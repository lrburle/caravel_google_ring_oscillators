magic
tech sky130A
magscale 1 2
timestamp 1696005323
<< error_p >>
rect 55 469 64 478
rect 102 469 111 478
rect 1319 469 1328 478
rect 1366 469 1375 478
rect 1711 469 1720 478
rect 1758 469 1767 478
rect 1911 469 1920 478
rect 1958 469 1967 478
rect 46 460 55 469
rect 111 460 120 469
rect 1310 460 1319 469
rect 1025 450 1031 456
rect 1071 450 1077 456
rect 1333 455 1345 463
rect 1355 455 1367 463
rect 1375 460 1384 469
rect 1434 463 1450 464
rect 1329 452 1331 455
rect 1369 452 1371 455
rect 1428 451 1439 463
rect 1702 460 1711 469
rect 1767 463 1776 469
rect 1708 457 1711 459
rect 1715 457 1721 463
rect 1761 460 1776 463
rect 1902 460 1911 469
rect 1967 462 1976 469
rect 1761 457 1767 460
rect 1019 444 1025 450
rect 1077 444 1083 450
rect 1310 443 1316 449
rect 1321 443 1329 451
rect 1332 449 1367 451
rect 1332 448 1333 449
rect 1365 448 1367 449
rect 47 438 55 442
rect 38 435 77 438
rect 1079 435 1118 440
rect 1304 437 1310 443
rect 1330 438 1332 447
rect 1333 443 1334 448
rect 1329 436 1330 438
rect 35 434 38 435
rect 47 434 55 435
rect 35 425 55 434
rect 57 425 69 434
rect 77 432 106 435
rect 106 426 110 432
rect 846 430 898 432
rect 1118 430 1132 435
rect 1328 432 1329 435
rect 793 428 898 430
rect 793 426 874 428
rect 110 425 111 426
rect 793 425 856 426
rect 31 423 35 425
rect 47 422 55 425
rect 759 423 789 425
rect 835 424 840 425
rect 23 410 31 422
rect 30 400 31 410
rect 35 419 69 422
rect 35 415 37 419
rect 35 408 36 415
rect 47 413 55 419
rect 66 417 69 419
rect 72 416 81 422
rect 34 406 36 408
rect 33 400 39 406
rect 44 400 47 413
rect 27 394 33 400
rect 30 388 31 394
rect 34 374 35 400
rect 67 394 69 416
rect 73 410 81 416
rect 111 413 120 422
rect 642 417 656 419
rect 668 417 759 423
rect 642 416 668 417
rect 642 415 656 416
rect 636 414 656 415
rect 677 414 682 417
rect 827 414 835 424
rect 874 417 891 426
rect 891 416 893 417
rect 79 400 85 406
rect 102 404 111 413
rect 627 409 651 414
rect 682 409 688 414
rect 826 413 827 414
rect 898 413 915 428
rect 1132 426 1142 430
rect 1327 428 1328 432
rect 1142 417 1164 426
rect 1325 424 1327 428
rect 1365 426 1369 448
rect 1371 439 1379 451
rect 1637 449 1649 457
rect 1698 453 1708 457
rect 1709 453 1715 457
rect 1673 449 1715 453
rect 1767 451 1773 457
rect 1920 456 1926 462
rect 1966 460 1976 462
rect 1929 456 1941 460
rect 1951 456 1963 460
rect 1966 456 1972 460
rect 1914 450 1920 456
rect 1972 450 1978 456
rect 1418 432 1428 448
rect 1449 446 1461 449
rect 1643 448 1649 449
rect 1695 448 1698 449
rect 1443 445 1463 446
rect 1637 445 1643 448
rect 1679 445 1709 448
rect 1443 443 1449 445
rect 1463 443 1493 445
rect 1440 437 1443 443
rect 1437 434 1443 437
rect 1495 436 1516 443
rect 1543 436 1549 442
rect 1164 416 1167 417
rect 85 394 91 400
rect 102 398 106 404
rect 614 401 627 409
rect 636 405 651 409
rect 100 386 101 391
rect 258 388 274 396
rect 441 388 457 401
rect 524 391 541 401
rect 600 393 614 401
rect 594 391 600 393
rect 541 390 594 391
rect 625 389 633 401
rect 637 399 642 401
rect 688 399 701 409
rect 258 386 315 388
rect 96 369 100 384
rect 258 380 303 386
rect 315 380 319 386
rect 34 356 41 369
rect 95 365 96 368
rect 94 361 95 364
rect 97 356 111 365
rect 242 364 258 380
rect 319 373 324 380
rect 506 364 512 370
rect 552 364 558 370
rect 625 368 633 379
rect 637 370 639 399
rect 887 396 889 413
rect 893 411 915 413
rect 893 401 901 411
rect 1019 398 1025 416
rect 1167 408 1188 416
rect 1322 414 1325 423
rect 1365 419 1367 426
rect 1356 417 1367 419
rect 1371 422 1379 429
rect 1371 417 1384 422
rect 1369 416 1370 417
rect 1370 413 1371 414
rect 1375 413 1384 417
rect 1418 414 1428 430
rect 1437 426 1440 434
rect 1491 430 1497 436
rect 1549 430 1555 436
rect 1625 433 1633 445
rect 1637 443 1671 445
rect 1637 442 1643 443
rect 1637 441 1640 442
rect 1437 425 1441 426
rect 1439 413 1441 425
rect 1077 407 1110 408
rect 1188 407 1190 408
rect 1112 405 1118 407
rect 1077 399 1083 404
rect 1118 403 1122 405
rect 1190 403 1200 407
rect 1320 403 1322 411
rect 1362 405 1375 413
rect 1437 410 1441 413
rect 1625 411 1633 423
rect 1637 414 1639 441
rect 1917 436 1920 448
rect 1972 444 1975 448
rect 1925 430 1929 444
rect 1972 433 1988 444
rect 1988 430 2004 433
rect 1714 419 1715 420
rect 1715 417 1716 418
rect 1637 413 1640 414
rect 1683 413 1711 414
rect 1637 411 1649 413
rect 1683 412 1709 413
rect 1367 404 1375 405
rect 1428 403 1432 408
rect 1437 403 1442 410
rect 1637 407 1641 411
rect 1683 410 1705 412
rect 1711 411 1715 413
rect 1683 408 1698 410
rect 1637 405 1643 407
rect 1683 406 1699 408
rect 1709 407 1715 411
rect 1718 409 1723 415
rect 1767 413 1776 422
rect 1902 413 1911 422
rect 1911 412 1917 413
rect 746 393 762 396
rect 764 393 780 396
rect 740 390 760 393
rect 881 391 893 396
rect 1017 391 1018 395
rect 1025 392 1031 398
rect 1035 395 1103 399
rect 1122 398 1134 403
rect 784 386 785 390
rect 742 384 834 386
rect 881 384 901 391
rect 1016 386 1017 391
rect 1035 389 1061 395
rect 1071 392 1077 395
rect 1103 389 1116 395
rect 1134 390 1155 398
rect 1200 390 1234 403
rect 1366 400 1367 402
rect 1304 391 1310 397
rect 1320 395 1321 399
rect 1363 397 1366 398
rect 1015 384 1016 386
rect 1053 384 1061 389
rect 646 375 742 384
rect 784 381 785 384
rect 743 375 755 377
rect 646 372 743 375
rect 637 369 641 370
rect 646 369 742 372
rect 637 368 646 369
rect 620 367 644 368
rect 648 367 671 368
rect 620 365 639 367
rect 688 366 703 369
rect 613 364 620 365
rect 633 364 634 365
rect 249 356 258 364
rect 500 358 506 364
rect 558 358 564 364
rect 594 361 613 364
rect 681 363 688 366
rect 637 362 648 363
rect 679 362 681 363
rect 572 358 594 361
rect 564 357 586 358
rect 27 348 33 354
rect 33 342 39 348
rect 41 346 66 356
rect 81 348 97 356
rect 79 346 97 348
rect 245 347 249 356
rect 637 355 649 362
rect 252 352 258 353
rect 252 351 294 352
rect 298 351 304 353
rect 252 348 263 351
rect 252 347 258 348
rect 294 347 304 351
rect 245 346 252 347
rect 72 341 75 346
rect 79 342 85 346
rect 68 335 72 341
rect 242 337 245 346
rect 246 341 252 346
rect 304 341 310 347
rect 311 345 323 353
rect 384 346 390 352
rect 430 346 436 352
rect 700 351 701 366
rect 730 364 740 369
rect 739 351 740 364
rect 785 364 796 380
rect 757 354 765 356
rect 747 352 757 354
rect 745 351 747 352
rect 325 344 327 345
rect 298 339 323 341
rect 63 326 68 335
rect 156 334 186 336
rect 236 334 242 337
rect 61 319 63 326
rect 29 307 30 317
rect 59 308 61 319
rect 132 318 156 334
rect 186 328 236 334
rect 321 327 323 339
rect 327 329 335 341
rect 372 338 384 346
rect 436 340 442 346
rect 558 338 561 342
rect 687 339 745 351
rect 785 350 789 364
rect 826 359 827 380
rect 834 377 906 384
rect 830 375 906 377
rect 834 368 906 375
rect 915 374 916 380
rect 909 368 916 374
rect 955 368 961 374
rect 1010 368 1015 384
rect 877 367 918 368
rect 903 362 918 367
rect 961 362 967 368
rect 792 354 838 356
rect 838 352 846 354
rect 846 351 849 352
rect 757 342 769 350
rect 779 342 791 350
rect 682 338 687 339
rect 441 334 443 336
rect 321 318 324 327
rect 360 322 368 334
rect 372 332 390 334
rect 372 328 374 332
rect 443 328 450 334
rect 58 303 59 307
rect 57 300 58 303
rect 57 283 58 287
rect 108 280 132 318
rect 321 309 323 318
rect 298 307 323 309
rect 327 307 335 319
rect 371 318 374 328
rect 450 326 453 328
rect 561 326 575 338
rect 668 335 682 338
rect 691 336 700 339
rect 789 338 791 342
rect 849 339 896 351
rect 909 347 918 362
rect 1008 361 1010 368
rect 1026 364 1035 380
rect 1044 367 1053 384
rect 1116 380 1133 389
rect 1155 380 1194 390
rect 1006 355 1008 361
rect 911 346 916 347
rect 961 345 967 348
rect 896 338 901 339
rect 909 338 911 345
rect 967 342 974 345
rect 984 342 996 350
rect 1004 349 1006 354
rect 1026 349 1035 362
rect 1040 355 1044 367
rect 1086 366 1115 376
rect 1133 375 1194 380
rect 1133 369 1155 375
rect 1194 372 1204 375
rect 1079 357 1115 366
rect 1126 364 1135 366
rect 1038 349 1040 354
rect 997 338 1004 349
rect 1026 346 1038 349
rect 1070 348 1079 357
rect 1086 356 1115 357
rect 1116 357 1135 364
rect 1155 362 1176 369
rect 1204 366 1219 372
rect 1234 368 1291 390
rect 1310 385 1316 391
rect 1321 389 1322 395
rect 1362 391 1368 397
rect 1322 384 1323 389
rect 1356 386 1362 391
rect 1363 386 1366 391
rect 1356 385 1363 386
rect 1362 384 1363 385
rect 1320 380 1323 384
rect 1371 383 1373 403
rect 1432 397 1438 403
rect 1443 400 1444 402
rect 1445 398 1448 399
rect 1448 397 1453 398
rect 1432 396 1488 397
rect 1637 396 1648 405
rect 1683 402 1695 406
rect 1709 405 1723 407
rect 1767 405 1773 411
rect 1911 410 1918 412
rect 1920 410 1929 430
rect 2004 413 2081 430
rect 2081 410 2091 413
rect 1711 404 1721 405
rect 1758 404 1767 405
rect 1911 404 1929 410
rect 1972 404 1978 410
rect 2091 404 2136 410
rect 2231 406 2249 407
rect 2219 404 2231 406
rect 1683 398 1701 402
rect 1715 399 1721 404
rect 1761 399 1767 404
rect 1920 403 1926 404
rect 1920 401 1927 403
rect 1928 402 1929 404
rect 1958 403 1961 404
rect 1920 398 1926 401
rect 1928 399 1932 400
rect 1947 399 1958 403
rect 1963 398 1972 404
rect 2091 400 2219 404
rect 1432 395 1497 396
rect 1641 395 1649 396
rect 1449 393 1497 395
rect 1449 391 1461 393
rect 1643 390 1659 395
rect 1664 393 1665 396
rect 1491 384 1497 390
rect 1549 384 1555 390
rect 1320 379 1325 380
rect 1361 379 1362 383
rect 1311 370 1325 379
rect 1291 367 1310 368
rect 1311 367 1323 370
rect 1219 363 1226 366
rect 1291 363 1323 367
rect 1325 363 1326 369
rect 1226 362 1228 363
rect 1116 356 1128 357
rect 1086 355 1093 356
rect 1135 355 1144 357
rect 1086 354 1091 355
rect 1086 353 1088 354
rect 1086 352 1132 353
rect 1133 352 1144 355
rect 1082 351 1087 352
rect 1094 351 1128 352
rect 1082 350 1128 351
rect 1082 349 1094 350
rect 1031 338 1038 346
rect 1081 343 1094 349
rect 1125 348 1128 350
rect 1132 349 1144 352
rect 1176 349 1278 362
rect 1291 361 1311 363
rect 1314 361 1330 362
rect 1303 360 1330 361
rect 1303 357 1311 360
rect 1314 355 1341 360
rect 1355 355 1361 379
rect 1373 363 1375 380
rect 1497 378 1503 384
rect 1506 379 1509 384
rect 1375 361 1380 362
rect 1368 355 1380 361
rect 1509 355 1518 379
rect 1543 378 1555 384
rect 1648 380 1659 390
rect 1683 392 1702 398
rect 1683 385 1720 392
rect 1844 388 1860 396
rect 1922 394 1925 398
rect 1921 388 1922 393
rect 1665 380 1669 384
rect 1549 357 1555 378
rect 1659 365 1671 380
rect 1687 377 1720 385
rect 1804 380 1807 388
rect 1845 387 1860 388
rect 1920 382 1921 387
rect 1963 381 1966 398
rect 1975 384 2076 389
rect 2076 381 2087 384
rect 2118 381 2219 400
rect 2249 392 2271 406
rect 1665 356 1669 365
rect 1671 363 1673 365
rect 1126 343 1128 348
rect 1139 343 1145 349
rect 1176 346 1310 349
rect 1314 346 1330 355
rect 1341 346 1405 355
rect 1673 354 1693 363
rect 1702 360 1720 377
rect 1800 369 1804 380
rect 1795 367 1800 369
rect 1757 362 1758 365
rect 1506 348 1588 354
rect 1489 346 1506 348
rect 1082 342 1094 343
rect 659 333 668 335
rect 647 332 659 333
rect 686 332 691 336
rect 600 327 686 332
rect 588 326 600 327
rect 628 326 647 327
rect 745 326 753 338
rect 757 336 791 338
rect 453 325 583 326
rect 561 321 575 325
rect 617 323 628 326
rect 610 319 616 323
rect 360 311 368 312
rect 370 311 371 318
rect 246 298 252 301
rect 294 298 323 307
rect 326 304 327 306
rect 360 300 370 311
rect 372 302 374 318
rect 500 312 506 318
rect 506 306 512 312
rect 534 304 547 312
rect 577 304 588 319
rect 602 312 607 316
rect 739 313 748 325
rect 757 313 759 336
rect 372 300 390 302
rect 534 301 543 304
rect 547 303 549 304
rect 589 301 591 303
rect 599 301 608 310
rect 748 304 759 313
rect 789 304 791 336
rect 795 326 803 338
rect 901 336 911 338
rect 968 336 996 338
rect 997 336 1008 338
rect 901 335 909 336
rect 906 333 909 335
rect 961 333 962 336
rect 994 333 1008 336
rect 827 319 841 333
rect 896 322 906 333
rect 960 329 961 333
rect 896 319 909 322
rect 959 319 960 328
rect 994 327 996 333
rect 997 327 1008 333
rect 1031 336 1039 338
rect 1031 327 1038 336
rect 1039 333 1043 336
rect 1042 330 1048 333
rect 1043 328 1048 330
rect 994 323 997 327
rect 999 326 1008 327
rect 999 324 1000 326
rect 841 318 896 319
rect 903 316 909 319
rect 958 316 959 318
rect 961 316 967 322
rect 994 318 996 323
rect 1000 319 1002 324
rect 1002 318 1003 319
rect 993 316 996 318
rect 1003 316 1004 318
rect 909 310 915 316
rect 951 314 954 316
rect 955 314 961 316
rect 950 310 961 314
rect 992 313 993 316
rect 950 304 957 310
rect 991 309 992 312
rect 989 306 991 307
rect 994 306 996 316
rect 962 304 996 306
rect 1000 313 1008 316
rect 1000 304 1014 313
rect 989 303 991 304
rect 1014 302 1017 304
rect 367 299 370 300
rect 173 282 294 298
rect 304 295 310 298
rect 311 295 323 298
rect 169 280 173 282
rect 260 280 262 282
rect 295 280 296 291
rect 298 289 304 295
rect 364 287 367 298
rect 368 296 370 299
rect 378 296 384 300
rect 372 294 384 296
rect 372 288 390 294
rect 403 291 406 300
rect 436 294 442 300
rect 402 287 403 291
rect 430 288 441 294
rect 543 292 552 301
rect 589 300 599 301
rect 987 300 989 301
rect 590 299 599 300
rect 590 292 610 299
rect 792 297 793 300
rect 753 294 754 296
rect 962 292 974 300
rect 984 294 996 300
rect 1017 296 1019 302
rect 1021 297 1031 327
rect 1048 324 1061 328
rect 1061 319 1073 324
rect 1076 318 1078 319
rect 1087 318 1094 342
rect 1139 340 1140 343
rect 1262 331 1310 346
rect 1330 344 1405 346
rect 1422 345 1473 346
rect 1475 345 1486 346
rect 1422 344 1483 345
rect 1330 342 1422 344
rect 1078 316 1083 318
rect 1087 316 1139 318
rect 1083 311 1139 316
rect 1070 301 1079 310
rect 1087 308 1156 311
rect 1087 303 1144 308
rect 1156 304 1181 308
rect 1278 306 1286 331
rect 1310 328 1317 331
rect 1330 330 1346 342
rect 1348 330 1364 342
rect 1469 341 1484 344
rect 1465 339 1469 341
rect 1449 334 1465 339
rect 1475 338 1484 341
rect 1518 338 1525 348
rect 1478 332 1483 334
rect 1296 312 1300 328
rect 1317 326 1348 328
rect 1349 326 1351 330
rect 1317 321 1349 326
rect 1340 319 1357 321
rect 1340 314 1349 319
rect 1357 318 1361 319
rect 1300 308 1301 311
rect 1320 310 1340 314
rect 1081 301 1145 303
rect 1181 302 1193 304
rect 1277 302 1278 305
rect 1079 297 1145 301
rect 982 292 996 294
rect 360 282 364 287
rect 359 281 360 282
rect 400 281 402 287
rect 354 280 359 281
rect 89 274 108 280
rect 160 274 169 280
rect 85 268 89 274
rect 153 269 160 274
rect 152 268 153 269
rect 83 253 85 268
rect 149 261 152 268
rect 151 250 160 254
rect 198 250 207 254
rect 210 250 226 266
rect 228 250 244 266
rect 262 250 266 279
rect 293 259 295 279
rect 340 276 354 280
rect 396 276 397 279
rect 399 276 400 281
rect 436 279 441 288
rect 553 287 556 292
rect 597 291 610 292
rect 337 274 340 276
rect 331 269 337 274
rect 330 268 331 269
rect 320 266 330 268
rect 306 261 330 266
rect 306 250 320 261
rect 393 250 399 276
rect 441 263 446 279
rect 556 272 563 287
rect 595 285 610 287
rect 446 259 451 263
rect 451 257 466 259
rect 79 216 83 250
rect 148 245 160 250
rect 194 245 210 250
rect 244 249 260 250
rect 251 246 260 249
rect 142 244 155 245
rect 194 244 216 245
rect 140 243 149 244
rect 140 223 142 243
rect 143 238 149 243
rect 139 222 142 223
rect 140 216 142 222
rect 148 232 149 238
rect 186 236 216 244
rect 186 234 210 236
rect 255 235 260 246
rect 290 244 306 250
rect 388 245 393 249
rect 395 245 397 250
rect 436 249 448 257
rect 458 253 471 257
rect 458 249 470 253
rect 471 250 472 253
rect 506 250 522 266
rect 524 250 540 266
rect 563 254 572 272
rect 564 253 572 254
rect 576 257 577 274
rect 576 255 580 257
rect 608 256 610 285
rect 611 281 622 287
rect 614 276 622 281
rect 614 275 627 276
rect 618 266 627 275
rect 754 272 758 291
rect 791 278 792 292
rect 873 279 879 285
rect 919 279 925 285
rect 958 280 959 281
rect 982 279 987 292
rect 1006 281 1021 296
rect 1079 292 1098 297
rect 867 273 873 279
rect 925 273 931 279
rect 980 272 982 279
rect 1006 278 1022 281
rect 618 265 636 266
rect 607 255 610 256
rect 576 253 610 255
rect 614 262 636 265
rect 678 265 736 270
rect 678 264 688 265
rect 736 264 737 265
rect 758 264 759 270
rect 792 266 793 270
rect 737 262 740 264
rect 614 253 622 262
rect 627 252 636 262
rect 472 249 479 250
rect 490 249 503 250
rect 429 245 432 247
rect 436 245 495 249
rect 386 244 395 245
rect 424 244 429 245
rect 265 235 266 240
rect 290 237 428 244
rect 436 243 470 245
rect 276 235 306 237
rect 386 236 395 237
rect 255 234 276 235
rect 290 234 306 235
rect 186 233 201 234
rect 238 233 259 234
rect 209 232 229 233
rect 148 216 164 232
rect 194 216 210 232
rect 220 227 244 229
rect 254 224 255 229
rect 83 211 102 216
rect 113 211 148 216
rect 83 209 113 211
rect 132 200 149 211
rect 210 209 213 215
rect 210 200 220 209
rect 140 198 149 200
rect 213 198 222 200
rect 265 199 266 234
rect 293 232 298 234
rect 290 216 306 232
rect 388 230 393 236
rect 387 225 388 229
rect 385 224 387 225
rect 381 221 385 224
rect 378 217 381 221
rect 342 216 378 217
rect 293 201 298 216
rect 306 215 342 216
rect 306 205 322 215
rect 324 205 340 215
rect 419 213 429 214
rect 468 213 470 243
rect 472 236 482 245
rect 540 236 556 250
rect 610 249 614 252
rect 634 250 636 252
rect 658 250 664 256
rect 704 251 710 256
rect 700 250 712 251
rect 759 250 762 262
rect 794 253 810 266
rect 865 264 873 270
rect 863 262 873 264
rect 977 263 980 272
rect 926 260 936 262
rect 936 258 942 260
rect 975 259 977 263
rect 853 256 867 258
rect 942 256 949 258
rect 793 252 810 253
rect 793 250 797 252
rect 576 241 588 249
rect 598 241 610 249
rect 636 244 716 250
rect 740 244 748 250
rect 762 244 763 249
rect 576 240 577 241
rect 474 233 572 236
rect 479 225 572 233
rect 577 230 579 240
rect 636 236 652 244
rect 658 243 712 244
rect 658 239 710 243
rect 653 236 657 237
rect 579 226 581 230
rect 602 225 653 236
rect 396 211 419 213
rect 424 211 432 213
rect 384 210 396 211
rect 361 207 384 210
rect 432 207 434 210
rect 342 205 361 207
rect 303 201 342 205
rect 436 203 470 213
rect 474 211 482 223
rect 540 216 556 225
rect 572 224 600 225
rect 581 221 582 224
rect 582 217 583 221
rect 539 215 540 216
rect 538 211 540 215
rect 583 211 584 215
rect 472 207 474 210
rect 533 203 540 211
rect 584 204 586 211
rect 658 205 678 239
rect 704 237 712 239
rect 710 207 712 237
rect 716 227 724 239
rect 739 234 748 244
rect 739 231 740 234
rect 739 221 748 231
rect 763 226 766 241
rect 778 234 797 250
rect 831 245 840 254
rect 853 253 873 256
rect 949 255 953 256
rect 953 254 958 255
rect 974 254 975 256
rect 970 253 981 254
rect 1006 253 1021 278
rect 1022 266 1025 277
rect 1087 272 1098 292
rect 1129 292 1139 297
rect 1129 272 1130 292
rect 1133 291 1139 292
rect 1193 291 1260 302
rect 1275 293 1277 301
rect 1301 293 1305 308
rect 1315 303 1320 310
rect 1361 304 1418 318
rect 1418 303 1421 304
rect 1312 293 1314 301
rect 1421 300 1435 303
rect 1481 302 1483 332
rect 1487 322 1495 334
rect 1525 314 1535 338
rect 1555 322 1562 348
rect 1588 346 1592 348
rect 1669 347 1670 354
rect 1592 345 1593 346
rect 1593 339 1596 345
rect 1596 334 1599 339
rect 1599 331 1601 334
rect 1601 328 1602 331
rect 1452 300 1483 302
rect 1487 300 1495 312
rect 1535 311 1536 314
rect 1562 312 1564 322
rect 1602 314 1609 328
rect 1670 322 1674 347
rect 1693 346 1709 354
rect 1720 347 1721 354
rect 1707 345 1713 346
rect 1707 344 1715 345
rect 1721 344 1722 347
rect 1757 346 1772 362
rect 1795 360 1807 367
rect 1794 359 1807 360
rect 1817 359 1829 367
rect 1860 364 1876 380
rect 1791 357 1800 359
rect 1790 355 1791 357
rect 1794 355 1800 357
rect 1833 355 1834 357
rect 1840 355 1846 360
rect 1783 354 1790 355
rect 1794 354 1829 355
rect 1833 354 1846 355
rect 1783 349 1794 354
rect 1795 353 1829 354
rect 1777 344 1787 349
rect 1788 348 1794 349
rect 1828 348 1829 353
rect 1846 348 1852 354
rect 1860 346 1876 362
rect 1912 346 1920 380
rect 1966 368 1967 380
rect 1971 377 1972 381
rect 2087 380 2106 381
rect 2114 380 2118 381
rect 2078 376 2114 380
rect 2164 377 2168 381
rect 1715 343 1756 344
rect 1721 330 1738 343
rect 1740 338 1756 343
rect 1774 342 1777 344
rect 1767 338 1774 342
rect 1859 339 1860 343
rect 1740 330 1767 338
rect 1858 332 1860 339
rect 1910 334 1912 344
rect 1921 334 1929 346
rect 1933 334 1935 368
rect 1971 363 1972 376
rect 2078 372 2126 376
rect 2069 366 2078 372
rect 1966 360 1967 363
rect 1972 348 1973 360
rect 2058 348 2069 366
rect 2107 361 2126 372
rect 2126 360 2128 361
rect 2168 360 2173 377
rect 2271 373 2274 392
rect 2274 366 2275 372
rect 2053 346 2069 348
rect 1973 340 1979 346
rect 1974 334 1979 340
rect 2053 340 2065 346
rect 2075 340 2087 348
rect 2128 346 2147 360
rect 2173 346 2178 360
rect 2275 346 2278 366
rect 2147 344 2148 346
rect 2148 340 2149 342
rect 2178 341 2180 346
rect 2053 336 2058 340
rect 2091 338 2092 340
rect 2093 336 2096 337
rect 1857 331 1860 332
rect 1721 317 1722 330
rect 1749 328 1767 330
rect 1856 330 1860 331
rect 1856 328 1857 330
rect 1909 328 1910 331
rect 1929 328 1930 333
rect 1743 324 1749 328
rect 1852 321 1856 328
rect 1908 321 1909 328
rect 1930 324 1932 328
rect 1960 325 1967 334
rect 1974 328 1975 334
rect 1953 323 1960 325
rect 1971 323 1975 328
rect 2041 324 2049 336
rect 2053 334 2087 336
rect 2053 333 2056 334
rect 1933 322 1971 323
rect 1722 314 1723 316
rect 1609 311 1611 314
rect 1564 306 1565 311
rect 1611 308 1612 311
rect 1435 297 1446 300
rect 1449 297 1488 300
rect 1446 296 1488 297
rect 1261 284 1268 291
rect 1269 281 1275 293
rect 1268 277 1275 281
rect 1269 272 1275 277
rect 1299 278 1312 293
rect 1449 291 1488 296
rect 1537 293 1539 301
rect 1471 288 1483 291
rect 1488 286 1510 291
rect 1524 284 1529 286
rect 1539 284 1546 293
rect 1529 278 1546 284
rect 1098 266 1099 272
rect 1268 266 1271 272
rect 1022 264 1028 266
rect 1025 253 1028 264
rect 1090 261 1106 266
rect 1089 260 1103 261
rect 1108 260 1124 266
rect 1081 253 1089 260
rect 1103 254 1126 260
rect 853 250 867 253
rect 973 251 974 253
rect 981 252 1021 253
rect 1027 252 1028 253
rect 1079 252 1081 253
rect 1006 251 1054 252
rect 1077 250 1079 252
rect 1093 251 1105 254
rect 1186 253 1202 266
rect 1204 253 1220 266
rect 1266 259 1268 265
rect 1269 264 1271 266
rect 1299 264 1317 278
rect 1539 275 1555 278
rect 1502 264 1516 266
rect 1126 252 1127 253
rect 1179 252 1180 253
rect 1098 250 1105 251
rect 847 246 861 250
rect 847 245 858 246
rect 822 236 831 245
rect 793 232 797 234
rect 778 226 797 232
rect 766 221 767 224
rect 704 206 712 207
rect 716 206 724 217
rect 738 216 748 221
rect 767 211 769 220
rect 778 216 794 226
rect 853 224 861 236
rect 865 226 867 250
rect 970 244 973 250
rect 925 227 931 233
rect 959 230 977 244
rect 919 226 925 227
rect 964 226 966 230
rect 865 224 899 226
rect 908 224 967 226
rect 977 225 983 230
rect 978 224 984 225
rect 797 220 798 224
rect 889 223 899 224
rect 888 221 899 223
rect 903 222 908 224
rect 880 220 898 221
rect 900 220 903 222
rect 919 221 925 224
rect 798 216 799 220
rect 865 217 877 220
rect 880 217 899 220
rect 865 216 878 217
rect 734 206 738 211
rect 794 206 802 216
rect 825 212 877 216
rect 887 212 899 217
rect 704 205 734 206
rect 794 205 804 206
rect 658 204 710 205
rect 716 204 732 205
rect 794 204 806 205
rect 280 199 303 201
rect 306 200 322 201
rect 324 200 340 201
rect 436 199 448 203
rect 458 201 523 203
rect 532 201 540 203
rect 586 201 592 204
rect 458 200 540 201
rect 458 199 532 200
rect 29 167 30 195
rect 58 184 59 195
rect 142 192 149 198
rect 207 197 223 198
rect 264 197 280 199
rect 207 195 254 197
rect 258 195 266 197
rect 201 194 229 195
rect 258 194 264 195
rect 186 192 229 194
rect 142 189 155 192
rect 195 189 201 192
rect 207 191 229 192
rect 256 191 258 194
rect 207 189 216 191
rect 149 186 188 189
rect 195 186 207 189
rect 59 171 67 184
rect 151 180 188 186
rect 198 180 207 186
rect 242 183 254 191
rect 264 180 265 189
rect 59 167 70 171
rect 30 161 31 167
rect 67 165 70 167
rect 68 162 73 165
rect 42 159 71 160
rect 74 159 75 161
rect 24 125 31 137
rect 36 128 37 159
rect 65 157 70 159
rect 69 128 70 157
rect 71 150 82 159
rect 298 152 302 194
rect 386 189 395 198
rect 470 196 532 199
rect 592 196 599 201
rect 652 200 732 204
rect 770 202 771 204
rect 794 201 815 204
rect 794 200 809 201
rect 630 198 716 200
rect 804 198 809 200
rect 815 199 820 201
rect 820 198 824 199
rect 825 198 876 212
rect 888 205 898 212
rect 950 205 964 223
rect 967 222 975 224
rect 978 222 989 224
rect 997 223 1006 250
rect 1028 234 1044 250
rect 1068 244 1076 250
rect 975 220 997 222
rect 1028 220 1044 232
rect 1097 223 1099 250
rect 1100 249 1105 250
rect 1102 248 1105 249
rect 1127 250 1128 252
rect 1177 250 1179 252
rect 1103 246 1107 248
rect 1108 244 1109 246
rect 1127 244 1140 250
rect 1101 240 1105 242
rect 978 216 1044 220
rect 982 212 1028 216
rect 1068 213 1069 216
rect 887 202 888 205
rect 948 202 950 205
rect 599 195 600 196
rect 601 195 634 198
rect 635 195 636 197
rect 451 194 590 195
rect 451 189 460 194
rect 601 191 607 195
rect 632 191 635 195
rect 658 192 664 198
rect 700 193 712 198
rect 820 197 831 198
rect 822 195 831 197
rect 822 194 834 195
rect 704 192 710 193
rect 770 191 771 193
rect 607 189 612 191
rect 631 189 632 191
rect 395 180 404 189
rect 442 180 451 189
rect 607 188 631 189
rect 767 184 770 191
rect 822 189 831 194
rect 837 191 840 193
rect 840 189 859 191
rect 887 189 896 198
rect 918 194 924 200
rect 945 198 948 202
rect 982 200 1010 212
rect 1012 207 1053 212
rect 1069 210 1071 213
rect 1095 210 1097 222
rect 1103 210 1105 240
rect 1109 230 1117 242
rect 1126 234 1140 244
rect 1170 248 1179 250
rect 1232 249 1236 253
rect 1264 251 1266 259
rect 1299 250 1312 264
rect 1317 260 1320 264
rect 1447 254 1453 256
rect 1447 250 1461 254
rect 1493 250 1499 256
rect 1500 250 1516 264
rect 1539 250 1546 275
rect 1555 265 1558 275
rect 1558 250 1563 264
rect 1565 250 1581 302
rect 1612 300 1616 308
rect 1720 302 1723 308
rect 1729 303 1740 320
rect 1795 315 1807 321
rect 1907 320 1908 321
rect 1836 315 1852 320
rect 1906 315 1907 320
rect 1953 315 1960 322
rect 1807 314 1836 315
rect 1905 308 1906 311
rect 1788 302 1794 308
rect 1846 302 1852 308
rect 1616 286 1624 300
rect 1718 297 1720 301
rect 1726 298 1729 302
rect 1624 275 1629 286
rect 1629 271 1631 275
rect 1655 266 1674 297
rect 1701 293 1718 297
rect 1794 296 1800 302
rect 1804 299 1805 302
rect 1814 298 1821 302
rect 1701 286 1724 293
rect 1689 278 1718 286
rect 1687 275 1689 278
rect 1685 271 1687 275
rect 1701 271 1718 278
rect 1683 268 1685 271
rect 1681 266 1683 268
rect 1655 263 1683 266
rect 1655 251 1681 263
rect 1655 250 1675 251
rect 1170 234 1177 248
rect 1194 238 1206 244
rect 1191 237 1250 238
rect 1251 237 1264 250
rect 1191 235 1199 237
rect 1250 235 1264 237
rect 1271 235 1274 250
rect 1126 232 1129 234
rect 1190 233 1191 235
rect 1069 208 1105 210
rect 1109 208 1117 220
rect 1126 216 1140 232
rect 1182 228 1190 232
rect 1194 230 1201 232
rect 1182 220 1188 228
rect 1194 226 1195 230
rect 1251 228 1279 235
rect 1286 228 1299 249
rect 1320 234 1332 250
rect 1441 244 1447 250
rect 1445 242 1447 244
rect 1449 242 1482 250
rect 1499 244 1505 250
rect 1516 244 1532 250
rect 1546 244 1547 250
rect 1499 242 1532 244
rect 1563 242 1581 250
rect 1631 242 1632 250
rect 1655 242 1674 250
rect 1688 242 1701 271
rect 1718 258 1725 270
rect 1730 260 1731 292
rect 1797 288 1803 291
rect 1794 286 1797 288
rect 1785 281 1794 286
rect 1778 272 1779 275
rect 1805 272 1810 297
rect 1811 296 1813 297
rect 1840 296 1864 302
rect 1903 300 1905 308
rect 1773 260 1778 272
rect 1730 259 1735 260
rect 1730 258 1764 259
rect 1771 258 1776 260
rect 1725 256 1726 258
rect 1770 256 1771 258
rect 1767 254 1769 255
rect 1730 246 1742 253
rect 1752 246 1764 253
rect 1810 242 1821 271
rect 1842 250 1864 296
rect 1901 286 1903 300
rect 1898 275 1901 286
rect 1897 268 1898 271
rect 1935 268 1953 315
rect 2041 302 2049 314
rect 2053 302 2055 333
rect 2086 332 2087 334
rect 2093 324 2099 336
rect 2149 325 2151 337
rect 2180 336 2196 340
rect 2266 337 2275 346
rect 2258 336 2266 337
rect 2180 325 2258 336
rect 2093 323 2096 324
rect 2096 315 2101 322
rect 2134 317 2196 325
rect 2128 315 2134 317
rect 2087 302 2128 315
rect 2096 300 2101 302
rect 2151 301 2153 317
rect 2049 298 2052 300
rect 2101 298 2102 300
rect 2153 297 2154 300
rect 2052 296 2054 297
rect 2053 295 2055 296
rect 2053 291 2056 295
rect 2102 292 2103 294
rect 2053 290 2057 291
rect 2056 288 2057 290
rect 2103 288 2104 292
rect 2154 288 2155 291
rect 2180 290 2196 317
rect 2057 281 2060 286
rect 1995 273 1996 274
rect 1874 263 1890 266
rect 1894 263 1897 268
rect 1933 263 1935 268
rect 1976 266 1988 267
rect 1874 255 1894 263
rect 1930 255 1933 263
rect 1970 261 1988 266
rect 1998 261 2010 267
rect 2060 261 2067 281
rect 2086 261 2100 266
rect 1970 260 2067 261
rect 1970 255 2061 260
rect 2067 256 2068 259
rect 2084 255 2100 261
rect 1872 251 1875 255
rect 1928 251 1930 255
rect 1964 254 2010 255
rect 1964 252 1968 254
rect 1970 253 2010 254
rect 1957 251 1967 252
rect 1970 251 1976 253
rect 1951 250 1956 251
rect 1970 250 1971 251
rect 1842 242 1872 250
rect 1925 248 1928 250
rect 1947 249 1951 250
rect 1938 248 1944 249
rect 1925 246 1938 248
rect 1915 245 1919 246
rect 1909 244 1915 245
rect 1896 242 1909 244
rect 1925 243 1928 246
rect 1437 239 1445 242
rect 1449 240 1452 242
rect 1436 233 1446 239
rect 1125 214 1126 216
rect 1012 200 1028 207
rect 1053 205 1064 207
rect 1071 206 1078 208
rect 1078 205 1084 206
rect 1095 205 1097 208
rect 1064 204 1069 205
rect 1084 204 1104 205
rect 1107 204 1109 207
rect 1124 206 1125 208
rect 964 194 970 200
rect 982 198 997 200
rect 1084 198 1105 204
rect 1121 201 1124 205
rect 1127 202 1129 216
rect 1106 200 1124 201
rect 1106 198 1121 200
rect 1177 198 1178 200
rect 1182 198 1188 210
rect 1236 201 1237 213
rect 1251 202 1264 228
rect 1266 224 1274 228
rect 1266 216 1275 224
rect 1279 219 1311 228
rect 1320 219 1332 232
rect 1412 219 1436 233
rect 1437 230 1445 233
rect 1275 213 1276 215
rect 1286 213 1299 219
rect 1311 216 1332 219
rect 1276 209 1304 213
rect 1311 209 1330 216
rect 1398 211 1412 219
rect 1276 208 1330 209
rect 1391 208 1398 211
rect 1437 208 1445 220
rect 1449 208 1451 240
rect 1517 234 1746 242
rect 1517 232 1519 234
rect 1520 232 1746 234
rect 1517 226 1746 232
rect 1774 226 1896 242
rect 1919 230 1925 243
rect 1954 234 1970 250
rect 1917 227 1924 230
rect 1517 224 1774 226
rect 1519 216 1532 224
rect 1549 219 1551 224
rect 1519 215 1520 216
rect 1520 213 1521 214
rect 1517 208 1520 213
rect 1550 211 1551 219
rect 1562 216 1574 224
rect 1574 215 1575 216
rect 1579 215 1581 220
rect 1598 215 1677 224
rect 1575 214 1677 215
rect 1578 211 1594 214
rect 1195 199 1197 200
rect 1194 198 1200 199
rect 976 194 982 198
rect 1093 196 1105 198
rect 831 184 859 189
rect 760 171 767 184
rect 831 180 840 184
rect 878 180 887 189
rect 912 188 918 194
rect 970 188 982 194
rect 1094 188 1095 193
rect 970 178 974 185
rect 1126 184 1127 198
rect 1178 195 1179 198
rect 1189 196 1191 197
rect 1235 196 1236 200
rect 1250 199 1251 202
rect 1276 201 1320 208
rect 1330 207 1332 208
rect 1332 204 1339 207
rect 1389 205 1391 208
rect 1488 207 1516 208
rect 1339 201 1343 204
rect 1276 200 1298 201
rect 1300 200 1316 201
rect 1343 200 1345 201
rect 1385 200 1389 205
rect 1502 204 1516 207
rect 1546 205 1550 211
rect 1257 199 1264 200
rect 1272 199 1286 200
rect 1345 199 1348 200
rect 1249 198 1257 199
rect 1244 197 1257 198
rect 1276 197 1286 199
rect 1441 198 1447 204
rect 1499 203 1516 204
rect 1543 203 1546 205
rect 1499 201 1555 203
rect 1576 201 1594 211
rect 1596 208 1677 214
rect 1688 212 1701 224
rect 1764 216 1765 219
rect 1499 200 1516 201
rect 1543 200 1546 201
rect 1555 200 1594 201
rect 1598 200 1677 208
rect 1499 198 1505 200
rect 1241 196 1250 197
rect 1179 192 1191 195
rect 1194 192 1195 193
rect 1203 192 1241 196
rect 1179 191 1238 192
rect 1194 186 1206 191
rect 1125 175 1127 184
rect 1244 175 1250 196
rect 1276 196 1290 197
rect 750 168 767 171
rect 1091 168 1094 175
rect 750 166 760 168
rect 1090 166 1091 168
rect 750 165 754 166
rect 739 161 781 165
rect 739 160 766 161
rect 737 159 739 160
rect 781 159 784 161
rect 723 157 737 159
rect 255 150 261 152
rect 298 151 307 152
rect 75 147 93 150
rect 82 137 93 147
rect 255 146 267 150
rect 301 146 307 151
rect 690 150 723 157
rect 684 149 689 150
rect 249 140 255 146
rect 307 141 313 146
rect 661 145 684 149
rect 738 147 746 159
rect 750 158 755 159
rect 655 143 661 145
rect 271 140 402 141
rect 255 138 271 140
rect 307 139 610 140
rect 637 139 643 141
rect 402 138 403 139
rect 610 138 643 139
rect 646 138 651 143
rect 36 126 40 128
rect 67 126 70 128
rect 36 125 70 126
rect 75 125 93 137
rect 243 126 251 138
rect 255 136 261 138
rect 31 123 32 125
rect 32 120 37 123
rect 70 120 75 123
rect 36 119 48 120
rect 35 113 48 119
rect 58 113 70 120
rect 82 119 93 125
rect 35 106 37 113
rect 93 102 100 119
rect 243 104 251 116
rect 255 106 257 136
rect 404 131 408 138
rect 610 135 645 138
rect 683 135 689 141
rect 408 120 415 131
rect 631 129 637 135
rect 638 131 645 135
rect 689 131 695 135
rect 738 131 746 137
rect 750 131 752 158
rect 1079 156 1085 162
rect 1087 156 1090 166
rect 1125 162 1126 175
rect 1231 169 1237 174
rect 1243 169 1244 174
rect 1276 170 1286 196
rect 1290 195 1294 196
rect 1349 195 1355 198
rect 1384 195 1385 198
rect 1447 196 1461 198
rect 1447 195 1453 196
rect 1485 195 1489 196
rect 1356 193 1358 194
rect 1358 192 1361 193
rect 1374 192 1384 195
rect 1303 187 1309 191
rect 1309 184 1314 187
rect 1361 184 1384 192
rect 1315 178 1339 184
rect 1374 181 1406 184
rect 1412 181 1485 195
rect 1493 192 1499 198
rect 1500 196 1501 197
rect 1541 196 1543 200
rect 1576 195 1579 200
rect 1585 199 1677 200
rect 1649 198 1677 199
rect 1626 197 1677 198
rect 1685 197 1688 211
rect 1763 209 1764 213
rect 1810 212 1821 226
rect 1842 216 1874 226
rect 1911 219 1924 227
rect 1908 217 1924 219
rect 1954 217 1970 232
rect 2008 223 2010 253
rect 2014 243 2022 255
rect 2061 250 2101 255
rect 2104 254 2111 286
rect 2146 252 2154 264
rect 2158 254 2160 286
rect 2190 269 2195 286
rect 2190 254 2192 269
rect 2195 264 2196 268
rect 2158 252 2192 254
rect 2196 252 2204 264
rect 2111 250 2112 252
rect 2198 250 2200 252
rect 2101 249 2116 250
rect 2158 249 2159 250
rect 2110 248 2116 249
rect 2155 248 2157 249
rect 1992 221 2010 223
rect 2014 221 2022 233
rect 2071 217 2081 248
rect 2110 244 2125 248
rect 2113 220 2125 244
rect 2158 240 2170 248
rect 2180 240 2192 248
rect 2198 240 2212 250
rect 2159 232 2161 240
rect 2112 219 2125 220
rect 1897 216 2010 217
rect 1762 203 1763 208
rect 1761 200 1762 203
rect 1821 201 1824 211
rect 1842 206 1864 216
rect 1874 215 2010 216
rect 1874 207 1890 215
rect 1892 211 2010 215
rect 2081 213 2085 217
rect 2111 216 2125 219
rect 2146 227 2161 232
rect 2200 234 2212 240
rect 2200 232 2202 234
rect 2146 216 2162 227
rect 2200 217 2212 232
rect 2202 216 2212 217
rect 2110 215 2111 216
rect 2109 213 2110 214
rect 2057 211 2100 213
rect 1892 208 2057 211
rect 2081 208 2100 211
rect 1894 207 1998 208
rect 2081 207 2085 208
rect 1874 206 1908 207
rect 1842 204 1890 206
rect 1835 201 1864 204
rect 1750 197 1761 200
rect 1810 199 1835 201
rect 1797 198 1810 199
rect 1793 197 1797 198
rect 1652 196 1655 197
rect 1673 196 1761 197
rect 1673 195 1750 196
rect 1766 195 1793 197
rect 1821 196 1824 199
rect 1495 191 1496 192
rect 1533 181 1541 195
rect 1575 190 1576 195
rect 1651 193 1652 195
rect 1674 194 1676 195
rect 1650 190 1651 193
rect 1676 192 1679 194
rect 1684 193 1685 195
rect 1742 194 1766 195
rect 1731 191 1742 194
rect 1679 190 1682 191
rect 1231 168 1249 169
rect 1277 168 1283 170
rect 1225 162 1289 168
rect 1314 165 1344 178
rect 1374 175 1412 181
rect 1530 175 1533 181
rect 1374 171 1406 175
rect 1314 162 1350 165
rect 1371 164 1374 170
rect 1375 167 1406 171
rect 1403 166 1405 167
rect 1406 166 1409 167
rect 1525 166 1530 175
rect 1402 164 1403 166
rect 1409 163 1414 166
rect 1524 164 1525 166
rect 1125 156 1131 162
rect 1231 157 1283 162
rect 1035 154 1079 156
rect 884 153 918 154
rect 1035 153 1041 154
rect 847 152 884 153
rect 824 151 847 152
rect 821 149 824 151
rect 1073 150 1079 154
rect 1131 150 1137 156
rect 796 135 821 149
rect 912 142 918 148
rect 970 143 976 148
rect 1225 145 1237 157
rect 1271 147 1276 157
rect 1001 143 1037 145
rect 918 136 924 142
rect 942 141 1001 143
rect 1037 141 1043 143
rect 940 138 942 141
rect 791 132 796 135
rect 689 129 771 131
rect 692 128 771 129
rect 788 128 796 132
rect 738 125 746 128
rect 750 127 752 128
rect 771 127 800 128
rect 750 125 784 127
rect 781 121 784 125
rect 788 125 796 127
rect 800 126 828 127
rect 788 123 791 125
rect 785 121 788 123
rect 828 122 842 126
rect 934 125 940 138
rect 964 136 970 141
rect 1043 138 1054 141
rect 1231 138 1237 145
rect 1033 134 1035 135
rect 1054 134 1065 138
rect 1230 135 1237 138
rect 1065 133 1067 134
rect 1067 132 1071 133
rect 415 119 416 120
rect 637 119 638 120
rect 750 113 762 121
rect 772 113 784 121
rect 842 117 848 122
rect 932 120 934 125
rect 931 119 932 120
rect 848 115 859 117
rect 476 109 610 112
rect 776 110 780 113
rect 859 111 872 115
rect 872 110 877 111
rect 352 107 476 109
rect 610 107 616 109
rect 255 104 261 106
rect 330 104 352 107
rect 37 100 38 102
rect 251 100 253 103
rect 254 100 255 102
rect 307 101 330 104
rect 616 101 628 107
rect 760 102 776 110
rect 877 106 893 110
rect 893 104 909 106
rect 909 103 918 104
rect 924 103 931 118
rect 628 100 631 101
rect 635 100 637 102
rect 38 81 48 100
rect 249 94 255 100
rect 307 94 313 100
rect 631 98 637 100
rect 254 92 267 94
rect 254 88 261 92
rect 301 88 307 94
rect 635 89 637 98
rect 737 93 760 102
rect 918 101 940 103
rect 737 91 807 93
rect 48 70 58 81
rect 50 68 64 70
rect 100 68 116 84
rect 254 80 255 88
rect 631 83 637 89
rect 689 90 760 91
rect 689 88 753 90
rect 807 88 816 91
rect 689 83 695 88
rect 254 68 266 80
rect 634 77 643 83
rect 683 77 689 83
rect 634 74 637 77
rect 718 74 737 88
rect 816 87 820 88
rect 820 84 822 87
rect 824 79 825 81
rect 634 70 636 74
rect 714 71 718 74
rect 825 72 840 79
rect 924 74 930 101
rect 940 98 975 101
rect 1025 98 1033 110
rect 1037 98 1039 132
rect 1225 123 1237 135
rect 1276 123 1278 138
rect 1314 135 1344 162
rect 1370 161 1371 163
rect 1414 162 1416 163
rect 1354 158 1356 159
rect 1368 157 1370 161
rect 1357 149 1371 157
rect 1399 156 1401 161
rect 1419 159 1422 161
rect 1422 158 1424 159
rect 1424 155 1428 158
rect 1448 155 1460 161
rect 1519 156 1522 161
rect 1554 156 1575 190
rect 1641 168 1650 190
rect 1679 188 1684 190
rect 1685 188 1731 191
rect 1824 190 1825 193
rect 1679 187 1731 188
rect 1679 168 1684 187
rect 1825 184 1829 190
rect 1825 168 1832 184
rect 1842 168 1864 201
rect 1874 200 1890 204
rect 1894 200 1908 206
rect 1970 200 1986 207
rect 2086 206 2100 208
rect 2085 204 2100 206
rect 2086 200 2100 204
rect 2087 199 2088 200
rect 2088 195 2089 197
rect 2090 184 2093 191
rect 2113 190 2125 216
rect 2162 211 2163 214
rect 2162 208 2164 211
rect 2200 208 2202 212
rect 2162 203 2170 208
rect 2197 203 2200 208
rect 2162 200 2178 203
rect 2180 200 2196 203
rect 1636 157 1641 168
rect 1676 156 1679 168
rect 1829 162 1832 168
rect 1829 156 1836 162
rect 1864 156 1866 168
rect 1894 163 1906 171
rect 1916 163 1928 171
rect 2093 167 2098 184
rect 2125 182 2129 190
rect 1876 159 1882 162
rect 1930 161 1932 162
rect 1883 159 1889 161
rect 1876 158 1889 159
rect 1875 156 1883 158
rect 1894 157 1930 159
rect 1932 157 1940 159
rect 1364 146 1365 149
rect 1371 146 1375 149
rect 1363 144 1364 146
rect 1375 144 1379 146
rect 1360 137 1363 143
rect 1379 141 1383 144
rect 1393 141 1399 155
rect 1428 153 1460 155
rect 1456 152 1461 153
rect 1463 149 1466 151
rect 1516 150 1519 156
rect 1550 149 1554 156
rect 1425 148 1426 149
rect 1455 146 1465 149
rect 1466 146 1472 149
rect 1478 146 1484 149
rect 1460 144 1465 146
rect 1355 123 1360 136
rect 1383 124 1411 141
rect 1424 138 1425 143
rect 1465 139 1469 144
rect 1471 143 1484 146
rect 1507 143 1513 146
rect 1524 143 1530 149
rect 1614 146 1620 152
rect 1633 150 1636 156
rect 1651 152 1663 154
rect 1632 146 1633 148
rect 1651 146 1666 152
rect 1675 149 1676 154
rect 1824 150 1830 156
rect 1882 150 1888 156
rect 1894 155 1896 157
rect 1674 146 1675 149
rect 1469 138 1471 139
rect 1472 138 1478 143
rect 1226 122 1230 123
rect 1231 122 1283 123
rect 1225 118 1289 122
rect 1220 116 1289 118
rect 1352 116 1355 123
rect 1079 110 1085 111
rect 1093 110 1131 111
rect 1073 107 1085 110
rect 1089 107 1137 110
rect 1073 104 1079 107
rect 1089 105 1127 107
rect 1080 104 1127 105
rect 1131 104 1137 107
rect 1079 98 1085 104
rect 1115 103 1119 104
rect 1109 101 1115 103
rect 1097 98 1109 101
rect 1125 98 1131 104
rect 1220 102 1225 116
rect 1231 111 1249 116
rect 1231 110 1237 111
rect 1277 110 1283 116
rect 1350 111 1352 116
rect 1278 108 1279 110
rect 1348 107 1350 110
rect 1384 107 1393 124
rect 1412 121 1415 123
rect 1420 121 1424 138
rect 1471 129 1481 138
rect 1530 137 1536 143
rect 1543 137 1548 146
rect 1608 144 1672 146
rect 1608 142 1666 144
rect 1667 142 1672 144
rect 1673 142 1674 145
rect 1608 140 1664 142
rect 1541 133 1542 136
rect 1481 121 1483 129
rect 1535 123 1541 133
rect 1415 120 1417 121
rect 1414 119 1418 120
rect 1414 115 1420 119
rect 1426 117 1427 119
rect 1426 115 1443 117
rect 1345 106 1348 107
rect 975 96 994 98
rect 1070 96 1071 98
rect 1092 96 1097 98
rect 994 95 1002 96
rect 1002 93 1023 95
rect 1033 93 1035 96
rect 1023 91 1037 93
rect 1033 90 1035 91
rect 1037 90 1058 91
rect 1070 90 1092 96
rect 1216 91 1220 101
rect 1279 98 1281 102
rect 1335 101 1345 106
rect 1331 100 1335 101
rect 1381 100 1384 107
rect 1417 102 1420 115
rect 1423 111 1425 112
rect 1426 108 1450 111
rect 1426 103 1438 108
rect 1450 105 1464 108
rect 1464 103 1476 105
rect 1483 103 1485 118
rect 1530 114 1535 123
rect 1614 108 1629 140
rect 1661 138 1664 140
rect 1667 138 1675 142
rect 1661 136 1663 138
rect 1662 112 1663 136
rect 1664 130 1675 138
rect 1664 126 1668 130
rect 1664 122 1667 126
rect 1670 124 1672 130
rect 1926 127 1928 157
rect 1930 154 1940 157
rect 2100 155 2102 161
rect 2110 155 2116 161
rect 2129 158 2152 182
rect 2156 155 2162 161
rect 2104 154 2110 155
rect 1932 150 1940 154
rect 1932 147 1950 150
rect 1940 143 1950 147
rect 2102 143 2110 154
rect 2115 150 2116 154
rect 2148 151 2154 154
rect 2113 143 2115 150
rect 2149 149 2154 151
rect 2162 149 2168 155
rect 1900 126 1928 127
rect 1895 125 1928 126
rect 1932 125 1940 137
rect 1950 133 1956 143
rect 2102 133 2113 143
rect 2094 132 2113 133
rect 2094 124 2103 132
rect 1669 122 1670 123
rect 1667 119 1671 122
rect 1929 121 1932 123
rect 1903 120 1906 121
rect 1666 114 1671 119
rect 1891 118 1901 120
rect 1882 116 1891 118
rect 1661 108 1663 111
rect 1476 102 1478 103
rect 1304 98 1331 100
rect 1380 98 1381 100
rect 1279 96 1311 98
rect 1269 95 1311 96
rect 1242 93 1311 95
rect 1224 91 1311 93
rect 1377 91 1380 96
rect 1036 88 1067 90
rect 1068 89 1071 90
rect 1197 89 1311 91
rect 1070 88 1071 89
rect 1037 86 1049 88
rect 1051 87 1070 88
rect 1175 87 1197 89
rect 1203 88 1311 89
rect 1216 87 1220 88
rect 1051 83 1078 87
rect 1127 83 1175 87
rect 1051 82 1089 83
rect 1116 82 1159 83
rect 1051 76 1159 82
rect 1053 74 1063 76
rect 1216 74 1217 87
rect 1281 84 1283 87
rect 1374 85 1377 91
rect 930 72 931 74
rect 1044 72 1053 74
rect 712 70 714 71
rect 414 68 416 69
rect 634 68 635 70
rect 710 68 712 70
rect 66 52 82 68
rect 84 52 100 68
rect 267 65 269 68
rect 407 65 413 68
rect 636 65 639 68
rect 706 65 710 68
rect 269 63 271 65
rect 406 64 407 65
rect 704 64 706 65
rect 404 63 406 64
rect 271 61 347 63
rect 399 61 404 63
rect 639 61 643 64
rect 702 62 704 64
rect 692 61 702 62
rect 354 60 398 61
rect 650 52 666 61
rect 667 60 668 61
rect 840 56 1064 72
rect 1281 71 1284 84
rect 1413 78 1417 101
rect 1476 97 1483 102
rect 1614 100 1666 108
rect 1667 104 1671 114
rect 1824 104 1830 110
rect 1882 104 1888 110
rect 1671 100 1673 102
rect 1472 91 1483 97
rect 1530 91 1536 97
rect 1608 94 1673 100
rect 1830 98 1836 104
rect 1876 98 1882 104
rect 1894 102 1895 118
rect 1916 113 1928 121
rect 2107 119 2113 132
rect 2150 129 2154 149
rect 2106 118 2107 119
rect 2102 109 2106 118
rect 2154 109 2156 129
rect 2102 103 2110 109
rect 2162 103 2168 109
rect 2102 102 2106 103
rect 1895 98 1897 102
rect 1476 85 1484 91
rect 1524 85 1530 91
rect 1614 88 1620 94
rect 1660 88 1666 94
rect 1476 78 1483 85
rect 1616 84 1619 88
rect 1217 68 1218 70
rect 1282 69 1284 71
rect 1280 68 1284 69
rect 1218 66 1221 68
rect 1279 66 1280 68
rect 1314 66 1344 75
rect 1348 66 1361 72
rect 1413 71 1415 78
rect 1476 77 1484 78
rect 1162 56 1348 66
rect 1415 65 1417 71
rect 1473 68 1484 77
rect 1610 72 1619 84
rect 1672 84 1673 94
rect 1610 68 1616 72
rect 1672 68 1676 84
rect 1888 72 1897 98
rect 2096 86 2102 102
rect 2110 97 2116 103
rect 2156 97 2162 103
rect 2156 86 2159 97
rect 1472 65 1473 67
rect 1615 66 1616 68
rect 946 52 962 56
rect 1064 53 1075 56
rect 1115 53 1162 56
rect 1075 52 1115 53
rect 1252 52 1268 56
rect 1314 48 1344 56
rect 1452 52 1468 65
rect 1615 56 1625 66
rect 1888 64 1901 72
rect 1956 68 1972 84
rect 2094 77 2103 86
rect 2156 79 2168 86
rect 2159 77 2168 79
rect 2096 68 2097 77
rect 2103 68 2112 77
rect 2150 68 2164 77
rect 1923 64 1956 68
rect 2156 64 2159 68
rect 1903 63 1922 64
rect 1671 57 1672 63
rect 1626 52 1642 56
rect 1644 52 1660 56
rect 1940 52 1956 64
rect 2097 57 2107 64
rect 2151 58 2156 64
rect 2145 57 2151 58
rect 2107 56 2148 57
rect 2132 52 2148 56
rect 1645 51 1646 52
<< nwell >>
rect -48 262 2440 583
<< pwell >>
rect 33 -17 67 17
rect 425 -17 459 17
rect 913 -17 947 17
rect 1401 -17 1435 17
rect 1793 -17 1827 17
<< nmos >>
rect 116 48 146 178
rect 212 48 242 178
rect 308 48 338 178
rect 508 48 538 178
rect 604 48 634 178
rect 700 48 730 178
rect 796 48 826 178
rect 996 48 1026 178
rect 1092 48 1122 178
rect 1188 48 1218 178
rect 1284 48 1314 178
rect 1484 48 1514 178
rect 1580 48 1610 178
rect 1676 48 1706 178
rect 1876 48 1906 178
rect 1972 48 2002 178
rect 2068 48 2098 178
rect 2164 48 2194 178
<< pmos >>
rect 116 298 146 498
rect 212 298 242 498
rect 308 298 338 498
rect 508 298 538 498
rect 604 298 634 498
rect 700 298 730 498
rect 796 298 826 498
rect 996 298 1026 498
rect 1092 298 1122 498
rect 1188 298 1218 498
rect 1284 298 1314 498
rect 1484 298 1514 498
rect 1580 298 1610 498
rect 1676 298 1706 498
rect 1876 298 1906 498
rect 1972 298 2002 498
rect 2068 298 2098 498
rect 2164 298 2194 498
<< ndiff >>
rect 58 102 116 178
rect 58 68 66 102
rect 100 68 116 102
rect 58 48 116 68
rect 146 102 212 178
rect 146 68 162 102
rect 196 68 212 102
rect 146 48 212 68
rect 242 48 308 178
rect 338 102 396 178
rect 338 68 354 102
rect 388 68 396 102
rect 338 48 396 68
rect 450 102 508 178
rect 450 68 458 102
rect 492 68 508 102
rect 450 48 508 68
rect 538 48 604 178
rect 634 102 700 178
rect 634 68 650 102
rect 684 68 700 102
rect 634 48 700 68
rect 730 48 796 178
rect 826 102 884 178
rect 826 68 842 102
rect 876 68 884 102
rect 826 48 884 68
rect 938 102 996 178
rect 938 68 946 102
rect 980 68 996 102
rect 938 48 996 68
rect 1026 48 1092 178
rect 1122 102 1188 178
rect 1122 68 1138 102
rect 1172 68 1188 102
rect 1122 48 1188 68
rect 1218 102 1284 178
rect 1218 68 1234 102
rect 1268 68 1284 102
rect 1218 48 1284 68
rect 1314 102 1372 178
rect 1314 68 1330 102
rect 1364 68 1372 102
rect 1314 48 1372 68
rect 1426 102 1484 178
rect 1426 68 1434 102
rect 1468 68 1484 102
rect 1426 48 1484 68
rect 1514 102 1580 178
rect 1514 68 1530 102
rect 1564 68 1580 102
rect 1514 48 1580 68
rect 1610 102 1676 178
rect 1610 68 1626 102
rect 1660 68 1676 102
rect 1610 48 1676 68
rect 1706 102 1764 178
rect 1706 68 1722 102
rect 1756 68 1764 102
rect 1706 48 1764 68
rect 1818 102 1876 178
rect 1818 68 1826 102
rect 1860 68 1876 102
rect 1818 48 1876 68
rect 1906 102 1972 178
rect 1906 68 1922 102
rect 1956 68 1972 102
rect 1906 48 1972 68
rect 2002 102 2068 178
rect 2002 68 2018 102
rect 2052 68 2068 102
rect 2002 48 2068 68
rect 2098 102 2164 178
rect 2098 68 2114 102
rect 2148 68 2164 102
rect 2098 48 2164 68
rect 2194 102 2252 178
rect 2194 68 2210 102
rect 2244 68 2252 102
rect 2194 48 2252 68
<< pdiff >>
rect 58 408 116 498
rect 58 374 66 408
rect 100 374 116 408
rect 58 298 116 374
rect 146 478 212 498
rect 146 444 162 478
rect 196 444 212 478
rect 146 298 212 444
rect 242 380 308 498
rect 242 346 258 380
rect 292 346 308 380
rect 242 298 308 346
rect 338 478 396 498
rect 338 444 354 478
rect 388 444 396 478
rect 338 298 396 444
rect 450 380 508 498
rect 450 346 458 380
rect 492 346 508 380
rect 450 298 508 346
rect 538 478 604 498
rect 538 444 554 478
rect 588 444 604 478
rect 538 298 604 444
rect 634 380 700 498
rect 634 346 650 380
rect 684 346 700 380
rect 634 298 700 346
rect 730 380 796 498
rect 730 346 746 380
rect 780 346 796 380
rect 730 298 796 346
rect 826 380 884 498
rect 826 346 842 380
rect 876 346 884 380
rect 826 298 884 346
rect 938 478 996 498
rect 938 444 946 478
rect 980 444 996 478
rect 938 298 996 444
rect 1026 380 1092 498
rect 1026 346 1042 380
rect 1076 346 1092 380
rect 1026 298 1092 346
rect 1122 478 1188 498
rect 1122 444 1138 478
rect 1172 444 1188 478
rect 1122 298 1188 444
rect 1218 298 1284 498
rect 1314 380 1372 498
rect 1314 346 1330 380
rect 1364 346 1372 380
rect 1314 298 1372 346
rect 1426 448 1484 498
rect 1426 414 1434 448
rect 1468 414 1484 448
rect 1426 298 1484 414
rect 1514 478 1580 498
rect 1514 444 1530 478
rect 1564 444 1580 478
rect 1514 298 1580 444
rect 1610 298 1676 498
rect 1706 380 1764 498
rect 1706 346 1722 380
rect 1756 346 1764 380
rect 1706 298 1764 346
rect 1818 380 1876 498
rect 1818 346 1826 380
rect 1860 346 1876 380
rect 1818 298 1876 346
rect 1906 298 1972 498
rect 2002 478 2068 498
rect 2002 444 2018 478
rect 2052 444 2068 478
rect 2002 298 2068 444
rect 2098 298 2164 498
rect 2194 380 2252 498
rect 2194 346 2210 380
rect 2244 346 2252 380
rect 2194 298 2252 346
<< ndiffc >>
rect 66 68 100 102
rect 162 68 196 102
rect 354 68 388 102
rect 458 68 492 102
rect 650 68 684 102
rect 842 68 876 102
rect 946 68 980 102
rect 1138 68 1172 102
rect 1234 68 1268 102
rect 1330 68 1364 102
rect 1434 68 1468 102
rect 1530 68 1564 102
rect 1626 68 1660 102
rect 1722 68 1756 102
rect 1826 68 1860 102
rect 1922 68 1956 102
rect 2018 68 2052 102
rect 2114 68 2148 102
rect 2210 68 2244 102
<< pdiffc >>
rect 66 374 100 408
rect 162 444 196 478
rect 258 346 292 380
rect 354 444 388 478
rect 458 346 492 380
rect 554 444 588 478
rect 650 346 684 380
rect 746 346 780 380
rect 842 346 876 380
rect 946 444 980 478
rect 1042 346 1076 380
rect 1138 444 1172 478
rect 1330 346 1364 380
rect 1434 414 1468 448
rect 1530 444 1564 478
rect 1722 346 1756 380
rect 1826 346 1860 380
rect 2018 444 2052 478
rect 2210 346 2244 380
<< poly >>
rect 116 498 146 524
rect 212 498 242 524
rect 308 498 338 524
rect 508 498 538 524
rect 604 498 634 524
rect 700 498 730 524
rect 796 498 826 524
rect 996 498 1026 524
rect 1092 498 1122 524
rect 1188 498 1218 524
rect 1284 498 1314 524
rect 1484 498 1514 524
rect 1580 498 1610 524
rect 1676 498 1706 524
rect 1876 498 1906 524
rect 1972 498 2002 524
rect 2068 498 2098 524
rect 2164 498 2194 524
rect 116 266 146 298
rect 212 266 242 298
rect 308 266 338 298
rect 508 266 538 298
rect 604 266 634 298
rect 700 266 730 298
rect 796 266 826 298
rect 996 266 1026 298
rect 1092 266 1122 298
rect 1188 266 1218 298
rect 1284 266 1314 298
rect 1484 266 1514 298
rect 1580 266 1610 298
rect 1676 266 1706 298
rect 1876 266 1906 298
rect 1972 266 2002 298
rect 2068 266 2098 298
rect 2164 266 2194 298
rect 104 250 158 266
rect 104 216 114 250
rect 148 216 158 250
rect 104 200 158 216
rect 200 250 254 266
rect 200 216 210 250
rect 244 216 254 250
rect 200 200 254 216
rect 296 250 350 266
rect 296 216 306 250
rect 340 216 350 250
rect 296 200 350 216
rect 496 250 550 266
rect 496 216 506 250
rect 540 216 550 250
rect 496 200 550 216
rect 592 250 646 266
rect 592 216 602 250
rect 636 216 646 250
rect 592 200 646 216
rect 688 250 742 266
rect 688 216 698 250
rect 732 216 742 250
rect 688 200 742 216
rect 784 250 838 266
rect 784 216 794 250
rect 828 216 838 250
rect 784 200 838 216
rect 984 250 1038 266
rect 984 216 994 250
rect 1028 216 1038 250
rect 984 200 1038 216
rect 1080 250 1134 266
rect 1080 216 1090 250
rect 1124 216 1134 250
rect 1080 200 1134 216
rect 1176 250 1230 266
rect 1176 216 1186 250
rect 1220 216 1230 250
rect 1176 200 1230 216
rect 1272 250 1326 266
rect 1272 216 1282 250
rect 1316 216 1326 250
rect 1272 200 1326 216
rect 1472 250 1526 266
rect 1472 216 1482 250
rect 1516 216 1526 250
rect 1472 200 1526 216
rect 1568 250 1622 266
rect 1568 216 1578 250
rect 1612 216 1622 250
rect 1568 200 1622 216
rect 1664 250 1718 266
rect 1664 216 1674 250
rect 1708 216 1718 250
rect 1664 200 1718 216
rect 1864 250 1918 266
rect 1864 216 1874 250
rect 1908 216 1918 250
rect 1864 200 1918 216
rect 1960 250 2014 266
rect 1960 216 1970 250
rect 2004 216 2014 250
rect 1960 200 2014 216
rect 2056 250 2110 266
rect 2056 216 2066 250
rect 2100 216 2110 250
rect 2056 200 2110 216
rect 2152 250 2206 266
rect 2152 216 2162 250
rect 2196 216 2206 250
rect 2152 200 2206 216
rect 116 178 146 200
rect 212 178 242 200
rect 308 178 338 200
rect 508 178 538 200
rect 604 178 634 200
rect 700 178 730 200
rect 796 178 826 200
rect 996 178 1026 200
rect 1092 178 1122 200
rect 1188 178 1218 200
rect 1284 178 1314 200
rect 1484 178 1514 200
rect 1580 178 1610 200
rect 1676 178 1706 200
rect 1876 178 1906 200
rect 1972 178 2002 200
rect 2068 178 2098 200
rect 2164 178 2194 200
rect 116 22 146 48
rect 212 22 242 48
rect 308 22 338 48
rect 508 22 538 48
rect 604 22 634 48
rect 700 22 730 48
rect 796 22 826 48
rect 996 22 1026 48
rect 1092 22 1122 48
rect 1188 22 1218 48
rect 1284 22 1314 48
rect 1484 22 1514 48
rect 1580 22 1610 48
rect 1676 22 1706 48
rect 1876 22 1906 48
rect 1972 22 2002 48
rect 2068 22 2098 48
rect 2164 22 2194 48
<< polycont >>
rect 114 216 148 250
rect 210 216 244 250
rect 306 216 340 250
rect 506 216 540 250
rect 602 216 636 250
rect 698 216 732 250
rect 794 216 828 250
rect 994 216 1028 250
rect 1090 216 1124 250
rect 1186 216 1220 250
rect 1282 216 1316 250
rect 1482 216 1516 250
rect 1578 216 1612 250
rect 1674 216 1708 250
rect 1874 216 1908 250
rect 1970 216 2004 250
rect 2066 216 2100 250
rect 2162 216 2196 250
<< locali >>
rect 0 528 29 562
rect 63 528 121 562
rect 155 528 213 562
rect 247 528 305 562
rect 339 528 397 562
rect 431 528 489 562
rect 523 528 581 562
rect 615 528 673 562
rect 707 528 765 562
rect 799 528 857 562
rect 891 528 949 562
rect 983 528 1041 562
rect 1075 528 1133 562
rect 1167 528 1225 562
rect 1259 528 1317 562
rect 1351 528 1409 562
rect 1443 528 1501 562
rect 1535 528 1593 562
rect 1627 528 1685 562
rect 1719 528 1777 562
rect 1811 528 1869 562
rect 1903 528 1961 562
rect 1995 528 2053 562
rect 2087 528 2145 562
rect 2179 528 2237 562
rect 2271 528 2329 562
rect 2363 528 2392 562
rect 162 478 196 528
tri 38 435 53 438 se
tri 53 435 77 438 sw
tri 35 426 38 435 se
rect 38 432 77 435
tri 77 432 106 435 sw
rect 38 426 106 432
tri 106 426 110 432 sw
rect 162 428 196 444
rect 354 478 388 528
rect 354 428 388 444
rect 554 478 588 528
rect 554 428 588 444
rect 946 478 980 528
tri 846 428 855 432 se
tri 855 428 898 432 sw
rect 946 428 980 444
rect 1138 478 1172 528
rect 1530 478 1564 528
tri 1428 451 1439 463 se
rect 1439 451 1488 463
tri 1332 448 1333 451 se
rect 1138 428 1172 444
tri 1330 438 1332 447 se
rect 1332 438 1333 448
tri 1329 436 1330 438 se
rect 1330 436 1333 438
tri 1328 432 1329 435 se
rect 1329 432 1333 436
tri 1327 428 1328 432 se
rect 1328 428 1333 432
tri 840 426 846 428 se
rect 846 426 898 428
rect 35 425 110 426
tri 110 425 111 426 sw
rect 35 422 111 425
tri 835 424 840 426 se
rect 840 424 898 426
rect 69 408 111 422
tri 642 414 656 419 se
rect 656 414 677 419
tri 677 414 682 419 sw
tri 827 414 835 424 se
rect 835 414 898 424
tri 627 409 642 414 se
rect 642 409 682 414
tri 682 409 688 414 sw
tri 826 413 827 414 se
rect 827 413 898 414
tri 34 374 35 408 se
rect 35 374 66 388
rect 100 374 111 408
tri 614 401 627 409 se
rect 627 401 688 409
tri 441 388 457 401 se
rect 457 391 524 401
tri 524 391 541 401 sw
tri 600 393 614 401 se
rect 614 393 637 401
tri 594 391 600 393 se
rect 600 391 637 393
rect 457 390 541 391
tri 541 390 590 391 sw
tri 590 390 594 391 se
rect 594 390 637 391
rect 457 388 637 390
tri 260 380 303 388 se
tri 303 386 315 388 sw
rect 303 380 315 386
tri 315 380 319 386 sw
rect 441 380 637 388
rect 671 399 688 401
tri 688 399 701 409 sw
rect 671 380 701 399
tri 740 390 760 393 se
rect 760 390 784 393
rect 740 381 784 390
tri 784 381 785 390 sw
rect 740 380 785 381
rect 826 380 855 413
rect 889 411 898 413
tri 898 411 915 428 sw
tri 1325 424 1327 428 se
rect 1327 424 1333 428
tri 1322 414 1325 423 se
rect 1325 417 1333 424
rect 1428 448 1488 451
tri 1367 426 1369 448 sw
rect 1367 417 1369 426
rect 1325 416 1369 417
tri 1369 416 1370 417 sw
rect 1325 414 1370 416
rect 1428 414 1434 448
rect 1468 437 1488 448
rect 34 369 111 374
tri 34 356 41 369 ne
rect 41 365 111 369
rect 41 356 97 365
tri 97 356 111 365 nw
tri 249 356 258 380 se
tri 41 346 66 356 ne
rect 66 346 81 356
tri 81 346 97 356 nw
tri 245 346 249 356 se
rect 249 346 258 356
rect 292 373 319 380
tri 319 373 324 380 sw
rect 292 346 324 373
tri 242 337 245 346 se
rect 245 341 324 346
rect 245 337 289 341
tri 156 334 168 336 se
tri 168 334 186 336 sw
tri 236 334 242 337 se
rect 242 334 289 337
tri 132 318 156 334 se
rect 156 328 186 334
tri 186 328 229 334 sw
tri 229 328 236 334 se
rect 236 328 289 334
rect 156 318 289 328
tri 108 280 132 318 se
rect 132 307 289 318
rect 323 327 324 341
rect 441 346 458 380
rect 492 367 637 380
rect 492 346 650 367
rect 684 346 700 380
tri 700 346 701 380 nw
tri 739 346 740 380 se
rect 740 346 746 380
rect 780 347 785 380
tri 785 347 789 380 sw
tri 826 359 827 380 ne
rect 780 346 789 347
rect 827 346 842 380
rect 889 379 915 411
tri 1320 403 1322 411 se
rect 1322 405 1370 414
tri 1370 405 1371 414 sw
rect 1322 403 1371 405
rect 1428 408 1449 414
tri 1428 403 1432 408 ne
rect 1432 403 1449 408
rect 1483 403 1488 437
rect 2018 478 2052 528
tri 1679 445 1709 448 se
rect 1709 445 1717 448
rect 1530 428 1564 444
rect 1671 414 1717 445
rect 1751 414 1758 448
rect 1671 411 1758 414
tri 1637 405 1641 411 ne
rect 1641 405 1758 411
tri 1925 406 1929 444 se
rect 2018 428 2052 444
rect 1929 406 1963 414
tri 2231 406 2235 407 se
tri 2235 406 2249 407 sw
rect 1320 399 1371 403
tri 1035 389 1059 399 se
tri 1059 395 1103 399 sw
tri 1320 395 1321 399 ne
rect 1321 395 1371 399
rect 1059 389 1103 395
tri 1103 389 1116 395 sw
tri 1321 389 1322 395 ne
rect 1322 389 1371 395
rect 1035 380 1116 389
tri 1116 380 1133 389 sw
tri 1322 382 1323 389 ne
rect 1323 383 1371 389
tri 1371 383 1373 403 sw
tri 1432 395 1438 403 ne
rect 1438 397 1488 403
tri 1438 395 1488 397 nw
tri 1641 395 1648 405 ne
rect 1648 395 1758 405
rect 1323 380 1373 383
tri 1648 380 1659 395 ne
rect 1659 380 1758 395
tri 1922 394 1925 406 se
rect 1925 394 1963 406
tri 2219 404 2231 406 se
rect 2231 404 2249 406
tri 1921 388 1922 393 se
rect 1922 388 1963 394
tri 1804 380 1807 388 se
rect 1807 387 1845 388
tri 1845 387 1860 388 sw
rect 1807 380 1860 387
tri 1920 382 1921 387 se
rect 1921 382 1963 388
rect 1920 381 1963 382
tri 1963 381 1966 404 sw
tri 2118 381 2219 404 se
rect 2219 392 2249 404
tri 2249 392 2271 406 sw
rect 2219 381 2271 392
rect 876 369 915 379
tri 915 369 916 380 sw
rect 876 346 911 369
tri 911 346 916 369 nw
rect 1035 346 1042 380
rect 1076 369 1133 380
tri 1133 369 1155 380 sw
tri 1323 370 1325 380 ne
rect 1325 369 1330 380
rect 1076 362 1155 369
tri 1155 362 1176 369 sw
tri 1325 363 1326 369 ne
rect 1326 362 1330 369
rect 1076 352 1176 362
rect 1076 346 1094 352
rect 441 343 700 346
rect 441 336 691 343
tri 691 336 700 343 nw
rect 739 338 789 346
tri 789 338 791 346 sw
tri 441 334 443 336 ne
rect 443 334 686 336
tri 323 318 324 327 nw
tri 371 318 372 328 se
tri 370 311 371 318 se
rect 371 311 372 318
rect 132 298 294 307
tri 294 298 323 307 nw
tri 367 299 370 311 se
rect 370 300 372 311
tri 443 328 450 334 ne
rect 450 332 686 334
tri 686 332 691 336 nw
rect 450 328 600 332
tri 450 326 453 328 ne
rect 453 327 600 328
tri 600 327 686 332 nw
rect 453 326 588 327
tri 588 326 600 327 nw
tri 453 325 556 326 ne
tri 556 325 583 326 nw
rect 739 325 757 338
tri 739 313 748 325 ne
rect 748 313 757 325
tri 748 304 757 313 ne
rect 827 345 911 346
rect 827 336 909 345
tri 909 336 911 345 nw
rect 1035 341 1094 346
tri 1035 338 1038 341 ne
rect 1038 338 1094 341
rect 827 333 906 336
tri 906 333 909 336 nw
tri 961 333 962 336 se
tri 827 319 841 333 ne
rect 841 319 896 333
tri 896 319 906 333 nw
tri 960 329 961 333 se
rect 961 329 962 333
tri 959 319 960 328 se
rect 960 319 962 329
tri 841 318 879 319 ne
tri 879 318 896 319 nw
tri 958 316 959 318 se
rect 959 316 962 319
rect 958 304 962 316
tri 1038 336 1039 338 ne
rect 1039 336 1094 338
tri 996 333 997 336 sw
tri 1039 333 1043 336 ne
rect 1043 333 1094 336
rect 996 328 997 333
tri 997 328 999 333 sw
tri 1043 328 1048 333 ne
rect 1048 328 1094 333
rect 996 324 999 328
tri 999 324 1000 328 sw
tri 1048 324 1061 328 ne
rect 1061 324 1094 328
rect 996 319 1000 324
tri 1000 319 1002 324 sw
tri 1061 319 1073 324 ne
rect 1073 319 1094 324
rect 996 318 1002 319
tri 1002 318 1003 319 sw
tri 1076 318 1078 319 ne
rect 1078 318 1094 319
rect 1128 346 1176 352
tri 1176 346 1278 362 sw
tri 1326 346 1330 362 ne
rect 1364 363 1373 380
tri 1373 363 1375 380 sw
tri 1659 365 1671 380 ne
rect 1671 365 1722 380
tri 1671 363 1673 365 ne
rect 1673 363 1722 365
rect 1364 361 1375 363
rect 1364 346 1368 361
tri 1368 346 1375 361 nw
tri 1673 354 1693 363 ne
rect 1693 354 1722 363
tri 1506 348 1577 354 se
tri 1577 348 1588 354 sw
tri 1489 346 1506 348 se
rect 1506 346 1588 348
tri 1588 346 1592 348 sw
tri 1693 346 1709 354 ne
rect 1709 346 1722 354
rect 1756 365 1758 380
tri 1800 369 1804 380 se
rect 1804 369 1826 380
rect 1756 346 1757 365
tri 1757 346 1758 365 nw
tri 1795 355 1800 369 se
rect 1800 355 1826 369
rect 1128 331 1278 346
tri 1278 331 1296 346 sw
tri 1479 345 1486 346 se
rect 1486 345 1592 346
tri 1592 345 1593 346 sw
tri 1709 345 1713 346 ne
rect 1713 345 1757 346
tri 1469 341 1479 345 se
rect 1479 341 1593 345
tri 1465 339 1469 341 se
rect 1469 339 1593 341
tri 1593 339 1596 345 sw
tri 1713 344 1715 345 ne
rect 1715 344 1757 345
tri 1715 343 1732 344 ne
tri 1732 343 1741 344 nw
rect 1128 318 1296 331
tri 1449 334 1465 339 se
rect 1465 334 1596 339
tri 1596 334 1599 339 sw
rect 996 316 1003 318
tri 1003 316 1004 318 sw
tri 1078 316 1083 318 ne
rect 1083 316 1296 318
rect 996 313 1004 316
tri 1004 313 1005 316 sw
rect 996 304 1005 313
tri 1005 304 1014 313 sw
tri 1083 311 1098 316 ne
rect 1098 312 1296 316
tri 1296 312 1300 328 sw
rect 1098 311 1300 312
tri 1098 308 1156 311 ne
rect 1156 308 1300 311
tri 1300 308 1301 311 sw
tri 1156 304 1181 308 ne
rect 1181 304 1301 308
rect 370 299 403 300
rect 132 282 173 298
tri 173 282 294 298 nw
tri 364 287 367 298 se
rect 367 291 403 299
tri 403 291 406 300 nw
rect 958 302 1014 304
tri 1014 302 1017 304 sw
tri 1181 302 1193 304 ne
rect 1193 302 1301 304
rect 958 291 1017 302
tri 1017 291 1019 302 sw
tri 1193 291 1260 302 ne
rect 1260 291 1301 302
tri 1301 291 1305 308 sw
rect 1483 331 1599 334
tri 1599 331 1601 334 sw
rect 1483 328 1601 331
tri 1601 328 1602 331 sw
rect 1483 314 1602 328
tri 1602 314 1609 328 sw
rect 1829 343 1860 346
tri 1912 346 1920 380 se
rect 1920 368 1966 381
tri 2114 380 2118 381 se
rect 2118 380 2271 381
tri 1966 368 1967 380 sw
tri 2078 372 2114 380 se
rect 2114 372 2210 380
rect 1920 346 1933 368
rect 1829 339 1859 343
tri 1859 339 1860 343 nw
rect 1829 332 1858 339
tri 1858 334 1859 339 nw
tri 1910 334 1912 344 se
rect 1912 334 1933 346
tri 2069 366 2078 372 se
rect 2078 366 2210 372
tri 2058 346 2069 366 se
rect 2069 346 2210 366
rect 2244 373 2271 380
tri 2271 373 2274 392 sw
rect 2244 366 2274 373
tri 2274 366 2275 372 sw
rect 2244 346 2275 366
tri 2275 353 2278 366 sw
tri 2275 346 2278 353 nw
rect 1829 331 1857 332
tri 1857 331 1858 332 nw
rect 1829 328 1856 331
tri 1856 328 1857 331 nw
tri 1909 328 1910 331 se
rect 1910 328 1960 334
rect 1829 321 1852 328
tri 1852 321 1856 328 nw
tri 1908 321 1909 328 se
rect 1909 325 1960 328
tri 1960 325 1967 334 nw
tri 2053 336 2058 345 se
rect 2058 337 2266 346
tri 2266 337 2275 346 nw
rect 2058 336 2258 337
tri 2258 336 2266 337 nw
rect 1909 321 1953 325
tri 1795 315 1807 321 ne
rect 1807 320 1852 321
tri 1907 320 1908 321 se
rect 1908 320 1953 321
rect 1807 315 1836 320
tri 1836 315 1852 320 nw
tri 1906 315 1907 320 se
rect 1907 315 1953 320
tri 1953 315 1960 325 nw
tri 1807 314 1833 315 ne
tri 1833 314 1836 315 nw
rect 1483 311 1609 314
tri 1609 311 1611 314 sw
rect 1483 308 1611 311
tri 1611 308 1612 311 sw
tri 1905 308 1906 311 se
rect 1906 308 1935 315
rect 1483 300 1612 308
tri 1612 300 1616 308 sw
tri 1903 300 1905 308 se
rect 1905 300 1935 308
tri 1449 291 1488 300 ne
rect 1488 291 1616 300
rect 367 287 402 291
tri 402 287 403 291 nw
rect 958 288 1019 291
tri 1019 288 1020 291 sw
tri 360 282 364 287 se
rect 364 282 400 287
rect 132 280 169 282
tri 169 280 173 282 nw
tri 359 281 360 282 se
rect 360 281 400 282
tri 400 281 402 287 nw
tri 354 280 359 281 se
rect 359 280 399 281
tri 89 274 108 280 se
rect 108 274 160 280
tri 160 274 169 280 nw
tri 340 276 354 280 se
rect 354 276 399 280
tri 399 276 400 281 nw
tri 337 274 340 276 se
rect 340 274 393 276
tri 85 268 89 274 se
rect 89 269 153 274
tri 153 269 160 274 nw
tri 331 269 337 274 se
rect 337 269 393 274
rect 89 268 152 269
tri 152 268 153 269 nw
tri 330 268 331 269 se
rect 331 268 393 269
tri 83 253 85 268 se
rect 85 253 149 268
tri 149 261 152 268 nw
tri 320 261 330 268 se
rect 330 261 393 268
rect 83 250 149 253
tri 307 250 320 261 se
rect 320 250 393 261
tri 393 250 399 276 nw
rect 610 281 611 287
tri 611 281 614 287 sw
rect 958 284 1020 288
tri 1020 284 1021 287 sw
tri 1261 284 1268 291 ne
rect 1268 284 1305 291
tri 1305 284 1307 291 sw
tri 1488 286 1510 291 ne
rect 1510 286 1616 291
tri 1616 286 1624 300 sw
tri 1706 286 1724 293 se
rect 1724 292 1765 293
rect 1724 286 1730 292
tri 1524 284 1529 286 ne
rect 1529 284 1624 286
rect 958 281 1021 284
rect 1268 281 1307 284
rect 610 280 614 281
tri 614 280 615 281 sw
tri 958 280 959 281 ne
rect 610 276 615 280
tri 615 276 618 280 sw
rect 959 278 1021 281
tri 1021 278 1022 281 sw
rect 610 262 618 276
tri 618 262 627 276 sw
tri 678 264 688 270 se
tri 688 265 736 270 sw
rect 688 264 736 265
tri 736 264 737 265 sw
rect 959 264 1022 278
tri 1268 277 1269 281 ne
rect 1269 278 1307 281
tri 1307 278 1308 284 sw
tri 1529 278 1546 284 ne
rect 1546 278 1624 284
tri 1022 264 1025 277 sw
rect 1269 276 1308 278
tri 1269 264 1271 276 ne
rect 1271 264 1308 276
tri 1308 264 1317 278 sw
tri 1546 275 1555 278 ne
rect 1555 275 1624 278
tri 1624 275 1629 286 sw
tri 1689 278 1706 286 se
rect 1706 278 1730 286
tri 1687 275 1689 278 se
rect 1689 275 1730 278
tri 1555 265 1558 275 ne
rect 1558 271 1629 275
tri 1629 271 1631 275 sw
tri 1685 271 1687 275 se
rect 1687 271 1730 275
rect 1558 264 1631 271
tri 1683 268 1685 271 se
rect 1685 268 1730 271
rect 678 262 737 264
tri 737 262 740 264 sw
rect 610 253 627 262
rect 576 252 627 253
tri 627 252 634 262 sw
rect 576 250 634 252
tri 634 250 635 252 sw
rect 678 250 740 262
tri 855 252 865 258 se
tri 79 224 83 250 se
tri 79 216 83 224 ne
rect 83 216 114 250
tri 148 224 149 250 nw
tri 244 249 251 250 sw
rect 244 246 251 249
tri 251 246 255 249 sw
rect 244 229 255 246
tri 83 209 102 216 ne
rect 102 211 113 216
tri 113 211 148 216 nw
tri 254 224 255 229 nw
rect 210 215 220 216
tri 210 211 213 215 ne
tri 102 209 113 211 nw
rect 213 209 220 215
tri 213 195 220 209 ne
rect 340 249 393 250
tri 495 249 503 250 se
rect 503 249 506 250
rect 340 229 388 249
tri 388 230 393 249 nw
tri 436 245 495 249 se
rect 495 245 506 249
rect 340 225 387 229
tri 387 225 388 229 nw
rect 340 224 385 225
tri 385 224 387 225 nw
rect 340 221 381 224
tri 381 221 385 224 nw
rect 340 217 378 221
tri 378 217 381 221 nw
rect 340 216 342 217
tri 342 216 378 217 nw
tri 306 215 342 216 nw
rect 470 216 506 245
rect 576 244 602 250
tri 576 240 577 244 ne
rect 577 240 602 244
tri 577 230 579 240 ne
rect 579 230 602 240
tri 579 226 581 230 ne
rect 581 224 602 230
tri 581 221 582 224 ne
rect 582 221 602 224
tri 582 217 583 221 ne
rect 470 215 539 216
tri 539 215 540 216 nw
rect 583 216 602 221
rect 583 215 636 216
rect 470 211 538 215
tri 538 211 539 215 nw
tri 583 211 584 215 ne
rect 584 211 636 215
tri 436 203 470 211 ne
rect 470 203 533 211
tri 533 203 538 211 nw
tri 584 204 586 211 ne
rect 586 204 636 211
rect 678 239 698 250
rect 732 244 740 250
rect 732 221 739 244
tri 739 231 740 244 nw
rect 794 250 865 252
rect 732 216 738 221
tri 738 217 739 221 nw
rect 712 211 738 216
rect 712 206 734 211
tri 734 206 738 211 nw
rect 828 224 865 250
rect 959 253 1025 264
tri 1025 253 1027 264 sw
tri 1089 260 1097 261 se
tri 1097 260 1103 261 sw
rect 1271 260 1317 264
tri 1317 260 1320 264 sw
tri 1081 253 1089 260 se
rect 1089 254 1103 260
tri 1103 254 1126 260 sw
rect 1089 253 1126 254
rect 959 252 1027 253
tri 1027 252 1028 253 sw
tri 1079 252 1081 253 se
rect 1081 252 1126 253
tri 1126 252 1127 253 sw
tri 1179 252 1180 253 se
rect 1180 252 1232 253
rect 959 250 1028 252
tri 1077 250 1079 252 se
rect 1079 250 1127 252
tri 1127 250 1128 252 sw
rect 959 244 994 250
tri 959 230 977 244 ne
rect 977 230 994 244
tri 977 225 983 230 ne
rect 983 225 994 230
tri 983 224 984 225 ne
rect 984 224 994 225
rect 828 221 889 224
tri 889 221 899 224 nw
tri 984 221 989 224 ne
rect 989 221 994 224
rect 828 217 880 221
tri 880 217 889 221 nw
tri 989 217 993 221 ne
rect 993 217 994 221
rect 828 216 876 217
tri 876 216 878 217 nw
tri 1068 244 1076 250 se
rect 1076 244 1090 250
rect 1068 242 1090 244
rect 1124 248 1128 250
tri 1128 248 1130 250 sw
rect 1124 244 1129 248
tri 1129 244 1130 248 nw
tri 1177 248 1179 252 se
rect 1179 250 1232 252
rect 1179 248 1186 250
rect 1068 216 1071 242
rect 1124 216 1126 244
tri 1126 217 1129 244 nw
tri 794 206 802 216 ne
rect 802 206 825 216
tri 712 205 734 206 nw
tri 802 205 804 206 ne
tri 470 196 523 203 ne
rect 523 201 532 203
tri 532 201 533 203 nw
tri 586 201 592 204 ne
rect 592 201 636 204
tri 523 196 532 201 nw
tri 592 196 599 201 ne
rect 599 197 636 201
rect 804 204 825 206
tri 804 198 809 204 ne
rect 809 198 825 204
tri 825 198 876 216 nw
tri 1068 213 1069 216 ne
rect 1069 213 1071 216
tri 1069 208 1071 213 ne
rect 1105 208 1125 216
tri 1125 214 1126 216 nw
rect 1177 216 1186 248
rect 1220 249 1232 250
tri 1232 249 1236 253 sw
rect 1220 232 1236 249
tri 1071 206 1078 208 ne
rect 1078 206 1124 208
tri 1124 206 1125 208 nw
tri 1078 205 1084 206 ne
rect 1084 205 1124 206
tri 1084 198 1104 205 ne
rect 1104 201 1121 205
tri 1121 201 1124 205 nw
rect 1104 198 1106 201
tri 1106 198 1121 201 nw
rect 1177 200 1194 216
tri 1177 198 1178 200 ne
rect 1178 198 1194 200
rect 1228 200 1236 232
rect 1271 250 1320 260
tri 1558 250 1563 264 ne
rect 1563 250 1631 264
tri 1681 263 1683 268 se
rect 1683 263 1730 268
tri 1675 251 1681 263 se
rect 1681 258 1730 263
rect 1764 258 1765 292
tri 1901 286 1903 300 se
rect 1903 286 1935 300
tri 1898 275 1901 286 se
rect 1901 275 1935 286
tri 1897 268 1898 271 se
rect 1898 268 1935 275
tri 1935 268 1953 315 nw
rect 2087 325 2190 336
tri 2190 325 2258 336 nw
rect 2087 317 2134 325
tri 2134 317 2190 325 nw
rect 2087 315 2128 317
tri 2128 315 2134 317 nw
tri 2087 302 2128 315 nw
tri 1894 263 1897 268 se
rect 1897 263 1933 268
tri 1933 263 1935 268 nw
rect 1681 251 1765 258
tri 1875 255 1894 263 se
rect 1894 255 1930 263
tri 1930 255 1933 263 nw
tri 1978 255 2019 261 se
tri 2019 255 2061 261 sw
tri 1674 250 1675 251 se
rect 1675 250 1765 251
tri 1872 251 1875 255 se
rect 1875 251 1928 255
tri 1928 251 1930 255 nw
tri 1971 251 1976 255 se
rect 1872 250 1928 251
tri 1271 230 1274 250 ne
rect 1274 224 1282 250
tri 1274 221 1275 224 ne
rect 1275 216 1282 224
rect 1316 216 1320 250
rect 1275 215 1320 216
tri 1275 213 1276 215 ne
rect 1276 213 1320 215
tri 1236 204 1237 213 sw
tri 1236 201 1237 204 nw
tri 1276 201 1304 213 ne
rect 1304 209 1320 213
tri 1304 201 1320 209 nw
tri 1449 242 1482 250 se
tri 1516 242 1517 250 sw
tri 1563 242 1566 250 ne
rect 1566 242 1578 250
rect 1516 224 1517 242
tri 1517 224 1519 242 sw
rect 1516 216 1519 224
tri 1566 218 1574 242 ne
rect 1574 216 1578 242
rect 1612 220 1631 250
tri 1631 220 1632 250 sw
rect 1612 216 1627 220
tri 1627 216 1632 220 nw
tri 1673 216 1674 235 se
rect 1708 219 1765 250
rect 1708 216 1764 219
tri 1764 216 1765 219 nw
tri 1871 227 1872 250 se
rect 1872 227 1874 250
tri 1871 216 1874 227 ne
rect 1908 243 1925 250
tri 1925 243 1928 250 nw
tri 1970 250 1971 251 se
rect 1971 250 1976 251
rect 2010 250 2061 255
tri 2061 250 2101 255 sw
tri 2192 269 2195 286 sw
rect 2192 264 2195 269
tri 2195 264 2196 268 sw
rect 2192 256 2196 264
tri 2196 256 2198 263 sw
rect 2192 252 2198 256
rect 2158 250 2198 252
rect 1908 230 1919 243
tri 1919 230 1925 243 nw
rect 1908 227 1917 230
tri 1917 227 1919 230 nw
rect 1908 219 1911 227
tri 1911 219 1917 227 nw
rect 2010 221 2066 250
tri 1908 216 1911 219 nw
rect 2004 216 2066 221
rect 2100 249 2101 250
tri 2101 249 2110 250 sw
tri 2158 249 2159 250 ne
rect 2100 244 2110 249
tri 2110 244 2113 249 sw
rect 2100 243 2113 244
tri 2113 243 2114 244 sw
rect 2100 222 2114 243
rect 2159 243 2162 250
tri 2159 230 2161 243 ne
rect 2100 220 2113 222
tri 2113 220 2114 222 nw
rect 2161 227 2162 243
tri 2161 220 2162 227 ne
rect 2100 219 2112 220
tri 2112 219 2113 220 nw
rect 2100 216 2111 219
tri 2111 216 2112 219 nw
rect 2196 240 2198 250
tri 2198 240 2200 252 sw
rect 2196 217 2200 240
tri 2200 217 2202 240 sw
rect 2196 216 2202 217
rect 1483 215 1519 216
tri 1519 215 1520 216 sw
tri 1574 215 1575 216 ne
rect 1575 215 1625 216
rect 1483 213 1520 215
tri 1575 214 1625 215 ne
tri 1625 214 1627 216 nw
tri 1520 213 1521 214 nw
rect 1673 213 1764 216
tri 1874 215 1882 216 ne
tri 1882 215 1898 216 nw
tri 1971 215 1973 216 ne
rect 1973 215 2110 216
tri 2110 215 2111 216 nw
tri 1974 214 1976 215 ne
rect 1976 214 2110 215
tri 1976 213 1980 214 ne
rect 1980 213 2109 214
tri 2109 213 2110 214 nw
rect 2162 214 2202 216
tri 2162 213 2163 214 ne
rect 1483 208 1517 213
tri 1517 208 1520 213 nw
rect 1673 208 1763 213
tri 1763 209 1764 213 nw
tri 1981 209 1996 213 ne
rect 1996 211 2057 213
tri 2057 211 2100 213 nw
rect 2163 212 2202 214
rect 2163 211 2200 212
rect 1996 209 1998 211
tri 1996 208 1998 209 ne
tri 1998 208 2057 211 nw
tri 2163 208 2164 211 ne
rect 2164 208 2200 211
tri 2200 208 2202 212 nw
tri 1488 207 1516 208 ne
rect 1673 203 1762 208
tri 1762 203 1763 208 nw
tri 2164 203 2170 208 ne
rect 2170 203 2197 208
tri 2197 203 2200 208 nw
rect 1228 198 1235 200
rect 599 196 635 197
tri 599 195 600 196 ne
rect 600 195 635 196
tri 635 195 636 197 nw
tri 1178 195 1179 198 ne
rect 1179 195 1235 198
tri 1235 195 1236 200 nw
rect 1673 200 1761 203
tri 1761 200 1762 203 nw
rect 1673 196 1750 200
tri 1750 196 1761 200 nw
tri 1673 195 1674 196 ne
rect 1674 195 1742 196
tri 601 191 607 195 ne
rect 607 191 632 195
tri 632 191 635 195 nw
tri 1179 191 1191 195 ne
rect 1191 194 1235 195
tri 1674 194 1676 195 ne
rect 1676 194 1742 195
tri 1742 194 1750 196 nw
rect 1191 192 1209 194
tri 1209 192 1235 194 nw
tri 1676 192 1679 194 ne
tri 1191 191 1209 192 nw
rect 1679 191 1731 194
tri 1731 191 1742 194 nw
tri 607 188 612 191 ne
rect 612 189 631 191
tri 631 189 632 191 nw
tri 1679 189 1682 191 ne
rect 1682 189 1685 191
tri 612 188 631 189 nw
tri 1682 188 1683 189 ne
rect 1683 188 1685 189
tri 1683 187 1685 188 ne
tri 1685 187 1731 191 nw
tri 739 160 766 165 se
tri 766 161 781 165 sw
rect 766 160 781 161
rect 35 159 42 160
tri 42 159 71 160 sw
tri 737 159 739 160 se
rect 739 159 781 160
tri 781 159 784 161 sw
rect 35 125 36 159
rect 70 150 71 159
tri 71 150 82 159 sw
tri 723 157 737 159 se
rect 737 157 750 159
tri 690 150 723 157 se
rect 723 150 750 157
rect 70 125 82 150
rect 35 119 82 125
tri 82 119 93 150 sw
tri 684 149 689 150 se
rect 689 149 750 150
tri 661 145 684 149 se
rect 684 145 750 149
tri 655 143 661 145 se
rect 661 143 750 145
tri 271 140 402 141 se
tri 255 138 271 140 se
rect 271 138 402 140
tri 402 138 403 140 sw
tri 646 138 651 143 se
rect 651 138 750 143
tri 35 106 37 119 ne
rect 37 102 93 119
tri 93 102 100 119 sw
tri 37 100 38 102 ne
rect 38 100 66 102
tri 38 81 48 100 ne
rect 48 81 66 100
tri 48 70 58 81 ne
rect 58 70 66 81
tri 58 68 64 70 ne
rect 64 68 66 70
rect 162 102 196 118
rect 289 131 404 138
tri 404 131 408 138 sw
tri 638 131 645 138 se
rect 645 131 750 138
rect 289 120 408 131
tri 408 120 415 131 sw
rect 638 125 750 131
tri 1235 150 1237 157 se
tri 1233 145 1235 149 se
rect 1235 145 1237 150
tri 1001 143 1033 145 se
tri 1033 143 1037 145 sw
tri 942 141 1001 143 se
rect 1001 141 1037 143
tri 1037 141 1043 143 sw
tri 1232 141 1233 143 se
rect 1233 141 1237 145
tri 940 138 942 141 se
rect 942 138 1043 141
tri 1043 138 1054 141 sw
tri 1231 138 1232 141 se
rect 1232 138 1237 141
tri 934 125 940 138 se
rect 940 134 1054 138
tri 1054 134 1065 138 sw
tri 1230 134 1231 138 se
rect 1231 134 1237 138
rect 940 133 1065 134
tri 1065 133 1067 134 sw
rect 940 132 1067 133
tri 1067 132 1071 133 sw
rect 940 125 1037 132
rect 638 120 781 125
tri 781 120 784 125 nw
tri 932 120 934 125 se
rect 934 120 1037 125
rect 289 119 415 120
tri 415 119 416 120 sw
rect 289 104 416 119
tri 637 119 638 120 se
rect 638 119 780 120
tri 780 119 781 120 nw
tri 931 119 932 120 se
rect 932 119 1037 120
rect 637 118 780 119
rect 255 102 416 104
tri 254 80 255 102 se
rect 255 80 354 102
tri 254 68 266 80 ne
rect 266 68 354 80
rect 388 69 416 102
rect 388 68 414 69
tri 414 68 416 69 nw
rect 458 102 492 118
rect 637 110 776 118
tri 776 110 780 118 nw
rect 637 102 760 110
tri 760 102 776 110 nw
rect 842 102 876 118
tri 636 74 637 102 se
rect 637 74 650 102
tri 635 70 636 73 se
rect 636 70 650 74
rect 635 68 650 70
rect 684 90 737 102
tri 737 90 760 102 nw
rect 684 74 718 90
tri 718 74 737 90 nw
rect 684 71 714 74
tri 714 71 718 74 nw
rect 684 70 712 71
tri 712 70 714 71 nw
rect 684 68 710 70
tri 710 68 712 70 nw
tri 924 103 931 118 se
rect 931 103 1037 119
rect 924 102 1037 103
tri 924 74 930 102 ne
rect 930 74 946 102
tri 930 70 931 74 ne
rect 931 70 946 74
tri 931 68 932 70 ne
rect 932 68 946 70
rect 980 98 1037 102
tri 1226 120 1230 132 se
rect 1230 123 1237 134
tri 1271 147 1276 157 sw
rect 1271 123 1276 147
tri 1425 148 1426 149 se
tri 1424 138 1425 143 se
rect 1425 138 1426 148
rect 1230 122 1276 123
tri 1276 122 1278 138 sw
rect 1230 120 1278 122
tri 1225 118 1226 119 se
rect 1226 118 1278 120
tri 1420 121 1424 138 se
rect 1424 121 1426 138
rect 980 88 1070 98
tri 1070 88 1071 98 nw
rect 1138 102 1172 118
rect 980 78 1063 88
tri 1063 78 1070 88 nw
rect 980 74 1053 78
tri 1053 74 1063 78 nw
rect 980 70 1044 74
tri 1044 70 1053 74 nw
rect 980 68 1040 70
tri 1040 68 1044 70 nw
tri 1220 102 1225 118 se
rect 1225 108 1278 118
tri 1278 108 1279 118 sw
rect 1225 102 1279 108
rect 1330 102 1364 118
tri 1216 87 1220 101 se
rect 1220 87 1234 102
tri 1216 74 1217 87 ne
rect 1217 70 1234 87
tri 1217 68 1218 70 ne
rect 1218 68 1234 70
rect 1268 88 1279 102
tri 1279 88 1281 102 sw
rect 1268 71 1281 88
tri 1281 71 1283 87 sw
rect 1268 69 1282 71
tri 1282 70 1283 71 nw
rect 1268 68 1280 69
tri 1280 68 1282 69 nw
tri 1417 102 1420 118 se
rect 1420 115 1426 121
tri 1460 144 1465 149 sw
rect 1460 139 1465 144
tri 1465 139 1469 144 sw
tri 1622 139 1626 144 se
tri 1626 143 1657 144 sw
rect 1626 142 1657 143
tri 1657 142 1663 143 sw
rect 1626 139 1629 142
rect 1460 138 1469 139
tri 1469 138 1471 139 sw
tri 1621 138 1622 139 se
rect 1622 138 1629 139
rect 1460 129 1471 138
tri 1471 129 1481 138 sw
tri 1620 129 1621 138 se
rect 1621 129 1629 138
rect 1460 121 1481 129
tri 1481 121 1483 129 sw
rect 1460 115 1483 121
rect 1420 102 1483 115
tri 1483 110 1485 118 sw
tri 1483 103 1485 110 nw
tri 1413 78 1417 101 se
rect 1417 78 1434 102
tri 1413 71 1415 78 ne
rect 1415 71 1434 78
rect 162 18 196 68
tri 267 65 269 68 ne
rect 269 65 407 68
tri 407 65 413 68 nw
tri 269 63 271 65 ne
rect 271 64 406 65
tri 406 64 407 65 nw
rect 271 63 404 64
tri 404 63 406 64 nw
tri 271 61 347 63 ne
rect 347 61 399 63
tri 399 61 404 63 nw
tri 354 60 396 61 ne
tri 396 60 398 61 nw
rect 458 18 492 68
tri 636 65 639 68 ne
rect 639 65 706 68
tri 706 65 710 68 nw
rect 639 64 704 65
tri 704 64 706 65 nw
tri 639 61 643 64 ne
rect 643 62 702 64
tri 702 62 704 64 nw
rect 643 61 692 62
tri 692 61 702 62 nw
rect 842 18 876 68
rect 932 65 1035 68
tri 1035 65 1040 68 nw
rect 932 64 1030 65
tri 1030 64 1031 65 nw
rect 932 63 1023 64
tri 1023 63 1028 64 nw
tri 932 59 934 63 ne
rect 934 59 998 63
tri 998 59 1023 63 nw
rect 1138 18 1172 68
tri 1218 65 1221 68 ne
rect 1221 65 1279 68
tri 1279 65 1280 68 nw
rect 1221 64 1278 65
tri 1278 64 1279 65 nw
tri 1221 63 1222 64 ne
rect 1222 63 1278 64
tri 1222 57 1227 63 ne
rect 1227 62 1277 63
tri 1277 62 1278 63 nw
rect 1227 57 1264 62
tri 1264 57 1277 62 nw
tri 1227 56 1228 57 ne
rect 1228 56 1262 57
tri 1262 56 1264 57 nw
rect 1330 18 1364 68
tri 1415 65 1417 71 ne
rect 1417 68 1434 71
rect 1468 77 1476 102
tri 1476 78 1483 102 nw
rect 1530 102 1564 118
tri 1619 107 1620 118 se
rect 1620 108 1629 129
tri 1663 138 1664 142 sw
rect 1663 122 1664 138
tri 1664 122 1667 138 sw
tri 1928 157 1930 159 sw
rect 1928 154 1930 157
tri 1930 154 1935 157 sw
rect 1928 150 1935 154
tri 1935 150 1940 154 sw
tri 2115 150 2116 154 se
rect 1928 143 1940 150
tri 1940 143 1950 150 sw
tri 2113 143 2115 150 se
rect 2115 143 2116 150
rect 1928 133 1950 143
tri 1950 133 1956 143 sw
rect 1928 125 1956 133
rect 1663 108 1667 122
rect 1620 107 1667 108
rect 1619 104 1667 107
tri 1667 104 1671 122 sw
rect 1894 118 1956 125
tri 2107 119 2113 143 se
rect 2113 120 2116 143
tri 2150 129 2154 154 sw
rect 2150 120 2154 129
rect 2113 119 2154 120
tri 2106 118 2107 119 se
rect 2107 118 2154 119
rect 1619 102 1671 104
rect 1722 102 1756 118
rect 1468 68 1473 77
tri 1473 68 1476 77 nw
tri 1616 72 1619 102 se
rect 1619 72 1626 102
rect 1616 68 1626 72
rect 1660 95 1671 102
tri 1671 95 1673 102 sw
rect 1660 68 1672 95
tri 1672 74 1673 95 nw
rect 1417 67 1473 68
rect 1417 65 1472 67
tri 1472 65 1473 67 nw
rect 1530 18 1564 68
tri 1615 66 1616 68 se
rect 1616 66 1672 68
tri 1615 56 1625 66 ne
rect 1625 63 1672 66
rect 1625 56 1671 63
tri 1671 57 1672 63 nw
rect 1722 18 1756 68
rect 1826 102 1860 118
tri 1894 102 1895 118 ne
rect 1895 102 1956 118
tri 1895 72 1897 102 ne
rect 1897 72 1922 102
rect 1826 18 1860 68
tri 1897 64 1901 72 ne
rect 1901 68 1922 72
rect 2018 102 2052 118
tri 2102 102 2106 118 se
rect 2106 109 2154 118
tri 2154 109 2156 129 sw
rect 2106 102 2156 109
rect 2210 102 2244 118
tri 2096 79 2102 102 se
rect 2102 79 2114 102
tri 2096 68 2097 79 ne
rect 2097 68 2114 79
rect 2148 79 2156 102
tri 2156 79 2159 102 sw
rect 2148 68 2159 79
tri 2159 70 2160 79 sw
tri 2159 69 2160 70 nw
rect 1901 64 1923 68
tri 1923 64 1954 68 nw
tri 1903 63 1914 64 ne
tri 1914 63 1922 64 nw
rect 2018 18 2052 68
rect 2097 64 2156 68
tri 2156 64 2159 68 nw
tri 2097 57 2107 64 ne
rect 2107 58 2151 64
tri 2151 58 2156 64 nw
rect 2107 57 2145 58
tri 2145 57 2151 58 nw
tri 2107 56 2138 57 ne
tri 2138 56 2145 57 nw
rect 2210 18 2244 68
rect 0 -16 29 18
rect 63 -16 121 18
rect 155 -16 213 18
rect 247 -16 305 18
rect 339 -16 397 18
rect 431 -16 489 18
rect 523 -16 581 18
rect 615 -16 673 18
rect 707 -16 765 18
rect 799 -16 857 18
rect 891 -16 949 18
rect 983 -16 1041 18
rect 1075 -16 1133 18
rect 1167 -16 1225 18
rect 1259 -16 1317 18
rect 1351 -16 1409 18
rect 1443 -16 1501 18
rect 1535 -16 1593 18
rect 1627 -16 1685 18
rect 1719 -16 1777 18
rect 1811 -16 1869 18
rect 1903 -16 1961 18
rect 1995 -16 2053 18
rect 2087 -16 2145 18
rect 2179 -16 2237 18
rect 2271 -16 2329 18
rect 2363 -16 2392 18
<< viali >>
rect 29 528 63 562
rect 121 528 155 562
rect 213 528 247 562
rect 305 528 339 562
rect 397 528 431 562
rect 489 528 523 562
rect 581 528 615 562
rect 673 528 707 562
rect 765 528 799 562
rect 857 528 891 562
rect 949 528 983 562
rect 1041 528 1075 562
rect 1133 528 1167 562
rect 1225 528 1259 562
rect 1317 528 1351 562
rect 1409 528 1443 562
rect 1501 528 1535 562
rect 1593 528 1627 562
rect 1685 528 1719 562
rect 1777 528 1811 562
rect 1869 528 1903 562
rect 1961 528 1995 562
rect 2053 528 2087 562
rect 2145 528 2179 562
rect 2237 528 2271 562
rect 2329 528 2363 562
rect 35 408 69 422
rect 35 388 66 408
rect 66 388 69 408
rect 637 380 671 401
rect 855 380 889 413
rect 1333 417 1367 451
rect 1449 414 1468 437
rect 1468 414 1483 437
rect 289 307 323 341
rect 637 367 650 380
rect 650 367 671 380
rect 855 379 876 380
rect 876 379 889 380
rect 1449 403 1483 414
rect 1637 411 1671 445
rect 1717 414 1751 448
rect 1929 414 1963 448
rect 372 300 406 334
rect 757 304 791 338
rect 962 304 996 338
rect 1094 318 1128 352
rect 1795 346 1826 355
rect 1826 346 1829 355
rect 1449 300 1483 334
rect 1795 321 1829 346
rect 1933 334 1967 368
rect 576 253 610 287
rect 220 216 244 229
rect 244 216 254 229
rect 220 195 254 216
rect 436 211 470 245
rect 678 216 698 239
rect 698 216 712 239
rect 678 205 712 216
rect 865 224 899 258
rect 1071 216 1090 242
rect 1090 216 1105 242
rect 1071 208 1105 216
rect 1194 216 1220 232
rect 1220 216 1228 232
rect 1194 198 1228 216
rect 1730 258 1764 292
rect 2053 302 2087 336
rect 1449 216 1482 242
rect 1482 216 1483 242
rect 1976 250 2010 255
rect 2158 252 2192 286
rect 1976 221 2004 250
rect 2004 221 2010 250
rect 1449 208 1483 216
rect 36 125 70 159
rect 255 104 289 138
rect 750 125 784 159
rect 1037 98 1071 132
rect 1237 123 1271 157
rect 1426 115 1460 149
rect 1629 108 1663 142
rect 1894 125 1928 159
rect 2116 120 2150 154
rect 29 -16 63 18
rect 121 -16 155 18
rect 213 -16 247 18
rect 305 -16 339 18
rect 397 -16 431 18
rect 489 -16 523 18
rect 581 -16 615 18
rect 673 -16 707 18
rect 765 -16 799 18
rect 857 -16 891 18
rect 949 -16 983 18
rect 1041 -16 1075 18
rect 1133 -16 1167 18
rect 1225 -16 1259 18
rect 1317 -16 1351 18
rect 1409 -16 1443 18
rect 1501 -16 1535 18
rect 1593 -16 1627 18
rect 1685 -16 1719 18
rect 1777 -16 1811 18
rect 1869 -16 1903 18
rect 1961 -16 1995 18
rect 2053 -16 2087 18
rect 2145 -16 2179 18
rect 2237 -16 2271 18
rect 2329 -16 2363 18
<< metal1 >>
rect 0 562 2392 593
rect 0 528 29 562
rect 63 528 121 562
rect 155 528 213 562
rect 247 528 305 562
rect 339 528 397 562
rect 431 528 489 562
rect 523 528 581 562
rect 615 528 673 562
rect 707 528 765 562
rect 799 528 857 562
rect 891 528 949 562
rect 983 528 1041 562
rect 1075 528 1133 562
rect 1167 528 1225 562
rect 1259 528 1317 562
rect 1351 528 1409 562
rect 1443 528 1501 562
rect 1535 528 1593 562
rect 1627 528 1685 562
rect 1719 528 1777 562
rect 1811 528 1869 562
rect 1903 528 1961 562
rect 1995 528 2053 562
rect 2087 528 2145 562
rect 2179 528 2237 562
rect 2271 528 2329 562
rect 2363 528 2392 562
rect 0 497 2392 528
tri 1329 452 1331 455 se
rect 1331 452 1369 455
tri 1369 452 1371 455 sw
rect 1329 451 1371 452
tri 793 425 856 430 se
tri 856 426 874 430 sw
rect 856 425 874 426
tri 31 423 35 425 se
rect 35 423 70 425
tri 70 423 72 425 sw
tri 759 423 789 425 se
rect 789 423 874 425
rect 31 422 72 423
tri 30 388 31 415 se
rect 31 400 35 422
rect 69 416 72 422
tri 668 417 759 423 se
rect 759 417 874 423
tri 874 417 891 426 sw
tri 72 416 73 417 sw
tri 653 416 668 417 se
rect 668 416 891 417
tri 891 416 893 417 sw
rect 69 400 73 416
tri 651 415 653 416 se
rect 653 415 893 416
tri 636 405 651 415 se
rect 651 413 893 415
rect 651 405 855 413
tri 633 403 635 405 se
rect 635 403 855 405
rect 633 401 855 403
rect 31 388 33 400
rect 30 348 33 388
rect 633 367 637 401
rect 671 379 855 401
rect 889 379 893 413
tri 1326 443 1329 450 se
rect 1329 443 1333 451
rect 1077 435 1079 440
tri 1079 435 1118 440 sw
rect 1077 430 1118 435
tri 1118 430 1132 435 sw
rect 1077 426 1132 430
tri 1132 426 1142 430 sw
rect 1077 417 1142 426
tri 1142 417 1164 426 sw
rect 1367 417 1371 451
tri 1673 449 1715 453 se
tri 1634 447 1636 449 se
rect 1636 448 1715 449
rect 1636 447 1643 448
tri 1443 443 1449 446 se
tri 1449 445 1463 446 sw
rect 1633 445 1643 447
rect 1449 443 1463 445
tri 1463 443 1493 445 sw
tri 1440 434 1443 443 se
rect 1443 437 1495 443
rect 1443 434 1449 437
rect 1077 416 1164 417
tri 1164 416 1167 417 sw
rect 1077 408 1167 416
tri 1167 408 1188 416 sw
tri 1077 407 1110 408 ne
rect 1110 407 1188 408
tri 1188 407 1190 408 sw
tri 1112 405 1118 407 ne
rect 1118 405 1190 407
tri 1118 403 1122 405 ne
rect 1122 403 1190 405
tri 1190 403 1200 407 sw
tri 1122 398 1134 403 ne
rect 1134 398 1200 403
tri 1134 390 1155 398 ne
rect 1155 390 1200 398
tri 1200 390 1234 403 sw
rect 1362 415 1371 417
rect 1362 413 1369 415
tri 1369 413 1371 415 nw
tri 1439 426 1440 434 se
rect 1440 426 1449 434
tri 1439 413 1441 426 ne
rect 1441 410 1449 426
tri 1441 409 1442 410 ne
rect 1442 403 1449 410
rect 1483 436 1495 437
tri 1495 436 1516 443 sw
rect 1483 403 1497 436
tri 1442 402 1443 403 ne
rect 1443 402 1497 403
tri 1443 400 1444 402 ne
rect 1444 400 1497 402
tri 1444 399 1445 400 ne
rect 1445 399 1497 400
tri 1445 398 1448 399 ne
rect 1448 398 1497 399
tri 1448 396 1453 398 ne
rect 1453 396 1497 398
tri 1453 393 1497 396 ne
rect 671 377 890 379
rect 671 375 743 377
tri 743 375 755 377 nw
tri 830 375 853 377 ne
rect 853 375 890 377
tri 890 375 893 379 nw
tri 1155 375 1194 390 ne
rect 1194 375 1234 390
rect 671 372 703 375
tri 703 372 743 375 nw
tri 1194 372 1204 375 ne
rect 1204 372 1234 375
rect 671 367 688 372
rect 633 366 688 367
tri 688 366 703 372 nw
tri 633 364 634 366 ne
rect 634 364 681 366
rect 30 346 75 348
rect 30 341 72 346
tri 72 341 75 346 nw
rect 304 344 325 345
tri 325 344 327 345 sw
rect 304 341 327 344
rect 30 335 68 341
tri 68 335 72 341 nw
rect 30 326 63 335
tri 63 326 68 335 nw
rect 30 319 61 326
tri 61 319 63 326 nw
tri 29 307 30 317 se
rect 30 307 59 319
tri 59 308 61 319 nw
rect 29 303 58 307
tri 58 303 59 307 nw
rect 323 307 327 341
rect 29 283 57 303
tri 57 300 58 303 nw
rect 304 306 327 307
rect 304 304 326 306
tri 326 304 327 306 nw
tri 368 336 370 338 se
rect 370 336 384 338
rect 368 334 384 336
rect 304 303 325 304
tri 325 303 326 304 nw
rect 368 300 372 334
rect 635 363 681 364
tri 681 363 688 366 nw
tri 638 362 648 363 ne
rect 648 362 679 363
tri 679 362 681 363 nw
tri 558 338 561 342 sw
tri 753 340 755 342 se
rect 755 340 793 342
tri 793 340 795 342 sw
rect 753 338 795 340
rect 558 321 561 338
tri 561 321 575 338 sw
rect 558 319 575 321
tri 575 319 577 321 sw
rect 558 312 577 319
tri 534 304 547 312 ne
rect 547 304 577 312
tri 577 304 588 319 sw
rect 753 304 757 338
rect 791 304 795 338
tri 1204 366 1219 372 ne
rect 1219 368 1234 372
tri 1234 368 1291 390 sw
rect 1633 411 1637 445
rect 1633 410 1643 411
tri 1633 407 1636 410 ne
rect 1636 407 1643 410
rect 1695 408 1715 448
tri 1695 406 1699 408 nw
tri 1972 433 1988 444 sw
rect 1972 430 1988 433
tri 1988 430 2004 433 sw
rect 1972 413 2004 430
tri 2004 413 2081 430 sw
rect 1972 410 2081 413
tri 2081 410 2091 413 sw
rect 1972 404 2091 410
rect 1928 403 2091 404
tri 1928 402 1929 403 ne
rect 1929 402 2091 403
rect 1928 400 2091 402
tri 2091 400 2136 410 sw
rect 1929 396 2136 400
tri 2136 396 2157 400 sw
rect 1929 393 2157 396
tri 2157 393 2159 396 sw
rect 1929 389 2159 393
rect 1929 384 1975 389
tri 1975 384 2054 389 nw
tri 2054 384 2076 389 ne
rect 2076 388 2159 389
tri 2159 388 2164 393 sw
rect 2076 384 2164 388
rect 1929 381 1972 384
tri 1972 381 1975 384 nw
tri 2076 381 2087 384 ne
rect 2087 381 2164 384
rect 1929 368 1971 381
tri 1971 377 1972 381 nw
tri 2087 377 2106 381 ne
rect 2106 377 2164 381
tri 2164 377 2168 388 sw
rect 2107 376 2168 377
rect 1219 366 1291 368
tri 1219 363 1226 366 ne
rect 1226 363 1291 366
tri 1226 362 1228 363 ne
rect 1228 362 1291 363
tri 1229 361 1231 362 ne
rect 1231 361 1291 362
tri 1291 361 1310 368 sw
tri 1231 358 1240 361 ne
rect 1240 360 1310 361
tri 1310 360 1317 361 sw
rect 1240 358 1317 360
tri 1240 357 1241 358 ne
rect 1241 357 1317 358
tri 1243 356 1244 357 ne
rect 1244 356 1317 357
tri 1091 355 1093 356 se
rect 1093 355 1130 356
tri 1244 355 1246 356 ne
rect 1246 355 1317 356
tri 1317 355 1341 360 sw
tri 1791 357 1794 359 se
rect 1794 357 1831 359
tri 1831 357 1833 359 sw
tri 1790 355 1791 357 se
rect 1791 355 1833 357
tri 1088 354 1091 355 se
rect 1091 354 1130 355
tri 1130 354 1131 355 sw
tri 1087 353 1088 354 se
rect 1088 353 1132 354
rect 1087 352 1132 353
tri 1086 351 1087 352 se
rect 1087 351 1094 352
rect 1086 349 1094 351
rect 1128 349 1132 352
tri 1246 351 1258 355 ne
rect 1258 351 1341 355
tri 1258 349 1262 351 ne
rect 1262 349 1341 351
rect 1086 348 1087 349
tri 961 345 967 348 sw
rect 961 342 967 345
tri 967 342 974 345 sw
rect 961 339 998 342
tri 998 339 1000 342 sw
rect 961 338 1000 339
rect 961 316 962 338
tri 951 314 954 316 ne
rect 954 314 962 316
tri 954 312 955 314 ne
rect 955 311 962 314
tri 955 304 957 311 ne
rect 957 304 962 311
rect 996 304 1000 338
tri 547 303 549 304 ne
rect 549 303 588 304
tri 588 303 589 304 sw
tri 549 302 550 303 ne
rect 368 299 384 300
tri 368 296 370 299 ne
rect 370 296 384 299
rect 550 300 589 303
tri 589 300 591 303 sw
rect 753 302 795 304
tri 957 303 958 304 ne
rect 753 300 793 302
tri 793 300 795 302 nw
rect 958 302 1000 304
tri 958 300 960 302 ne
rect 960 300 998 302
tri 998 300 1000 302 nw
tri 1262 331 1310 349 ne
rect 1310 342 1341 349
tri 1341 342 1405 355 sw
tri 1787 349 1790 355 se
rect 1790 354 1795 355
rect 1829 354 1833 355
tri 1833 354 1834 357 sw
rect 1790 349 1794 354
tri 1422 344 1473 346 se
tri 1473 344 1475 346 sw
tri 1777 344 1787 349 se
rect 1787 344 1794 349
tri 1405 342 1422 344 se
rect 1422 342 1475 344
rect 1310 338 1475 342
tri 1475 338 1484 344 sw
tri 1774 342 1777 344 se
rect 1777 342 1794 344
tri 1767 338 1774 342 se
rect 1774 338 1794 342
rect 1310 336 1485 338
tri 1485 336 1487 338 sw
rect 1310 334 1487 336
rect 1310 331 1449 334
tri 1310 328 1317 331 ne
rect 1317 328 1449 331
tri 1317 321 1348 328 ne
rect 1348 321 1449 328
tri 1348 319 1357 321 ne
rect 1357 319 1449 321
tri 1357 318 1361 319 ne
rect 1361 318 1449 319
tri 550 299 551 300 ne
rect 551 299 591 300
tri 551 296 552 299 ne
rect 552 294 591 299
rect 553 293 591 294
tri 591 293 597 300 sw
rect 753 297 792 300
tri 792 297 793 300 nw
tri 1361 304 1418 318 ne
rect 1418 304 1449 318
tri 1418 303 1421 304 ne
rect 1421 303 1449 304
tri 1421 300 1435 303 ne
rect 1435 300 1449 303
rect 1483 300 1487 334
tri 1749 328 1767 338 se
rect 1767 328 1794 338
tri 1743 324 1749 328 se
rect 1749 324 1794 328
tri 1740 321 1743 324 se
rect 1743 321 1794 324
rect 1929 334 1933 368
rect 1967 363 1971 368
tri 1971 363 1972 376 sw
rect 1967 348 1972 363
tri 2107 361 2126 376 ne
rect 2126 361 2168 376
tri 2126 360 2128 361 ne
rect 2128 360 2168 361
tri 2168 360 2173 377 sw
tri 1972 348 1973 360 sw
rect 1967 340 1973 348
tri 2128 346 2147 360 ne
rect 2147 346 2173 360
tri 2173 346 2178 360 sw
tri 2147 344 2148 346 ne
rect 2148 342 2178 346
tri 2148 340 2149 342 ne
rect 2149 341 2178 342
tri 2178 341 2180 346 sw
rect 1967 334 1974 340
tri 2049 337 2052 340 se
rect 2052 338 2091 340
tri 2091 338 2092 340 sw
rect 2052 337 2093 338
rect 2149 337 2180 341
rect 2049 336 2093 337
rect 1929 333 1974 334
tri 1929 328 1930 333 ne
rect 1930 328 1974 333
tri 1974 328 1975 336 sw
tri 1930 324 1932 328 ne
rect 1932 324 1971 328
tri 1932 323 1933 324 ne
rect 1933 323 1971 324
tri 1971 323 1975 328 nw
tri 1933 322 1935 323 ne
tri 1935 322 1971 323 nw
tri 1729 303 1740 320 se
rect 1740 303 1794 321
rect 1729 302 1794 303
rect 2049 302 2053 336
rect 2087 323 2093 336
tri 2093 323 2096 337 sw
tri 2149 324 2151 337 ne
rect 2087 302 2096 323
rect 2151 322 2180 337
tri 1435 297 1446 300 ne
rect 1446 298 1487 300
rect 1446 297 1485 298
rect 753 296 791 297
tri 791 296 792 297 nw
tri 1446 296 1452 297 ne
rect 1452 296 1485 297
tri 1485 296 1487 298 nw
tri 1726 298 1729 302 se
rect 1729 298 1814 302
tri 1814 298 1821 302 nw
rect 2049 300 2096 302
tri 2096 300 2101 322 sw
tri 2151 301 2153 322 ne
rect 2153 300 2180 322
tri 2049 298 2052 300 ne
rect 2052 298 2101 300
tri 2101 298 2102 300 sw
rect 1726 297 1813 298
tri 1813 297 1814 298 nw
rect 2052 297 2102 298
tri 2153 297 2154 300 ne
tri 1725 296 1726 297 se
rect 1726 296 1811 297
tri 1811 296 1813 297 nw
tri 2052 296 2054 297 ne
rect 2054 296 2102 297
tri 753 294 754 296 ne
rect 553 292 597 293
tri 553 287 556 292 ne
rect 556 291 597 292
tri 597 291 601 293 sw
rect 754 291 791 296
rect 1725 295 1810 296
rect 1725 294 1807 295
tri 1807 294 1810 295 nw
rect 2055 295 2102 296
tri 2055 294 2056 295 ne
rect 1725 292 1805 294
tri 1805 292 1807 294 nw
rect 2056 292 2102 295
tri 2102 292 2103 294 sw
rect 556 289 612 291
tri 612 289 614 291 sw
rect 556 287 614 289
tri 57 283 58 287 sw
rect 29 195 58 283
tri 556 272 563 287 ne
rect 563 272 576 287
tri 563 254 572 272 ne
rect 572 253 576 272
rect 610 253 614 287
tri 754 272 758 291 ne
rect 758 278 791 291
tri 791 278 792 292 sw
rect 758 270 792 278
tri 758 264 759 270 ne
rect 759 266 792 270
tri 792 266 793 270 sw
tri 572 249 576 253 ne
rect 576 252 614 253
rect 576 249 610 252
tri 610 249 614 252 nw
rect 759 262 793 266
tri 863 262 873 264 se
tri 759 250 762 262 ne
tri 432 247 434 249 se
rect 434 247 472 249
tri 472 247 474 249 sw
tri 429 245 432 247 se
rect 432 245 474 247
tri 428 244 429 245 se
rect 429 244 436 245
tri 29 167 30 195 ne
rect 30 184 58 195
tri 58 184 59 195 sw
tri 301 237 428 244 se
rect 428 237 436 244
tri 276 235 301 237 se
rect 301 235 436 237
tri 259 234 276 235 se
rect 276 234 436 235
tri 238 233 259 234 se
rect 259 233 436 234
tri 209 232 214 233 se
rect 214 232 436 233
tri 201 231 203 232 sw
tri 203 231 209 232 se
rect 209 231 436 232
rect 201 229 436 231
rect 201 195 220 229
rect 254 214 436 229
rect 254 213 419 214
tri 419 213 426 214 nw
tri 426 213 429 214 ne
rect 429 213 436 214
rect 254 211 396 213
tri 396 211 419 213 nw
rect 254 210 384 211
tri 384 210 396 211 nw
tri 429 210 432 213 ne
rect 432 211 436 213
rect 470 211 474 245
rect 432 210 474 211
rect 254 207 361 210
tri 361 207 384 210 nw
tri 432 207 434 210 ne
rect 434 207 472 210
tri 472 207 474 210 nw
rect 762 249 793 262
tri 861 260 863 262 se
rect 863 260 873 262
rect 861 258 873 260
rect 925 260 926 262
tri 926 260 936 262 sw
rect 925 258 936 260
tri 936 258 942 260 sw
rect 1725 258 1730 292
rect 1764 291 1803 292
tri 1803 291 1804 292 nw
rect 2056 291 2103 292
rect 1764 288 1797 291
tri 1797 288 1803 291 nw
tri 2056 288 2057 291 ne
rect 2057 288 2103 291
tri 2103 288 2104 292 sw
rect 1764 286 1794 288
tri 1794 286 1797 288 nw
rect 2057 286 2104 288
rect 2154 291 2180 300
tri 2154 288 2155 291 ne
rect 2155 290 2180 291
tri 2180 290 2196 340 sw
tri 2154 287 2155 288 se
rect 2155 287 2196 290
rect 2154 286 2196 287
rect 1764 281 1785 286
tri 1785 281 1794 286 nw
tri 2057 281 2060 286 ne
rect 2060 281 2104 286
rect 1764 275 1779 281
tri 1779 275 1785 281 nw
rect 1764 272 1778 275
tri 1778 272 1779 275 nw
rect 1764 260 1773 272
tri 1773 260 1778 272 nw
tri 2060 260 2067 281 ne
rect 1764 258 1771 260
tri 1771 258 1773 260 nw
rect 2067 259 2104 281
tri 1972 258 1975 259 se
rect 1975 258 2012 259
tri 762 244 763 249 ne
rect 710 241 714 243
tri 714 241 716 243 sw
rect 710 239 716 241
rect 254 205 342 207
tri 342 205 361 207 nw
rect 712 205 716 239
rect 763 241 793 249
tri 763 226 766 241 ne
rect 766 226 793 241
tri 793 226 797 253 sw
rect 766 224 797 226
rect 861 224 865 258
rect 925 256 942 258
tri 942 256 949 258 sw
tri 1725 256 1726 258 ne
rect 1726 256 1770 258
tri 1770 256 1771 258 nw
rect 925 255 949 256
tri 949 255 953 256 sw
rect 925 254 953 255
tri 953 254 958 255 sw
tri 1726 254 1728 256 ne
rect 1728 255 1769 256
tri 1769 255 1770 256 nw
rect 1728 254 1767 255
tri 1767 254 1769 255 nw
tri 1968 254 1972 258 se
rect 1972 257 2012 258
tri 2012 257 2014 259 sw
rect 1972 255 2014 257
tri 2067 256 2068 259 ne
rect 2068 255 2104 259
rect 1972 254 1976 255
rect 925 253 970 254
tri 970 253 981 254 sw
rect 1729 253 1766 254
tri 1766 253 1767 254 nw
rect 925 252 981 253
tri 981 252 1009 253 sw
tri 1967 252 1968 253 se
rect 1968 252 1976 254
rect 925 251 1009 252
tri 1009 251 1054 252 sw
tri 1957 251 1967 252 se
rect 1967 251 1976 252
rect 925 250 1098 251
tri 1098 250 1100 251 sw
tri 1951 250 1956 251 se
rect 1956 250 1976 251
rect 925 249 1100 250
tri 1100 249 1101 250 sw
rect 925 248 1102 249
tri 1102 248 1103 249 sw
rect 925 246 1103 248
tri 1103 246 1107 248 sw
rect 925 244 1108 246
tri 1108 244 1109 246 sw
rect 925 242 1109 244
rect 925 227 1071 242
rect 899 226 1071 227
rect 899 224 908 226
tri 908 224 957 226 nw
tri 957 224 967 226 ne
rect 967 224 1071 226
tri 766 221 767 224 ne
rect 767 220 797 224
tri 797 220 798 224 sw
rect 861 222 903 224
tri 903 222 908 224 nw
tri 967 222 975 224 ne
rect 975 222 1071 224
tri 861 220 863 222 ne
rect 863 220 900 222
tri 900 220 903 222 nw
tri 975 220 987 222 ne
rect 987 220 1071 222
tri 767 211 769 220 ne
rect 769 212 798 220
tri 798 212 799 220 sw
tri 987 212 1028 220 ne
rect 1028 212 1071 220
rect 769 208 799 212
tri 799 208 801 212 sw
tri 769 207 770 208 ne
rect 254 201 303 205
tri 303 201 342 205 nw
rect 254 199 280 201
tri 280 199 303 201 nw
rect 254 197 264 199
tri 264 197 280 199 nw
rect 710 203 716 205
rect 710 201 714 203
tri 714 201 716 203 nw
rect 770 205 801 208
tri 801 205 804 208 sw
tri 1028 207 1053 212 ne
rect 1053 208 1071 212
rect 1105 208 1109 242
tri 1445 242 1447 246 se
tri 1947 249 1951 250 se
rect 1951 249 1976 250
tri 1938 248 1944 249 se
rect 1944 248 1976 249
tri 1925 246 1938 248 se
rect 1938 246 1976 248
tri 1915 245 1919 246 se
rect 1919 245 1976 246
tri 1909 244 1915 245 se
rect 1915 244 1976 245
tri 1499 242 1520 244 sw
tri 1896 242 1909 244 se
rect 1909 242 1976 244
tri 1191 235 1199 238 se
tri 1199 237 1250 238 sw
rect 1199 235 1250 237
tri 1250 235 1255 237 sw
tri 1190 233 1191 235 se
rect 1191 233 1255 235
rect 1190 232 1255 233
rect 1053 207 1109 208
tri 1053 205 1064 207 ne
rect 1064 205 1107 207
rect 770 204 804 205
tri 804 204 806 205 sw
tri 1064 204 1069 205 ne
rect 1069 204 1107 205
tri 1107 204 1109 207 nw
tri 1188 228 1190 232 se
rect 1190 228 1194 232
tri 770 202 771 204 ne
rect 771 201 806 204
tri 806 201 815 204 sw
rect 771 199 815 201
tri 815 199 820 201 sw
rect 771 197 820 199
tri 820 197 824 199 sw
rect 1188 198 1194 228
rect 1228 228 1255 232
tri 1255 228 1279 235 sw
rect 1228 219 1279 228
tri 1279 219 1311 228 sw
rect 1228 208 1311 219
tri 1311 208 1330 219 sw
rect 1228 207 1330 208
tri 1330 207 1332 208 sw
rect 1228 204 1332 207
tri 1332 204 1339 207 sw
rect 1445 206 1447 242
rect 1499 224 1520 242
tri 1520 224 1746 242 sw
tri 1774 226 1896 242 se
rect 1896 226 1976 242
tri 1746 224 1774 226 se
rect 1774 224 1976 226
rect 1499 221 1976 224
rect 2010 221 2014 255
tri 2014 254 2015 255 nw
tri 2068 254 2069 255 ne
rect 2069 254 2104 255
tri 2104 254 2111 286 sw
rect 2069 252 2111 254
rect 2154 252 2158 286
rect 2192 252 2196 286
tri 2069 250 2070 252 ne
rect 2070 250 2111 252
tri 2111 250 2112 252 sw
tri 2070 249 2071 250 ne
rect 1499 219 2014 221
rect 1499 217 2012 219
tri 2012 217 2014 219 nw
rect 2071 248 2112 250
rect 2154 250 2196 252
tri 2154 249 2155 250 ne
rect 2155 249 2194 250
tri 2112 248 2113 249 sw
tri 2155 248 2157 249 ne
rect 2157 248 2194 249
tri 2194 248 2196 250 nw
tri 2071 217 2081 248 ne
rect 2081 217 2113 248
tri 1445 204 1447 206 ne
rect 1228 201 1339 204
tri 1339 201 1343 204 sw
rect 1228 200 1343 201
tri 1343 200 1345 201 sw
rect 1228 199 1257 200
tri 1257 199 1264 200 nw
tri 1272 199 1278 200 ne
rect 1278 199 1345 200
tri 1345 199 1348 200 sw
rect 1228 198 1249 199
tri 1188 197 1189 198 ne
rect 1189 197 1249 198
tri 1249 197 1257 199 nw
tri 1278 197 1284 199 ne
rect 1284 198 1348 199
tri 1348 198 1349 199 sw
rect 1499 207 1897 217
tri 1897 207 1998 217 nw
tri 2081 207 2085 217 ne
rect 1499 206 1882 207
tri 1882 206 1897 207 nw
rect 2085 206 2113 217
rect 1499 204 1859 206
tri 1859 204 1882 206 nw
tri 2085 204 2086 206 ne
rect 2086 204 2113 206
rect 1499 203 1835 204
tri 1499 201 1555 203 ne
rect 1555 201 1835 203
tri 1835 201 1859 204 nw
tri 2086 201 2087 204 ne
rect 2087 201 2113 204
tri 1555 200 1585 201 ne
rect 1585 200 1810 201
tri 1585 199 1626 200 ne
rect 1626 199 1810 200
tri 1810 199 1835 201 nw
tri 2087 199 2088 201 ne
rect 1649 198 1797 199
tri 1797 198 1810 199 nw
rect 1284 197 1349 198
rect 254 195 258 197
tri 213 194 214 195 ne
rect 214 194 258 195
tri 258 194 264 197 nw
rect 771 196 824 197
tri 824 196 829 197 sw
tri 1189 196 1191 197 ne
rect 1191 196 1241 197
tri 1241 196 1249 197 nw
tri 1284 196 1290 197 ne
rect 1290 196 1349 197
rect 771 195 829 196
tri 829 195 831 196 sw
rect 771 194 831 195
tri 831 194 834 195 sw
tri 1191 194 1193 196 ne
rect 1193 195 1241 196
tri 1290 195 1294 196 ne
rect 1294 195 1349 196
tri 1349 195 1355 198 sw
tri 1626 197 1649 198 ne
tri 1649 197 1673 198 ne
rect 1673 197 1793 198
tri 1793 197 1797 198 nw
rect 2088 197 2113 201
tri 1673 195 1750 197 ne
rect 1750 195 1766 197
tri 1766 195 1793 197 nw
tri 2088 195 2089 197 ne
tri 216 191 219 194 ne
rect 219 191 256 194
tri 256 191 258 194 nw
rect 771 193 834 194
tri 770 191 771 193 se
rect 771 191 837 193
tri 837 191 840 193 sw
tri 767 184 770 191 se
rect 770 184 840 191
tri 840 184 859 191 sw
rect 30 167 59 184
tri 59 167 67 184 sw
tri 760 168 767 184 se
rect 767 168 918 184
tri 30 161 31 167 ne
rect 31 165 67 167
tri 67 165 68 167 sw
tri 754 166 760 168 se
rect 760 166 918 168
tri 753 165 754 166 se
rect 754 165 918 166
rect 31 162 68 165
tri 68 162 73 165 sw
tri 748 163 753 165 se
rect 753 163 918 165
rect 31 161 73 162
tri 73 161 74 162 sw
tri 746 161 748 163 se
rect 748 161 918 163
rect 31 159 74 161
tri 74 159 75 161 sw
rect 31 125 36 159
rect 70 125 75 159
rect 746 159 918 161
tri 31 123 32 125 ne
rect 32 123 75 125
tri 32 120 37 123 ne
rect 37 120 70 123
tri 70 120 75 123 nw
tri 251 140 253 142 se
rect 253 140 255 142
rect 251 103 255 140
tri 307 139 605 140 se
tri 605 139 610 140 sw
rect 307 135 610 139
tri 610 135 639 139 sw
rect 307 112 637 135
rect 307 109 476 112
tri 476 109 600 112 nw
tri 600 109 610 112 ne
rect 610 109 637 112
rect 307 107 352 109
tri 352 107 476 109 nw
tri 610 107 616 109 ne
rect 616 107 637 109
rect 307 104 330 107
tri 330 104 352 107 nw
tri 251 100 253 103 ne
rect 253 100 255 103
tri 307 101 330 104 nw
tri 616 101 628 107 ne
rect 628 101 637 107
tri 628 100 631 101 ne
rect 631 100 637 101
tri 631 98 636 100 ne
rect 636 98 637 100
rect 746 125 750 159
rect 784 154 918 159
rect 784 153 884 154
tri 884 153 918 154 nw
rect 784 152 847 153
tri 847 152 884 153 nw
rect 784 151 824 152
tri 824 151 847 152 nw
rect 784 149 821 151
tri 821 149 824 151 nw
rect 784 135 796 149
tri 796 135 821 149 nw
rect 1193 193 1238 195
tri 1194 191 1195 193 ne
rect 1195 191 1238 193
tri 1238 192 1241 195 nw
tri 1294 194 1295 195 ne
rect 1295 194 1355 195
tri 1355 194 1356 195 sw
tri 1750 194 1762 195 ne
tri 1762 194 1766 195 nw
tri 1298 193 1299 194 ne
rect 1299 193 1356 194
tri 1356 193 1358 194 sw
rect 2089 193 2113 197
tri 1301 191 1303 193 ne
rect 1303 192 1358 193
tri 1358 192 1361 193 sw
tri 2089 192 2090 193 ne
rect 1303 191 1361 192
tri 1303 187 1309 191 ne
rect 1309 187 1361 191
tri 1309 184 1314 187 ne
rect 1314 184 1361 187
tri 1361 184 1375 192 sw
rect 2090 191 2113 193
tri 2090 184 2093 191 ne
rect 2093 190 2113 191
tri 2113 190 2125 248 sw
rect 2093 184 2125 190
tri 1315 168 1339 184 ne
rect 1339 168 1375 184
tri 1339 167 1341 168 ne
rect 1341 167 1375 168
tri 1375 167 1406 184 sw
tri 2093 167 2098 184 ne
rect 2098 182 2125 184
tri 2125 182 2129 190 sw
rect 2098 167 2129 182
tri 1342 166 1344 167 ne
rect 1344 166 1406 167
tri 1406 166 1409 167 sw
tri 2098 166 2099 167 ne
rect 1344 165 1409 166
tri 1344 162 1350 165 ne
rect 1350 163 1409 165
tri 1409 163 1414 166 sw
rect 2099 163 2129 167
rect 1350 162 1414 163
tri 1414 162 1416 163 sw
tri 1350 161 1351 162 ne
rect 1351 161 1416 162
tri 1416 161 1417 162 sw
tri 1890 161 1892 163 se
rect 1892 162 1929 163
tri 1929 162 1930 163 sw
tri 2099 162 2100 163 ne
rect 1892 161 1930 162
tri 1930 161 1932 162 sw
tri 1352 159 1354 161 ne
rect 1354 159 1419 161
tri 1419 159 1422 161 sw
tri 1354 158 1356 159 ne
rect 1356 158 1422 159
tri 1422 158 1424 159 sw
tri 1883 158 1889 161 se
rect 1889 159 1932 161
rect 1889 158 1894 159
tri 1356 157 1357 158 ne
rect 1357 157 1424 158
tri 1035 153 1041 156 se
tri 1041 154 1079 156 sw
rect 1041 153 1079 154
rect 784 132 791 135
tri 791 133 796 135 nw
tri 1033 134 1035 135 se
rect 1035 134 1079 153
rect 784 125 788 132
rect 746 123 788 125
tri 788 123 791 132 nw
rect 1033 132 1079 134
tri 746 121 748 123 ne
rect 748 121 785 123
tri 785 121 788 123 nw
rect 1033 98 1037 132
rect 1071 104 1079 132
tri 1357 149 1371 157 ne
rect 1371 155 1424 157
tri 1424 155 1428 158 sw
tri 1875 156 1883 158 se
rect 1883 156 1894 158
rect 1371 153 1428 155
tri 1428 153 1456 155 sw
rect 1371 152 1456 153
tri 1456 152 1461 153 sw
rect 1371 151 1462 152
tri 1462 151 1463 152 sw
rect 1371 149 1463 151
tri 1463 149 1466 151 sw
tri 1371 146 1375 149 ne
rect 1375 146 1426 149
tri 1375 144 1379 146 ne
rect 1379 144 1426 146
tri 1379 141 1383 144 ne
rect 1383 141 1426 144
tri 1383 124 1411 141 ne
rect 1411 124 1426 141
tri 1411 123 1412 124 ne
rect 1412 123 1426 124
tri 1412 121 1415 123 ne
rect 1415 121 1426 123
tri 1415 120 1417 121 ne
rect 1417 120 1426 121
tri 1417 119 1418 120 ne
rect 1418 119 1426 120
tri 1418 116 1420 119 ne
rect 1420 115 1426 119
rect 1460 146 1466 149
tri 1466 146 1471 149 sw
rect 1460 143 1471 146
tri 1471 143 1480 146 sw
rect 1460 115 1478 143
tri 1420 112 1423 115 ne
rect 1423 112 1478 115
tri 1423 111 1425 112 ne
rect 1425 111 1478 112
tri 1437 108 1450 111 ne
rect 1450 108 1478 111
tri 1450 105 1464 108 ne
rect 1464 105 1478 108
rect 1071 103 1115 104
tri 1115 103 1119 104 nw
tri 1464 103 1476 105 ne
rect 1476 103 1478 105
rect 1071 101 1109 103
tri 1109 101 1115 103 nw
tri 1476 102 1478 103 ne
rect 1071 98 1097 101
tri 1097 98 1109 101 nw
rect 1033 96 1092 98
tri 1092 96 1097 98 nw
tri 1033 90 1035 96 ne
rect 1035 90 1071 96
tri 1071 90 1092 96 nw
tri 1666 144 1667 145 sw
rect 1666 126 1667 144
tri 1667 126 1668 136 sw
rect 1666 112 1668 126
rect 1666 106 1667 112
tri 1667 111 1668 112 nw
tri 1666 105 1667 106 nw
rect 1882 125 1894 156
rect 1928 125 1932 159
rect 2100 161 2129 163
tri 2100 155 2102 161 ne
rect 2102 158 2129 161
tri 2129 158 2152 182 sw
rect 2102 155 2152 158
tri 2152 155 2155 158 sw
rect 2102 154 2110 155
tri 2102 132 2110 154 ne
rect 1882 123 1932 125
rect 1882 121 1929 123
tri 1929 121 1932 123 nw
rect 1882 120 1903 121
tri 1903 120 1906 121 nw
rect 1882 118 1891 120
tri 1891 118 1901 120 nw
tri 1882 116 1891 118 nw
tri 1036 88 1067 90 ne
rect 1067 89 1068 90
tri 1068 89 1071 90 nw
tri 1067 88 1068 89 nw
rect 0 18 2392 49
rect 0 -16 29 18
rect 63 -16 121 18
rect 155 -16 213 18
rect 247 -16 305 18
rect 339 -16 397 18
rect 431 -16 489 18
rect 523 -16 581 18
rect 615 -16 673 18
rect 707 -16 765 18
rect 799 -16 857 18
rect 891 -16 949 18
rect 983 -16 1041 18
rect 1075 -16 1133 18
rect 1167 -16 1225 18
rect 1259 -16 1317 18
rect 1351 -16 1409 18
rect 1443 -16 1501 18
rect 1535 -16 1593 18
rect 1627 -16 1685 18
rect 1719 -16 1777 18
rect 1811 -16 1869 18
rect 1903 -16 1961 18
rect 1995 -16 2053 18
rect 2087 -16 2145 18
rect 2179 -16 2237 18
rect 2271 -16 2329 18
rect 2363 -16 2392 18
rect 0 -47 2392 -16
<< via1 >>
rect 33 388 35 400
rect 35 388 69 400
rect 69 388 85 400
rect 33 348 85 388
rect 1025 398 1077 450
rect 1310 417 1333 443
rect 1333 417 1362 443
rect 1715 448 1767 457
rect 1643 445 1695 448
rect 1310 391 1362 417
rect 252 341 304 347
rect 252 307 289 341
rect 289 307 304 341
rect 252 295 304 307
rect 384 334 436 346
rect 384 300 406 334
rect 406 300 436 334
rect 506 312 558 364
rect 909 316 961 368
rect 1497 384 1549 436
rect 1643 411 1671 445
rect 1671 411 1695 445
rect 1643 396 1695 411
rect 1715 414 1717 448
rect 1717 414 1751 448
rect 1751 414 1767 448
rect 1715 405 1767 414
rect 1920 448 1972 456
rect 1920 414 1929 448
rect 1929 414 1963 448
rect 1963 414 1972 448
rect 1920 404 1972 414
rect 384 294 436 300
rect 1087 318 1094 349
rect 1094 318 1128 349
rect 1128 318 1139 349
rect 1087 297 1139 318
rect 1794 321 1795 354
rect 1795 321 1829 354
rect 1829 321 1846 354
rect 1794 302 1846 321
rect 149 192 201 244
rect 658 239 710 250
rect 873 258 925 279
rect 658 205 678 239
rect 678 205 710 239
rect 873 227 899 258
rect 899 227 925 258
rect 658 198 710 205
rect 1447 242 1499 250
rect 1447 208 1449 242
rect 1449 208 1483 242
rect 1483 208 1499 242
rect 1447 198 1499 208
rect 255 138 307 146
rect 255 104 289 138
rect 289 104 307 138
rect 255 94 307 104
rect 637 83 689 135
rect 918 142 970 194
rect 1231 157 1283 168
rect 1079 104 1131 156
rect 1231 123 1237 157
rect 1237 123 1271 157
rect 1271 123 1283 157
rect 1231 116 1283 123
rect 1478 91 1530 143
rect 1614 142 1666 146
rect 1614 108 1629 142
rect 1629 108 1663 142
rect 1663 108 1666 142
rect 1614 94 1666 108
rect 1830 104 1882 156
rect 2110 154 2162 155
rect 2110 120 2116 154
rect 2116 120 2150 154
rect 2150 120 2162 154
rect 2110 103 2162 120
<< metal2 >>
tri 47 413 55 442 se
tri 44 400 47 413 se
rect 47 400 102 413
rect 85 396 102 400
tri 102 398 106 413 nw
tri 1019 398 1025 416 se
tri 1708 457 1711 459 se
tri 1698 450 1708 457 se
rect 1708 450 1711 457
tri 1695 448 1698 450 se
rect 1698 448 1711 450
rect 85 391 101 396
tri 101 395 102 396 nw
tri 1018 395 1019 396 se
rect 1019 395 1053 398
tri 1017 391 1018 395 se
rect 1018 391 1053 395
rect 85 384 100 391
tri 100 386 101 391 nw
tri 1016 386 1017 391 se
rect 1017 386 1053 391
tri 742 384 755 386 se
tri 755 384 834 386 sw
tri 1015 384 1016 386 se
rect 1016 384 1053 386
tri 1053 384 1061 398 nw
rect 1362 402 1367 413
tri 1367 405 1369 413 nw
rect 1362 398 1366 402
tri 1366 400 1367 402 nw
rect 1362 391 1363 398
rect 1323 386 1363 391
tri 1363 386 1366 398 nw
tri 1322 384 1323 386 se
rect 1323 384 1362 386
tri 1362 384 1363 386 nw
rect 1695 414 1711 448
rect 1695 413 1709 414
tri 1709 413 1711 414 nw
rect 1695 412 1705 413
tri 1705 412 1709 413 nw
rect 1695 410 1698 412
tri 1698 410 1705 412 nw
tri 1695 407 1698 410 nw
rect 1917 412 1920 413
tri 1917 410 1918 412 ne
rect 1918 410 1920 412
tri 1918 406 1919 410 ne
rect 1919 404 1920 410
rect 1919 403 1958 404
tri 1958 403 1961 404 nw
tri 1921 401 1927 403 ne
rect 1927 401 1947 403
tri 1695 400 1696 401 sw
tri 1927 400 1928 401 ne
rect 1928 400 1947 401
rect 1695 398 1696 400
tri 1928 399 1932 400 ne
rect 1932 399 1947 400
tri 1947 399 1958 403 nw
tri 1696 398 1697 399 sw
rect 1695 396 1697 398
tri 1664 393 1665 396 ne
rect 1665 392 1697 396
tri 1697 392 1702 398 sw
rect 1665 384 1702 392
rect 85 368 96 384
tri 96 369 100 384 nw
tri 646 369 742 384 se
rect 742 369 834 384
tri 639 368 646 369 se
rect 646 368 834 369
tri 834 368 906 384 sw
tri 1010 368 1015 384 se
rect 1015 368 1044 384
rect 85 364 95 368
tri 95 365 96 368 nw
tri 620 365 639 368 se
rect 639 367 906 368
tri 906 367 909 368 sw
rect 639 365 909 367
tri 613 364 620 365 se
rect 620 364 909 365
rect 85 361 94 364
tri 94 361 95 364 nw
rect 85 355 88 361
tri 88 355 94 361 nw
tri 594 361 613 364 se
rect 613 361 909 364
tri 572 358 594 361 se
rect 594 358 909 361
tri 564 357 572 358 se
rect 572 357 909 358
tri 258 348 263 352 se
tri 263 351 294 352 sw
rect 263 348 294 351
tri 257 347 258 348 se
rect 258 347 294 348
tri 294 347 299 351 sw
rect 260 294 296 295
rect 599 356 909 357
rect 599 354 757 356
tri 757 354 765 356 nw
tri 792 354 838 356 ne
rect 838 354 909 356
rect 599 352 747 354
tri 747 352 757 354 nw
tri 838 352 846 354 ne
rect 846 352 909 354
rect 599 351 745 352
tri 745 351 747 352 nw
tri 846 351 849 352 ne
rect 849 351 909 352
rect 599 339 687 351
tri 687 339 745 351 nw
tri 849 339 896 351 ne
rect 896 339 909 351
rect 599 338 682 339
tri 682 338 687 339 nw
tri 896 338 901 339 ne
rect 901 338 909 339
rect 599 335 668 338
tri 668 335 682 338 nw
tri 901 335 909 338 ne
rect 599 333 659 335
tri 659 333 668 335 nw
rect 599 330 647 333
tri 647 330 659 333 nw
rect 599 326 628 330
tri 628 326 647 330 nw
rect 599 323 617 326
tri 617 323 628 326 nw
rect 599 319 610 323
tri 610 319 616 323 nw
rect 599 316 607 319
tri 607 316 610 319 nw
tri 1008 361 1010 368 se
rect 1010 367 1044 368
tri 1044 367 1053 384 nw
tri 1320 379 1322 384 se
rect 1322 383 1362 384
rect 1322 379 1361 383
tri 1361 379 1362 383 nw
tri 1506 379 1509 384 ne
rect 1509 379 1549 384
tri 1311 367 1320 379 se
rect 1320 367 1355 379
rect 1010 361 1040 367
tri 1006 355 1008 361 se
rect 1008 355 1040 361
tri 1040 355 1044 367 nw
tri 1303 357 1311 367 se
rect 1311 357 1355 367
rect 1006 354 1040 355
tri 1004 349 1006 354 se
rect 1006 349 1038 354
tri 1038 349 1040 354 nw
tri 1296 350 1303 357 se
rect 1303 354 1355 357
tri 1355 354 1361 379 nw
tri 1509 355 1518 379 ne
rect 1518 357 1549 379
tri 1549 357 1555 384 sw
rect 1518 354 1555 357
tri 1665 356 1669 384 ne
rect 1669 360 1702 384
tri 1702 360 1720 392 sw
rect 1669 354 1720 360
rect 1303 350 1351 354
tri 997 327 1004 349 se
rect 1004 327 1031 349
tri 1031 327 1038 349 nw
tri 996 323 997 327 se
rect 997 323 1021 327
tri 994 319 996 323 se
rect 996 319 1021 323
tri 993 316 994 318 se
rect 994 316 1021 319
rect 599 312 602 316
tri 602 312 607 316 nw
tri 992 313 993 316 se
rect 993 313 1021 316
tri 537 309 543 312 ne
tri 599 309 602 312 nw
tri 991 309 992 312 se
rect 992 309 1021 313
tri 989 303 991 307 se
rect 991 303 1021 309
tri 987 297 989 301 se
rect 989 297 1021 303
tri 1021 297 1031 327 nw
tri 1290 343 1296 349 se
rect 1296 343 1351 350
tri 1286 338 1290 343 se
rect 1290 338 1351 343
tri 1351 338 1355 354 nw
tri 1518 338 1525 354 ne
rect 1525 338 1555 354
tri 1278 306 1286 338 se
rect 1286 326 1349 338
tri 1349 326 1351 338 nw
rect 1286 314 1340 326
tri 1340 314 1349 326 nw
tri 1525 314 1535 338 ne
rect 1535 322 1555 338
tri 1555 322 1562 354 sw
tri 1669 347 1670 354 ne
rect 1670 347 1720 354
tri 1720 347 1721 354 sw
tri 1670 322 1674 347 ne
rect 1535 314 1562 322
rect 1286 310 1320 314
tri 1320 310 1340 314 nw
tri 1535 311 1536 314 ne
rect 1536 312 1562 314
tri 1562 312 1564 322 sw
rect 1286 306 1315 310
tri 1277 302 1278 305 se
rect 1278 302 1315 306
tri 1315 303 1320 310 nw
rect 1536 306 1564 312
rect 1674 317 1721 347
tri 1721 317 1722 347 sw
rect 1674 314 1722 317
tri 1722 314 1723 316 sw
tri 1564 306 1565 311 sw
rect 1536 303 1565 306
tri 1536 302 1537 303 ne
rect 1277 301 1314 302
tri 1314 301 1315 302 nw
rect 1537 301 1565 303
rect 1674 308 1723 314
tri 1085 297 1087 301 ne
rect 987 296 1021 297
tri 260 280 262 294 ne
rect 262 291 296 294
rect 262 279 295 291
tri 295 280 296 291 nw
tri 262 250 266 279 ne
tri 140 211 142 244 se
tri 142 243 149 244 sw
rect 142 211 149 243
tri 140 198 149 211 ne
tri 265 198 266 240 se
rect 266 199 293 279
tri 293 259 295 279 nw
rect 396 279 436 294
tri 436 279 441 294 sw
tri 982 279 987 294 se
rect 987 279 1006 296
tri 396 262 397 279 ne
rect 397 263 441 279
tri 441 263 446 279 sw
rect 397 259 446 263
tri 446 259 451 263 sw
rect 397 257 451 259
tri 451 257 466 259 sw
rect 397 253 466 257
tri 466 253 471 257 sw
tri 865 253 873 256 se
rect 397 250 471 253
tri 471 250 472 253 sw
tri 858 250 865 253 se
rect 865 250 873 253
tri 293 199 298 250 sw
rect 397 245 472 250
rect 266 198 298 199
tri 155 180 162 189 ne
tri 162 180 188 189 nw
tri 264 180 265 189 se
rect 265 180 298 198
rect 264 151 298 180
tri 298 151 302 194 sw
rect 451 236 472 245
tri 472 236 479 250 sw
tri 653 236 657 237 se
rect 657 236 658 237
rect 451 225 479 236
tri 479 225 572 236 sw
tri 602 225 653 236 se
rect 653 225 658 236
rect 451 224 572 225
tri 572 224 583 225 sw
tri 583 224 600 225 se
rect 600 224 658 225
rect 451 200 658 224
rect 451 198 634 200
tri 634 198 655 200 nw
tri 847 245 858 250 se
rect 858 245 873 250
tri 980 272 982 279 se
rect 982 272 1006 279
tri 977 263 980 272 se
rect 980 263 1006 272
tri 975 259 977 263 se
rect 977 259 1006 263
tri 974 253 975 256 se
rect 975 253 1006 259
tri 973 251 974 253 se
rect 974 251 1006 253
tri 1006 251 1021 296 nw
tri 1087 272 1098 297 ne
rect 1098 272 1129 297
tri 1129 272 1130 297 nw
tri 1275 293 1277 301 se
rect 1277 293 1312 301
tri 1312 293 1314 301 nw
tri 1537 293 1539 301 ne
rect 1539 293 1565 301
tri 1269 272 1275 293 se
rect 1275 272 1299 293
tri 1098 266 1099 272 ne
rect 973 250 1006 251
rect 1099 250 1129 272
tri 1268 266 1269 272 se
rect 1269 266 1299 272
tri 1266 259 1268 265 se
rect 1268 259 1299 266
tri 1264 251 1266 259 se
rect 1266 251 1299 259
tri 970 243 973 250 se
rect 973 243 997 250
tri 968 234 970 243 se
rect 970 234 997 243
tri 966 230 968 234 se
rect 968 230 997 234
rect 451 195 601 198
tri 601 195 634 198 nw
tri 451 194 590 195 nw
rect 887 223 898 227
tri 898 224 901 227 nw
tri 964 224 966 230 se
rect 966 224 997 230
rect 887 205 888 223
tri 888 205 898 223 nw
tri 950 205 964 223 se
rect 964 222 997 224
tri 997 223 1006 250 nw
tri 1097 223 1099 250 se
rect 1099 223 1127 250
rect 964 205 982 222
tri 887 202 888 205 nw
tri 948 202 950 205 se
rect 950 202 982 205
tri 945 198 948 202 se
rect 948 198 982 202
tri 982 198 997 222 nw
tri 1095 198 1097 222 se
rect 1097 198 1127 223
tri 1127 202 1129 250 nw
tri 1251 202 1264 250 se
rect 1264 249 1299 251
tri 1299 250 1312 293 nw
tri 1539 250 1546 293 ne
rect 1546 250 1565 293
rect 1264 205 1286 249
tri 1286 205 1299 249 nw
tri 1436 233 1446 239 se
rect 1446 233 1447 239
tri 1412 219 1436 233 se
rect 1436 219 1447 233
tri 1398 211 1412 219 se
rect 1412 211 1447 219
tri 1391 208 1398 211 se
rect 1398 208 1447 211
tri 1389 205 1391 208 se
rect 1391 205 1447 208
rect 1264 202 1276 205
tri 1250 198 1251 202 se
rect 1251 198 1276 202
tri 943 196 945 198 se
rect 945 196 976 198
rect 943 195 976 196
rect 942 194 976 195
rect 264 146 302 151
rect 970 187 976 194
tri 976 188 982 198 nw
tri 1094 188 1095 193 se
rect 1095 188 1126 198
rect 970 185 974 187
tri 974 185 976 187 nw
tri 970 178 974 185 nw
tri 1091 168 1094 175 se
rect 1094 168 1126 188
tri 1126 175 1127 198 nw
tri 1244 175 1250 198 se
rect 1250 175 1276 198
tri 1243 169 1244 174 se
rect 1244 169 1276 175
tri 1276 170 1286 205 nw
tri 1385 200 1389 205 se
rect 1389 200 1447 205
rect 1385 198 1447 200
tri 1546 244 1547 250 ne
rect 1547 241 1565 250
tri 1547 233 1549 241 ne
rect 1549 233 1565 241
tri 1549 219 1551 233 ne
rect 1551 229 1565 233
tri 1565 229 1581 302 sw
rect 1674 301 1720 308
tri 1720 302 1723 308 nw
rect 1674 297 1718 301
tri 1718 297 1720 301 nw
tri 1804 299 1805 302 ne
rect 1805 297 1842 302
rect 1551 220 1581 229
tri 1550 211 1551 219 se
rect 1551 211 1579 220
tri 1579 211 1581 220 nw
tri 1655 211 1674 297 se
rect 1674 271 1701 297
tri 1701 271 1718 297 nw
tri 1805 272 1810 297 ne
rect 1810 271 1842 297
rect 1674 211 1688 271
tri 1688 212 1701 271 nw
tri 1810 212 1821 271 ne
tri 1546 205 1550 211 se
rect 1550 205 1576 211
tri 1543 200 1546 205 se
rect 1546 200 1576 205
tri 1384 195 1385 198 se
rect 1385 196 1489 198
tri 1489 196 1491 198 nw
tri 1541 196 1543 200 se
rect 1543 196 1576 200
rect 1385 195 1485 196
tri 1485 195 1489 196 nw
rect 1541 195 1576 196
tri 1576 195 1579 211 nw
tri 1652 196 1655 211 se
rect 1655 196 1685 211
tri 1685 196 1688 211 nw
rect 1821 211 1842 271
tri 1821 196 1824 211 ne
rect 1652 195 1685 196
tri 1374 171 1384 195 se
rect 1384 181 1412 195
tri 1412 181 1485 195 nw
tri 1533 181 1541 195 se
rect 1541 190 1575 195
tri 1575 190 1576 195 nw
tri 1651 193 1652 195 se
rect 1652 193 1684 195
tri 1684 193 1685 195 nw
rect 1824 193 1842 211
tri 1650 190 1651 193 se
rect 1651 190 1684 193
tri 1824 190 1825 193 ne
rect 1825 190 1842 193
rect 1541 181 1554 190
rect 1384 175 1405 181
tri 1405 175 1412 181 nw
tri 1530 175 1533 181 se
rect 1533 175 1554 181
rect 1384 171 1403 175
rect 1243 168 1276 169
tri 1090 166 1091 168 se
rect 1091 166 1125 168
tri 1087 156 1090 166 se
rect 1090 156 1125 166
tri 1125 156 1126 168 nw
rect 689 128 692 131
tri 692 128 771 131 sw
rect 689 127 771 128
tri 771 127 800 128 sw
rect 689 126 800 127
tri 800 126 828 127 sw
rect 689 122 828 126
tri 828 122 842 126 sw
rect 689 117 842 122
tri 842 117 848 122 sw
rect 689 115 848 117
tri 848 115 859 117 sw
rect 689 111 859 115
tri 859 111 872 115 sw
rect 689 110 872 111
tri 872 110 877 111 sw
rect 689 106 877 110
tri 877 106 893 110 sw
rect 689 104 893 106
tri 893 104 909 106 sw
tri 1371 164 1374 170 se
rect 1374 166 1403 171
tri 1403 166 1405 175 nw
tri 1525 166 1530 175 se
rect 1530 166 1554 175
rect 1374 164 1402 166
tri 1402 164 1403 166 nw
tri 1524 164 1525 166 se
rect 1525 164 1554 166
rect 1371 163 1402 164
tri 1370 161 1371 163 se
rect 1371 161 1401 163
tri 1401 162 1402 163 nw
tri 1523 163 1524 164 se
rect 1524 163 1554 164
tri 1522 161 1523 162 se
rect 1523 161 1554 163
tri 1368 156 1370 161 se
rect 1370 156 1399 161
tri 1399 156 1401 161 nw
tri 1519 156 1522 161 se
rect 1522 156 1554 161
tri 1554 156 1575 190 nw
tri 1641 168 1650 190 se
rect 1650 168 1679 190
tri 1679 168 1684 190 nw
tri 1825 168 1829 190 ne
rect 1829 168 1842 190
tri 1842 168 1864 302 sw
tri 1636 157 1641 168 se
rect 1641 157 1676 168
tri 1365 149 1368 156 se
rect 1368 155 1399 156
rect 1368 149 1393 155
tri 1364 146 1365 149 se
rect 1365 146 1393 149
tri 1363 144 1364 146 se
rect 1364 144 1393 146
tri 1360 137 1363 143 se
rect 1363 137 1393 144
tri 1393 137 1399 155 nw
tri 1516 150 1519 156 se
rect 1519 150 1550 156
tri 1513 146 1516 149 se
rect 1516 148 1550 150
tri 1550 149 1554 156 nw
tri 1633 150 1636 156 se
rect 1636 154 1676 157
tri 1676 156 1679 168 nw
tri 1829 156 1832 168 ne
rect 1832 156 1864 168
tri 1864 156 1866 168 sw
rect 1636 150 1675 154
rect 1633 149 1675 150
tri 1675 149 1676 154 nw
rect 1516 146 1548 148
tri 1548 146 1550 148 nw
tri 1632 146 1633 148 se
rect 1633 146 1674 149
tri 1674 146 1675 149 nw
tri 1507 143 1513 146 se
rect 1513 143 1543 146
rect 1360 136 1393 137
tri 1355 123 1360 136 se
rect 1360 123 1384 136
tri 1352 116 1355 123 se
rect 1355 116 1384 123
tri 1350 111 1352 116 se
rect 1352 111 1384 116
tri 1348 107 1350 110 se
rect 1350 107 1384 111
tri 1384 107 1393 136 nw
tri 1345 106 1348 107 se
rect 1348 106 1381 107
rect 689 103 909 104
tri 909 103 918 104 sw
rect 689 101 918 103
tri 918 101 940 103 sw
tri 1335 101 1345 106 se
rect 1345 101 1381 106
rect 689 98 940 101
tri 940 98 975 101 sw
tri 1331 100 1335 101 se
rect 1335 100 1381 101
tri 1381 100 1384 107 nw
tri 1304 98 1331 100 se
rect 1331 98 1380 100
tri 1380 98 1381 100 nw
rect 689 96 975 98
tri 975 96 994 98 sw
tri 1279 96 1304 98 se
rect 1304 96 1380 98
rect 689 95 994 96
tri 994 95 1002 96 sw
tri 1269 95 1279 96 se
rect 1279 95 1377 96
rect 689 93 1002 95
tri 1002 93 1023 95 sw
tri 1242 93 1269 95 se
rect 1269 93 1377 95
rect 689 91 753 93
tri 753 91 787 93 nw
tri 787 91 807 93 ne
rect 807 91 1023 93
tri 1023 91 1037 93 sw
tri 1224 91 1242 93 se
rect 1242 91 1377 93
tri 1377 91 1380 96 nw
rect 1530 136 1543 143
tri 1543 137 1548 146 nw
rect 1530 133 1541 136
tri 1541 133 1542 136 nw
rect 1530 123 1535 133
tri 1535 123 1541 133 nw
tri 1530 114 1535 123 nw
rect 1666 145 1674 146
rect 1666 139 1673 145
tri 1673 140 1674 145 nw
rect 1666 133 1672 139
tri 1672 137 1673 139 nw
rect 1666 123 1670 133
tri 1670 124 1672 133 nw
rect 1666 119 1669 123
tri 1669 119 1670 123 nw
tri 1666 114 1669 119 nw
tri 2109 144 2110 145 se
tri 2108 133 2109 144 se
rect 2109 133 2110 144
tri 689 88 753 91 nw
tri 807 88 816 91 ne
rect 816 89 1037 91
tri 1037 89 1058 91 sw
tri 1197 89 1224 91 se
rect 1224 89 1374 91
rect 816 88 1058 89
tri 816 87 820 88 ne
rect 820 87 1058 88
tri 1058 87 1064 89 sw
tri 1175 87 1197 89 se
rect 1197 87 1374 89
tri 820 84 822 87 ne
rect 822 83 1064 87
tri 1064 83 1078 87 sw
tri 1127 83 1175 87 se
rect 1175 85 1374 87
tri 1374 85 1377 91 nw
rect 1175 83 1361 85
tri 822 81 824 83 ne
rect 824 82 1078 83
tri 1078 82 1089 83 sw
tri 1116 82 1121 83 se
rect 1121 82 1361 83
rect 824 81 1361 82
tri 824 79 825 81 ne
rect 825 79 1361 81
tri 825 72 840 79 ne
rect 840 72 1361 79
tri 1361 72 1374 85 nw
tri 840 56 1064 72 ne
rect 1064 66 1348 72
tri 1348 66 1361 72 nw
rect 1064 56 1162 66
tri 1162 56 1348 66 nw
tri 1064 53 1075 56 ne
rect 1075 53 1115 56
tri 1115 53 1162 56 nw
tri 1075 52 1105 53 ne
tri 1105 52 1115 53 nw
<< via2 >>
rect 55 413 111 469
rect 1319 443 1375 469
rect 1711 457 1767 469
rect 1319 413 1362 443
rect 1362 413 1375 443
rect 1711 413 1715 457
rect 1715 413 1767 457
rect 1911 456 1967 469
rect 1911 413 1920 456
rect 1920 413 1967 456
rect 543 312 558 357
rect 558 312 599 357
rect 1079 349 1135 357
rect 543 301 599 312
rect 1079 301 1087 349
rect 1087 301 1135 349
rect 151 244 207 245
rect 151 192 201 244
rect 201 192 207 244
rect 151 189 207 192
rect 395 189 451 245
rect 831 227 873 245
rect 873 227 887 245
rect 831 189 887 227
rect 2103 103 2110 133
rect 2110 103 2159 133
rect 2103 77 2159 103
<< metal3 >>
rect 50 469 196 474
rect 50 413 55 469
rect 111 413 196 469
rect 50 408 196 413
rect 1314 469 1460 474
rect 1314 413 1319 469
rect 1375 413 1460 469
rect 1314 408 1460 413
rect 1654 469 1800 474
rect 1654 413 1711 469
rect 1767 413 1800 469
rect 1654 408 1800 413
rect 1861 469 1972 474
rect 1861 413 1911 469
rect 1967 413 1972 469
rect 1861 408 1972 413
rect 538 357 684 362
rect 538 301 543 357
rect 599 301 684 357
rect 538 296 684 301
rect 1074 357 1185 362
rect 1074 301 1079 357
rect 1135 301 1185 357
rect 1074 296 1185 301
rect 116 245 262 250
rect 116 189 151 245
rect 207 189 262 245
rect 116 184 262 189
rect 323 245 469 250
rect 323 189 395 245
rect 451 189 469 245
rect 323 184 469 189
rect 826 245 972 250
rect 826 189 831 245
rect 887 189 972 245
rect 826 184 972 189
rect 1125 135 1185 296
rect 1284 135 1314 178
rect 1861 135 1921 408
rect 1125 75 1921 135
rect 2098 133 2244 138
rect 2098 77 2103 133
rect 2159 77 2244 133
rect 1284 48 1314 75
rect 2098 72 2244 77
<< labels >>
flabel nwell s 33 528 67 562 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 425 528 459 562 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 913 528 947 562 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 1401 528 1435 562 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 1793 528 1827 562 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel pwell s 33 -16 67 18 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 425 -16 459 18 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 913 -16 947 18 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 1401 -16 1435 18 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 1793 -16 1827 18 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel comment s 0 1 0 1 0 FreeSans 100 0 0 0 mul2
flabel metal3 s 826 184 972 250 0 FreeSans 100 0 0 0 A1
port 3 nsew
flabel metal3 s 2098 72 2244 138 0 FreeSans 100 0 0 0 R3
port 4 nsew
flabel metal3 s 50 408 196 474 0 FreeSans 100 0 0 0 R0
port 5 nsew
flabel metal3 s 1314 408 1460 474 0 FreeSans 100 0 0 0 R2
port 6 nsew
flabel metal3 s 1654 408 1800 474 0 FreeSans 100 0 0 0 R1
port 7 nsew
flabel metal3 s 538 296 684 362 0 FreeSans 100 0 0 0 B1
port 8 nsew
flabel metal3 s 116 184 262 250 0 FreeSans 100 0 0 0 A0
port 9 nsew
flabel metal3 s 323 184 469 250 0 FreeSans 100 0 0 0 B0
port 10 nsew
flabel metal1 s 31 -16 65 18 0 FreeSans 100 0 0 0 vgnd
port 11 nsew
flabel metal1 s 31 528 65 562 0 FreeSans 100 0 0 0 vpwr
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 2392 544
<< end >>
