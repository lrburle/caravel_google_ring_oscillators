magic
tech sky130A
magscale 1 2
timestamp 1708622636
<< error_s >>
rect 3119 2104 3120 2115
rect 3309 2104 3310 2115
rect 3395 2104 3396 2115
rect 4618 2104 4619 2115
rect 4808 2104 4809 2115
rect 4894 2104 4895 2115
rect 5745 2104 5746 2115
rect 5935 2104 5936 2115
rect 6021 2104 6022 2115
rect 6294 2104 6295 2115
rect 6492 2104 6493 2115
rect 7670 2104 7671 2115
rect 7860 2104 7861 2115
rect 7946 2104 7947 2115
rect 8797 2104 8798 2115
rect 8987 2104 8988 2115
rect 9073 2104 9074 2115
rect 9346 2104 9347 2115
rect 9544 2104 9545 2115
rect 10722 2104 10723 2115
rect 10912 2104 10913 2115
rect 10998 2104 10999 2115
rect 11849 2104 11850 2115
rect 12039 2104 12040 2115
rect 12125 2104 12126 2115
rect 12398 2104 12399 2115
rect 12596 2104 12597 2115
rect 13774 2104 13775 2115
rect 13964 2104 13965 2115
rect 14050 2104 14051 2115
rect 14901 2104 14902 2115
rect 15091 2104 15092 2115
rect 15177 2104 15178 2115
rect 15450 2104 15451 2115
rect 15648 2104 15649 2115
rect 16826 2104 16827 2115
rect 17016 2104 17017 2115
rect 17102 2104 17103 2115
rect 17953 2104 17954 2115
rect 18143 2104 18144 2115
rect 18229 2104 18230 2115
rect 18502 2104 18503 2115
rect 18700 2104 18701 2115
rect 3130 2064 3131 2104
rect 3320 2064 3321 2104
rect 3406 2064 3407 2104
rect 4629 2064 4630 2104
rect 4819 2064 4820 2104
rect 4905 2064 4906 2104
rect 5756 2064 5757 2104
rect 5946 2064 5947 2104
rect 6032 2064 6033 2104
rect 6305 2064 6306 2104
rect 6503 2064 6504 2104
rect 7681 2064 7682 2104
rect 7871 2064 7872 2104
rect 7957 2064 7958 2104
rect 8808 2064 8809 2104
rect 8998 2064 8999 2104
rect 9084 2064 9085 2104
rect 9357 2064 9358 2104
rect 9555 2064 9556 2104
rect 10733 2064 10734 2104
rect 10923 2064 10924 2104
rect 11009 2064 11010 2104
rect 11860 2064 11861 2104
rect 12050 2064 12051 2104
rect 12136 2064 12137 2104
rect 12409 2064 12410 2104
rect 12607 2064 12608 2104
rect 13785 2064 13786 2104
rect 13975 2064 13976 2104
rect 14061 2064 14062 2104
rect 14912 2064 14913 2104
rect 15102 2064 15103 2104
rect 15188 2064 15189 2104
rect 15461 2064 15462 2104
rect 15659 2064 15660 2104
rect 16837 2064 16838 2104
rect 17027 2064 17028 2104
rect 17113 2064 17114 2104
rect 17964 2064 17965 2104
rect 18154 2064 18155 2104
rect 18240 2064 18241 2104
rect 18513 2064 18514 2104
rect 18711 2064 18712 2104
rect 5953 1937 5980 1944
rect 9005 1937 9032 1944
rect 12057 1937 12084 1944
rect 15109 1937 15136 1944
rect 18161 1937 18188 1944
rect 5953 1916 6021 1937
rect 9005 1916 9073 1937
rect 12057 1916 12125 1937
rect 15109 1916 15177 1937
rect 18161 1916 18229 1937
rect 5953 1910 6008 1916
rect 9005 1910 9060 1916
rect 12057 1910 12112 1916
rect 15109 1910 15164 1916
rect 18161 1910 18216 1916
rect 5992 1909 5993 1910
rect 9044 1909 9045 1910
rect 12096 1909 12097 1910
rect 15148 1909 15149 1910
rect 18200 1909 18201 1910
rect 5965 1903 6020 1909
rect 9017 1903 9072 1909
rect 12069 1903 12124 1909
rect 15121 1903 15176 1909
rect 18173 1903 18228 1909
rect 5992 1881 5993 1903
rect 9044 1881 9045 1903
rect 12096 1881 12097 1903
rect 15148 1881 15149 1903
rect 18200 1881 18201 1903
rect 3119 1674 3120 1685
rect 3309 1674 3310 1685
rect 3395 1674 3396 1685
rect 4618 1674 4619 1685
rect 4808 1674 4809 1685
rect 4894 1674 4895 1685
rect 5745 1674 5746 1685
rect 5935 1674 5936 1685
rect 6021 1674 6022 1685
rect 6294 1674 6295 1685
rect 6492 1674 6493 1685
rect 7670 1674 7671 1685
rect 7860 1674 7861 1685
rect 7946 1674 7947 1685
rect 8797 1674 8798 1685
rect 8987 1674 8988 1685
rect 9073 1674 9074 1685
rect 9346 1674 9347 1685
rect 9544 1674 9545 1685
rect 10722 1674 10723 1685
rect 10912 1674 10913 1685
rect 10998 1674 10999 1685
rect 11849 1674 11850 1685
rect 12039 1674 12040 1685
rect 12125 1674 12126 1685
rect 12398 1674 12399 1685
rect 12596 1674 12597 1685
rect 13774 1674 13775 1685
rect 13964 1674 13965 1685
rect 14050 1674 14051 1685
rect 14901 1674 14902 1685
rect 15091 1674 15092 1685
rect 15177 1674 15178 1685
rect 15450 1674 15451 1685
rect 15648 1674 15649 1685
rect 16826 1674 16827 1685
rect 17016 1674 17017 1685
rect 17102 1674 17103 1685
rect 17953 1674 17954 1685
rect 18143 1674 18144 1685
rect 18229 1674 18230 1685
rect 18502 1674 18503 1685
rect 18700 1674 18701 1685
rect 3130 1478 3131 1674
rect 3320 1478 3321 1674
rect 3406 1478 3407 1674
rect 4629 1478 4630 1674
rect 4819 1478 4820 1674
rect 4905 1478 4906 1674
rect 5756 1478 5757 1674
rect 5946 1478 5947 1674
rect 6032 1478 6033 1674
rect 6305 1478 6306 1674
rect 6503 1478 6504 1674
rect 7681 1478 7682 1674
rect 7871 1478 7872 1674
rect 7957 1478 7958 1674
rect 8808 1478 8809 1674
rect 8998 1478 8999 1674
rect 9084 1478 9085 1674
rect 9357 1478 9358 1674
rect 9555 1478 9556 1674
rect 10733 1478 10734 1674
rect 10923 1478 10924 1674
rect 11009 1478 11010 1674
rect 11860 1478 11861 1674
rect 12050 1478 12051 1674
rect 12136 1478 12137 1674
rect 12409 1478 12410 1674
rect 12607 1478 12608 1674
rect 13785 1478 13786 1674
rect 13975 1478 13976 1674
rect 14061 1478 14062 1674
rect 14912 1478 14913 1674
rect 15102 1478 15103 1674
rect 15188 1478 15189 1674
rect 15461 1478 15462 1674
rect 15659 1478 15660 1674
rect 16837 1478 16838 1674
rect 17027 1478 17028 1674
rect 17113 1478 17114 1674
rect 17964 1478 17965 1674
rect 18154 1478 18155 1674
rect 18240 1478 18241 1674
rect 18513 1478 18514 1674
rect 18711 1478 18712 1674
rect 3444 1374 3468 1408
rect 4943 1374 4967 1408
rect 6070 1374 6094 1408
rect 7995 1374 8019 1408
rect 9122 1374 9146 1408
rect 11047 1374 11071 1408
rect 12174 1374 12198 1408
rect 14099 1374 14123 1408
rect 15226 1374 15250 1408
rect 17151 1374 17175 1408
rect 18278 1374 18302 1408
rect 6070 1085 6094 1119
rect 9122 1085 9146 1119
rect 12174 1085 12198 1119
rect 15226 1085 15250 1119
rect 18278 1085 18302 1119
rect 4790 1054 4799 1055
rect 7842 1054 7851 1055
rect 10894 1054 10903 1055
rect 13946 1054 13955 1055
rect 16998 1054 17007 1055
rect 4710 1049 4790 1054
rect 4799 1050 4835 1054
rect 4835 1049 4837 1050
rect 7762 1049 7842 1054
rect 7851 1050 7887 1054
rect 7887 1049 7889 1050
rect 10814 1049 10894 1054
rect 10903 1050 10939 1054
rect 10939 1049 10941 1050
rect 13866 1049 13946 1054
rect 13955 1050 13991 1054
rect 16982 1053 16998 1054
rect 13991 1049 13993 1050
rect 16918 1049 16982 1053
rect 17007 1050 17043 1054
rect 17043 1049 17045 1050
rect 4442 1041 4710 1049
rect 4837 1041 4854 1049
rect 7494 1041 7762 1049
rect 7889 1041 7906 1049
rect 10546 1041 10814 1049
rect 10941 1041 10958 1049
rect 13598 1041 13866 1049
rect 13993 1041 14010 1049
rect 16650 1041 16918 1049
rect 17045 1041 17062 1049
rect 4431 1040 4442 1041
rect 4411 1038 4442 1040
rect 4855 1038 4859 1041
rect 7483 1040 7494 1041
rect 7463 1038 7494 1040
rect 7907 1038 7911 1041
rect 10535 1040 10546 1041
rect 10515 1038 10546 1040
rect 10959 1038 10963 1041
rect 13587 1040 13598 1041
rect 13567 1038 13598 1040
rect 14011 1038 14015 1041
rect 16639 1040 16650 1041
rect 16619 1038 16650 1040
rect 17063 1038 17067 1041
rect 4393 1027 4431 1038
rect 4861 1030 4867 1036
rect 4060 1025 4099 1026
rect 4060 1024 4097 1025
rect 4099 1024 4100 1025
rect 4058 1022 4060 1024
rect 4086 1016 4098 1024
rect 4100 1022 4101 1024
rect 4360 1022 4393 1027
rect 4765 1025 4821 1027
rect 4101 1016 4107 1022
rect 4348 1020 4393 1022
rect 4660 1021 4765 1025
rect 4821 1021 4831 1025
rect 4348 1016 4404 1020
rect 4049 1015 4101 1016
rect 4048 1012 4049 1015
rect 4107 1013 4108 1016
rect 4104 1012 4108 1013
rect 4348 1014 4364 1016
rect 4392 1015 4404 1016
rect 4366 1014 4388 1015
rect 4400 1014 4404 1015
rect 4348 1012 4409 1014
rect 4440 1012 4660 1021
rect 4831 1017 4842 1021
rect 4831 1014 4849 1017
rect 4852 1014 4917 1030
rect 4831 1012 4917 1014
rect 4038 1005 4044 1011
rect 4047 1008 4048 1012
rect 4046 1005 4047 1008
rect 4084 1005 4090 1011
rect 4032 999 4038 1005
rect 4090 999 4096 1005
rect 4058 990 4059 997
rect 4097 995 4098 1012
rect 4103 1001 4110 1012
rect 4348 1011 4406 1012
rect 4339 1008 4345 1011
rect 4346 1009 4348 1011
rect 4350 1010 4355 1011
rect 4349 1009 4355 1010
rect 4409 1009 4410 1011
rect 4431 1010 4439 1012
rect 4837 1011 4846 1012
rect 4831 1010 4844 1011
rect 4852 1010 4917 1012
rect 4346 1008 4353 1009
rect 4411 1008 4431 1010
rect 4339 1006 4347 1008
rect 4332 1005 4347 1006
rect 4349 1005 4353 1008
rect 4329 1001 4347 1005
rect 4401 1001 4404 1008
rect 4103 998 4104 1001
rect 4102 997 4103 998
rect 4096 990 4098 994
rect 4099 990 4103 997
rect 4311 994 4329 1001
rect 4332 997 4347 1001
rect 4058 989 4075 990
rect 4059 988 4075 989
rect 4044 978 4075 988
rect 4079 978 4110 990
rect 4289 986 4311 994
rect 4332 990 4348 997
rect 4402 996 4403 1000
rect 4407 998 4431 1008
rect 4831 1009 4843 1010
rect 4844 1009 4917 1010
rect 4933 1009 5014 1030
rect 7445 1027 7483 1038
rect 7913 1030 7919 1036
rect 5745 1015 5746 1026
rect 5935 1015 5936 1026
rect 6021 1015 6022 1026
rect 6294 1015 6295 1026
rect 6491 1015 6492 1026
rect 7112 1025 7151 1026
rect 7112 1024 7149 1025
rect 7151 1024 7152 1025
rect 7110 1022 7112 1024
rect 7138 1016 7150 1024
rect 7152 1022 7153 1024
rect 7412 1022 7445 1027
rect 7817 1025 7873 1027
rect 7153 1016 7159 1022
rect 7400 1020 7445 1022
rect 7712 1021 7817 1025
rect 7873 1021 7883 1025
rect 7400 1016 7456 1020
rect 7101 1015 7153 1016
rect 4831 1005 4852 1009
rect 4407 996 4416 998
rect 4402 995 4404 996
rect 4407 995 4411 996
rect 4347 988 4348 990
rect 4270 979 4289 986
rect 4044 972 4110 978
rect 4256 974 4270 979
rect 4005 967 4011 968
rect 3766 965 3768 967
rect 3821 964 3822 967
rect 3998 964 4002 967
rect 4011 964 4018 967
rect 3822 962 3824 964
rect 3985 956 3998 964
rect 4018 963 4023 964
rect 4023 959 4034 963
rect 4060 961 4076 972
rect 4078 966 4098 972
rect 4248 971 4254 973
rect 4332 972 4348 988
rect 4392 992 4407 995
rect 4413 993 4415 996
rect 4392 986 4408 992
rect 4414 988 4415 993
rect 4413 986 4414 988
rect 4557 986 4578 1002
rect 4824 1001 4831 1005
rect 4837 1001 4852 1005
rect 4810 994 4824 1001
rect 4844 998 4852 1001
rect 4870 1005 4880 1009
rect 5014 1005 5031 1009
rect 4870 1003 4883 1005
rect 4852 995 4853 998
rect 4392 985 4416 986
rect 4771 985 4777 991
rect 4795 986 4810 994
rect 4793 985 4795 986
rect 4817 985 4823 991
rect 4853 985 4860 995
rect 4391 983 4392 985
rect 4396 974 4416 985
rect 4591 974 4603 982
rect 4613 974 4625 982
rect 4765 979 4771 985
rect 4823 979 4829 985
rect 4855 980 4863 985
rect 4855 979 4864 980
rect 4855 978 4865 979
rect 4855 975 4867 978
rect 4243 970 4248 971
rect 4240 969 4243 970
rect 4348 968 4366 971
rect 4396 970 4408 974
rect 4855 973 4869 975
rect 4870 973 4871 1003
rect 4876 993 4897 1003
rect 5031 999 5053 1005
rect 5053 997 5055 999
rect 4880 983 4897 993
rect 5055 992 5061 997
rect 5061 986 5065 992
rect 4855 971 4871 973
rect 4876 972 4897 983
rect 5065 982 5068 986
rect 5068 975 5072 982
rect 5072 973 5073 975
rect 4876 971 4998 972
rect 5073 971 5074 972
rect 4585 970 4587 971
rect 4627 970 4664 971
rect 4396 969 4405 970
rect 4140 967 4144 968
rect 4146 967 4151 968
rect 4078 961 4094 966
rect 4132 965 4140 967
rect 4130 964 4132 965
rect 4151 964 4154 967
rect 4232 966 4239 968
rect 4228 964 4232 966
rect 4127 963 4130 964
rect 4126 962 4127 963
rect 4154 962 4157 964
rect 4224 963 4228 964
rect 4046 959 4094 961
rect 4023 958 4038 959
rect 4046 958 4096 959
rect 4119 958 4128 962
rect 4157 959 4161 962
rect 4204 961 4224 963
rect 4026 956 4040 958
rect 4041 957 4096 958
rect 3982 954 3985 956
rect 4026 954 4043 956
rect 4046 954 4096 957
rect 4115 956 4128 958
rect 4161 956 4164 959
rect 4212 958 4218 961
rect 4111 954 4128 956
rect 4164 954 4167 956
rect 4201 954 4209 957
rect 4333 956 4339 959
rect 4348 956 4364 968
rect 4366 967 4373 968
rect 4396 967 4404 969
rect 4373 965 4384 967
rect 4392 966 4404 967
rect 4391 965 4404 966
rect 4384 964 4404 965
rect 4424 964 4430 970
rect 4470 966 4476 970
rect 4579 969 4585 970
rect 4460 964 4476 966
rect 4392 962 4404 964
rect 4311 954 4339 956
rect 3822 946 3823 949
rect 3821 945 3860 946
rect 3819 944 3821 945
rect 3804 934 3819 944
rect 3780 920 3804 934
rect 3777 918 3780 920
rect 3770 913 3777 918
rect 3822 913 3823 945
rect 3860 944 3887 945
rect 3964 944 3982 954
rect 4026 953 4096 954
rect 4026 951 4048 953
rect 4077 951 4078 953
rect 4084 951 4090 953
rect 4104 951 4128 954
rect 4026 948 4128 951
rect 4026 947 4081 948
rect 4084 947 4090 948
rect 4026 946 4060 947
rect 4062 946 4081 947
rect 4093 946 4128 948
rect 4026 944 4081 946
rect 4091 945 4128 946
rect 4090 944 4128 945
rect 4167 953 4190 954
rect 4198 953 4201 954
rect 4311 953 4329 954
rect 4333 953 4359 954
rect 4391 953 4397 959
rect 4418 958 4482 964
rect 4529 963 4535 969
rect 4575 968 4581 969
rect 4570 966 4581 968
rect 4564 964 4569 966
rect 4560 963 4564 964
rect 4575 963 4581 966
rect 4591 968 4625 970
rect 4629 969 4637 970
rect 4424 954 4476 958
rect 4523 957 4529 963
rect 4581 957 4587 963
rect 4167 946 4198 953
rect 4284 946 4323 953
rect 4339 947 4345 953
rect 4385 947 4391 953
rect 4167 944 4190 946
rect 4278 945 4284 946
rect 4273 944 4278 945
rect 3887 938 4128 944
rect 4157 938 4172 944
rect 4180 939 4190 944
rect 4186 938 4190 939
rect 4239 938 4273 944
rect 4424 938 4438 954
rect 3948 922 3964 938
rect 4010 937 4033 938
rect 4010 934 4038 937
rect 4010 933 4046 934
rect 4048 933 4056 935
rect 4077 934 4078 938
rect 4152 937 4157 938
rect 4143 935 4151 936
rect 4079 934 4126 935
rect 4138 934 4143 935
rect 4063 933 4126 934
rect 4190 933 4206 938
rect 4233 936 4239 938
rect 4424 936 4439 938
rect 4229 935 4232 936
rect 4224 933 4228 934
rect 4010 925 4118 933
rect 4077 924 4078 925
rect 4016 922 4033 924
rect 3948 916 3964 920
rect 3999 917 4014 922
rect 4037 920 4062 922
rect 3850 913 3891 916
rect 3895 913 3964 916
rect 3767 911 3770 913
rect 3822 911 3850 913
rect 3948 911 3992 913
rect 3998 911 4014 917
rect 4035 917 4062 920
rect 4081 918 4140 922
rect 4188 920 4224 933
rect 4422 931 4439 936
rect 4418 928 4422 931
rect 4411 924 4418 928
rect 4403 920 4411 924
rect 4424 920 4439 931
rect 4470 920 4472 954
rect 4476 950 4489 954
rect 4591 953 4612 968
rect 4622 967 4625 968
rect 4630 963 4637 969
rect 4665 968 4668 970
rect 4855 969 4869 971
rect 4870 970 4998 971
rect 4880 969 4897 970
rect 4901 969 4998 970
rect 4668 967 4670 968
rect 4670 966 4672 967
rect 4633 960 4635 963
rect 4851 960 4854 961
rect 4638 954 4645 957
rect 4770 953 4771 957
rect 4832 954 4851 960
rect 4855 957 4874 969
rect 4832 953 4856 954
rect 4590 952 4612 953
rect 4590 950 4591 952
rect 4476 942 4484 950
rect 4589 938 4590 949
rect 4646 946 4658 953
rect 4829 952 4832 953
rect 4659 944 4661 945
rect 4661 940 4668 944
rect 4476 920 4484 932
rect 4183 918 4188 920
rect 4063 917 4140 918
rect 4035 915 4047 917
rect 4107 916 4118 917
rect 4055 914 4067 916
rect 4106 915 4108 916
rect 3763 909 3767 911
rect 3821 910 3823 911
rect 3820 909 3824 910
rect 3819 906 3824 909
rect 3766 903 3767 904
rect 3818 903 3824 906
rect 3948 904 3964 911
rect 3992 910 4017 911
rect 3983 908 4014 910
rect 4017 909 4028 910
rect 4028 908 4035 909
rect 3973 906 4014 908
rect 4035 907 4048 908
rect 4056 906 4063 907
rect 3983 905 4014 906
rect 3998 904 4014 905
rect 3757 894 3758 899
rect 3811 896 3812 900
rect 3817 899 3824 903
rect 3816 895 3817 899
rect 3810 876 3812 895
rect 3964 888 3980 904
rect 3982 888 3998 904
rect 4075 888 4077 911
rect 4140 909 4156 917
rect 4172 913 4183 918
rect 4167 911 4171 913
rect 4161 909 4167 911
rect 4190 909 4206 920
rect 4390 912 4403 920
rect 4422 918 4476 920
rect 4487 918 4489 926
rect 4526 920 4529 937
rect 4668 935 4677 940
rect 4764 939 4770 952
rect 4774 946 4795 949
rect 4811 946 4812 949
rect 4823 948 4829 952
rect 4840 946 4856 953
rect 4764 936 4771 939
rect 4772 938 4774 946
rect 4795 939 4856 946
rect 4869 942 4874 957
rect 4897 968 4998 969
rect 5075 968 5076 970
rect 4803 938 4856 939
rect 4822 937 4872 938
rect 4589 925 4592 929
rect 4678 928 4688 934
rect 4764 933 4772 936
rect 4822 933 4829 937
rect 4418 912 4488 918
rect 4523 917 4525 919
rect 4592 918 4607 925
rect 4688 923 4692 928
rect 4692 920 4693 923
rect 4607 917 4630 918
rect 4523 916 4529 917
rect 4521 912 4529 916
rect 4388 911 4390 912
rect 4422 911 4437 912
rect 4438 911 4439 912
rect 4140 908 4206 909
rect 4126 907 4206 908
rect 4382 907 4388 911
rect 4422 907 4443 911
rect 4460 908 4476 912
rect 4084 906 4107 907
rect 4140 904 4206 907
rect 4174 888 4190 904
rect 4368 900 4382 907
rect 4422 904 4437 907
rect 4438 904 4439 907
rect 4470 906 4476 908
rect 4479 904 4488 912
rect 4523 911 4529 912
rect 4581 916 4630 917
rect 4581 911 4587 916
rect 4598 914 4630 916
rect 4607 913 4631 914
rect 4607 911 4630 913
rect 4633 911 4658 913
rect 4672 911 4686 920
rect 4693 918 4694 920
rect 4759 918 4764 933
rect 4770 927 4777 933
rect 4770 925 4772 927
rect 4694 913 4696 918
rect 4696 911 4697 913
rect 4757 911 4759 915
rect 4518 907 4520 911
rect 4423 900 4436 904
rect 4477 900 4479 903
rect 4514 900 4518 907
rect 4529 905 4535 911
rect 4348 888 4371 900
rect 4418 897 4423 900
rect 4402 888 4418 897
rect 4435 896 4438 899
rect 4472 896 4477 899
rect 4512 897 4514 900
rect 4438 888 4454 896
rect 4456 888 4472 896
rect 4506 888 4512 897
rect 3816 875 3824 888
rect 4012 880 4142 888
rect 4345 883 4348 888
rect 4394 883 4402 888
rect 4503 883 4506 888
rect 4260 880 4308 883
rect 3990 875 4032 880
rect 3810 873 3816 875
rect 3979 873 4032 875
rect 3767 870 3771 873
rect 3800 871 3810 873
rect 3813 872 3816 873
rect 3800 870 3812 871
rect 3960 870 4032 873
rect 4075 870 4077 880
rect 4119 879 4260 880
rect 4122 875 4260 879
rect 4308 875 4309 880
rect 4341 875 4345 883
rect 4380 876 4394 883
rect 4498 876 4503 883
rect 4374 875 4380 876
rect 4541 875 4565 910
rect 4575 905 4581 911
rect 4607 909 4686 911
rect 4697 909 4698 911
rect 4620 904 4686 909
rect 4698 904 4700 908
rect 4636 888 4652 904
rect 4654 893 4670 904
rect 4700 899 4702 903
rect 4702 893 4704 899
rect 4745 898 4757 910
rect 4766 909 4770 925
rect 4803 916 4811 933
rect 4817 927 4823 933
rect 4765 904 4766 909
rect 4783 905 4803 915
rect 4770 903 4782 905
rect 4783 903 4804 905
rect 4822 904 4823 927
rect 4856 922 4872 937
rect 4874 936 4875 941
rect 4897 938 4918 968
rect 4938 967 4998 968
rect 5076 967 5077 968
rect 4947 965 4998 967
rect 5077 965 5080 967
rect 4967 963 4998 965
rect 5080 963 5082 965
rect 4976 961 4998 963
rect 5082 961 5086 963
rect 4930 938 4946 954
rect 4948 938 4964 954
rect 4988 949 5016 961
rect 5086 954 5095 961
rect 4974 938 4975 949
rect 5016 947 5020 949
rect 5095 947 5103 954
rect 5020 946 5021 947
rect 5021 944 5022 946
rect 5103 944 5105 947
rect 5291 944 5292 949
rect 5320 944 5336 954
rect 5022 939 5028 944
rect 5105 940 5110 944
rect 5274 940 5341 944
rect 5110 939 5112 940
rect 5251 939 5274 940
rect 4897 936 4930 938
rect 4964 937 4980 938
rect 4944 936 4980 937
rect 5028 936 5030 938
rect 5112 936 5115 939
rect 5248 936 5251 939
rect 5291 938 5292 940
rect 5341 938 5342 939
rect 4875 916 4880 933
rect 4897 922 4929 936
rect 4944 935 4964 936
rect 4966 934 4980 936
rect 5030 934 5032 936
rect 5115 934 5119 936
rect 5245 934 5248 936
rect 4960 932 4980 934
rect 5032 932 5033 934
rect 5119 932 5121 934
rect 5244 932 5245 934
rect 4881 915 4887 921
rect 4897 919 4918 922
rect 4922 921 4929 922
rect 4918 915 4921 919
rect 4922 915 4933 921
rect 4875 909 4881 915
rect 4880 908 4881 909
rect 4922 906 4929 915
rect 4933 909 4939 915
rect 4971 904 5007 932
rect 5033 925 5040 932
rect 5121 925 5132 932
rect 5241 925 5244 932
rect 5040 924 5054 925
rect 5032 915 5054 924
rect 5132 919 5141 925
rect 5238 919 5241 925
rect 5141 916 5144 919
rect 5237 916 5238 919
rect 5040 907 5054 915
rect 5144 912 5149 916
rect 5235 912 5237 916
rect 5149 907 5153 912
rect 5232 910 5235 912
rect 5048 905 5057 907
rect 5054 904 5057 905
rect 5153 904 5155 907
rect 4979 903 4982 904
rect 5007 903 5008 904
rect 5057 903 5058 904
rect 4767 901 4807 903
rect 4764 900 4765 901
rect 4763 899 4764 900
rect 4767 899 4803 901
rect 4807 899 4808 901
rect 4762 898 4767 899
rect 4745 896 4767 898
rect 4705 893 4757 896
rect 4762 893 4767 896
rect 4654 888 4673 893
rect 4704 888 4757 893
rect 4601 877 4610 881
rect 4648 877 4657 881
rect 4667 879 4673 888
rect 4699 886 4711 888
rect 4694 883 4699 886
rect 4704 883 4711 886
rect 4693 882 4711 883
rect 4685 880 4711 882
rect 4682 879 4711 880
rect 4667 877 4711 879
rect 4593 875 4711 877
rect 4122 870 4224 875
rect 4262 874 4416 875
rect 4262 872 4409 874
rect 4235 871 4262 872
rect 4341 871 4345 872
rect 4374 871 4380 872
rect 4416 871 4430 874
rect 4496 871 4498 875
rect 4535 872 4593 875
rect 4601 872 4704 875
rect 4227 870 4235 871
rect 4430 870 4434 871
rect 4535 870 4601 872
rect 4602 870 4704 872
rect 4711 870 4713 875
rect 4745 872 4757 888
rect 4758 881 4763 893
rect 4762 880 4763 881
rect 4783 871 4803 899
rect 4808 893 4811 899
rect 4811 881 4816 893
rect 4919 887 4922 903
rect 4975 902 4979 903
rect 4974 899 4975 901
rect 5008 899 5014 903
rect 4967 893 4974 899
rect 4979 897 4980 899
rect 5013 893 5014 899
rect 5049 893 5056 898
rect 5058 893 5072 903
rect 4967 887 4973 893
rect 4811 877 4815 881
rect 4922 877 4947 887
rect 5056 885 5068 893
rect 5072 887 5081 893
rect 5155 887 5168 903
rect 5228 902 5240 910
rect 5250 902 5262 910
rect 5302 904 5303 938
rect 5341 934 5352 938
rect 5342 922 5352 934
rect 5342 903 5343 922
rect 5228 898 5231 902
rect 5264 899 5266 902
rect 5216 886 5224 898
rect 5228 896 5262 898
rect 5228 895 5231 896
rect 4815 873 4816 875
rect 4947 870 4965 877
rect 4967 875 4973 877
rect 5068 876 5075 885
rect 5081 879 5087 886
rect 5168 879 5173 886
rect 5087 877 5089 879
rect 5173 877 5175 879
rect 4967 870 4974 875
rect 4979 870 4980 872
rect 5089 871 5092 877
rect 5175 870 5179 877
rect 3771 869 3800 870
rect 3808 867 3812 870
rect 3956 869 3960 870
rect 4222 869 4227 870
rect 4310 869 4311 870
rect 3807 866 3812 867
rect 3943 866 3956 869
rect 4213 868 4222 869
rect 4205 866 4213 868
rect 4311 867 4312 869
rect 3755 859 3756 866
rect 3805 864 3812 866
rect 3921 865 3955 866
rect 4200 865 4205 866
rect 3805 859 3807 864
rect 3921 862 3943 865
rect 3920 859 3943 862
rect 3955 859 3962 865
rect 4167 859 4200 865
rect 3804 855 3805 859
rect 3916 855 3921 859
rect 3924 854 3943 859
rect 3962 857 3965 859
rect 4161 858 4167 859
rect 4154 857 4161 858
rect 4138 854 4153 857
rect 4312 854 4317 866
rect 4339 863 4341 870
rect 4371 863 4374 870
rect 4434 868 4446 870
rect 4338 860 4339 863
rect 4370 860 4371 863
rect 4446 859 4484 868
rect 4489 863 4494 870
rect 4524 869 4535 870
rect 4512 868 4524 869
rect 4510 866 4512 868
rect 4507 864 4510 866
rect 4537 864 4540 869
rect 4487 860 4489 863
rect 3803 851 3804 854
rect 3914 851 3916 854
rect 3923 850 3924 854
rect 3754 838 3755 850
rect 3799 838 3803 850
rect 3907 838 3914 850
rect 3753 816 3754 837
rect 3792 816 3799 838
rect 3907 835 3913 838
rect 3901 829 3907 835
rect 3915 828 3920 842
rect 3953 835 3959 841
rect 3965 839 3966 854
rect 4042 850 4138 854
rect 4317 850 4318 854
rect 4336 853 4338 859
rect 4367 853 4370 859
rect 4479 858 4489 859
rect 4479 853 4486 858
rect 4489 857 4495 858
rect 4504 857 4507 864
rect 4592 863 4601 870
rect 4657 863 4666 870
rect 4675 868 4676 870
rect 4713 868 4714 870
rect 4535 860 4537 863
rect 4676 861 4678 868
rect 4714 860 4717 868
rect 4743 864 4744 866
rect 4742 861 4743 863
rect 4758 859 4764 870
rect 4780 864 4783 870
rect 4816 866 4818 870
rect 4965 869 4975 870
rect 4855 868 4856 869
rect 4854 867 4855 868
rect 4853 865 4854 866
rect 4846 864 4853 865
rect 4770 859 4772 861
rect 4495 855 4518 857
rect 4533 856 4535 859
rect 4495 854 4508 855
rect 4528 854 4533 856
rect 4479 852 4482 853
rect 4479 851 4481 852
rect 4503 851 4504 854
rect 4508 851 4549 854
rect 4594 851 4600 857
rect 4640 851 4646 857
rect 4679 855 4680 857
rect 4718 854 4719 857
rect 4740 856 4741 859
rect 4766 856 4774 859
rect 4727 854 4766 856
rect 4776 855 4780 863
rect 4804 859 4846 864
rect 4875 863 4881 869
rect 4933 863 4939 869
rect 4967 867 4975 869
rect 5075 868 5076 870
rect 5092 869 5093 870
rect 4976 867 4985 868
rect 4967 866 4988 867
rect 4967 865 4975 866
rect 4976 865 4988 866
rect 5048 865 5050 868
rect 5093 867 5094 869
rect 5179 867 5181 869
rect 5228 868 5230 895
rect 5094 865 5095 866
rect 4976 863 4985 865
rect 4775 854 4776 855
rect 4650 851 4727 854
rect 4739 853 4740 854
rect 4768 853 4781 854
rect 3982 843 4043 850
rect 3981 841 3982 842
rect 3959 832 3965 835
rect 3966 832 3967 838
rect 3959 829 3967 832
rect 3975 829 3981 841
rect 3985 840 3996 842
rect 4042 840 4043 843
rect 4053 843 4243 850
rect 4318 846 4321 850
rect 4328 846 4336 851
rect 4359 847 4367 851
rect 4354 846 4415 847
rect 4265 843 4347 846
rect 4053 839 4138 843
rect 4231 842 4249 843
rect 4318 842 4321 843
rect 4213 839 4231 842
rect 4249 841 4261 842
rect 4264 839 4267 841
rect 4051 838 4053 839
rect 4046 835 4050 838
rect 4040 830 4046 835
rect 4073 831 4075 839
rect 4205 838 4213 839
rect 4189 835 4205 838
rect 3963 828 3967 829
rect 4039 828 4040 830
rect 3752 810 3753 816
rect 3791 811 3792 816
rect 3820 811 3836 824
rect 3914 813 3915 828
rect 3959 826 3961 827
rect 3963 826 3975 828
rect 3961 816 3983 826
rect 4012 817 4028 824
rect 3959 812 3983 816
rect 4002 812 4028 817
rect 3959 811 3961 812
rect 3789 807 3791 810
rect 3965 808 3967 811
rect 3751 800 3752 805
rect 3786 800 3788 805
rect 3785 798 3786 800
rect 3781 790 3785 798
rect 3804 792 3815 808
rect 3964 806 3965 808
rect 3983 807 3992 812
rect 4000 809 4028 812
rect 3998 808 4009 809
rect 4012 808 4028 809
rect 4030 808 4046 824
rect 4069 818 4075 831
rect 4155 830 4189 835
rect 4113 823 4155 830
rect 4267 829 4269 839
rect 4321 829 4326 842
rect 4328 828 4336 843
rect 4105 822 4113 823
rect 4080 818 4105 822
rect 4069 816 4080 818
rect 4065 812 4075 816
rect 3996 807 4012 808
rect 3992 806 4012 807
rect 3992 805 4009 806
rect 4046 805 4062 808
rect 3914 790 3915 805
rect 3779 786 3781 790
rect 3900 787 3915 790
rect 3953 789 3964 805
rect 3990 803 4023 805
rect 3990 794 4018 803
rect 4040 797 4062 805
rect 3990 793 4012 794
rect 3996 792 4012 793
rect 4002 790 4012 792
rect 4036 792 4062 797
rect 4036 791 4046 792
rect 3953 787 3965 789
rect 3750 782 3751 786
rect 3900 783 3965 787
rect 3996 787 4012 790
rect 4029 790 4046 791
rect 4029 787 4062 790
rect 3996 783 4062 787
rect 3900 782 3964 783
rect 3749 771 3750 781
rect 3778 773 3779 782
rect 3900 774 3966 782
rect 3990 774 4062 783
rect 4069 777 4073 812
rect 4097 803 4106 812
rect 4126 808 4142 823
rect 4144 803 4153 812
rect 4204 808 4220 824
rect 4222 808 4238 824
rect 4269 813 4273 828
rect 4326 825 4336 828
rect 4359 825 4367 846
rect 4416 843 4429 846
rect 4433 842 4435 843
rect 4437 842 4479 851
rect 4435 839 4479 842
rect 4437 835 4479 839
rect 4495 846 4549 851
rect 4588 850 4594 851
rect 4646 850 4727 851
rect 4554 846 4652 850
rect 4681 849 4683 850
rect 4692 849 4701 850
rect 4678 847 4688 849
rect 4693 848 4701 849
rect 4495 835 4525 846
rect 4549 845 4652 846
rect 4549 843 4561 845
rect 4576 843 4594 845
rect 4548 842 4549 843
rect 4683 842 4684 845
rect 4437 830 4525 835
rect 4537 831 4548 842
rect 4719 840 4725 850
rect 4437 825 4479 830
rect 4489 828 4513 830
rect 4536 828 4537 831
rect 4685 830 4688 838
rect 4726 830 4729 838
rect 4732 830 4738 850
rect 4759 839 4781 853
rect 4820 840 4825 858
rect 4881 857 4887 863
rect 4881 841 4886 857
rect 4923 841 4925 863
rect 4927 857 4933 863
rect 4975 862 4985 863
rect 4976 861 4985 862
rect 4976 859 4991 861
rect 5048 859 5054 865
rect 5095 864 5096 865
rect 4979 856 5004 859
rect 4979 853 4994 856
rect 4996 853 5002 856
rect 5032 854 5041 859
rect 5042 854 5048 859
rect 5078 857 5079 861
rect 5096 859 5098 864
rect 5098 856 5100 859
rect 5100 854 5101 856
rect 5181 854 5189 866
rect 5228 864 5231 868
rect 5260 864 5262 896
rect 5266 889 5274 898
rect 5266 879 5293 889
rect 5340 881 5343 885
rect 5333 879 5340 881
rect 5266 870 5333 879
rect 5287 869 5291 870
rect 5273 866 5287 869
rect 5268 865 5273 866
rect 5264 864 5268 865
rect 5224 856 5225 861
rect 5223 854 5225 856
rect 4985 850 4994 853
rect 5032 850 5051 854
rect 5040 846 5051 850
rect 5051 842 5052 846
rect 5079 842 5082 854
rect 5101 850 5103 854
rect 5189 851 5191 854
rect 5103 845 5107 850
rect 5107 843 5109 845
rect 5191 844 5196 850
rect 5109 842 5110 843
rect 5110 841 5112 842
rect 4881 839 4914 841
rect 4688 828 4689 830
rect 4489 825 4498 828
rect 4272 808 4273 813
rect 4324 824 4331 825
rect 4324 814 4334 824
rect 4324 812 4328 814
rect 4331 812 4334 814
rect 4356 813 4358 824
rect 4396 814 4412 824
rect 4389 813 4412 814
rect 4414 813 4437 824
rect 4481 820 4489 825
rect 4493 824 4498 825
rect 4157 803 4158 808
rect 4088 794 4101 803
rect 4153 794 4162 803
rect 4097 787 4101 794
rect 4157 792 4158 794
rect 4188 792 4204 808
rect 4239 807 4254 808
rect 4323 807 4324 811
rect 4332 808 4334 812
rect 4240 799 4254 807
rect 4273 800 4274 807
rect 4322 804 4323 807
rect 4321 800 4322 803
rect 4334 800 4350 808
rect 4355 807 4356 812
rect 4389 808 4430 813
rect 4380 806 4401 808
rect 4412 807 4418 808
rect 4354 800 4355 806
rect 4380 802 4396 806
rect 4406 802 4412 807
rect 4377 801 4423 802
rect 4377 800 4418 801
rect 4194 790 4200 792
rect 4203 791 4204 792
rect 4231 792 4254 799
rect 4274 797 4276 800
rect 4231 791 4246 792
rect 4202 790 4204 791
rect 4188 787 4204 790
rect 4205 789 4207 790
rect 4240 789 4246 791
rect 4205 787 4246 789
rect 4276 787 4286 797
rect 4318 787 4321 797
rect 4334 792 4354 800
rect 4349 790 4354 792
rect 4377 792 4396 800
rect 4430 792 4446 808
rect 4458 807 4464 813
rect 4471 812 4481 820
rect 4492 813 4498 824
rect 4513 823 4539 828
rect 4503 822 4546 823
rect 4503 821 4544 822
rect 4533 813 4536 821
rect 4546 818 4553 822
rect 4553 816 4554 818
rect 4465 807 4471 812
rect 4492 809 4493 813
rect 4554 812 4557 816
rect 4588 813 4604 824
rect 4606 813 4622 824
rect 4657 816 4666 825
rect 4689 824 4690 828
rect 4646 815 4657 816
rect 4579 812 4581 813
rect 4619 812 4623 813
rect 4532 809 4533 811
rect 4579 810 4623 812
rect 4579 808 4613 810
rect 4464 801 4470 807
rect 4476 792 4492 808
rect 4377 790 4387 792
rect 4389 790 4396 792
rect 4188 785 4243 787
rect 4099 777 4100 785
rect 4161 777 4167 783
rect 4188 781 4211 785
rect 3779 768 3780 771
rect 3916 767 3932 774
rect 3934 767 3950 774
rect 3990 771 3998 774
rect 4002 771 4048 774
rect 3998 767 4001 769
rect 4012 767 4028 771
rect 4030 767 4046 771
rect 3748 743 3749 767
rect 3780 742 3783 767
rect 3916 759 3950 767
rect 4002 759 4046 767
rect 3916 758 3932 759
rect 3934 758 3953 759
rect 4012 758 4028 759
rect 4030 758 4046 759
rect 4069 763 4072 777
rect 4074 763 4080 771
rect 3938 753 3953 758
rect 4069 757 4080 763
rect 4009 753 4018 756
rect 4063 754 4080 757
rect 4097 756 4100 777
rect 4045 753 4080 754
rect 3882 740 4080 753
rect 4088 747 4100 756
rect 4166 771 4173 777
rect 4188 774 4209 781
rect 3953 738 3962 740
rect 3968 737 4074 740
rect 4097 738 4106 747
rect 4108 741 4115 747
rect 3783 733 3784 737
rect 3784 724 3785 731
rect 4046 730 4048 737
rect 4069 730 4075 737
rect 4166 731 4167 771
rect 4194 753 4209 774
rect 4241 778 4242 785
rect 4246 778 4255 787
rect 4241 756 4243 778
rect 4247 775 4255 778
rect 4284 782 4299 787
rect 4316 782 4318 787
rect 4334 782 4354 790
rect 4284 778 4354 782
rect 4380 780 4396 790
rect 4284 774 4359 778
rect 4300 772 4316 774
rect 4318 772 4334 774
rect 4349 772 4359 774
rect 4377 774 4396 780
rect 4430 774 4446 790
rect 4476 780 4492 790
rect 4527 789 4532 808
rect 4562 803 4564 806
rect 4572 805 4588 808
rect 4623 807 4638 808
rect 4648 807 4657 815
rect 4684 810 4700 824
rect 4702 810 4718 824
rect 4729 823 4732 830
rect 4729 818 4734 823
rect 4728 816 4729 818
rect 4732 816 4734 818
rect 4759 816 4775 839
rect 4782 830 4789 838
rect 4825 830 4828 839
rect 4876 835 4887 839
rect 4876 831 4881 835
rect 4789 824 4792 830
rect 4828 828 4829 830
rect 4874 828 4876 831
rect 4885 828 4887 835
rect 4780 816 4796 824
rect 4724 813 4727 815
rect 4676 808 4719 810
rect 4734 808 4738 816
rect 4757 812 4759 816
rect 4668 807 4679 808
rect 4693 807 4695 808
rect 4719 807 4738 808
rect 4572 799 4594 805
rect 4572 798 4588 799
rect 4568 792 4588 798
rect 4594 793 4600 799
rect 4568 789 4575 792
rect 4579 789 4588 792
rect 4622 792 4638 807
rect 4646 799 4652 805
rect 4640 793 4646 799
rect 4622 790 4623 792
rect 4527 780 4542 789
rect 4572 788 4588 789
rect 4476 774 4542 780
rect 4567 778 4588 788
rect 4617 787 4619 790
rect 4622 787 4638 790
rect 4611 778 4613 787
rect 4567 776 4613 778
rect 4617 776 4638 787
rect 4655 785 4676 807
rect 4696 803 4697 805
rect 4709 799 4715 804
rect 4698 795 4699 797
rect 4719 795 4734 807
rect 4754 806 4757 812
rect 4780 811 4801 816
rect 4829 813 4834 828
rect 4867 817 4874 828
rect 4880 818 4881 828
rect 4867 816 4880 817
rect 4864 815 4867 816
rect 4849 814 4861 815
rect 4847 813 4849 814
rect 4825 812 4839 813
rect 4813 811 4825 812
rect 4780 810 4813 811
rect 4780 808 4801 810
rect 4829 808 4834 812
rect 4738 801 4740 805
rect 4745 795 4754 806
rect 4689 787 4705 795
rect 4719 792 4745 795
rect 4764 792 4780 808
rect 4796 806 4801 808
rect 4873 806 4880 816
rect 4885 809 4886 828
rect 4885 806 4888 809
rect 4917 807 4919 839
rect 5052 836 5054 841
rect 5082 836 5083 841
rect 5112 839 5136 841
rect 4873 805 4881 806
rect 4909 805 4919 807
rect 4923 805 4931 817
rect 4972 815 4988 824
rect 4990 815 5006 824
rect 4972 814 5006 815
rect 5054 814 5056 836
rect 5083 824 5089 836
rect 5114 830 5128 839
rect 5196 836 5198 842
rect 5221 841 5225 854
rect 5220 836 5225 841
rect 5213 834 5225 836
rect 5237 860 5265 861
rect 5237 855 5264 860
rect 5128 828 5136 830
rect 5129 825 5132 828
rect 4972 813 5007 814
rect 4970 811 4972 813
rect 5005 812 5006 813
rect 4970 808 5006 811
rect 5068 809 5102 824
rect 5132 815 5136 825
rect 5136 811 5137 814
rect 5137 809 5138 811
rect 5198 809 5199 811
rect 5065 808 5102 809
rect 5138 808 5139 809
rect 4801 801 4803 805
rect 4834 800 4836 805
rect 4881 802 4885 805
rect 4885 801 4909 802
rect 4917 801 4919 805
rect 4956 801 4982 808
rect 4992 801 5004 808
rect 4836 797 4837 800
rect 4805 795 4806 797
rect 4733 790 4745 792
rect 4806 791 4809 795
rect 4572 774 4583 776
rect 4618 774 4638 776
rect 4300 766 4365 772
rect 4377 768 4387 774
rect 4389 771 4423 774
rect 4426 771 4430 774
rect 4389 768 4430 771
rect 4300 758 4359 766
rect 4385 764 4387 768
rect 4396 764 4412 768
rect 4240 753 4243 756
rect 4246 753 4249 754
rect 4194 744 4249 753
rect 4307 749 4359 758
rect 4389 758 4412 764
rect 4414 758 4430 768
rect 4492 761 4508 774
rect 4389 756 4401 758
rect 4406 755 4412 758
rect 4464 755 4470 761
rect 4489 758 4508 761
rect 4510 758 4526 774
rect 4588 772 4604 774
rect 4606 772 4622 774
rect 4541 761 4547 767
rect 4579 764 4622 772
rect 4652 768 4656 785
rect 4689 780 4706 787
rect 4676 768 4682 773
rect 4702 772 4706 780
rect 4719 780 4749 790
rect 4719 774 4734 780
rect 4745 779 4749 780
rect 4728 773 4733 774
rect 4706 771 4707 772
rect 4489 755 4495 758
rect 4547 755 4553 761
rect 4588 758 4604 764
rect 4606 758 4622 764
rect 4412 749 4418 755
rect 4458 749 4464 755
rect 4491 754 4495 755
rect 4650 754 4656 768
rect 4698 767 4719 771
rect 4723 767 4728 773
rect 4664 757 4666 758
rect 4663 755 4664 757
rect 4488 750 4492 754
rect 4659 752 4663 755
rect 4698 753 4723 767
rect 4749 763 4760 779
rect 4764 774 4780 790
rect 4809 779 4814 790
rect 4814 776 4822 779
rect 4837 778 4853 797
rect 4885 793 4897 801
rect 4907 793 4919 801
rect 4950 797 4972 801
rect 4996 797 5002 801
rect 4950 795 5004 797
rect 5006 795 5022 808
rect 5052 795 5065 808
rect 5083 806 5089 808
rect 5089 802 5090 806
rect 4915 778 4919 793
rect 4944 789 4972 795
rect 4837 776 4875 778
rect 4814 775 4853 776
rect 4814 774 4830 775
rect 4760 754 4766 763
rect 4780 758 4796 774
rect 4798 763 4822 774
rect 4837 764 4853 775
rect 4860 775 4875 776
rect 4860 774 4876 775
rect 4876 763 4878 774
rect 4915 763 4917 778
rect 4798 758 4814 763
rect 4822 753 4827 763
rect 4853 754 4858 763
rect 4876 758 4881 763
rect 4916 761 4917 763
rect 4950 774 4972 789
rect 5002 792 5022 795
rect 5002 790 5016 792
rect 5002 789 5022 790
rect 5002 781 5004 789
rect 5003 774 5004 781
rect 5006 774 5022 789
rect 5045 784 5055 795
rect 5057 787 5058 795
rect 5090 786 5093 800
rect 5102 792 5118 808
rect 5043 780 5045 784
rect 5058 782 5059 786
rect 5093 781 5094 786
rect 5041 774 5043 780
rect 5094 778 5095 781
rect 5095 774 5097 778
rect 5102 774 5118 790
rect 5139 786 5147 808
rect 5213 806 5220 834
rect 5237 826 5258 855
rect 5212 802 5213 806
rect 5225 803 5234 812
rect 5237 808 5248 826
rect 5274 824 5284 847
rect 5260 818 5294 824
rect 5756 819 5757 1015
rect 5946 819 5947 1015
rect 6032 819 6033 1015
rect 6305 819 6306 1015
rect 6502 819 6503 1015
rect 7100 1012 7101 1015
rect 7159 1013 7160 1016
rect 7156 1012 7160 1013
rect 7400 1014 7416 1016
rect 7444 1015 7456 1016
rect 7418 1014 7440 1015
rect 7452 1014 7456 1015
rect 7400 1012 7461 1014
rect 7492 1012 7712 1021
rect 7883 1017 7894 1021
rect 7883 1014 7901 1017
rect 7904 1014 7969 1030
rect 7883 1012 7969 1014
rect 7090 1005 7096 1011
rect 7099 1008 7100 1012
rect 7098 1005 7099 1008
rect 7136 1005 7142 1011
rect 7084 999 7090 1005
rect 7142 999 7148 1005
rect 7110 990 7111 997
rect 7149 995 7150 1012
rect 7155 1001 7162 1012
rect 7400 1011 7458 1012
rect 7391 1008 7397 1011
rect 7398 1009 7400 1011
rect 7402 1010 7407 1011
rect 7401 1009 7407 1010
rect 7461 1009 7462 1011
rect 7483 1010 7491 1012
rect 7889 1011 7898 1012
rect 7883 1010 7896 1011
rect 7904 1010 7969 1012
rect 7398 1008 7405 1009
rect 7463 1008 7483 1010
rect 7391 1006 7399 1008
rect 7384 1005 7399 1006
rect 7401 1005 7405 1008
rect 7381 1001 7399 1005
rect 7453 1001 7456 1008
rect 7155 998 7156 1001
rect 7154 997 7155 998
rect 7148 990 7150 994
rect 7151 990 7155 997
rect 7363 994 7381 1001
rect 7384 997 7399 1001
rect 7110 989 7127 990
rect 7111 988 7127 989
rect 7096 978 7127 988
rect 7131 978 7162 990
rect 7341 986 7363 994
rect 7384 990 7400 997
rect 7454 996 7455 1000
rect 7459 998 7483 1008
rect 7883 1009 7895 1010
rect 7896 1009 7969 1010
rect 7985 1009 8066 1030
rect 10497 1027 10535 1038
rect 10965 1030 10971 1036
rect 8797 1015 8798 1026
rect 8987 1015 8988 1026
rect 9073 1015 9074 1026
rect 9346 1015 9347 1026
rect 9543 1015 9544 1026
rect 10164 1025 10203 1026
rect 10164 1024 10201 1025
rect 10203 1024 10204 1025
rect 10162 1022 10164 1024
rect 10190 1016 10202 1024
rect 10204 1022 10205 1024
rect 10464 1022 10497 1027
rect 10869 1025 10925 1027
rect 10205 1016 10211 1022
rect 10452 1020 10497 1022
rect 10764 1021 10869 1025
rect 10925 1021 10935 1025
rect 10452 1016 10508 1020
rect 10153 1015 10205 1016
rect 7883 1005 7904 1009
rect 7459 996 7468 998
rect 7454 995 7456 996
rect 7459 995 7463 996
rect 7399 988 7400 990
rect 7322 979 7341 986
rect 7096 972 7162 978
rect 7308 974 7322 979
rect 7057 967 7063 968
rect 6818 965 6820 967
rect 6873 964 6874 967
rect 7050 964 7054 967
rect 7063 964 7070 967
rect 6874 962 6876 964
rect 7037 956 7050 964
rect 7070 963 7075 964
rect 7075 959 7086 963
rect 7112 961 7128 972
rect 7130 966 7150 972
rect 7300 971 7306 973
rect 7384 972 7400 988
rect 7444 992 7459 995
rect 7465 993 7467 996
rect 7444 986 7460 992
rect 7466 988 7467 993
rect 7465 986 7466 988
rect 7609 986 7630 1002
rect 7876 1001 7883 1005
rect 7889 1001 7904 1005
rect 7862 994 7876 1001
rect 7896 998 7904 1001
rect 7922 1005 7932 1009
rect 8066 1005 8083 1009
rect 7922 1003 7935 1005
rect 7904 995 7905 998
rect 7444 985 7468 986
rect 7823 985 7829 991
rect 7847 986 7862 994
rect 7845 985 7847 986
rect 7869 985 7875 991
rect 7905 985 7912 995
rect 7443 983 7444 985
rect 7448 974 7468 985
rect 7643 974 7655 982
rect 7665 974 7677 982
rect 7817 979 7823 985
rect 7875 979 7881 985
rect 7907 980 7915 985
rect 7907 979 7916 980
rect 7907 978 7917 979
rect 7907 975 7919 978
rect 7295 970 7300 971
rect 7292 969 7295 970
rect 7400 968 7418 971
rect 7448 970 7460 974
rect 7907 973 7921 975
rect 7922 973 7923 1003
rect 7928 993 7949 1003
rect 8083 999 8105 1005
rect 8105 997 8107 999
rect 7932 983 7949 993
rect 8107 992 8113 997
rect 8113 986 8117 992
rect 7907 971 7923 973
rect 7928 972 7949 983
rect 8117 982 8120 986
rect 8120 975 8124 982
rect 8124 973 8125 975
rect 7928 971 8050 972
rect 8125 971 8126 972
rect 7637 970 7639 971
rect 7679 970 7716 971
rect 7448 969 7457 970
rect 7192 967 7196 968
rect 7198 967 7203 968
rect 7130 961 7146 966
rect 7184 965 7192 967
rect 7182 964 7184 965
rect 7203 964 7206 967
rect 7284 966 7291 968
rect 7280 964 7284 966
rect 7179 963 7182 964
rect 7178 962 7179 963
rect 7206 962 7209 964
rect 7276 963 7280 964
rect 7098 959 7146 961
rect 7075 958 7090 959
rect 7098 958 7148 959
rect 7171 958 7180 962
rect 7209 959 7213 962
rect 7256 961 7276 963
rect 7078 956 7092 958
rect 7093 957 7148 958
rect 7034 954 7037 956
rect 7078 954 7095 956
rect 7098 954 7148 957
rect 7167 956 7180 958
rect 7213 956 7216 959
rect 7264 958 7270 961
rect 7163 954 7180 956
rect 7216 954 7219 956
rect 7253 954 7261 957
rect 7385 956 7391 959
rect 7400 956 7416 968
rect 7418 967 7425 968
rect 7448 967 7456 969
rect 7425 965 7436 967
rect 7444 966 7456 967
rect 7443 965 7456 966
rect 7436 964 7456 965
rect 7476 964 7482 970
rect 7522 966 7528 970
rect 7631 969 7637 970
rect 7512 964 7528 966
rect 7444 962 7456 964
rect 7363 954 7391 956
rect 6874 946 6875 949
rect 6873 945 6912 946
rect 6871 944 6873 945
rect 6856 934 6871 944
rect 6832 920 6856 934
rect 6829 918 6832 920
rect 6822 913 6829 918
rect 6874 913 6875 945
rect 6912 944 6939 945
rect 7016 944 7034 954
rect 7078 953 7148 954
rect 7078 951 7100 953
rect 7129 951 7130 953
rect 7136 951 7142 953
rect 7156 951 7180 954
rect 7078 948 7180 951
rect 7078 947 7133 948
rect 7136 947 7142 948
rect 7078 946 7112 947
rect 7114 946 7133 947
rect 7145 946 7180 948
rect 7078 944 7133 946
rect 7143 945 7180 946
rect 7142 944 7180 945
rect 7219 953 7242 954
rect 7250 953 7253 954
rect 7363 953 7381 954
rect 7385 953 7411 954
rect 7443 953 7449 959
rect 7470 958 7534 964
rect 7581 963 7587 969
rect 7627 968 7633 969
rect 7622 966 7633 968
rect 7616 964 7621 966
rect 7612 963 7616 964
rect 7627 963 7633 966
rect 7643 968 7677 970
rect 7681 969 7689 970
rect 7476 954 7528 958
rect 7575 957 7581 963
rect 7633 957 7639 963
rect 7219 946 7250 953
rect 7336 946 7375 953
rect 7391 947 7397 953
rect 7437 947 7443 953
rect 7219 944 7242 946
rect 7330 945 7336 946
rect 7325 944 7330 945
rect 6939 938 7180 944
rect 7209 938 7224 944
rect 7232 939 7242 944
rect 7238 938 7242 939
rect 7291 938 7325 944
rect 7476 938 7490 954
rect 7000 922 7016 938
rect 7062 937 7085 938
rect 7062 934 7090 937
rect 7062 933 7098 934
rect 7100 933 7108 935
rect 7129 934 7130 938
rect 7204 937 7209 938
rect 7195 935 7203 936
rect 7131 934 7178 935
rect 7190 934 7195 935
rect 7115 933 7178 934
rect 7242 933 7258 938
rect 7285 936 7291 938
rect 7476 936 7491 938
rect 7281 935 7284 936
rect 7276 933 7280 934
rect 7062 925 7170 933
rect 7129 924 7130 925
rect 7068 922 7085 924
rect 7000 916 7016 920
rect 7051 917 7066 922
rect 7089 920 7114 922
rect 6902 913 6943 916
rect 6947 913 7016 916
rect 6819 911 6822 913
rect 6874 911 6902 913
rect 7000 911 7044 913
rect 7050 911 7066 917
rect 7087 917 7114 920
rect 7133 918 7192 922
rect 7240 920 7276 933
rect 7474 931 7491 936
rect 7470 928 7474 931
rect 7463 924 7470 928
rect 7455 920 7463 924
rect 7476 920 7491 931
rect 7522 920 7524 954
rect 7528 950 7541 954
rect 7643 953 7664 968
rect 7674 967 7677 968
rect 7682 963 7689 969
rect 7717 968 7720 970
rect 7907 969 7921 971
rect 7922 970 8050 971
rect 7932 969 7949 970
rect 7953 969 8050 970
rect 7720 967 7722 968
rect 7722 966 7724 967
rect 7685 960 7687 963
rect 7903 960 7906 961
rect 7690 954 7697 957
rect 7822 953 7823 957
rect 7884 954 7903 960
rect 7907 957 7926 969
rect 7884 953 7908 954
rect 7642 952 7664 953
rect 7642 950 7643 952
rect 7528 942 7536 950
rect 7641 938 7642 949
rect 7698 946 7710 953
rect 7881 952 7884 953
rect 7711 944 7713 945
rect 7713 940 7720 944
rect 7528 920 7536 932
rect 7235 918 7240 920
rect 7115 917 7192 918
rect 7087 915 7099 917
rect 7159 916 7170 917
rect 7107 914 7119 916
rect 7158 915 7160 916
rect 6815 909 6819 911
rect 6873 910 6875 911
rect 6872 909 6876 910
rect 6871 906 6876 909
rect 6818 903 6819 904
rect 6870 903 6876 906
rect 7000 904 7016 911
rect 7044 910 7069 911
rect 7035 908 7066 910
rect 7069 909 7080 910
rect 7080 908 7087 909
rect 7025 906 7066 908
rect 7087 907 7100 908
rect 7108 906 7115 907
rect 7035 905 7066 906
rect 7050 904 7066 905
rect 6809 894 6810 899
rect 6863 896 6864 900
rect 6869 899 6876 903
rect 6868 895 6869 899
rect 6862 876 6864 895
rect 7016 888 7032 904
rect 7034 888 7050 904
rect 7127 888 7129 911
rect 7192 909 7208 917
rect 7224 913 7235 918
rect 7219 911 7223 913
rect 7213 909 7219 911
rect 7242 909 7258 920
rect 7442 912 7455 920
rect 7474 918 7528 920
rect 7539 918 7541 926
rect 7578 920 7581 937
rect 7720 935 7729 940
rect 7816 939 7822 952
rect 7826 946 7847 949
rect 7863 946 7864 949
rect 7875 948 7881 952
rect 7892 946 7908 953
rect 7816 936 7823 939
rect 7824 938 7826 946
rect 7847 939 7908 946
rect 7921 942 7926 957
rect 7949 968 8050 969
rect 8127 968 8128 970
rect 7855 938 7908 939
rect 7874 937 7924 938
rect 7641 925 7644 929
rect 7730 928 7740 934
rect 7816 933 7824 936
rect 7874 933 7881 937
rect 7470 912 7540 918
rect 7575 917 7577 919
rect 7644 918 7659 925
rect 7740 923 7744 928
rect 7744 920 7745 923
rect 7659 917 7682 918
rect 7575 916 7581 917
rect 7573 912 7581 916
rect 7440 911 7442 912
rect 7474 911 7489 912
rect 7490 911 7491 912
rect 7192 908 7258 909
rect 7178 907 7258 908
rect 7434 907 7440 911
rect 7474 907 7495 911
rect 7512 908 7528 912
rect 7136 906 7159 907
rect 7192 904 7258 907
rect 7226 888 7242 904
rect 7420 900 7434 907
rect 7474 904 7489 907
rect 7490 904 7491 907
rect 7522 906 7528 908
rect 7531 904 7540 912
rect 7575 911 7581 912
rect 7633 916 7682 917
rect 7633 911 7639 916
rect 7650 914 7682 916
rect 7659 913 7683 914
rect 7659 911 7682 913
rect 7685 911 7710 913
rect 7724 911 7738 920
rect 7745 918 7746 920
rect 7811 918 7816 933
rect 7822 927 7829 933
rect 7822 925 7824 927
rect 7746 913 7748 918
rect 7748 911 7749 913
rect 7809 911 7811 915
rect 7570 907 7572 911
rect 7475 900 7488 904
rect 7529 900 7531 903
rect 7566 900 7570 907
rect 7581 905 7587 911
rect 7400 888 7423 900
rect 7470 897 7475 900
rect 7454 888 7470 897
rect 7487 896 7490 899
rect 7524 896 7529 899
rect 7564 897 7566 900
rect 7490 888 7506 896
rect 7508 888 7524 896
rect 7558 888 7564 897
rect 6868 875 6876 888
rect 7064 880 7194 888
rect 7397 883 7400 888
rect 7446 883 7454 888
rect 7555 883 7558 888
rect 7312 880 7360 883
rect 7042 875 7084 880
rect 6862 873 6868 875
rect 7031 873 7084 875
rect 6819 870 6823 873
rect 6852 871 6862 873
rect 6865 872 6868 873
rect 6852 870 6864 871
rect 7012 870 7084 873
rect 7127 870 7129 880
rect 7171 879 7312 880
rect 7174 875 7312 879
rect 7360 875 7361 880
rect 7393 875 7397 883
rect 7432 876 7446 883
rect 7550 876 7555 883
rect 7426 875 7432 876
rect 7593 875 7617 910
rect 7627 905 7633 911
rect 7659 909 7738 911
rect 7749 909 7750 911
rect 7672 904 7738 909
rect 7750 904 7752 908
rect 7688 888 7704 904
rect 7706 893 7722 904
rect 7752 899 7754 903
rect 7754 893 7756 899
rect 7797 898 7809 910
rect 7818 909 7822 925
rect 7855 916 7863 933
rect 7869 927 7875 933
rect 7817 904 7818 909
rect 7835 905 7855 915
rect 7822 903 7834 905
rect 7835 903 7856 905
rect 7874 904 7875 927
rect 7908 922 7924 937
rect 7926 936 7927 941
rect 7949 938 7970 968
rect 7990 967 8050 968
rect 8128 967 8129 968
rect 7999 965 8050 967
rect 8129 965 8132 967
rect 8019 963 8050 965
rect 8132 963 8134 965
rect 8028 961 8050 963
rect 8134 961 8138 963
rect 7982 938 7998 954
rect 8000 938 8016 954
rect 8040 949 8068 961
rect 8138 954 8147 961
rect 8026 938 8027 949
rect 8068 947 8072 949
rect 8147 947 8155 954
rect 8072 946 8073 947
rect 8073 944 8074 946
rect 8155 944 8157 947
rect 8343 944 8344 949
rect 8372 944 8388 954
rect 8074 939 8080 944
rect 8157 940 8162 944
rect 8326 940 8393 944
rect 8162 939 8164 940
rect 8303 939 8326 940
rect 7949 936 7982 938
rect 8016 937 8032 938
rect 7996 936 8032 937
rect 8080 936 8082 938
rect 8164 936 8167 939
rect 8300 936 8303 939
rect 8343 938 8344 940
rect 8393 938 8394 939
rect 7927 916 7932 933
rect 7949 922 7981 936
rect 7996 935 8016 936
rect 8018 934 8032 936
rect 8082 934 8084 936
rect 8167 934 8171 936
rect 8297 934 8300 936
rect 8012 932 8032 934
rect 8084 932 8085 934
rect 8171 932 8173 934
rect 8296 932 8297 934
rect 7933 915 7939 921
rect 7949 919 7970 922
rect 7974 921 7981 922
rect 7970 915 7973 919
rect 7974 915 7985 921
rect 7927 909 7933 915
rect 7932 908 7933 909
rect 7974 906 7981 915
rect 7985 909 7991 915
rect 8023 904 8059 932
rect 8085 925 8092 932
rect 8173 925 8184 932
rect 8293 925 8296 932
rect 8092 924 8106 925
rect 8084 915 8106 924
rect 8184 919 8193 925
rect 8290 919 8293 925
rect 8193 916 8196 919
rect 8289 916 8290 919
rect 8092 907 8106 915
rect 8196 912 8201 916
rect 8287 912 8289 916
rect 8201 907 8205 912
rect 8284 910 8287 912
rect 8100 905 8109 907
rect 8106 904 8109 905
rect 8205 904 8207 907
rect 8031 903 8034 904
rect 8059 903 8060 904
rect 8109 903 8110 904
rect 7819 901 7859 903
rect 7816 900 7817 901
rect 7815 899 7816 900
rect 7819 899 7855 901
rect 7859 899 7860 901
rect 7814 898 7819 899
rect 7797 896 7819 898
rect 7757 893 7809 896
rect 7814 893 7819 896
rect 7706 888 7725 893
rect 7756 888 7809 893
rect 7653 877 7662 881
rect 7700 877 7709 881
rect 7719 879 7725 888
rect 7751 886 7763 888
rect 7746 883 7751 886
rect 7756 883 7763 886
rect 7745 882 7763 883
rect 7737 880 7763 882
rect 7734 879 7763 880
rect 7719 877 7763 879
rect 7645 875 7763 877
rect 7174 870 7276 875
rect 7314 874 7468 875
rect 7314 872 7461 874
rect 7287 871 7314 872
rect 7393 871 7397 872
rect 7426 871 7432 872
rect 7468 871 7482 874
rect 7548 871 7550 875
rect 7587 872 7645 875
rect 7653 872 7756 875
rect 7279 870 7287 871
rect 7482 870 7486 871
rect 7587 870 7653 872
rect 7654 870 7756 872
rect 7763 870 7765 875
rect 7797 872 7809 888
rect 7810 881 7815 893
rect 7814 880 7815 881
rect 7835 871 7855 899
rect 7860 893 7863 899
rect 7863 881 7868 893
rect 7971 887 7974 903
rect 8027 902 8031 903
rect 8026 899 8027 901
rect 8060 899 8066 903
rect 8019 893 8026 899
rect 8031 897 8032 899
rect 8065 893 8066 899
rect 8101 893 8108 898
rect 8110 893 8124 903
rect 8019 887 8025 893
rect 7863 877 7867 881
rect 7974 877 7999 887
rect 8108 885 8120 893
rect 8124 887 8133 893
rect 8207 887 8220 903
rect 8280 902 8292 910
rect 8302 902 8314 910
rect 8354 904 8355 938
rect 8393 934 8404 938
rect 8394 922 8404 934
rect 8394 903 8395 922
rect 8280 898 8283 902
rect 8316 899 8318 902
rect 8268 886 8276 898
rect 8280 896 8314 898
rect 8280 895 8283 896
rect 7867 873 7868 875
rect 7999 870 8017 877
rect 8019 875 8025 877
rect 8120 876 8127 885
rect 8133 879 8139 886
rect 8220 879 8225 886
rect 8139 877 8141 879
rect 8225 877 8227 879
rect 8019 870 8026 875
rect 8031 870 8032 872
rect 8141 871 8144 877
rect 8227 870 8231 877
rect 6823 869 6852 870
rect 6860 867 6864 870
rect 7008 869 7012 870
rect 7274 869 7279 870
rect 7362 869 7363 870
rect 6859 866 6864 867
rect 6995 866 7008 869
rect 7265 868 7274 869
rect 7257 866 7265 868
rect 7363 867 7364 869
rect 6807 859 6808 866
rect 6857 864 6864 866
rect 6973 865 7007 866
rect 7252 865 7257 866
rect 6857 859 6859 864
rect 6973 862 6995 865
rect 6972 859 6995 862
rect 7007 859 7014 865
rect 7219 859 7252 865
rect 6856 855 6857 859
rect 6968 855 6973 859
rect 6976 854 6995 859
rect 7014 857 7017 859
rect 7213 858 7219 859
rect 7206 857 7213 858
rect 7190 854 7205 857
rect 7364 854 7369 866
rect 7391 863 7393 870
rect 7423 863 7426 870
rect 7486 868 7498 870
rect 7390 860 7391 863
rect 7422 860 7423 863
rect 7498 859 7536 868
rect 7541 863 7546 870
rect 7576 869 7587 870
rect 7564 868 7576 869
rect 7562 866 7564 868
rect 7559 864 7562 866
rect 7589 864 7592 869
rect 7539 860 7541 863
rect 6855 851 6856 854
rect 6966 851 6968 854
rect 6975 850 6976 854
rect 6806 838 6807 850
rect 6851 838 6855 850
rect 6959 838 6966 850
rect 5260 812 5276 818
rect 5278 812 5294 818
rect 6805 816 6806 837
rect 6844 816 6851 838
rect 6959 835 6965 838
rect 6953 829 6959 835
rect 6967 828 6972 842
rect 7005 835 7011 841
rect 7017 839 7018 854
rect 7094 850 7190 854
rect 7369 850 7370 854
rect 7388 853 7390 859
rect 7419 853 7422 859
rect 7531 858 7541 859
rect 7531 853 7538 858
rect 7541 857 7547 858
rect 7556 857 7559 864
rect 7644 863 7653 870
rect 7709 863 7718 870
rect 7727 868 7728 870
rect 7765 868 7766 870
rect 7587 860 7589 863
rect 7728 861 7730 868
rect 7766 860 7769 868
rect 7795 864 7796 866
rect 7794 861 7795 863
rect 7810 859 7816 870
rect 7832 864 7835 870
rect 7868 866 7870 870
rect 8017 869 8027 870
rect 7907 868 7908 869
rect 7906 867 7907 868
rect 7905 865 7906 866
rect 7898 864 7905 865
rect 7822 859 7824 861
rect 7547 855 7570 857
rect 7585 856 7587 859
rect 7547 854 7560 855
rect 7580 854 7585 856
rect 7531 852 7534 853
rect 7531 851 7533 852
rect 7555 851 7556 854
rect 7560 851 7601 854
rect 7646 851 7652 857
rect 7692 851 7698 857
rect 7731 855 7732 857
rect 7770 854 7771 857
rect 7792 856 7793 859
rect 7818 856 7826 859
rect 7779 854 7818 856
rect 7828 855 7832 863
rect 7856 859 7898 864
rect 7927 863 7933 869
rect 7985 863 7991 869
rect 8019 867 8027 869
rect 8127 868 8128 870
rect 8144 869 8145 870
rect 8028 867 8037 868
rect 8019 866 8040 867
rect 8019 865 8027 866
rect 8028 865 8040 866
rect 8100 865 8102 868
rect 8145 867 8146 869
rect 8231 867 8233 869
rect 8280 868 8282 895
rect 8146 865 8147 866
rect 8028 863 8037 865
rect 7827 854 7828 855
rect 7702 851 7779 854
rect 7791 853 7792 854
rect 7820 853 7833 854
rect 7034 843 7095 850
rect 7033 841 7034 842
rect 7011 832 7017 835
rect 7018 832 7019 838
rect 7011 829 7019 832
rect 7027 829 7033 841
rect 7037 840 7048 842
rect 7094 840 7095 843
rect 7105 843 7295 850
rect 7370 846 7373 850
rect 7380 846 7388 851
rect 7411 847 7419 851
rect 7406 846 7467 847
rect 7317 843 7399 846
rect 7105 839 7190 843
rect 7283 842 7301 843
rect 7370 842 7373 843
rect 7265 839 7283 842
rect 7301 841 7313 842
rect 7316 839 7319 841
rect 7103 838 7105 839
rect 7098 835 7102 838
rect 7092 830 7098 835
rect 7125 831 7127 839
rect 7257 838 7265 839
rect 7241 835 7257 838
rect 7015 828 7019 829
rect 7091 828 7092 830
rect 5260 809 5294 812
rect 6804 810 6805 816
rect 6843 811 6844 816
rect 6872 811 6888 824
rect 6966 813 6967 828
rect 7011 826 7013 827
rect 7015 826 7027 828
rect 7013 816 7035 826
rect 7064 817 7080 824
rect 7011 812 7035 816
rect 7054 812 7080 817
rect 7011 811 7013 812
rect 5260 808 5306 809
rect 5209 790 5212 800
rect 5216 794 5225 803
rect 5237 792 5260 808
rect 5272 803 5281 808
rect 5306 805 5311 808
rect 6841 807 6843 810
rect 7017 808 7019 811
rect 5281 794 5290 803
rect 5199 787 5214 790
rect 5147 779 5153 786
rect 5172 780 5214 787
rect 5220 786 5224 792
rect 5237 790 5247 792
rect 5237 787 5260 790
rect 5216 780 5218 784
rect 5237 781 5274 787
rect 5148 774 5164 779
rect 5172 774 5216 780
rect 5244 774 5274 781
rect 5311 774 5327 805
rect 6803 800 6804 805
rect 6838 800 6840 805
rect 6837 798 6838 800
rect 6833 790 6837 798
rect 6856 792 6867 808
rect 7016 806 7017 808
rect 7035 807 7044 812
rect 7052 809 7080 812
rect 7050 808 7061 809
rect 7064 808 7080 809
rect 7082 808 7098 824
rect 7121 818 7127 831
rect 7207 830 7241 835
rect 7165 823 7207 830
rect 7319 829 7321 839
rect 7373 829 7378 842
rect 7380 828 7388 843
rect 7157 822 7165 823
rect 7132 818 7157 822
rect 7121 816 7132 818
rect 7117 812 7127 816
rect 7048 807 7064 808
rect 7044 806 7064 807
rect 7044 805 7061 806
rect 7098 805 7114 808
rect 6966 790 6967 805
rect 6831 786 6833 790
rect 6952 787 6967 790
rect 7005 789 7016 805
rect 7042 803 7075 805
rect 7042 794 7070 803
rect 7092 797 7114 805
rect 7042 793 7064 794
rect 7048 792 7064 793
rect 7054 790 7064 792
rect 7088 792 7114 797
rect 7088 791 7098 792
rect 7005 787 7017 789
rect 6802 782 6803 786
rect 6952 783 7017 787
rect 7048 787 7064 790
rect 7081 790 7098 791
rect 7081 787 7114 790
rect 7048 783 7114 787
rect 6952 782 7016 783
rect 4950 761 5006 774
rect 5008 763 5016 774
rect 5038 763 5041 774
rect 5059 764 5060 770
rect 4878 753 4881 758
rect 4917 758 5006 761
rect 5037 760 5040 763
rect 5091 760 5102 774
rect 4307 745 4366 749
rect 4488 746 4495 750
rect 4649 748 4659 752
rect 4696 749 4698 753
rect 4527 746 4624 748
rect 4647 746 4659 748
rect 4695 746 4696 748
rect 4487 745 4495 746
rect 4498 745 4633 746
rect 4644 745 4646 746
rect 4649 745 4659 746
rect 4194 741 4246 744
rect 4249 742 4250 744
rect 4188 736 4252 741
rect 4307 740 4446 745
rect 4487 744 4659 745
rect 4188 735 4254 736
rect 4109 730 4115 731
rect 4030 727 4132 730
rect 4030 724 4157 727
rect 4166 725 4173 731
rect 4194 729 4200 735
rect 4209 727 4212 732
rect 4240 729 4246 735
rect 4251 727 4254 735
rect 4213 725 4214 727
rect 4254 725 4255 727
rect 4307 726 4315 740
rect 4359 736 4446 740
rect 4361 730 4446 736
rect 4479 743 4659 744
rect 4691 743 4695 745
rect 4705 744 4723 753
rect 4827 750 4829 753
rect 4858 750 4860 753
rect 4728 744 4768 745
rect 4769 744 4780 750
rect 4479 740 4656 743
rect 4479 732 4493 740
rect 4691 735 4705 743
rect 4368 729 4369 730
rect 4369 727 4370 729
rect 3746 713 3747 724
rect 3785 717 3786 724
rect 4030 720 4079 724
rect 4030 717 4086 720
rect 4115 719 4121 724
rect 4030 716 4038 717
rect 4030 715 4037 716
rect 3786 711 3787 713
rect 4049 712 4051 717
rect 4079 710 4086 717
rect 3745 707 3746 710
rect 3930 707 4013 710
rect 4051 696 4054 709
rect 4086 708 4096 709
rect 4064 700 4076 708
rect 4086 700 4098 708
rect 4055 698 4060 700
rect 4062 698 4107 700
rect 4055 697 4107 698
rect 4133 697 4135 722
rect 4161 719 4167 725
rect 4214 723 4215 725
rect 4255 720 4256 722
rect 4301 720 4317 726
rect 4217 715 4219 719
rect 4256 716 4257 719
rect 4303 716 4317 720
rect 4321 716 4324 719
rect 4347 718 4349 726
rect 4359 720 4365 726
rect 4446 725 4455 730
rect 4371 723 4372 725
rect 4346 716 4349 718
rect 4353 716 4361 720
rect 4219 709 4223 715
rect 4257 710 4259 715
rect 4303 714 4313 716
rect 4303 713 4312 714
rect 4315 713 4336 716
rect 4346 713 4348 716
rect 4351 713 4361 716
rect 4312 710 4313 713
rect 4324 710 4327 713
rect 4340 712 4344 713
rect 4344 711 4349 712
rect 4351 711 4353 713
rect 4336 710 4351 711
rect 4372 710 4379 722
rect 4455 713 4460 724
rect 4487 722 4493 732
rect 4616 723 4622 729
rect 4632 727 4638 732
rect 4627 723 4632 727
rect 4662 723 4668 729
rect 4688 727 4691 735
rect 4692 727 4705 735
rect 4688 725 4692 727
rect 4713 726 4721 744
rect 4728 740 4780 744
rect 4726 735 4762 740
rect 4768 737 4780 740
rect 4829 747 4832 750
rect 4768 735 4785 737
rect 4726 731 4728 735
rect 4769 734 4785 735
rect 4829 734 4834 747
rect 4779 731 4785 734
rect 4780 730 4785 731
rect 4783 729 4787 730
rect 4832 729 4834 734
rect 4785 726 4789 729
rect 4479 719 4493 722
rect 4479 716 4495 719
rect 4547 716 4548 719
rect 4610 717 4616 723
rect 4668 717 4674 723
rect 4684 722 4688 724
rect 4689 723 4692 725
rect 4715 724 4716 726
rect 4787 725 4789 726
rect 4833 725 4834 729
rect 4721 724 4722 725
rect 4224 698 4230 708
rect 4260 698 4262 708
rect 4315 701 4327 710
rect 4328 698 4334 708
rect 4337 701 4349 710
rect 4351 709 4416 710
rect 4358 707 4416 709
rect 4365 706 4416 707
rect 4373 703 4416 706
rect 4379 700 4385 703
rect 4387 702 4416 703
rect 4388 701 4416 702
rect 4379 698 4393 700
rect 4230 697 4234 698
rect 4055 696 4234 697
rect 3744 692 3745 696
rect 4051 695 4060 696
rect 4052 694 4060 695
rect 4064 694 4234 696
rect 4262 694 4266 698
rect 3749 690 3750 692
rect 3747 676 3750 690
rect 3744 670 3747 676
rect 3737 663 3747 670
rect 3749 663 3750 676
rect 3782 690 3783 692
rect 3784 690 3794 692
rect 3782 687 3809 690
rect 4049 688 4055 694
rect 3782 673 3813 687
rect 4052 684 4055 688
rect 4064 692 4160 694
rect 4064 690 4192 692
rect 4230 691 4289 694
rect 4230 690 4234 691
rect 4262 690 4266 691
rect 4289 690 4293 691
rect 4334 690 4335 696
rect 4385 695 4393 698
rect 4395 697 4416 701
rect 4457 709 4461 713
rect 4479 712 4497 716
rect 4522 712 4525 713
rect 4479 711 4495 712
rect 4479 710 4493 711
rect 4487 709 4495 710
rect 4497 709 4499 711
rect 4500 710 4525 712
rect 4540 710 4542 712
rect 4547 710 4553 715
rect 4601 710 4616 716
rect 4683 715 4688 722
rect 4676 711 4682 714
rect 4684 711 4688 715
rect 4710 716 4727 724
rect 4506 709 4608 710
rect 4457 707 4462 709
rect 4487 707 4493 709
rect 4528 707 4608 709
rect 4457 706 4463 707
rect 4490 706 4528 707
rect 4457 702 4464 706
rect 4457 701 4465 702
rect 4428 698 4438 699
rect 4457 698 4467 701
rect 4490 698 4503 706
rect 4541 703 4547 707
rect 4552 706 4608 707
rect 4676 709 4684 711
rect 4676 706 4682 709
rect 4710 708 4732 716
rect 4724 706 4732 708
rect 4743 706 4749 712
rect 4552 705 4621 706
rect 4668 705 4676 706
rect 4552 703 4676 705
rect 4552 700 4589 703
rect 4421 697 4425 698
rect 4403 695 4421 697
rect 4379 694 4421 695
rect 4439 696 4467 698
rect 4385 692 4416 694
rect 4385 691 4404 692
rect 4382 690 4390 691
rect 4064 688 4113 690
rect 4064 683 4098 688
rect 4064 682 4072 683
rect 4064 681 4071 682
rect 3964 673 3998 676
rect 3782 663 3783 673
rect 3788 663 3795 670
rect 3737 658 3795 663
rect 3812 660 3813 673
rect 3743 657 3788 658
rect 3743 653 3744 657
rect 3747 654 3785 657
rect 3749 646 3761 654
rect 3771 646 3783 654
rect 3743 630 3752 644
rect 3822 642 3823 671
rect 4105 663 4107 688
rect 4133 663 4135 690
rect 4196 688 4199 690
rect 4235 687 4236 690
rect 4293 688 4297 690
rect 4375 688 4382 690
rect 4236 678 4242 687
rect 4269 678 4276 687
rect 4285 685 4308 688
rect 4366 687 4375 688
rect 4285 684 4310 685
rect 4285 683 4331 684
rect 4335 683 4337 687
rect 4361 685 4366 687
rect 4358 684 4361 685
rect 4356 683 4358 684
rect 4285 682 4356 683
rect 4393 682 4402 691
rect 4409 690 4416 692
rect 4439 692 4469 696
rect 4439 691 4470 692
rect 4488 691 4490 698
rect 4552 691 4585 700
rect 4668 695 4676 703
rect 4710 693 4732 706
rect 4737 700 4743 706
rect 4783 700 4785 725
rect 4787 713 4797 725
rect 4833 719 4839 725
rect 4860 719 4875 750
rect 4881 749 4882 753
rect 4917 751 5004 758
rect 5032 753 5038 760
rect 5082 758 5102 760
rect 5164 758 5180 774
rect 5182 770 5198 774
rect 5200 771 5207 774
rect 5211 773 5216 774
rect 5200 770 5206 771
rect 5209 770 5211 773
rect 5246 770 5252 774
rect 5182 764 5200 770
rect 5252 764 5258 770
rect 5182 758 5198 764
rect 5260 760 5274 774
rect 5327 761 5335 774
rect 6801 771 6802 781
rect 6830 773 6831 782
rect 6952 774 7018 782
rect 7042 774 7114 783
rect 7121 777 7125 812
rect 7149 803 7158 812
rect 7178 808 7194 823
rect 7196 803 7205 812
rect 7256 808 7272 824
rect 7274 808 7290 824
rect 7321 813 7325 828
rect 7378 825 7388 828
rect 7411 825 7419 846
rect 7468 843 7481 846
rect 7485 842 7487 843
rect 7489 842 7531 851
rect 7487 839 7531 842
rect 7489 835 7531 839
rect 7547 846 7601 851
rect 7640 850 7646 851
rect 7698 850 7779 851
rect 7606 846 7704 850
rect 7733 849 7735 850
rect 7744 849 7753 850
rect 7730 847 7740 849
rect 7745 848 7753 849
rect 7547 835 7577 846
rect 7601 845 7704 846
rect 7601 843 7613 845
rect 7628 843 7646 845
rect 7600 842 7601 843
rect 7735 842 7736 845
rect 7489 830 7577 835
rect 7589 831 7600 842
rect 7771 840 7777 850
rect 7489 825 7531 830
rect 7541 828 7565 830
rect 7588 828 7589 831
rect 7737 830 7740 838
rect 7778 830 7781 838
rect 7784 830 7790 850
rect 7811 839 7833 853
rect 7872 840 7877 858
rect 7933 857 7939 863
rect 7933 841 7938 857
rect 7975 841 7977 863
rect 7979 857 7985 863
rect 8027 862 8037 863
rect 8028 861 8037 862
rect 8028 859 8043 861
rect 8100 859 8106 865
rect 8147 864 8148 865
rect 8031 856 8056 859
rect 8031 853 8046 856
rect 8048 853 8054 856
rect 8084 854 8093 859
rect 8094 854 8100 859
rect 8130 857 8131 861
rect 8148 859 8150 864
rect 8150 856 8152 859
rect 8152 854 8153 856
rect 8233 854 8241 866
rect 8280 864 8283 868
rect 8312 864 8314 896
rect 8318 889 8326 898
rect 8318 879 8345 889
rect 8392 881 8395 885
rect 8385 879 8392 881
rect 8318 870 8385 879
rect 8339 869 8343 870
rect 8325 866 8339 869
rect 8320 865 8325 866
rect 8316 864 8320 865
rect 8276 856 8277 861
rect 8275 854 8277 856
rect 8037 850 8046 853
rect 8084 850 8103 854
rect 8092 846 8103 850
rect 8103 842 8104 846
rect 8131 842 8134 854
rect 8153 850 8155 854
rect 8241 851 8243 854
rect 8155 845 8159 850
rect 8159 843 8161 845
rect 8243 844 8248 850
rect 8161 842 8162 843
rect 8162 841 8164 842
rect 7933 839 7966 841
rect 7740 828 7741 830
rect 7541 825 7550 828
rect 7324 808 7325 813
rect 7376 824 7383 825
rect 7376 814 7386 824
rect 7376 812 7380 814
rect 7383 812 7386 814
rect 7408 813 7410 824
rect 7448 814 7464 824
rect 7441 813 7464 814
rect 7466 813 7489 824
rect 7533 820 7541 825
rect 7545 824 7550 825
rect 7209 803 7210 808
rect 7140 794 7153 803
rect 7205 794 7214 803
rect 7149 787 7153 794
rect 7209 792 7210 794
rect 7240 792 7256 808
rect 7291 807 7306 808
rect 7375 807 7376 811
rect 7384 808 7386 812
rect 7292 799 7306 807
rect 7325 800 7326 807
rect 7374 804 7375 807
rect 7373 800 7374 803
rect 7386 800 7402 808
rect 7407 807 7408 812
rect 7441 808 7482 813
rect 7432 806 7453 808
rect 7464 807 7470 808
rect 7406 800 7407 806
rect 7432 802 7448 806
rect 7458 802 7464 807
rect 7429 801 7475 802
rect 7429 800 7470 801
rect 7246 790 7252 792
rect 7255 791 7256 792
rect 7283 792 7306 799
rect 7326 797 7328 800
rect 7283 791 7298 792
rect 7254 790 7256 791
rect 7240 787 7256 790
rect 7257 789 7259 790
rect 7292 789 7298 791
rect 7257 787 7298 789
rect 7328 787 7338 797
rect 7370 787 7373 797
rect 7386 792 7406 800
rect 7401 790 7406 792
rect 7429 792 7448 800
rect 7482 792 7498 808
rect 7510 807 7516 813
rect 7523 812 7533 820
rect 7544 813 7550 824
rect 7565 823 7591 828
rect 7555 822 7598 823
rect 7555 821 7596 822
rect 7585 813 7588 821
rect 7598 818 7605 822
rect 7605 816 7606 818
rect 7517 807 7523 812
rect 7544 809 7545 813
rect 7606 812 7609 816
rect 7640 813 7656 824
rect 7658 813 7674 824
rect 7709 816 7718 825
rect 7741 824 7742 828
rect 7698 815 7709 816
rect 7631 812 7633 813
rect 7671 812 7675 813
rect 7584 809 7585 811
rect 7631 810 7675 812
rect 7631 808 7665 810
rect 7516 801 7522 807
rect 7528 792 7544 808
rect 7429 790 7439 792
rect 7441 790 7448 792
rect 7240 785 7295 787
rect 7151 777 7152 785
rect 7213 777 7219 783
rect 7240 781 7263 785
rect 6831 768 6832 771
rect 6968 767 6984 774
rect 6986 767 7002 774
rect 7042 771 7050 774
rect 7054 771 7100 774
rect 7050 767 7053 769
rect 7064 767 7080 771
rect 7082 767 7098 771
rect 5260 758 5277 760
rect 5082 753 5091 758
rect 5099 755 5100 757
rect 5271 753 5277 758
rect 5307 753 5319 761
rect 5327 756 5341 761
rect 5329 753 5341 756
rect 4917 749 5002 751
rect 5027 750 5040 753
rect 4882 746 4883 748
rect 4917 745 5008 749
rect 5020 748 5040 750
rect 5076 748 5082 753
rect 5020 746 5038 748
rect 5075 746 5076 748
rect 5024 745 5038 746
rect 4883 735 4885 744
rect 4936 743 5038 745
rect 4936 740 4968 743
rect 4984 740 5038 743
rect 4885 732 4886 735
rect 4886 730 4887 731
rect 4887 726 4888 730
rect 4936 729 5038 740
rect 5061 732 5063 743
rect 5070 740 5075 746
rect 5100 742 5103 753
rect 5067 736 5070 740
rect 5066 735 5067 736
rect 5064 732 5066 735
rect 5059 730 5064 732
rect 4947 727 4951 729
rect 4988 728 4992 729
rect 4946 725 4951 727
rect 4987 725 4988 727
rect 5049 725 5059 730
rect 4879 719 4885 725
rect 4888 721 4892 724
rect 4945 722 4951 725
rect 5007 724 5059 725
rect 4944 721 4951 722
rect 4985 721 4986 722
rect 5007 721 5049 724
rect 4827 713 4833 719
rect 4885 713 4891 719
rect 4892 717 4991 721
rect 5007 717 5042 721
rect 5061 720 5063 730
rect 5103 724 5104 742
rect 5206 740 5232 753
rect 5235 748 5240 753
rect 5277 748 5280 753
rect 5303 750 5304 752
rect 5335 749 5341 753
rect 5235 747 5241 748
rect 5235 740 5240 747
rect 5280 746 5282 748
rect 5295 746 5303 749
rect 5307 747 5341 749
rect 5338 746 5341 747
rect 5241 740 5242 746
rect 5282 740 5287 746
rect 5288 740 5301 746
rect 5104 719 5107 724
rect 5060 717 5061 719
rect 5194 718 5200 731
rect 5205 724 5206 730
rect 5242 726 5244 740
rect 5206 722 5208 724
rect 5206 721 5210 722
rect 5238 721 5240 724
rect 5206 719 5240 721
rect 5244 719 5246 726
rect 5264 725 5265 727
rect 5287 726 5301 740
rect 5252 722 5258 724
rect 5252 719 5262 722
rect 5288 720 5305 726
rect 5232 718 5262 719
rect 4787 712 4789 713
rect 4787 707 4795 712
rect 4892 707 5033 717
rect 5034 712 5042 717
rect 5200 716 5206 718
rect 5242 717 5252 718
rect 5242 716 5244 717
rect 5113 715 5115 716
rect 5200 715 5244 716
rect 5056 712 5058 715
rect 4789 706 4795 707
rect 4789 700 4801 706
rect 4412 687 4416 690
rect 4414 685 4416 687
rect 4415 683 4416 685
rect 4457 690 4470 691
rect 4457 687 4471 690
rect 4457 683 4479 687
rect 4335 678 4337 682
rect 4199 673 4200 676
rect 4197 668 4200 673
rect 4242 671 4246 678
rect 4276 671 4281 678
rect 4415 677 4419 683
rect 4457 679 4476 683
rect 4479 682 4481 683
rect 4484 682 4488 690
rect 4555 686 4575 691
rect 4549 683 4575 686
rect 4548 682 4575 683
rect 4585 682 4594 691
rect 4710 690 4727 693
rect 4732 691 4733 693
rect 4734 689 4738 690
rect 4789 689 4795 700
rect 4817 698 4826 700
rect 4817 691 4830 698
rect 4726 687 4738 689
rect 4787 688 4795 689
rect 4783 687 4787 688
rect 4726 685 4741 687
rect 4772 685 4783 687
rect 4726 683 4761 685
rect 4765 683 4772 685
rect 4481 681 4488 682
rect 4535 681 4575 682
rect 4481 680 4517 681
rect 4535 680 4547 681
rect 4484 679 4505 680
rect 4526 679 4558 680
rect 4457 678 4554 679
rect 4457 677 4476 678
rect 4348 675 4358 676
rect 4419 675 4420 676
rect 4476 675 4478 676
rect 4361 674 4369 675
rect 4366 671 4380 674
rect 4246 668 4248 671
rect 4190 667 4200 668
rect 4218 667 4229 668
rect 4173 664 4190 667
rect 4162 663 4173 664
rect 4055 662 4173 663
rect 4197 662 4200 667
rect 4229 666 4250 667
rect 4229 664 4252 666
rect 4249 663 4264 664
rect 4284 663 4289 668
rect 4380 667 4382 671
rect 4396 664 4407 667
rect 4391 663 4396 664
rect 4249 662 4396 663
rect 4055 659 4162 662
rect 4055 657 4141 659
rect 4196 657 4197 659
rect 4055 656 4129 657
rect 4055 655 4125 656
rect 4055 654 4118 655
rect 4055 653 4113 654
rect 4055 648 4107 653
rect 4049 642 4113 648
rect 3752 626 3756 630
rect 3812 626 3828 642
rect 4055 636 4061 642
rect 4071 638 4077 642
rect 4077 634 4082 638
rect 4101 636 4107 642
rect 4133 634 4135 657
rect 4192 642 4196 657
rect 4252 655 4256 660
rect 4264 659 4391 662
rect 4420 660 4427 675
rect 4477 671 4480 675
rect 4484 674 4488 678
rect 4610 675 4616 677
rect 4588 674 4616 675
rect 4483 672 4484 674
rect 4581 672 4589 674
rect 4610 671 4618 674
rect 4668 671 4674 677
rect 4726 674 4742 683
rect 4466 668 4483 671
rect 4434 664 4448 667
rect 4448 663 4454 664
rect 4461 663 4481 668
rect 4616 665 4622 671
rect 4662 665 4668 671
rect 4570 663 4573 664
rect 4789 663 4795 688
rect 4808 682 4823 691
rect 4936 689 4942 707
rect 4969 706 4984 707
rect 4969 705 4998 706
rect 4448 662 4573 663
rect 4454 660 4570 662
rect 4743 660 4795 663
rect 4461 659 4570 660
rect 4290 657 4379 659
rect 4290 654 4294 657
rect 4307 656 4372 657
rect 4311 655 4369 656
rect 4321 654 4363 655
rect 4256 652 4257 654
rect 4294 652 4295 654
rect 4327 653 4363 654
rect 4257 649 4259 652
rect 4260 642 4265 648
rect 4295 642 4304 652
rect 4337 644 4338 646
rect 4328 642 4343 644
rect 4192 634 4206 642
rect 4304 639 4306 642
rect 4328 639 4344 642
rect 4306 637 4307 639
rect 4328 637 4355 639
rect 4082 632 4149 634
rect 3756 624 3812 626
rect 3796 610 3812 624
rect 4133 614 4135 632
rect 4140 630 4152 632
rect 4191 630 4206 634
rect 4308 633 4311 637
rect 4328 635 4337 637
rect 4341 635 4386 637
rect 4393 635 4402 644
rect 4140 626 4156 630
rect 4190 626 4206 630
rect 4156 610 4172 626
rect 4174 610 4190 626
rect 4274 615 4291 633
rect 4309 625 4331 633
rect 4337 626 4346 635
rect 4384 626 4393 635
rect 4427 630 4442 659
rect 4464 657 4562 659
rect 4464 655 4470 657
rect 4475 656 4557 657
rect 4477 655 4557 656
rect 4479 652 4551 655
rect 4737 654 4801 660
rect 4458 650 4461 652
rect 4479 651 4538 652
rect 4479 650 4494 651
rect 4504 650 4510 651
rect 4451 645 4457 649
rect 4479 645 4502 650
rect 4513 645 4532 650
rect 4743 648 4749 654
rect 4758 652 4759 654
rect 4759 650 4760 652
rect 4479 644 4499 645
rect 4479 642 4481 644
rect 4483 642 4499 644
rect 4523 642 4532 645
rect 4760 644 4762 649
rect 4789 648 4795 654
rect 4444 639 4448 642
rect 4479 641 4499 642
rect 4479 634 4494 641
rect 4520 635 4532 642
rect 4585 635 4594 644
rect 4789 642 4790 648
rect 4817 645 4823 682
rect 4843 677 4846 683
rect 4879 676 4881 683
rect 4827 667 4833 673
rect 4834 667 4843 676
rect 4833 663 4843 667
rect 4847 663 4849 673
rect 4879 671 4882 676
rect 4931 674 4936 689
rect 4878 667 4882 671
rect 4885 667 4891 673
rect 4969 672 4984 705
rect 5015 704 5019 705
rect 5039 694 5049 705
rect 5115 694 5183 715
rect 5200 712 5218 715
rect 5205 708 5218 712
rect 5246 712 5252 717
rect 5285 715 5287 718
rect 5298 716 5305 720
rect 5305 715 5307 716
rect 5339 715 5341 746
rect 5345 737 5353 749
rect 6800 743 6801 767
rect 6832 742 6835 767
rect 6968 759 7002 767
rect 7054 759 7098 767
rect 6968 758 6984 759
rect 6986 758 7005 759
rect 7064 758 7080 759
rect 7082 758 7098 759
rect 7121 763 7124 777
rect 7126 763 7132 771
rect 6990 753 7005 758
rect 7121 757 7132 763
rect 7061 753 7070 756
rect 7115 754 7132 757
rect 7149 756 7152 777
rect 7097 753 7132 754
rect 6934 740 7132 753
rect 7140 747 7152 756
rect 7218 771 7225 777
rect 7240 774 7261 781
rect 7005 738 7014 740
rect 7020 737 7126 740
rect 7149 738 7158 747
rect 7160 741 7167 747
rect 6835 733 6836 737
rect 5345 715 5353 727
rect 6836 724 6837 731
rect 7098 730 7100 737
rect 7121 730 7127 737
rect 7218 731 7219 771
rect 7246 753 7261 774
rect 7293 778 7294 785
rect 7298 778 7307 787
rect 7293 756 7295 778
rect 7299 775 7307 778
rect 7336 782 7351 787
rect 7368 782 7370 787
rect 7386 782 7406 790
rect 7336 778 7406 782
rect 7432 780 7448 790
rect 7336 774 7411 778
rect 7352 772 7368 774
rect 7370 772 7386 774
rect 7401 772 7411 774
rect 7429 774 7448 780
rect 7482 774 7498 790
rect 7528 780 7544 790
rect 7579 789 7584 808
rect 7614 803 7616 806
rect 7624 805 7640 808
rect 7675 807 7690 808
rect 7700 807 7709 815
rect 7736 810 7752 824
rect 7754 810 7770 824
rect 7781 823 7784 830
rect 7781 818 7786 823
rect 7780 816 7781 818
rect 7784 816 7786 818
rect 7811 816 7827 839
rect 7834 830 7841 838
rect 7877 830 7880 839
rect 7928 835 7939 839
rect 7928 831 7933 835
rect 7841 824 7844 830
rect 7880 828 7881 830
rect 7926 828 7928 831
rect 7937 828 7939 835
rect 7832 816 7848 824
rect 7776 813 7779 815
rect 7728 808 7771 810
rect 7786 808 7790 816
rect 7809 812 7811 816
rect 7720 807 7731 808
rect 7745 807 7747 808
rect 7771 807 7790 808
rect 7624 799 7646 805
rect 7624 798 7640 799
rect 7620 792 7640 798
rect 7646 793 7652 799
rect 7620 789 7627 792
rect 7631 789 7640 792
rect 7674 792 7690 807
rect 7698 799 7704 805
rect 7692 793 7698 799
rect 7674 790 7675 792
rect 7579 780 7594 789
rect 7624 788 7640 789
rect 7528 774 7594 780
rect 7619 778 7640 788
rect 7669 787 7671 790
rect 7674 787 7690 790
rect 7663 778 7665 787
rect 7619 776 7665 778
rect 7669 776 7690 787
rect 7707 785 7728 807
rect 7748 803 7749 805
rect 7761 799 7767 804
rect 7750 795 7751 797
rect 7771 795 7786 807
rect 7806 806 7809 812
rect 7832 811 7853 816
rect 7881 813 7886 828
rect 7919 817 7926 828
rect 7932 818 7933 828
rect 7919 816 7932 817
rect 7916 815 7919 816
rect 7901 814 7913 815
rect 7899 813 7901 814
rect 7877 812 7891 813
rect 7865 811 7877 812
rect 7832 810 7865 811
rect 7832 808 7853 810
rect 7881 808 7886 812
rect 7790 801 7792 805
rect 7797 795 7806 806
rect 7741 787 7757 795
rect 7771 792 7797 795
rect 7816 792 7832 808
rect 7848 806 7853 808
rect 7925 806 7932 816
rect 7937 809 7938 828
rect 7937 806 7940 809
rect 7969 807 7971 839
rect 8104 836 8106 841
rect 8134 836 8135 841
rect 8164 839 8188 841
rect 7925 805 7933 806
rect 7961 805 7971 807
rect 7975 805 7983 817
rect 8024 815 8040 824
rect 8042 815 8058 824
rect 8024 814 8058 815
rect 8106 814 8108 836
rect 8135 824 8141 836
rect 8166 830 8180 839
rect 8248 836 8250 842
rect 8273 841 8277 854
rect 8272 836 8277 841
rect 8265 834 8277 836
rect 8289 860 8317 861
rect 8289 855 8316 860
rect 8180 828 8188 830
rect 8181 825 8184 828
rect 8024 813 8059 814
rect 8022 811 8024 813
rect 8057 812 8058 813
rect 8022 808 8058 811
rect 8120 809 8154 824
rect 8184 815 8188 825
rect 8188 811 8189 814
rect 8189 809 8190 811
rect 8250 809 8251 811
rect 8117 808 8154 809
rect 8190 808 8191 809
rect 7853 801 7855 805
rect 7886 800 7888 805
rect 7933 802 7937 805
rect 7937 801 7961 802
rect 7969 801 7971 805
rect 8008 801 8034 808
rect 8044 801 8056 808
rect 7888 797 7889 800
rect 7857 795 7858 797
rect 7785 790 7797 792
rect 7858 791 7861 795
rect 7624 774 7635 776
rect 7670 774 7690 776
rect 7352 766 7417 772
rect 7429 768 7439 774
rect 7441 771 7475 774
rect 7478 771 7482 774
rect 7441 768 7482 771
rect 7352 758 7411 766
rect 7437 764 7439 768
rect 7448 764 7464 768
rect 7292 753 7295 756
rect 7298 753 7301 754
rect 7246 744 7301 753
rect 7359 749 7411 758
rect 7441 758 7464 764
rect 7466 758 7482 768
rect 7544 761 7560 774
rect 7441 756 7453 758
rect 7458 755 7464 758
rect 7516 755 7522 761
rect 7541 758 7560 761
rect 7562 758 7578 774
rect 7640 772 7656 774
rect 7658 772 7674 774
rect 7593 761 7599 767
rect 7631 764 7674 772
rect 7704 768 7708 785
rect 7741 780 7758 787
rect 7728 768 7734 773
rect 7754 772 7758 780
rect 7771 780 7801 790
rect 7771 774 7786 780
rect 7797 779 7801 780
rect 7780 773 7785 774
rect 7758 771 7759 772
rect 7541 755 7547 758
rect 7599 755 7605 761
rect 7640 758 7656 764
rect 7658 758 7674 764
rect 7464 749 7470 755
rect 7510 749 7516 755
rect 7543 754 7547 755
rect 7702 754 7708 768
rect 7750 767 7771 771
rect 7775 767 7780 773
rect 7716 757 7718 758
rect 7715 755 7716 757
rect 7540 750 7544 754
rect 7711 752 7715 755
rect 7750 753 7775 767
rect 7801 763 7812 779
rect 7816 774 7832 790
rect 7861 779 7866 790
rect 7866 776 7874 779
rect 7889 778 7905 797
rect 7937 793 7949 801
rect 7959 793 7971 801
rect 8002 797 8024 801
rect 8048 797 8054 801
rect 8002 795 8056 797
rect 8058 795 8074 808
rect 8104 795 8117 808
rect 8135 806 8141 808
rect 8141 802 8142 806
rect 7967 778 7971 793
rect 7996 789 8024 795
rect 7889 776 7927 778
rect 7866 775 7905 776
rect 7866 774 7882 775
rect 7812 754 7818 763
rect 7832 758 7848 774
rect 7850 763 7874 774
rect 7889 764 7905 775
rect 7912 775 7927 776
rect 7912 774 7928 775
rect 7928 763 7930 774
rect 7967 763 7969 778
rect 7850 758 7866 763
rect 7874 753 7879 763
rect 7905 754 7910 763
rect 7928 758 7933 763
rect 7968 761 7969 763
rect 8002 774 8024 789
rect 8054 792 8074 795
rect 8054 790 8068 792
rect 8054 789 8074 790
rect 8054 781 8056 789
rect 8055 774 8056 781
rect 8058 774 8074 789
rect 8097 784 8107 795
rect 8109 787 8110 795
rect 8142 786 8145 800
rect 8154 792 8170 808
rect 8095 780 8097 784
rect 8110 782 8111 786
rect 8145 781 8146 786
rect 8093 774 8095 780
rect 8146 778 8147 781
rect 8147 774 8149 778
rect 8154 774 8170 790
rect 8191 786 8199 808
rect 8265 806 8272 834
rect 8289 826 8310 855
rect 8264 802 8265 806
rect 8277 803 8286 812
rect 8289 808 8300 826
rect 8326 824 8336 847
rect 8312 818 8346 824
rect 8808 819 8809 1015
rect 8998 819 8999 1015
rect 9084 819 9085 1015
rect 9357 819 9358 1015
rect 9554 819 9555 1015
rect 10152 1012 10153 1015
rect 10211 1013 10212 1016
rect 10208 1012 10212 1013
rect 10452 1014 10468 1016
rect 10496 1015 10508 1016
rect 10470 1014 10492 1015
rect 10504 1014 10508 1015
rect 10452 1012 10513 1014
rect 10544 1012 10764 1021
rect 10935 1017 10946 1021
rect 10935 1014 10953 1017
rect 10956 1014 11021 1030
rect 10935 1012 11021 1014
rect 10142 1005 10148 1011
rect 10151 1008 10152 1012
rect 10150 1005 10151 1008
rect 10188 1005 10194 1011
rect 10136 999 10142 1005
rect 10194 999 10200 1005
rect 10162 990 10163 997
rect 10201 995 10202 1012
rect 10207 1001 10214 1012
rect 10452 1011 10510 1012
rect 10443 1008 10449 1011
rect 10450 1009 10452 1011
rect 10454 1010 10459 1011
rect 10453 1009 10459 1010
rect 10513 1009 10514 1011
rect 10535 1010 10543 1012
rect 10941 1011 10950 1012
rect 10935 1010 10948 1011
rect 10956 1010 11021 1012
rect 10450 1008 10457 1009
rect 10515 1008 10535 1010
rect 10443 1006 10451 1008
rect 10436 1005 10451 1006
rect 10453 1005 10457 1008
rect 10433 1001 10451 1005
rect 10505 1001 10508 1008
rect 10207 998 10208 1001
rect 10206 997 10207 998
rect 10200 990 10202 994
rect 10203 990 10207 997
rect 10415 994 10433 1001
rect 10436 997 10451 1001
rect 10162 989 10179 990
rect 10163 988 10179 989
rect 10148 978 10179 988
rect 10183 978 10214 990
rect 10393 986 10415 994
rect 10436 990 10452 997
rect 10506 996 10507 1000
rect 10511 998 10535 1008
rect 10935 1009 10947 1010
rect 10948 1009 11021 1010
rect 11037 1009 11118 1030
rect 13549 1027 13587 1038
rect 14017 1030 14023 1036
rect 11849 1015 11850 1026
rect 12039 1015 12040 1026
rect 12125 1015 12126 1026
rect 12398 1015 12399 1026
rect 12595 1015 12596 1026
rect 13216 1025 13255 1026
rect 13216 1024 13253 1025
rect 13255 1024 13256 1025
rect 13214 1022 13216 1024
rect 13242 1016 13254 1024
rect 13256 1022 13257 1024
rect 13516 1022 13549 1027
rect 13921 1025 13977 1027
rect 13257 1016 13263 1022
rect 13504 1020 13549 1022
rect 13816 1021 13921 1025
rect 13977 1021 13987 1025
rect 13504 1016 13560 1020
rect 13205 1015 13257 1016
rect 10935 1005 10956 1009
rect 10511 996 10520 998
rect 10506 995 10508 996
rect 10511 995 10515 996
rect 10451 988 10452 990
rect 10374 979 10393 986
rect 10148 972 10214 978
rect 10360 974 10374 979
rect 10109 967 10115 968
rect 9870 965 9872 967
rect 9925 964 9926 967
rect 10102 964 10106 967
rect 10115 964 10122 967
rect 9926 962 9928 964
rect 10089 956 10102 964
rect 10122 963 10127 964
rect 10127 959 10138 963
rect 10164 961 10180 972
rect 10182 966 10202 972
rect 10352 971 10358 973
rect 10436 972 10452 988
rect 10496 992 10511 995
rect 10517 993 10519 996
rect 10496 986 10512 992
rect 10518 988 10519 993
rect 10517 986 10518 988
rect 10661 986 10682 1002
rect 10928 1001 10935 1005
rect 10941 1001 10956 1005
rect 10914 994 10928 1001
rect 10948 998 10956 1001
rect 10974 1005 10984 1009
rect 11118 1005 11135 1009
rect 10974 1003 10987 1005
rect 10956 995 10957 998
rect 10496 985 10520 986
rect 10875 985 10881 991
rect 10899 986 10914 994
rect 10897 985 10899 986
rect 10921 985 10927 991
rect 10957 985 10964 995
rect 10495 983 10496 985
rect 10500 974 10520 985
rect 10695 974 10707 982
rect 10717 974 10729 982
rect 10869 979 10875 985
rect 10927 979 10933 985
rect 10959 980 10967 985
rect 10959 979 10968 980
rect 10959 978 10969 979
rect 10959 975 10971 978
rect 10347 970 10352 971
rect 10344 969 10347 970
rect 10452 968 10470 971
rect 10500 970 10512 974
rect 10959 973 10973 975
rect 10974 973 10975 1003
rect 10980 993 11001 1003
rect 11135 999 11157 1005
rect 11157 997 11159 999
rect 10984 983 11001 993
rect 11159 992 11165 997
rect 11165 986 11169 992
rect 10959 971 10975 973
rect 10980 972 11001 983
rect 11169 982 11172 986
rect 11172 975 11176 982
rect 11176 973 11177 975
rect 10980 971 11102 972
rect 11177 971 11178 972
rect 10689 970 10691 971
rect 10731 970 10768 971
rect 10500 969 10509 970
rect 10244 967 10248 968
rect 10250 967 10255 968
rect 10182 961 10198 966
rect 10236 965 10244 967
rect 10234 964 10236 965
rect 10255 964 10258 967
rect 10336 966 10343 968
rect 10332 964 10336 966
rect 10231 963 10234 964
rect 10230 962 10231 963
rect 10258 962 10261 964
rect 10328 963 10332 964
rect 10150 959 10198 961
rect 10127 958 10142 959
rect 10150 958 10200 959
rect 10223 958 10232 962
rect 10261 959 10265 962
rect 10308 961 10328 963
rect 10130 956 10144 958
rect 10145 957 10200 958
rect 10086 954 10089 956
rect 10130 954 10147 956
rect 10150 954 10200 957
rect 10219 956 10232 958
rect 10265 956 10268 959
rect 10316 958 10322 961
rect 10215 954 10232 956
rect 10268 954 10271 956
rect 10305 954 10313 957
rect 10437 956 10443 959
rect 10452 956 10468 968
rect 10470 967 10477 968
rect 10500 967 10508 969
rect 10477 965 10488 967
rect 10496 966 10508 967
rect 10495 965 10508 966
rect 10488 964 10508 965
rect 10528 964 10534 970
rect 10574 966 10580 970
rect 10683 969 10689 970
rect 10564 964 10580 966
rect 10496 962 10508 964
rect 10415 954 10443 956
rect 9926 946 9927 949
rect 9925 945 9964 946
rect 9923 944 9925 945
rect 9908 934 9923 944
rect 9884 920 9908 934
rect 9881 918 9884 920
rect 9874 913 9881 918
rect 9926 913 9927 945
rect 9964 944 9991 945
rect 10068 944 10086 954
rect 10130 953 10200 954
rect 10130 951 10152 953
rect 10181 951 10182 953
rect 10188 951 10194 953
rect 10208 951 10232 954
rect 10130 948 10232 951
rect 10130 947 10185 948
rect 10188 947 10194 948
rect 10130 946 10164 947
rect 10166 946 10185 947
rect 10197 946 10232 948
rect 10130 944 10185 946
rect 10195 945 10232 946
rect 10194 944 10232 945
rect 10271 953 10294 954
rect 10302 953 10305 954
rect 10415 953 10433 954
rect 10437 953 10463 954
rect 10495 953 10501 959
rect 10522 958 10586 964
rect 10633 963 10639 969
rect 10679 968 10685 969
rect 10674 966 10685 968
rect 10668 964 10673 966
rect 10664 963 10668 964
rect 10679 963 10685 966
rect 10695 968 10729 970
rect 10733 969 10741 970
rect 10528 954 10580 958
rect 10627 957 10633 963
rect 10685 957 10691 963
rect 10271 946 10302 953
rect 10388 946 10427 953
rect 10443 947 10449 953
rect 10489 947 10495 953
rect 10271 944 10294 946
rect 10382 945 10388 946
rect 10377 944 10382 945
rect 9991 938 10232 944
rect 10261 938 10276 944
rect 10284 939 10294 944
rect 10290 938 10294 939
rect 10343 938 10377 944
rect 10528 938 10542 954
rect 10052 922 10068 938
rect 10114 937 10137 938
rect 10114 934 10142 937
rect 10114 933 10150 934
rect 10152 933 10160 935
rect 10181 934 10182 938
rect 10256 937 10261 938
rect 10247 935 10255 936
rect 10183 934 10230 935
rect 10242 934 10247 935
rect 10167 933 10230 934
rect 10294 933 10310 938
rect 10337 936 10343 938
rect 10528 936 10543 938
rect 10333 935 10336 936
rect 10328 933 10332 934
rect 10114 925 10222 933
rect 10181 924 10182 925
rect 10120 922 10137 924
rect 10052 916 10068 920
rect 10103 917 10118 922
rect 10141 920 10166 922
rect 9954 913 9995 916
rect 9999 913 10068 916
rect 9871 911 9874 913
rect 9926 911 9954 913
rect 10052 911 10096 913
rect 10102 911 10118 917
rect 10139 917 10166 920
rect 10185 918 10244 922
rect 10292 920 10328 933
rect 10526 931 10543 936
rect 10522 928 10526 931
rect 10515 924 10522 928
rect 10507 920 10515 924
rect 10528 920 10543 931
rect 10574 920 10576 954
rect 10580 950 10593 954
rect 10695 953 10716 968
rect 10726 967 10729 968
rect 10734 963 10741 969
rect 10769 968 10772 970
rect 10959 969 10973 971
rect 10974 970 11102 971
rect 10984 969 11001 970
rect 11005 969 11102 970
rect 10772 967 10774 968
rect 10774 966 10776 967
rect 10737 960 10739 963
rect 10955 960 10958 961
rect 10742 954 10749 957
rect 10874 953 10875 957
rect 10936 954 10955 960
rect 10959 957 10978 969
rect 10936 953 10960 954
rect 10694 952 10716 953
rect 10694 950 10695 952
rect 10580 942 10588 950
rect 10693 938 10694 949
rect 10750 946 10762 953
rect 10933 952 10936 953
rect 10763 944 10765 945
rect 10765 940 10772 944
rect 10580 920 10588 932
rect 10287 918 10292 920
rect 10167 917 10244 918
rect 10139 915 10151 917
rect 10211 916 10222 917
rect 10159 914 10171 916
rect 10210 915 10212 916
rect 9867 909 9871 911
rect 9925 910 9927 911
rect 9924 909 9928 910
rect 9923 906 9928 909
rect 9870 903 9871 904
rect 9922 903 9928 906
rect 10052 904 10068 911
rect 10096 910 10121 911
rect 10087 908 10118 910
rect 10121 909 10132 910
rect 10132 908 10139 909
rect 10077 906 10118 908
rect 10139 907 10152 908
rect 10160 906 10167 907
rect 10087 905 10118 906
rect 10102 904 10118 905
rect 9861 894 9862 899
rect 9915 896 9916 900
rect 9921 899 9928 903
rect 9920 895 9921 899
rect 9914 876 9916 895
rect 10068 888 10084 904
rect 10086 888 10102 904
rect 10179 888 10181 911
rect 10244 909 10260 917
rect 10276 913 10287 918
rect 10271 911 10275 913
rect 10265 909 10271 911
rect 10294 909 10310 920
rect 10494 912 10507 920
rect 10526 918 10580 920
rect 10591 918 10593 926
rect 10630 920 10633 937
rect 10772 935 10781 940
rect 10868 939 10874 952
rect 10878 946 10899 949
rect 10915 946 10916 949
rect 10927 948 10933 952
rect 10944 946 10960 953
rect 10868 936 10875 939
rect 10876 938 10878 946
rect 10899 939 10960 946
rect 10973 942 10978 957
rect 11001 968 11102 969
rect 11179 968 11180 970
rect 10907 938 10960 939
rect 10926 937 10976 938
rect 10693 925 10696 929
rect 10782 928 10792 934
rect 10868 933 10876 936
rect 10926 933 10933 937
rect 10522 912 10592 918
rect 10627 917 10629 919
rect 10696 918 10711 925
rect 10792 923 10796 928
rect 10796 920 10797 923
rect 10711 917 10734 918
rect 10627 916 10633 917
rect 10625 912 10633 916
rect 10492 911 10494 912
rect 10526 911 10541 912
rect 10542 911 10543 912
rect 10244 908 10310 909
rect 10230 907 10310 908
rect 10486 907 10492 911
rect 10526 907 10547 911
rect 10564 908 10580 912
rect 10188 906 10211 907
rect 10244 904 10310 907
rect 10278 888 10294 904
rect 10472 900 10486 907
rect 10526 904 10541 907
rect 10542 904 10543 907
rect 10574 906 10580 908
rect 10583 904 10592 912
rect 10627 911 10633 912
rect 10685 916 10734 917
rect 10685 911 10691 916
rect 10702 914 10734 916
rect 10711 913 10735 914
rect 10711 911 10734 913
rect 10737 911 10762 913
rect 10776 911 10790 920
rect 10797 918 10798 920
rect 10863 918 10868 933
rect 10874 927 10881 933
rect 10874 925 10876 927
rect 10798 913 10800 918
rect 10800 911 10801 913
rect 10861 911 10863 915
rect 10622 907 10624 911
rect 10527 900 10540 904
rect 10581 900 10583 903
rect 10618 900 10622 907
rect 10633 905 10639 911
rect 10452 888 10475 900
rect 10522 897 10527 900
rect 10506 888 10522 897
rect 10539 896 10542 899
rect 10576 896 10581 899
rect 10616 897 10618 900
rect 10542 888 10558 896
rect 10560 888 10576 896
rect 10610 888 10616 897
rect 9920 875 9928 888
rect 10116 880 10246 888
rect 10449 883 10452 888
rect 10498 883 10506 888
rect 10607 883 10610 888
rect 10364 880 10412 883
rect 10094 875 10136 880
rect 9914 873 9920 875
rect 10083 873 10136 875
rect 9871 870 9875 873
rect 9904 871 9914 873
rect 9917 872 9920 873
rect 9904 870 9916 871
rect 10064 870 10136 873
rect 10179 870 10181 880
rect 10223 879 10364 880
rect 10226 875 10364 879
rect 10412 875 10413 880
rect 10445 875 10449 883
rect 10484 876 10498 883
rect 10602 876 10607 883
rect 10478 875 10484 876
rect 10645 875 10669 910
rect 10679 905 10685 911
rect 10711 909 10790 911
rect 10801 909 10802 911
rect 10724 904 10790 909
rect 10802 904 10804 908
rect 10740 888 10756 904
rect 10758 893 10774 904
rect 10804 899 10806 903
rect 10806 893 10808 899
rect 10849 898 10861 910
rect 10870 909 10874 925
rect 10907 916 10915 933
rect 10921 927 10927 933
rect 10869 904 10870 909
rect 10887 905 10907 915
rect 10874 903 10886 905
rect 10887 903 10908 905
rect 10926 904 10927 927
rect 10960 922 10976 937
rect 10978 936 10979 941
rect 11001 938 11022 968
rect 11042 967 11102 968
rect 11180 967 11181 968
rect 11051 965 11102 967
rect 11181 965 11184 967
rect 11071 963 11102 965
rect 11184 963 11186 965
rect 11080 961 11102 963
rect 11186 961 11190 963
rect 11034 938 11050 954
rect 11052 938 11068 954
rect 11092 949 11120 961
rect 11190 954 11199 961
rect 11078 938 11079 949
rect 11120 947 11124 949
rect 11199 947 11207 954
rect 11124 946 11125 947
rect 11125 944 11126 946
rect 11207 944 11209 947
rect 11395 944 11396 949
rect 11424 944 11440 954
rect 11126 939 11132 944
rect 11209 940 11214 944
rect 11378 940 11445 944
rect 11214 939 11216 940
rect 11355 939 11378 940
rect 11001 936 11034 938
rect 11068 937 11084 938
rect 11048 936 11084 937
rect 11132 936 11134 938
rect 11216 936 11219 939
rect 11352 936 11355 939
rect 11395 938 11396 940
rect 11445 938 11446 939
rect 10979 916 10984 933
rect 11001 922 11033 936
rect 11048 935 11068 936
rect 11070 934 11084 936
rect 11134 934 11136 936
rect 11219 934 11223 936
rect 11349 934 11352 936
rect 11064 932 11084 934
rect 11136 932 11137 934
rect 11223 932 11225 934
rect 11348 932 11349 934
rect 10985 915 10991 921
rect 11001 919 11022 922
rect 11026 921 11033 922
rect 11022 915 11025 919
rect 11026 915 11037 921
rect 10979 909 10985 915
rect 10984 908 10985 909
rect 11026 906 11033 915
rect 11037 909 11043 915
rect 11075 904 11111 932
rect 11137 925 11144 932
rect 11225 925 11236 932
rect 11345 925 11348 932
rect 11144 924 11158 925
rect 11136 915 11158 924
rect 11236 919 11245 925
rect 11342 919 11345 925
rect 11245 916 11248 919
rect 11341 916 11342 919
rect 11144 907 11158 915
rect 11248 912 11253 916
rect 11339 912 11341 916
rect 11253 907 11257 912
rect 11336 910 11339 912
rect 11152 905 11161 907
rect 11158 904 11161 905
rect 11257 904 11259 907
rect 11083 903 11086 904
rect 11111 903 11112 904
rect 11161 903 11162 904
rect 10871 901 10911 903
rect 10868 900 10869 901
rect 10867 899 10868 900
rect 10871 899 10907 901
rect 10911 899 10912 901
rect 10866 898 10871 899
rect 10849 896 10871 898
rect 10809 893 10861 896
rect 10866 893 10871 896
rect 10758 888 10777 893
rect 10808 888 10861 893
rect 10705 877 10714 881
rect 10752 877 10761 881
rect 10771 879 10777 888
rect 10803 886 10815 888
rect 10798 883 10803 886
rect 10808 883 10815 886
rect 10797 882 10815 883
rect 10789 880 10815 882
rect 10786 879 10815 880
rect 10771 877 10815 879
rect 10697 875 10815 877
rect 10226 870 10328 875
rect 10366 874 10520 875
rect 10366 872 10513 874
rect 10339 871 10366 872
rect 10445 871 10449 872
rect 10478 871 10484 872
rect 10520 871 10534 874
rect 10600 871 10602 875
rect 10639 872 10697 875
rect 10705 872 10808 875
rect 10331 870 10339 871
rect 10534 870 10538 871
rect 10639 870 10705 872
rect 10706 870 10808 872
rect 10815 870 10817 875
rect 10849 872 10861 888
rect 10862 881 10867 893
rect 10866 880 10867 881
rect 10887 871 10907 899
rect 10912 893 10915 899
rect 10915 881 10920 893
rect 11023 887 11026 903
rect 11079 902 11083 903
rect 11078 899 11079 901
rect 11112 899 11118 903
rect 11071 893 11078 899
rect 11083 897 11084 899
rect 11117 893 11118 899
rect 11153 893 11160 898
rect 11162 893 11176 903
rect 11071 887 11077 893
rect 10915 877 10919 881
rect 11026 877 11051 887
rect 11160 885 11172 893
rect 11176 887 11185 893
rect 11259 887 11272 903
rect 11332 902 11344 910
rect 11354 902 11366 910
rect 11406 904 11407 938
rect 11445 934 11456 938
rect 11446 922 11456 934
rect 11446 903 11447 922
rect 11332 898 11335 902
rect 11368 899 11370 902
rect 11320 886 11328 898
rect 11332 896 11366 898
rect 11332 895 11335 896
rect 10919 873 10920 875
rect 11051 870 11069 877
rect 11071 875 11077 877
rect 11172 876 11179 885
rect 11185 879 11191 886
rect 11272 879 11277 886
rect 11191 877 11193 879
rect 11277 877 11279 879
rect 11071 870 11078 875
rect 11083 870 11084 872
rect 11193 871 11196 877
rect 11279 870 11283 877
rect 9875 869 9904 870
rect 9912 867 9916 870
rect 10060 869 10064 870
rect 10326 869 10331 870
rect 10414 869 10415 870
rect 9911 866 9916 867
rect 10047 866 10060 869
rect 10317 868 10326 869
rect 10309 866 10317 868
rect 10415 867 10416 869
rect 9859 859 9860 866
rect 9909 864 9916 866
rect 10025 865 10059 866
rect 10304 865 10309 866
rect 9909 859 9911 864
rect 10025 862 10047 865
rect 10024 859 10047 862
rect 10059 859 10066 865
rect 10271 859 10304 865
rect 9908 855 9909 859
rect 10020 855 10025 859
rect 10028 854 10047 859
rect 10066 857 10069 859
rect 10265 858 10271 859
rect 10258 857 10265 858
rect 10242 854 10257 857
rect 10416 854 10421 866
rect 10443 863 10445 870
rect 10475 863 10478 870
rect 10538 868 10550 870
rect 10442 860 10443 863
rect 10474 860 10475 863
rect 10550 859 10588 868
rect 10593 863 10598 870
rect 10628 869 10639 870
rect 10616 868 10628 869
rect 10614 866 10616 868
rect 10611 864 10614 866
rect 10641 864 10644 869
rect 10591 860 10593 863
rect 9907 851 9908 854
rect 10018 851 10020 854
rect 10027 850 10028 854
rect 9858 838 9859 850
rect 9903 838 9907 850
rect 10011 838 10018 850
rect 8312 812 8328 818
rect 8330 812 8346 818
rect 9857 816 9858 837
rect 9896 816 9903 838
rect 10011 835 10017 838
rect 10005 829 10011 835
rect 10019 828 10024 842
rect 10057 835 10063 841
rect 10069 839 10070 854
rect 10146 850 10242 854
rect 10421 850 10422 854
rect 10440 853 10442 859
rect 10471 853 10474 859
rect 10583 858 10593 859
rect 10583 853 10590 858
rect 10593 857 10599 858
rect 10608 857 10611 864
rect 10696 863 10705 870
rect 10761 863 10770 870
rect 10779 868 10780 870
rect 10817 868 10818 870
rect 10639 860 10641 863
rect 10780 861 10782 868
rect 10818 860 10821 868
rect 10847 864 10848 866
rect 10846 861 10847 863
rect 10862 859 10868 870
rect 10884 864 10887 870
rect 10920 866 10922 870
rect 11069 869 11079 870
rect 10959 868 10960 869
rect 10958 867 10959 868
rect 10957 865 10958 866
rect 10950 864 10957 865
rect 10874 859 10876 861
rect 10599 855 10622 857
rect 10637 856 10639 859
rect 10599 854 10612 855
rect 10632 854 10637 856
rect 10583 852 10586 853
rect 10583 851 10585 852
rect 10607 851 10608 854
rect 10612 851 10653 854
rect 10698 851 10704 857
rect 10744 851 10750 857
rect 10783 855 10784 857
rect 10822 854 10823 857
rect 10844 856 10845 859
rect 10870 856 10878 859
rect 10831 854 10870 856
rect 10880 855 10884 863
rect 10908 859 10950 864
rect 10979 863 10985 869
rect 11037 863 11043 869
rect 11071 867 11079 869
rect 11179 868 11180 870
rect 11196 869 11197 870
rect 11080 867 11089 868
rect 11071 866 11092 867
rect 11071 865 11079 866
rect 11080 865 11092 866
rect 11152 865 11154 868
rect 11197 867 11198 869
rect 11283 867 11285 869
rect 11332 868 11334 895
rect 11198 865 11199 866
rect 11080 863 11089 865
rect 10879 854 10880 855
rect 10754 851 10831 854
rect 10843 853 10844 854
rect 10872 853 10885 854
rect 10086 843 10147 850
rect 10085 841 10086 842
rect 10063 832 10069 835
rect 10070 832 10071 838
rect 10063 829 10071 832
rect 10079 829 10085 841
rect 10089 840 10100 842
rect 10146 840 10147 843
rect 10157 843 10347 850
rect 10422 846 10425 850
rect 10432 846 10440 851
rect 10463 847 10471 851
rect 10458 846 10519 847
rect 10369 843 10451 846
rect 10157 839 10242 843
rect 10335 842 10353 843
rect 10422 842 10425 843
rect 10317 839 10335 842
rect 10353 841 10365 842
rect 10368 839 10371 841
rect 10155 838 10157 839
rect 10150 835 10154 838
rect 10144 830 10150 835
rect 10177 831 10179 839
rect 10309 838 10317 839
rect 10293 835 10309 838
rect 10067 828 10071 829
rect 10143 828 10144 830
rect 8312 809 8346 812
rect 9856 810 9857 816
rect 9895 811 9896 816
rect 9924 811 9940 824
rect 10018 813 10019 828
rect 10063 826 10065 827
rect 10067 826 10079 828
rect 10065 816 10087 826
rect 10116 817 10132 824
rect 10063 812 10087 816
rect 10106 812 10132 817
rect 10063 811 10065 812
rect 8312 808 8358 809
rect 8261 790 8264 800
rect 8268 794 8277 803
rect 8289 792 8312 808
rect 8324 803 8333 808
rect 8358 805 8363 808
rect 9893 807 9895 810
rect 10069 808 10071 811
rect 8333 794 8342 803
rect 8251 787 8266 790
rect 8199 779 8205 786
rect 8224 780 8266 787
rect 8272 786 8276 792
rect 8289 790 8299 792
rect 8289 787 8312 790
rect 8268 780 8270 784
rect 8289 781 8326 787
rect 8200 774 8216 779
rect 8224 774 8268 780
rect 8296 774 8326 781
rect 8363 774 8379 805
rect 9855 800 9856 805
rect 9890 800 9892 805
rect 9889 798 9890 800
rect 9885 790 9889 798
rect 9908 792 9919 808
rect 10068 806 10069 808
rect 10087 807 10096 812
rect 10104 809 10132 812
rect 10102 808 10113 809
rect 10116 808 10132 809
rect 10134 808 10150 824
rect 10173 818 10179 831
rect 10259 830 10293 835
rect 10217 823 10259 830
rect 10371 829 10373 839
rect 10425 829 10430 842
rect 10432 828 10440 843
rect 10209 822 10217 823
rect 10184 818 10209 822
rect 10173 816 10184 818
rect 10169 812 10179 816
rect 10100 807 10116 808
rect 10096 806 10116 807
rect 10096 805 10113 806
rect 10150 805 10166 808
rect 10018 790 10019 805
rect 9883 786 9885 790
rect 10004 787 10019 790
rect 10057 789 10068 805
rect 10094 803 10127 805
rect 10094 794 10122 803
rect 10144 797 10166 805
rect 10094 793 10116 794
rect 10100 792 10116 793
rect 10106 790 10116 792
rect 10140 792 10166 797
rect 10140 791 10150 792
rect 10057 787 10069 789
rect 9854 782 9855 786
rect 10004 783 10069 787
rect 10100 787 10116 790
rect 10133 790 10150 791
rect 10133 787 10166 790
rect 10100 783 10166 787
rect 10004 782 10068 783
rect 8002 761 8058 774
rect 8060 763 8068 774
rect 8090 763 8093 774
rect 8111 764 8112 770
rect 7930 753 7933 758
rect 7969 758 8058 761
rect 8089 760 8092 763
rect 8143 760 8154 774
rect 7359 745 7418 749
rect 7540 746 7547 750
rect 7701 748 7711 752
rect 7748 749 7750 753
rect 7579 746 7676 748
rect 7699 746 7711 748
rect 7747 746 7748 748
rect 7539 745 7547 746
rect 7550 745 7685 746
rect 7696 745 7698 746
rect 7701 745 7711 746
rect 7246 741 7298 744
rect 7301 742 7302 744
rect 7240 736 7304 741
rect 7359 740 7498 745
rect 7539 744 7711 745
rect 7240 735 7306 736
rect 7161 730 7167 731
rect 7082 727 7184 730
rect 7082 724 7209 727
rect 7218 725 7225 731
rect 7246 729 7252 735
rect 7261 727 7264 732
rect 7292 729 7298 735
rect 7303 727 7306 735
rect 7265 725 7266 727
rect 7306 725 7307 727
rect 7359 726 7367 740
rect 7411 736 7498 740
rect 7413 730 7498 736
rect 7531 743 7711 744
rect 7743 743 7747 745
rect 7757 744 7775 753
rect 7879 750 7881 753
rect 7910 750 7912 753
rect 7780 744 7820 745
rect 7821 744 7832 750
rect 7531 740 7708 743
rect 7531 732 7545 740
rect 7743 735 7757 743
rect 7420 729 7421 730
rect 7421 727 7422 729
rect 5246 709 5247 712
rect 5206 707 5218 708
rect 5247 702 5248 703
rect 5206 698 5207 701
rect 5268 696 5285 714
rect 6798 713 6799 724
rect 6837 717 6838 724
rect 7082 720 7131 724
rect 7082 717 7138 720
rect 7167 719 7173 724
rect 7082 716 7090 717
rect 7082 715 7089 716
rect 5342 711 5345 713
rect 6838 711 6839 713
rect 7101 712 7103 717
rect 5335 710 5342 711
rect 7131 710 7138 717
rect 5329 708 5341 710
rect 5318 703 5341 708
rect 6797 707 6798 710
rect 6982 707 7065 710
rect 5318 696 5329 703
rect 7103 696 7106 709
rect 7138 708 7148 709
rect 7116 700 7128 708
rect 7138 700 7150 708
rect 7107 698 7112 700
rect 7114 698 7159 700
rect 7107 697 7159 698
rect 7185 697 7187 722
rect 7213 719 7219 725
rect 7266 723 7267 725
rect 7307 720 7308 722
rect 7353 720 7369 726
rect 7269 715 7271 719
rect 7308 716 7309 719
rect 7355 716 7369 720
rect 7373 716 7376 719
rect 7399 718 7401 726
rect 7411 720 7417 726
rect 7498 725 7507 730
rect 7423 723 7424 725
rect 7398 716 7401 718
rect 7405 716 7413 720
rect 7271 709 7275 715
rect 7309 710 7311 715
rect 7355 714 7365 716
rect 7355 713 7364 714
rect 7367 713 7388 716
rect 7398 713 7400 716
rect 7403 713 7413 716
rect 7364 710 7365 713
rect 7376 710 7379 713
rect 7392 712 7396 713
rect 7396 711 7401 712
rect 7403 711 7405 713
rect 7388 710 7403 711
rect 7424 710 7431 722
rect 7507 713 7512 724
rect 7539 722 7545 732
rect 7668 723 7674 729
rect 7684 727 7690 732
rect 7679 723 7684 727
rect 7714 723 7720 729
rect 7740 727 7743 735
rect 7744 727 7757 735
rect 7740 725 7744 727
rect 7765 726 7773 744
rect 7780 740 7832 744
rect 7778 735 7814 740
rect 7820 737 7832 740
rect 7881 747 7884 750
rect 7820 735 7837 737
rect 7778 731 7780 735
rect 7821 734 7837 735
rect 7881 734 7886 747
rect 7831 731 7837 734
rect 7832 730 7837 731
rect 7835 729 7839 730
rect 7884 729 7886 734
rect 7837 726 7841 729
rect 7531 719 7545 722
rect 7531 716 7547 719
rect 7599 716 7600 719
rect 7662 717 7668 723
rect 7720 717 7726 723
rect 7736 722 7740 724
rect 7741 723 7744 725
rect 7767 724 7768 726
rect 7839 725 7841 726
rect 7885 725 7886 729
rect 7773 724 7774 725
rect 7276 698 7282 708
rect 7312 698 7314 708
rect 7367 701 7379 710
rect 7380 698 7386 708
rect 7389 701 7401 710
rect 7403 709 7468 710
rect 7410 707 7468 709
rect 7417 706 7468 707
rect 7425 703 7468 706
rect 7431 700 7437 703
rect 7439 702 7468 703
rect 7440 701 7468 702
rect 7431 698 7445 700
rect 7282 697 7286 698
rect 7107 696 7286 697
rect 5248 695 5249 696
rect 5262 694 5280 696
rect 5030 690 5041 691
rect 5030 688 5039 690
rect 5030 687 5040 688
rect 5043 687 5044 690
rect 5046 688 5055 691
rect 5076 690 5078 691
rect 5183 688 5203 694
rect 5207 691 5208 692
rect 5239 690 5280 694
rect 6796 692 6797 696
rect 7103 695 7112 696
rect 7104 694 7112 695
rect 7116 694 7286 696
rect 7314 694 7318 698
rect 6801 690 6802 692
rect 5208 688 5210 690
rect 5239 688 5262 690
rect 5176 687 5270 688
rect 5027 685 5040 687
rect 5024 683 5027 685
rect 5013 677 5024 683
rect 5030 679 5038 685
rect 4929 667 4931 671
rect 4878 663 4885 667
rect 4833 661 4885 663
rect 4834 660 4893 661
rect 4817 644 4825 645
rect 4792 642 4799 643
rect 4763 637 4765 641
rect 4789 637 4799 642
rect 4808 642 4825 644
rect 4833 642 4834 659
rect 4835 649 4893 660
rect 4926 655 4929 667
rect 4925 652 4926 654
rect 4962 652 4969 672
rect 5009 668 5013 676
rect 5030 663 5038 669
rect 5042 663 5044 687
rect 5208 676 5210 687
rect 5249 682 5251 687
rect 5292 676 5302 680
rect 6799 676 6802 690
rect 5112 672 5132 673
rect 5096 664 5112 672
rect 5132 664 5184 672
rect 5092 663 5096 664
rect 5030 662 5096 663
rect 5184 663 5198 664
rect 5210 663 5212 676
rect 5286 674 5292 676
rect 5255 664 5286 674
rect 6796 670 6799 676
rect 5246 663 5255 664
rect 5184 662 5255 663
rect 4843 648 4885 649
rect 4843 645 4883 648
rect 4789 635 4796 637
rect 4808 635 4834 642
rect 4847 637 4859 645
rect 4869 644 4881 645
rect 4882 644 4883 645
rect 4869 642 4883 644
rect 4922 643 4924 647
rect 4960 645 4962 651
rect 4959 643 4960 645
rect 5007 642 5009 659
rect 5030 657 5091 662
rect 5198 661 5255 662
rect 6789 663 6799 670
rect 6801 663 6802 676
rect 6834 690 6835 692
rect 6836 690 6846 692
rect 6834 687 6861 690
rect 7101 688 7107 694
rect 6834 673 6865 687
rect 7104 684 7107 688
rect 7116 692 7212 694
rect 7116 690 7244 692
rect 7282 691 7341 694
rect 7282 690 7286 691
rect 7314 690 7318 691
rect 7341 690 7345 691
rect 7386 690 7387 696
rect 7437 695 7445 698
rect 7447 697 7468 701
rect 7509 709 7513 713
rect 7531 712 7549 716
rect 7574 712 7577 713
rect 7531 711 7547 712
rect 7531 710 7545 711
rect 7539 709 7547 710
rect 7549 709 7551 711
rect 7552 710 7577 712
rect 7592 710 7594 712
rect 7599 710 7605 715
rect 7653 710 7668 716
rect 7735 715 7740 722
rect 7728 711 7734 714
rect 7736 711 7740 715
rect 7762 716 7779 724
rect 7558 709 7660 710
rect 7509 707 7514 709
rect 7539 707 7545 709
rect 7580 707 7660 709
rect 7509 706 7515 707
rect 7542 706 7580 707
rect 7509 702 7516 706
rect 7509 701 7517 702
rect 7480 698 7490 699
rect 7509 698 7519 701
rect 7542 698 7555 706
rect 7593 703 7599 707
rect 7604 706 7660 707
rect 7728 709 7736 711
rect 7728 706 7734 709
rect 7762 708 7784 716
rect 7776 706 7784 708
rect 7795 706 7801 712
rect 7604 705 7673 706
rect 7720 705 7728 706
rect 7604 703 7728 705
rect 7604 700 7641 703
rect 7473 697 7477 698
rect 7455 695 7473 697
rect 7431 694 7473 695
rect 7491 696 7519 698
rect 7437 692 7468 694
rect 7437 691 7456 692
rect 7434 690 7442 691
rect 7116 688 7165 690
rect 7116 683 7150 688
rect 7116 682 7124 683
rect 7116 681 7123 682
rect 7016 673 7050 676
rect 6834 663 6835 673
rect 6840 663 6847 670
rect 5210 660 5212 661
rect 6789 658 6847 663
rect 6864 660 6865 673
rect 5038 656 5091 657
rect 6795 657 6840 658
rect 5038 655 5080 656
rect 5040 653 5078 655
rect 6795 653 6796 657
rect 6799 654 6837 657
rect 5042 645 5054 653
rect 5064 645 5076 653
rect 6801 646 6813 654
rect 6823 646 6835 654
rect 4869 641 4882 642
rect 4866 639 4882 641
rect 4869 637 4882 639
rect 4871 636 4882 637
rect 4861 635 4867 636
rect 4873 635 4882 636
rect 4426 626 4444 630
rect 4457 626 4494 634
rect 4529 626 4538 635
rect 4576 626 4585 635
rect 4766 630 4773 634
rect 4765 626 4773 630
rect 4426 625 4432 626
rect 4309 621 4324 625
rect 4421 621 4426 625
rect 4309 618 4331 621
rect 4417 618 4421 621
rect 4309 615 4332 618
rect 4413 615 4417 618
rect 4444 615 4481 626
rect 4766 615 4773 626
rect 4789 629 4799 635
rect 4817 630 4834 635
rect 4291 614 4332 615
rect 4291 609 4346 614
rect 4407 610 4412 614
rect 4444 610 4460 615
rect 4462 610 4478 615
rect 4773 610 4777 615
rect 4789 614 4813 629
rect 4817 626 4833 630
rect 4864 626 4873 635
rect 4878 626 4879 635
rect 4883 626 4884 642
rect 4919 641 4921 642
rect 4914 637 4919 641
rect 4894 635 4914 637
rect 4956 635 4959 642
rect 4894 632 4911 635
rect 4882 624 4884 626
rect 4889 627 4911 632
rect 4951 628 4956 635
rect 5004 630 5009 642
rect 4949 627 4951 628
rect 4889 625 4901 627
rect 4864 622 4882 624
rect 4833 620 4868 622
rect 4888 620 4901 625
rect 4789 612 4817 614
rect 4789 611 4831 612
rect 4834 611 4850 620
rect 4851 618 4868 620
rect 4852 614 4868 618
rect 4870 615 4901 620
rect 4932 616 4949 627
rect 5004 626 5007 630
rect 5078 626 5079 630
rect 5196 626 5212 642
rect 5251 630 5262 642
rect 6795 630 6804 644
rect 6874 642 6875 671
rect 7157 663 7159 688
rect 7185 663 7187 690
rect 7248 688 7251 690
rect 7287 687 7288 690
rect 7345 688 7349 690
rect 7427 688 7434 690
rect 7288 678 7294 687
rect 7321 678 7328 687
rect 7337 685 7360 688
rect 7418 687 7427 688
rect 7337 684 7362 685
rect 7337 683 7383 684
rect 7387 683 7389 687
rect 7413 685 7418 687
rect 7410 684 7413 685
rect 7408 683 7410 684
rect 7337 682 7408 683
rect 7445 682 7454 691
rect 7461 690 7468 692
rect 7491 692 7521 696
rect 7491 691 7522 692
rect 7540 691 7542 698
rect 7604 691 7637 700
rect 7720 695 7728 703
rect 7762 693 7784 706
rect 7789 700 7795 706
rect 7835 700 7837 725
rect 7839 713 7849 725
rect 7885 719 7891 725
rect 7912 719 7927 750
rect 7933 749 7934 753
rect 7969 751 8056 758
rect 8084 753 8090 760
rect 8134 758 8154 760
rect 8216 758 8232 774
rect 8234 770 8250 774
rect 8252 771 8259 774
rect 8263 773 8268 774
rect 8252 770 8258 771
rect 8261 770 8263 773
rect 8298 770 8304 774
rect 8234 764 8252 770
rect 8304 764 8310 770
rect 8234 758 8250 764
rect 8312 760 8326 774
rect 8379 761 8387 774
rect 9853 771 9854 781
rect 9882 773 9883 782
rect 10004 774 10070 782
rect 10094 774 10166 783
rect 10173 777 10177 812
rect 10201 803 10210 812
rect 10230 808 10246 823
rect 10248 803 10257 812
rect 10308 808 10324 824
rect 10326 808 10342 824
rect 10373 813 10377 828
rect 10430 825 10440 828
rect 10463 825 10471 846
rect 10520 843 10533 846
rect 10537 842 10539 843
rect 10541 842 10583 851
rect 10539 839 10583 842
rect 10541 835 10583 839
rect 10599 846 10653 851
rect 10692 850 10698 851
rect 10750 850 10831 851
rect 10658 846 10756 850
rect 10785 849 10787 850
rect 10796 849 10805 850
rect 10782 847 10792 849
rect 10797 848 10805 849
rect 10599 835 10629 846
rect 10653 845 10756 846
rect 10653 843 10665 845
rect 10680 843 10698 845
rect 10652 842 10653 843
rect 10787 842 10788 845
rect 10541 830 10629 835
rect 10641 831 10652 842
rect 10823 840 10829 850
rect 10541 825 10583 830
rect 10593 828 10617 830
rect 10640 828 10641 831
rect 10789 830 10792 838
rect 10830 830 10833 838
rect 10836 830 10842 850
rect 10863 839 10885 853
rect 10924 840 10929 858
rect 10985 857 10991 863
rect 10985 841 10990 857
rect 11027 841 11029 863
rect 11031 857 11037 863
rect 11079 862 11089 863
rect 11080 861 11089 862
rect 11080 859 11095 861
rect 11152 859 11158 865
rect 11199 864 11200 865
rect 11083 856 11108 859
rect 11083 853 11098 856
rect 11100 853 11106 856
rect 11136 854 11145 859
rect 11146 854 11152 859
rect 11182 857 11183 861
rect 11200 859 11202 864
rect 11202 856 11204 859
rect 11204 854 11205 856
rect 11285 854 11293 866
rect 11332 864 11335 868
rect 11364 864 11366 896
rect 11370 889 11378 898
rect 11370 879 11397 889
rect 11444 881 11447 885
rect 11437 879 11444 881
rect 11370 870 11437 879
rect 11391 869 11395 870
rect 11377 866 11391 869
rect 11372 865 11377 866
rect 11368 864 11372 865
rect 11328 856 11329 861
rect 11327 854 11329 856
rect 11089 850 11098 853
rect 11136 850 11155 854
rect 11144 846 11155 850
rect 11155 842 11156 846
rect 11183 842 11186 854
rect 11205 850 11207 854
rect 11293 851 11295 854
rect 11207 845 11211 850
rect 11211 843 11213 845
rect 11295 844 11300 850
rect 11213 842 11214 843
rect 11214 841 11216 842
rect 10985 839 11018 841
rect 10792 828 10793 830
rect 10593 825 10602 828
rect 10376 808 10377 813
rect 10428 824 10435 825
rect 10428 814 10438 824
rect 10428 812 10432 814
rect 10435 812 10438 814
rect 10460 813 10462 824
rect 10500 814 10516 824
rect 10493 813 10516 814
rect 10518 813 10541 824
rect 10585 820 10593 825
rect 10597 824 10602 825
rect 10261 803 10262 808
rect 10192 794 10205 803
rect 10257 794 10266 803
rect 10201 787 10205 794
rect 10261 792 10262 794
rect 10292 792 10308 808
rect 10343 807 10358 808
rect 10427 807 10428 811
rect 10436 808 10438 812
rect 10344 799 10358 807
rect 10377 800 10378 807
rect 10426 804 10427 807
rect 10425 800 10426 803
rect 10438 800 10454 808
rect 10459 807 10460 812
rect 10493 808 10534 813
rect 10484 806 10505 808
rect 10516 807 10522 808
rect 10458 800 10459 806
rect 10484 802 10500 806
rect 10510 802 10516 807
rect 10481 801 10527 802
rect 10481 800 10522 801
rect 10298 790 10304 792
rect 10307 791 10308 792
rect 10335 792 10358 799
rect 10378 797 10380 800
rect 10335 791 10350 792
rect 10306 790 10308 791
rect 10292 787 10308 790
rect 10309 789 10311 790
rect 10344 789 10350 791
rect 10309 787 10350 789
rect 10380 787 10390 797
rect 10422 787 10425 797
rect 10438 792 10458 800
rect 10453 790 10458 792
rect 10481 792 10500 800
rect 10534 792 10550 808
rect 10562 807 10568 813
rect 10575 812 10585 820
rect 10596 813 10602 824
rect 10617 823 10643 828
rect 10607 822 10650 823
rect 10607 821 10648 822
rect 10637 813 10640 821
rect 10650 818 10657 822
rect 10657 816 10658 818
rect 10569 807 10575 812
rect 10596 809 10597 813
rect 10658 812 10661 816
rect 10692 813 10708 824
rect 10710 813 10726 824
rect 10761 816 10770 825
rect 10793 824 10794 828
rect 10750 815 10761 816
rect 10683 812 10685 813
rect 10723 812 10727 813
rect 10636 809 10637 811
rect 10683 810 10727 812
rect 10683 808 10717 810
rect 10568 801 10574 807
rect 10580 792 10596 808
rect 10481 790 10491 792
rect 10493 790 10500 792
rect 10292 785 10347 787
rect 10203 777 10204 785
rect 10265 777 10271 783
rect 10292 781 10315 785
rect 9883 768 9884 771
rect 10020 767 10036 774
rect 10038 767 10054 774
rect 10094 771 10102 774
rect 10106 771 10152 774
rect 10102 767 10105 769
rect 10116 767 10132 771
rect 10134 767 10150 771
rect 8312 758 8329 760
rect 8134 753 8143 758
rect 8151 755 8152 757
rect 8323 753 8329 758
rect 8359 753 8371 761
rect 8379 756 8393 761
rect 8381 753 8393 756
rect 7969 749 8054 751
rect 8079 750 8092 753
rect 7934 746 7935 748
rect 7969 745 8060 749
rect 8072 748 8092 750
rect 8128 748 8134 753
rect 8072 746 8090 748
rect 8127 746 8128 748
rect 8076 745 8090 746
rect 7935 735 7937 744
rect 7988 743 8090 745
rect 7988 740 8020 743
rect 8036 740 8090 743
rect 7937 732 7938 735
rect 7938 730 7939 731
rect 7939 726 7940 730
rect 7988 729 8090 740
rect 8113 732 8115 743
rect 8122 740 8127 746
rect 8152 742 8155 753
rect 8119 736 8122 740
rect 8118 735 8119 736
rect 8116 732 8118 735
rect 8111 730 8116 732
rect 7999 727 8003 729
rect 8040 728 8044 729
rect 7998 725 8003 727
rect 8039 725 8040 727
rect 8101 725 8111 730
rect 7931 719 7937 725
rect 7940 721 7944 724
rect 7997 722 8003 725
rect 8059 724 8111 725
rect 7996 721 8003 722
rect 8037 721 8038 722
rect 8059 721 8101 724
rect 7879 713 7885 719
rect 7937 713 7943 719
rect 7944 717 8043 721
rect 8059 717 8094 721
rect 8113 720 8115 730
rect 8155 724 8156 742
rect 8258 740 8284 753
rect 8287 748 8292 753
rect 8329 748 8332 753
rect 8355 750 8356 752
rect 8387 749 8393 753
rect 8287 747 8293 748
rect 8287 740 8292 747
rect 8332 746 8334 748
rect 8347 746 8355 749
rect 8359 747 8393 749
rect 8390 746 8393 747
rect 8293 740 8294 746
rect 8334 740 8339 746
rect 8340 740 8353 746
rect 8156 719 8159 724
rect 8112 717 8113 719
rect 8246 718 8252 731
rect 8257 724 8258 730
rect 8294 726 8296 740
rect 8258 722 8260 724
rect 8258 721 8262 722
rect 8290 721 8292 724
rect 8258 719 8292 721
rect 8296 719 8298 726
rect 8316 725 8317 727
rect 8339 726 8353 740
rect 8304 722 8310 724
rect 8304 719 8314 722
rect 8340 720 8357 726
rect 8284 718 8314 719
rect 7839 712 7841 713
rect 7839 707 7847 712
rect 7944 707 8085 717
rect 8086 712 8094 717
rect 8252 716 8258 718
rect 8294 717 8304 718
rect 8294 716 8296 717
rect 8165 715 8167 716
rect 8252 715 8296 716
rect 8108 712 8110 715
rect 7841 706 7847 707
rect 7841 700 7853 706
rect 7464 687 7468 690
rect 7466 685 7468 687
rect 7467 683 7468 685
rect 7509 690 7522 691
rect 7509 687 7523 690
rect 7509 683 7531 687
rect 7387 678 7389 682
rect 7251 673 7252 676
rect 7249 668 7252 673
rect 7294 671 7298 678
rect 7328 671 7333 678
rect 7467 677 7471 683
rect 7509 679 7528 683
rect 7531 682 7533 683
rect 7536 682 7540 690
rect 7607 686 7627 691
rect 7601 683 7627 686
rect 7600 682 7627 683
rect 7637 682 7646 691
rect 7762 690 7779 693
rect 7784 691 7785 693
rect 7786 689 7790 690
rect 7841 689 7847 700
rect 7869 698 7878 700
rect 7869 691 7882 698
rect 7778 687 7790 689
rect 7839 688 7847 689
rect 7835 687 7839 688
rect 7778 685 7793 687
rect 7824 685 7835 687
rect 7778 683 7813 685
rect 7817 683 7824 685
rect 7533 681 7540 682
rect 7587 681 7627 682
rect 7533 680 7569 681
rect 7587 680 7599 681
rect 7536 679 7557 680
rect 7578 679 7610 680
rect 7509 678 7606 679
rect 7509 677 7528 678
rect 7400 675 7410 676
rect 7471 675 7472 676
rect 7528 675 7530 676
rect 7413 674 7421 675
rect 7418 671 7432 674
rect 7298 668 7300 671
rect 7242 667 7252 668
rect 7270 667 7281 668
rect 7225 664 7242 667
rect 7214 663 7225 664
rect 7107 662 7225 663
rect 7249 662 7252 667
rect 7281 666 7302 667
rect 7281 664 7304 666
rect 7301 663 7316 664
rect 7336 663 7341 668
rect 7432 667 7434 671
rect 7448 664 7459 667
rect 7443 663 7448 664
rect 7301 662 7448 663
rect 7107 659 7214 662
rect 7107 657 7193 659
rect 7248 657 7249 659
rect 7107 656 7181 657
rect 7107 655 7177 656
rect 7107 654 7170 655
rect 7107 653 7165 654
rect 7107 648 7159 653
rect 7101 642 7165 648
rect 5249 626 5262 630
rect 5077 624 5078 625
rect 5072 619 5077 624
rect 4882 614 4901 615
rect 4851 612 4901 614
rect 4852 611 4901 612
rect 4386 609 4407 610
rect 4789 609 4901 611
rect 4923 610 4932 616
rect 5007 615 5014 619
rect 5070 616 5072 619
rect 5067 615 5070 616
rect 5014 614 5067 615
rect 5020 610 5036 614
rect 5212 610 5228 626
rect 5230 610 5246 626
rect 5965 623 5992 629
rect 6804 626 6808 630
rect 6864 626 6880 642
rect 7107 636 7113 642
rect 7123 638 7129 642
rect 7129 634 7134 638
rect 7153 636 7159 642
rect 7185 634 7187 657
rect 7244 642 7248 657
rect 7304 655 7308 660
rect 7316 659 7443 662
rect 7472 660 7479 675
rect 7529 671 7532 675
rect 7536 674 7540 678
rect 7662 675 7668 677
rect 7640 674 7668 675
rect 7535 672 7536 674
rect 7633 672 7641 674
rect 7662 671 7670 674
rect 7720 671 7726 677
rect 7778 674 7794 683
rect 7518 668 7535 671
rect 7486 664 7500 667
rect 7500 663 7506 664
rect 7513 663 7533 668
rect 7668 665 7674 671
rect 7714 665 7720 671
rect 7622 663 7625 664
rect 7841 663 7847 688
rect 7860 682 7875 691
rect 7988 689 7994 707
rect 8021 706 8036 707
rect 8021 705 8050 706
rect 7500 662 7625 663
rect 7506 660 7622 662
rect 7795 660 7847 663
rect 7513 659 7622 660
rect 7342 657 7431 659
rect 7342 654 7346 657
rect 7359 656 7424 657
rect 7363 655 7421 656
rect 7373 654 7415 655
rect 7308 652 7309 654
rect 7346 652 7347 654
rect 7379 653 7415 654
rect 7309 649 7311 652
rect 7312 642 7317 648
rect 7347 642 7356 652
rect 7389 644 7390 646
rect 7380 642 7395 644
rect 7244 634 7258 642
rect 7356 639 7358 642
rect 7380 639 7396 642
rect 7358 637 7359 639
rect 7380 637 7407 639
rect 7134 632 7201 634
rect 6808 624 6864 626
rect 5993 623 6020 624
rect 6848 610 6864 624
rect 7185 614 7187 632
rect 7192 630 7204 632
rect 7243 630 7258 634
rect 7360 633 7363 637
rect 7380 635 7389 637
rect 7393 635 7438 637
rect 7445 635 7454 644
rect 7192 626 7208 630
rect 7242 626 7258 630
rect 7208 610 7224 626
rect 7226 610 7242 626
rect 7326 615 7343 633
rect 7361 625 7383 633
rect 7389 626 7398 635
rect 7436 626 7445 635
rect 7479 630 7494 659
rect 7516 657 7614 659
rect 7516 655 7522 657
rect 7527 656 7609 657
rect 7529 655 7609 656
rect 7531 652 7603 655
rect 7789 654 7853 660
rect 7510 650 7513 652
rect 7531 651 7590 652
rect 7531 650 7546 651
rect 7556 650 7562 651
rect 7503 645 7509 649
rect 7531 645 7554 650
rect 7565 645 7584 650
rect 7795 648 7801 654
rect 7810 652 7811 654
rect 7811 650 7812 652
rect 7531 644 7551 645
rect 7531 642 7533 644
rect 7535 642 7551 644
rect 7575 642 7584 645
rect 7812 644 7814 649
rect 7841 648 7847 654
rect 7496 639 7500 642
rect 7531 641 7551 642
rect 7531 634 7546 641
rect 7572 635 7584 642
rect 7637 635 7646 644
rect 7841 642 7842 648
rect 7869 645 7875 682
rect 7895 677 7898 683
rect 7931 676 7933 683
rect 7879 667 7885 673
rect 7886 667 7895 676
rect 7885 663 7895 667
rect 7899 663 7901 673
rect 7931 671 7934 676
rect 7983 674 7988 689
rect 7930 667 7934 671
rect 7937 667 7943 673
rect 8021 672 8036 705
rect 8067 704 8071 705
rect 8091 694 8101 705
rect 8167 694 8235 715
rect 8252 712 8270 715
rect 8257 708 8270 712
rect 8298 712 8304 717
rect 8337 715 8339 718
rect 8350 716 8357 720
rect 8357 715 8359 716
rect 8391 715 8393 746
rect 8397 737 8405 749
rect 9852 743 9853 767
rect 9884 742 9887 767
rect 10020 759 10054 767
rect 10106 759 10150 767
rect 10020 758 10036 759
rect 10038 758 10057 759
rect 10116 758 10132 759
rect 10134 758 10150 759
rect 10173 763 10176 777
rect 10178 763 10184 771
rect 10042 753 10057 758
rect 10173 757 10184 763
rect 10113 753 10122 756
rect 10167 754 10184 757
rect 10201 756 10204 777
rect 10149 753 10184 754
rect 9986 740 10184 753
rect 10192 747 10204 756
rect 10270 771 10277 777
rect 10292 774 10313 781
rect 10057 738 10066 740
rect 10072 737 10178 740
rect 10201 738 10210 747
rect 10212 741 10219 747
rect 9887 733 9888 737
rect 8397 715 8405 727
rect 9888 724 9889 731
rect 10150 730 10152 737
rect 10173 730 10179 737
rect 10270 731 10271 771
rect 10298 753 10313 774
rect 10345 778 10346 785
rect 10350 778 10359 787
rect 10345 756 10347 778
rect 10351 775 10359 778
rect 10388 782 10403 787
rect 10420 782 10422 787
rect 10438 782 10458 790
rect 10388 778 10458 782
rect 10484 780 10500 790
rect 10388 774 10463 778
rect 10404 772 10420 774
rect 10422 772 10438 774
rect 10453 772 10463 774
rect 10481 774 10500 780
rect 10534 774 10550 790
rect 10580 780 10596 790
rect 10631 789 10636 808
rect 10666 803 10668 806
rect 10676 805 10692 808
rect 10727 807 10742 808
rect 10752 807 10761 815
rect 10788 810 10804 824
rect 10806 810 10822 824
rect 10833 823 10836 830
rect 10833 818 10838 823
rect 10832 816 10833 818
rect 10836 816 10838 818
rect 10863 816 10879 839
rect 10886 830 10893 838
rect 10929 830 10932 839
rect 10980 835 10991 839
rect 10980 831 10985 835
rect 10893 824 10896 830
rect 10932 828 10933 830
rect 10978 828 10980 831
rect 10989 828 10991 835
rect 10884 816 10900 824
rect 10828 813 10831 815
rect 10780 808 10823 810
rect 10838 808 10842 816
rect 10861 812 10863 816
rect 10772 807 10783 808
rect 10797 807 10799 808
rect 10823 807 10842 808
rect 10676 799 10698 805
rect 10676 798 10692 799
rect 10672 792 10692 798
rect 10698 793 10704 799
rect 10672 789 10679 792
rect 10683 789 10692 792
rect 10726 792 10742 807
rect 10750 799 10756 805
rect 10744 793 10750 799
rect 10726 790 10727 792
rect 10631 780 10646 789
rect 10676 788 10692 789
rect 10580 774 10646 780
rect 10671 778 10692 788
rect 10721 787 10723 790
rect 10726 787 10742 790
rect 10715 778 10717 787
rect 10671 776 10717 778
rect 10721 776 10742 787
rect 10759 785 10780 807
rect 10800 803 10801 805
rect 10813 799 10819 804
rect 10802 795 10803 797
rect 10823 795 10838 807
rect 10858 806 10861 812
rect 10884 811 10905 816
rect 10933 813 10938 828
rect 10971 817 10978 828
rect 10984 818 10985 828
rect 10971 816 10984 817
rect 10968 815 10971 816
rect 10953 814 10965 815
rect 10951 813 10953 814
rect 10929 812 10943 813
rect 10917 811 10929 812
rect 10884 810 10917 811
rect 10884 808 10905 810
rect 10933 808 10938 812
rect 10842 801 10844 805
rect 10849 795 10858 806
rect 10793 787 10809 795
rect 10823 792 10849 795
rect 10868 792 10884 808
rect 10900 806 10905 808
rect 10977 806 10984 816
rect 10989 809 10990 828
rect 10989 806 10992 809
rect 11021 807 11023 839
rect 11156 836 11158 841
rect 11186 836 11187 841
rect 11216 839 11240 841
rect 10977 805 10985 806
rect 11013 805 11023 807
rect 11027 805 11035 817
rect 11076 815 11092 824
rect 11094 815 11110 824
rect 11076 814 11110 815
rect 11158 814 11160 836
rect 11187 824 11193 836
rect 11218 830 11232 839
rect 11300 836 11302 842
rect 11325 841 11329 854
rect 11324 836 11329 841
rect 11317 834 11329 836
rect 11341 860 11369 861
rect 11341 855 11368 860
rect 11232 828 11240 830
rect 11233 825 11236 828
rect 11076 813 11111 814
rect 11074 811 11076 813
rect 11109 812 11110 813
rect 11074 808 11110 811
rect 11172 809 11206 824
rect 11236 815 11240 825
rect 11240 811 11241 814
rect 11241 809 11242 811
rect 11302 809 11303 811
rect 11169 808 11206 809
rect 11242 808 11243 809
rect 10905 801 10907 805
rect 10938 800 10940 805
rect 10985 802 10989 805
rect 10989 801 11013 802
rect 11021 801 11023 805
rect 11060 801 11086 808
rect 11096 801 11108 808
rect 10940 797 10941 800
rect 10909 795 10910 797
rect 10837 790 10849 792
rect 10910 791 10913 795
rect 10676 774 10687 776
rect 10722 774 10742 776
rect 10404 766 10469 772
rect 10481 768 10491 774
rect 10493 771 10527 774
rect 10530 771 10534 774
rect 10493 768 10534 771
rect 10404 758 10463 766
rect 10489 764 10491 768
rect 10500 764 10516 768
rect 10344 753 10347 756
rect 10350 753 10353 754
rect 10298 744 10353 753
rect 10411 749 10463 758
rect 10493 758 10516 764
rect 10518 758 10534 768
rect 10596 761 10612 774
rect 10493 756 10505 758
rect 10510 755 10516 758
rect 10568 755 10574 761
rect 10593 758 10612 761
rect 10614 758 10630 774
rect 10692 772 10708 774
rect 10710 772 10726 774
rect 10645 761 10651 767
rect 10683 764 10726 772
rect 10756 768 10760 785
rect 10793 780 10810 787
rect 10780 768 10786 773
rect 10806 772 10810 780
rect 10823 780 10853 790
rect 10823 774 10838 780
rect 10849 779 10853 780
rect 10832 773 10837 774
rect 10810 771 10811 772
rect 10593 755 10599 758
rect 10651 755 10657 761
rect 10692 758 10708 764
rect 10710 758 10726 764
rect 10516 749 10522 755
rect 10562 749 10568 755
rect 10595 754 10599 755
rect 10754 754 10760 768
rect 10802 767 10823 771
rect 10827 767 10832 773
rect 10768 757 10770 758
rect 10767 755 10768 757
rect 10592 750 10596 754
rect 10763 752 10767 755
rect 10802 753 10827 767
rect 10853 763 10864 779
rect 10868 774 10884 790
rect 10913 779 10918 790
rect 10918 776 10926 779
rect 10941 778 10957 797
rect 10989 793 11001 801
rect 11011 793 11023 801
rect 11054 797 11076 801
rect 11100 797 11106 801
rect 11054 795 11108 797
rect 11110 795 11126 808
rect 11156 795 11169 808
rect 11187 806 11193 808
rect 11193 802 11194 806
rect 11019 778 11023 793
rect 11048 789 11076 795
rect 10941 776 10979 778
rect 10918 775 10957 776
rect 10918 774 10934 775
rect 10864 754 10870 763
rect 10884 758 10900 774
rect 10902 763 10926 774
rect 10941 764 10957 775
rect 10964 775 10979 776
rect 10964 774 10980 775
rect 10980 763 10982 774
rect 11019 763 11021 778
rect 10902 758 10918 763
rect 10926 753 10931 763
rect 10957 754 10962 763
rect 10980 758 10985 763
rect 11020 761 11021 763
rect 11054 774 11076 789
rect 11106 792 11126 795
rect 11106 790 11120 792
rect 11106 789 11126 790
rect 11106 781 11108 789
rect 11107 774 11108 781
rect 11110 774 11126 789
rect 11149 784 11159 795
rect 11161 787 11162 795
rect 11194 786 11197 800
rect 11206 792 11222 808
rect 11147 780 11149 784
rect 11162 782 11163 786
rect 11197 781 11198 786
rect 11145 774 11147 780
rect 11198 778 11199 781
rect 11199 774 11201 778
rect 11206 774 11222 790
rect 11243 786 11251 808
rect 11317 806 11324 834
rect 11341 826 11362 855
rect 11316 802 11317 806
rect 11329 803 11338 812
rect 11341 808 11352 826
rect 11378 824 11388 847
rect 11364 818 11398 824
rect 11860 819 11861 1015
rect 12050 819 12051 1015
rect 12136 819 12137 1015
rect 12409 819 12410 1015
rect 12606 819 12607 1015
rect 13204 1012 13205 1015
rect 13263 1013 13264 1016
rect 13260 1012 13264 1013
rect 13504 1014 13520 1016
rect 13548 1015 13560 1016
rect 13522 1014 13544 1015
rect 13556 1014 13560 1015
rect 13504 1012 13565 1014
rect 13596 1012 13816 1021
rect 13987 1017 13998 1021
rect 13987 1014 14005 1017
rect 14008 1014 14073 1030
rect 13987 1012 14073 1014
rect 13194 1005 13200 1011
rect 13203 1008 13204 1012
rect 13202 1005 13203 1008
rect 13240 1005 13246 1011
rect 13188 999 13194 1005
rect 13246 999 13252 1005
rect 13214 990 13215 997
rect 13253 995 13254 1012
rect 13259 1001 13266 1012
rect 13504 1011 13562 1012
rect 13495 1008 13501 1011
rect 13502 1009 13504 1011
rect 13506 1010 13511 1011
rect 13505 1009 13511 1010
rect 13565 1009 13566 1011
rect 13587 1010 13595 1012
rect 13993 1011 14002 1012
rect 13987 1010 14000 1011
rect 14008 1010 14073 1012
rect 13502 1008 13509 1009
rect 13567 1008 13587 1010
rect 13495 1006 13503 1008
rect 13488 1005 13503 1006
rect 13505 1005 13509 1008
rect 13485 1001 13503 1005
rect 13557 1001 13560 1008
rect 13259 998 13260 1001
rect 13258 997 13259 998
rect 13252 990 13254 994
rect 13255 990 13259 997
rect 13467 994 13485 1001
rect 13488 997 13503 1001
rect 13214 989 13231 990
rect 13215 988 13231 989
rect 13200 978 13231 988
rect 13235 978 13266 990
rect 13445 986 13467 994
rect 13488 990 13504 997
rect 13558 996 13559 1000
rect 13563 998 13587 1008
rect 13987 1009 13999 1010
rect 14000 1009 14073 1010
rect 14089 1009 14170 1030
rect 16601 1027 16639 1038
rect 17069 1030 17075 1036
rect 14901 1015 14902 1026
rect 15091 1015 15092 1026
rect 15177 1015 15178 1026
rect 15450 1015 15451 1026
rect 15647 1015 15648 1026
rect 16268 1025 16307 1026
rect 16268 1024 16305 1025
rect 16307 1024 16308 1025
rect 16266 1022 16268 1024
rect 16294 1016 16306 1024
rect 16308 1022 16309 1024
rect 16568 1022 16601 1027
rect 16973 1025 17029 1027
rect 16309 1016 16315 1022
rect 16556 1020 16601 1022
rect 16868 1021 16973 1025
rect 17029 1021 17039 1025
rect 16556 1016 16612 1020
rect 16257 1015 16309 1016
rect 13987 1005 14008 1009
rect 13563 996 13572 998
rect 13558 995 13560 996
rect 13563 995 13567 996
rect 13503 988 13504 990
rect 13426 979 13445 986
rect 13200 972 13266 978
rect 13412 974 13426 979
rect 13161 967 13167 968
rect 12922 965 12924 967
rect 12977 964 12978 967
rect 13154 964 13158 967
rect 13167 964 13174 967
rect 12978 962 12980 964
rect 13141 956 13154 964
rect 13174 963 13179 964
rect 13179 959 13190 963
rect 13216 961 13232 972
rect 13234 966 13254 972
rect 13404 971 13410 973
rect 13488 972 13504 988
rect 13548 992 13563 995
rect 13569 993 13571 996
rect 13548 986 13564 992
rect 13570 988 13571 993
rect 13567 986 13570 988
rect 13713 986 13734 1002
rect 13980 1001 13987 1005
rect 13993 1001 14008 1005
rect 13966 994 13980 1001
rect 14000 998 14008 1001
rect 14026 1005 14036 1009
rect 14170 1005 14187 1009
rect 14026 1003 14039 1005
rect 14008 995 14009 998
rect 13548 985 13572 986
rect 13927 985 13933 991
rect 13951 986 13966 994
rect 13949 985 13951 986
rect 13973 985 13979 991
rect 14009 985 14016 995
rect 13547 983 13548 985
rect 13552 974 13572 985
rect 13747 974 13759 982
rect 13769 974 13781 982
rect 13921 979 13927 985
rect 13979 979 13985 985
rect 14011 980 14019 985
rect 14011 979 14020 980
rect 14011 978 14021 979
rect 14011 975 14023 978
rect 13552 971 13564 974
rect 14011 973 14025 975
rect 14026 973 14027 1003
rect 14032 993 14053 1003
rect 14187 999 14209 1005
rect 14209 997 14211 999
rect 14036 983 14053 993
rect 14211 992 14217 997
rect 14217 986 14221 992
rect 14011 971 14027 973
rect 14032 972 14053 983
rect 14221 982 14224 986
rect 14224 975 14228 982
rect 14032 971 14154 972
rect 14228 971 14230 975
rect 13399 970 13404 971
rect 13396 969 13399 970
rect 13504 968 13522 971
rect 13548 970 13564 971
rect 13741 970 13743 971
rect 13783 970 13820 971
rect 13548 969 13561 970
rect 13296 967 13300 968
rect 13302 967 13307 968
rect 13234 961 13250 966
rect 13288 965 13296 967
rect 13286 964 13288 965
rect 13307 964 13310 967
rect 13388 966 13395 968
rect 13384 964 13388 966
rect 13283 963 13286 964
rect 13282 962 13283 963
rect 13310 962 13313 964
rect 13380 963 13384 964
rect 13202 959 13250 961
rect 13179 958 13194 959
rect 13202 958 13252 959
rect 13275 958 13284 962
rect 13313 959 13317 962
rect 13360 961 13380 963
rect 13182 956 13196 958
rect 13197 957 13252 958
rect 13138 954 13141 956
rect 13182 954 13199 956
rect 13202 954 13252 957
rect 13271 956 13284 958
rect 13317 956 13320 959
rect 13368 958 13374 961
rect 13267 954 13284 956
rect 13320 954 13323 956
rect 13357 954 13365 957
rect 13489 956 13495 959
rect 13504 956 13520 968
rect 13522 967 13529 968
rect 13529 965 13540 967
rect 13548 966 13560 969
rect 13547 965 13560 966
rect 13540 964 13560 965
rect 13580 964 13586 970
rect 13626 966 13632 970
rect 13735 969 13741 970
rect 13616 964 13632 966
rect 13548 962 13560 964
rect 13467 954 13495 956
rect 12978 946 12979 949
rect 12977 945 13016 946
rect 12975 944 12977 945
rect 12960 934 12975 944
rect 12936 920 12960 934
rect 12933 918 12936 920
rect 12926 913 12933 918
rect 12978 913 12979 945
rect 13016 944 13043 945
rect 13120 944 13138 954
rect 13182 953 13252 954
rect 13182 951 13204 953
rect 13233 951 13234 953
rect 13240 951 13246 953
rect 13260 951 13284 954
rect 13182 948 13284 951
rect 13182 947 13237 948
rect 13240 947 13246 948
rect 13182 946 13216 947
rect 13218 946 13237 947
rect 13249 946 13284 948
rect 13182 944 13237 946
rect 13247 945 13284 946
rect 13246 944 13284 945
rect 13323 953 13346 954
rect 13354 953 13357 954
rect 13323 946 13354 953
rect 13323 944 13346 946
rect 13043 938 13284 944
rect 13313 938 13328 944
rect 13336 939 13346 944
rect 13342 938 13346 939
rect 13395 938 13485 954
rect 13489 953 13515 954
rect 13547 953 13553 959
rect 13574 958 13638 964
rect 13685 963 13691 969
rect 13731 968 13737 969
rect 13726 966 13737 968
rect 13720 964 13725 966
rect 13716 963 13720 964
rect 13731 963 13737 966
rect 13747 968 13781 970
rect 13785 969 13793 970
rect 13580 954 13632 958
rect 13679 957 13685 963
rect 13737 957 13743 963
rect 13495 947 13501 953
rect 13541 947 13547 953
rect 13580 938 13594 954
rect 13104 922 13120 938
rect 13166 937 13189 938
rect 13166 934 13194 937
rect 13166 933 13202 934
rect 13204 933 13212 935
rect 13233 934 13234 938
rect 13308 937 13313 938
rect 13299 935 13307 936
rect 13235 934 13282 935
rect 13294 934 13299 935
rect 13219 933 13282 934
rect 13346 933 13362 938
rect 13389 936 13395 938
rect 13580 936 13595 938
rect 13385 935 13388 936
rect 13380 933 13384 934
rect 13166 925 13274 933
rect 13233 924 13234 925
rect 13172 922 13189 924
rect 13104 916 13120 920
rect 13155 917 13170 922
rect 13193 920 13218 922
rect 13006 913 13047 916
rect 13051 913 13120 916
rect 12923 911 12926 913
rect 12978 911 13006 913
rect 13104 911 13148 913
rect 13154 911 13170 917
rect 13191 917 13218 920
rect 13237 918 13296 922
rect 13344 920 13380 933
rect 13578 931 13595 936
rect 13574 928 13578 931
rect 13567 924 13574 928
rect 13559 920 13567 924
rect 13580 920 13595 931
rect 13626 920 13628 954
rect 13632 950 13645 954
rect 13747 953 13768 968
rect 13778 967 13781 968
rect 13786 963 13793 969
rect 13821 966 13828 970
rect 14011 969 14025 971
rect 14026 970 14154 971
rect 14036 969 14053 970
rect 14057 969 14154 970
rect 13789 960 13791 963
rect 14007 960 14010 961
rect 13794 954 13801 957
rect 13746 952 13768 953
rect 13746 950 13747 952
rect 13632 942 13640 950
rect 13745 938 13746 949
rect 13801 940 13824 954
rect 13926 953 13927 957
rect 13985 954 14007 960
rect 14011 957 14030 969
rect 13985 952 14012 954
rect 13632 920 13640 932
rect 13339 918 13344 920
rect 13219 917 13296 918
rect 13191 915 13203 917
rect 13263 916 13274 917
rect 13211 914 13223 916
rect 13262 915 13264 916
rect 12919 909 12923 911
rect 12977 910 12979 911
rect 12975 906 12980 910
rect 12922 903 12923 904
rect 12913 894 12914 899
rect 12967 896 12968 904
rect 12974 903 12980 906
rect 13104 904 13120 911
rect 13148 910 13173 911
rect 13139 908 13170 910
rect 13173 909 13184 910
rect 13184 908 13191 909
rect 13129 906 13170 908
rect 13191 907 13204 908
rect 13212 906 13219 907
rect 13139 905 13170 906
rect 13154 904 13170 905
rect 12972 899 12980 903
rect 12972 895 12974 899
rect 12966 876 12968 895
rect 13120 888 13136 904
rect 13138 888 13154 904
rect 13231 888 13233 911
rect 13296 909 13312 917
rect 13328 913 13339 918
rect 13323 911 13327 913
rect 13317 909 13323 911
rect 13346 909 13362 920
rect 13546 912 13559 920
rect 13578 918 13632 920
rect 13643 918 13645 926
rect 13682 920 13685 937
rect 13824 935 13833 940
rect 13920 939 13926 952
rect 13930 946 13951 949
rect 13967 946 13968 949
rect 13979 948 13985 952
rect 13996 946 14012 952
rect 13920 936 13927 939
rect 13928 938 13930 946
rect 13951 939 14012 946
rect 14025 942 14030 957
rect 14053 968 14154 969
rect 14231 968 14232 970
rect 13959 938 14012 939
rect 13978 937 14028 938
rect 13745 925 13748 929
rect 13833 928 13844 935
rect 13920 933 13928 936
rect 13978 933 13985 937
rect 13574 912 13644 918
rect 13679 917 13681 919
rect 13748 918 13763 925
rect 13844 923 13848 928
rect 13848 920 13849 923
rect 13763 917 13786 918
rect 13679 916 13685 917
rect 13677 912 13685 916
rect 13544 911 13546 912
rect 13578 911 13593 912
rect 13594 911 13595 912
rect 13296 908 13362 909
rect 13282 907 13362 908
rect 13538 907 13544 911
rect 13578 907 13599 911
rect 13616 908 13632 912
rect 13240 906 13263 907
rect 13296 904 13362 907
rect 13330 888 13346 904
rect 13524 900 13538 907
rect 13578 904 13593 907
rect 13594 904 13595 907
rect 13626 906 13632 908
rect 13635 904 13644 912
rect 13679 911 13685 912
rect 13737 916 13786 917
rect 13737 911 13743 916
rect 13754 914 13786 916
rect 13763 913 13787 914
rect 13763 911 13786 913
rect 13789 911 13814 913
rect 13828 911 13842 920
rect 13849 918 13850 920
rect 13915 918 13920 933
rect 13926 927 13933 933
rect 13926 925 13928 927
rect 13850 911 13853 918
rect 13913 911 13915 915
rect 13674 907 13676 911
rect 13579 900 13592 904
rect 13633 900 13635 904
rect 13670 900 13674 907
rect 13685 905 13691 911
rect 13504 888 13527 900
rect 13574 897 13579 900
rect 13558 888 13574 897
rect 13591 896 13594 899
rect 13628 896 13633 899
rect 13668 897 13670 900
rect 13594 888 13610 896
rect 13612 888 13628 896
rect 13662 888 13668 897
rect 12972 875 12980 888
rect 13168 880 13298 888
rect 13501 883 13504 888
rect 13550 883 13558 888
rect 13659 883 13662 888
rect 13416 880 13464 883
rect 13146 875 13188 880
rect 12966 873 12972 875
rect 13135 873 13188 875
rect 12923 870 12927 873
rect 12956 871 12966 873
rect 12969 872 12972 873
rect 12956 870 12968 871
rect 13116 870 13188 873
rect 13231 870 13233 880
rect 13275 879 13416 880
rect 13278 875 13416 879
rect 13464 875 13465 880
rect 13497 875 13501 883
rect 13536 876 13550 883
rect 13654 876 13659 883
rect 13530 875 13536 876
rect 13697 875 13721 910
rect 13731 905 13737 911
rect 13763 909 13842 911
rect 13853 909 13854 911
rect 13776 904 13842 909
rect 13854 904 13856 908
rect 13792 888 13808 904
rect 13810 893 13826 904
rect 13856 899 13858 903
rect 13858 893 13860 899
rect 13901 898 13913 910
rect 13922 909 13926 925
rect 13959 916 13967 933
rect 13973 927 13979 933
rect 13921 904 13922 909
rect 13939 905 13959 915
rect 13926 903 13938 905
rect 13939 903 13960 905
rect 13978 904 13979 927
rect 14012 922 14028 937
rect 14030 936 14031 941
rect 14053 938 14074 968
rect 14094 965 14154 968
rect 14232 967 14233 968
rect 14233 965 14236 967
rect 14123 963 14154 965
rect 14236 963 14238 965
rect 14132 961 14154 963
rect 14238 961 14242 963
rect 14086 938 14102 954
rect 14104 938 14120 954
rect 14144 949 14172 961
rect 14242 954 14251 961
rect 14130 938 14131 949
rect 14172 947 14176 949
rect 14251 947 14259 954
rect 14176 946 14177 947
rect 14177 944 14178 946
rect 14259 944 14261 947
rect 14447 944 14448 949
rect 14476 944 14492 954
rect 14178 939 14184 944
rect 14261 940 14266 944
rect 14430 940 14497 944
rect 14266 939 14268 940
rect 14407 939 14430 940
rect 14053 936 14086 938
rect 14091 936 14136 938
rect 14184 936 14186 938
rect 14268 936 14271 939
rect 14404 936 14407 939
rect 14447 938 14448 940
rect 14497 938 14498 939
rect 14031 916 14036 933
rect 14053 922 14085 936
rect 14122 934 14136 936
rect 14186 934 14188 936
rect 14271 934 14275 936
rect 14401 934 14404 936
rect 14116 932 14136 934
rect 14188 932 14189 934
rect 14275 932 14277 934
rect 14400 932 14401 934
rect 14037 915 14043 921
rect 14053 919 14074 922
rect 14078 921 14085 922
rect 14074 915 14077 919
rect 14078 915 14089 921
rect 14031 909 14037 915
rect 14036 908 14037 909
rect 14078 906 14085 915
rect 14089 909 14095 915
rect 14127 904 14163 932
rect 14189 925 14196 932
rect 14277 925 14288 932
rect 14397 925 14400 932
rect 14196 924 14210 925
rect 14188 915 14210 924
rect 14288 919 14297 925
rect 14394 919 14397 925
rect 14297 916 14300 919
rect 14393 916 14394 919
rect 14196 907 14210 915
rect 14300 912 14305 916
rect 14391 912 14393 916
rect 14305 907 14309 912
rect 14388 910 14391 912
rect 14204 905 14213 907
rect 14210 904 14213 905
rect 14309 904 14311 907
rect 13923 901 13963 903
rect 13920 900 13921 901
rect 13919 899 13920 900
rect 13923 899 13959 901
rect 13918 898 13923 899
rect 13901 896 13923 898
rect 13861 893 13913 896
rect 13918 893 13923 896
rect 13810 888 13829 893
rect 13860 888 13913 893
rect 13757 877 13766 881
rect 13804 877 13813 881
rect 13823 879 13829 888
rect 13855 886 13869 888
rect 13850 883 13855 886
rect 13860 883 13869 886
rect 13849 882 13869 883
rect 13841 880 13869 882
rect 13838 879 13869 880
rect 13823 877 13869 879
rect 13749 875 13869 877
rect 13278 870 13380 875
rect 13418 874 13572 875
rect 13418 872 13565 874
rect 13391 871 13418 872
rect 13383 870 13391 871
rect 12927 869 12956 870
rect 12964 867 12968 870
rect 13112 869 13116 870
rect 13378 869 13383 870
rect 12963 866 12968 867
rect 13099 866 13112 869
rect 13369 868 13378 869
rect 13361 866 13369 868
rect 13465 867 13468 872
rect 13497 871 13501 872
rect 13530 871 13536 872
rect 13572 871 13586 874
rect 13652 871 13654 875
rect 13668 872 13749 875
rect 13757 872 13869 875
rect 13901 872 13913 888
rect 13914 881 13919 893
rect 13918 880 13919 881
rect 13586 870 13590 871
rect 12911 859 12912 866
rect 12961 864 12968 866
rect 13077 865 13111 866
rect 13356 865 13361 866
rect 12961 859 12963 864
rect 13077 862 13099 865
rect 13076 859 13099 862
rect 13111 859 13118 865
rect 13323 859 13356 865
rect 12960 855 12961 859
rect 13072 855 13077 859
rect 13080 854 13099 859
rect 13118 857 13121 859
rect 13317 858 13323 859
rect 13310 857 13317 858
rect 13294 854 13309 857
rect 13468 854 13473 866
rect 13495 863 13497 870
rect 13527 863 13530 870
rect 13590 868 13602 870
rect 13494 860 13495 863
rect 13526 860 13527 863
rect 13602 859 13640 868
rect 13645 863 13650 870
rect 13668 868 13757 872
rect 13758 870 13869 872
rect 13939 871 13959 899
rect 13963 893 13967 901
rect 13967 873 13972 893
rect 14075 887 14078 904
rect 14135 903 14138 904
rect 14131 902 14135 903
rect 14130 899 14131 901
rect 14163 899 14170 904
rect 14123 887 14130 899
rect 14135 897 14136 899
rect 14169 893 14170 899
rect 14205 893 14212 898
rect 14213 893 14228 904
rect 14078 877 14103 887
rect 14129 877 14130 887
rect 14212 885 14224 893
rect 14228 887 14237 893
rect 14311 887 14324 904
rect 14384 902 14396 910
rect 14406 902 14418 910
rect 14458 904 14459 938
rect 14497 934 14508 938
rect 14498 922 14508 934
rect 14498 903 14499 922
rect 14384 898 14387 902
rect 14420 899 14422 902
rect 14372 886 14380 898
rect 14384 896 14418 898
rect 14384 895 14387 896
rect 14103 870 14130 877
rect 14224 876 14231 885
rect 14237 879 14243 886
rect 14324 879 14329 886
rect 14243 877 14245 879
rect 14329 877 14331 879
rect 14135 870 14136 872
rect 13666 866 13668 868
rect 13663 864 13666 866
rect 13693 864 13696 868
rect 13643 860 13645 863
rect 12959 851 12960 854
rect 13070 851 13072 854
rect 13079 850 13080 854
rect 12910 838 12911 850
rect 12955 838 12959 850
rect 13063 838 13070 850
rect 11364 812 11380 818
rect 11382 812 11398 818
rect 12909 816 12910 837
rect 12948 816 12955 838
rect 13063 835 13069 838
rect 13057 829 13063 835
rect 13071 828 13076 842
rect 13109 835 13115 841
rect 13121 839 13122 854
rect 13198 850 13294 854
rect 13473 850 13474 854
rect 13492 853 13494 859
rect 13523 853 13526 859
rect 13635 858 13645 859
rect 13635 853 13642 858
rect 13645 857 13651 858
rect 13660 857 13663 864
rect 13748 863 13757 868
rect 13813 863 13822 870
rect 13831 868 13832 870
rect 13869 868 13870 870
rect 13691 860 13693 863
rect 13832 861 13834 868
rect 13870 860 13873 868
rect 13899 864 13900 866
rect 13898 861 13899 863
rect 13914 859 13920 870
rect 13936 864 13939 870
rect 13972 866 13974 870
rect 14011 868 14012 869
rect 14009 865 14011 868
rect 14002 864 14009 865
rect 13926 859 13928 861
rect 13651 855 13674 857
rect 13689 856 13691 859
rect 13750 856 13756 857
rect 13796 856 13802 857
rect 13835 856 13836 857
rect 13874 856 13875 857
rect 13896 856 13897 859
rect 13922 856 13930 859
rect 13651 854 13664 855
rect 13684 854 13689 856
rect 13635 852 13638 853
rect 13635 851 13637 852
rect 13659 851 13660 854
rect 13664 851 13705 854
rect 13138 843 13199 850
rect 13137 841 13138 842
rect 13115 832 13121 835
rect 13122 832 13123 838
rect 13115 829 13123 832
rect 13131 829 13137 841
rect 13141 840 13152 842
rect 13198 840 13199 843
rect 13209 843 13399 850
rect 13474 846 13477 850
rect 13484 846 13492 851
rect 13515 847 13523 851
rect 13510 846 13571 847
rect 13421 843 13503 846
rect 13209 839 13294 843
rect 13387 842 13405 843
rect 13474 842 13477 843
rect 13369 839 13387 842
rect 13405 841 13417 842
rect 13420 839 13423 841
rect 13207 838 13209 839
rect 13202 835 13206 838
rect 13196 830 13202 835
rect 13229 831 13231 839
rect 13361 838 13369 839
rect 13345 835 13361 838
rect 13119 828 13123 829
rect 13195 828 13196 830
rect 11364 809 11398 812
rect 12908 810 12909 816
rect 12947 811 12948 816
rect 12976 811 12992 824
rect 13070 813 13071 828
rect 13115 826 13117 827
rect 13119 826 13131 828
rect 13117 816 13139 826
rect 13168 817 13184 824
rect 13115 812 13139 816
rect 13158 812 13184 817
rect 13115 811 13117 812
rect 11364 808 11410 809
rect 11313 790 11316 800
rect 11320 794 11329 803
rect 11341 792 11364 808
rect 11376 803 11385 808
rect 11410 805 11415 808
rect 12945 807 12947 810
rect 13121 808 13131 812
rect 11385 794 11394 803
rect 11303 787 11318 790
rect 11251 779 11257 786
rect 11276 780 11318 787
rect 11324 786 11328 792
rect 11341 790 11351 792
rect 11341 787 11364 790
rect 11320 780 11322 784
rect 11341 781 11378 787
rect 11252 774 11268 779
rect 11276 774 11320 780
rect 11348 774 11378 781
rect 11415 774 11431 805
rect 12907 800 12908 805
rect 12942 800 12944 805
rect 12941 798 12942 800
rect 12937 790 12941 798
rect 12960 792 12971 808
rect 13120 806 13121 808
rect 13139 807 13148 812
rect 13156 809 13184 812
rect 13154 808 13165 809
rect 13168 808 13184 809
rect 13186 808 13202 824
rect 13225 818 13231 831
rect 13311 830 13345 835
rect 13269 823 13311 830
rect 13423 829 13425 839
rect 13477 829 13482 842
rect 13484 828 13492 843
rect 13261 822 13269 823
rect 13236 818 13261 822
rect 13225 816 13236 818
rect 13221 812 13231 816
rect 13152 807 13168 808
rect 13148 806 13168 807
rect 13148 805 13165 806
rect 13202 805 13218 808
rect 13070 790 13071 805
rect 12935 786 12937 790
rect 13056 787 13071 790
rect 13109 789 13120 805
rect 13146 803 13179 805
rect 13146 794 13174 803
rect 13196 797 13218 805
rect 13146 793 13168 794
rect 13152 792 13168 793
rect 13158 790 13168 792
rect 13192 792 13218 797
rect 13192 791 13202 792
rect 13109 787 13121 789
rect 12906 782 12907 786
rect 13056 783 13121 787
rect 13152 787 13168 790
rect 13185 790 13202 791
rect 13185 787 13218 790
rect 13152 783 13218 787
rect 13056 782 13120 783
rect 11054 761 11110 774
rect 11112 763 11120 774
rect 11142 763 11145 774
rect 11163 764 11164 770
rect 10982 753 10985 758
rect 11021 758 11110 761
rect 11141 760 11144 763
rect 11195 760 11206 774
rect 10411 745 10470 749
rect 10592 746 10599 750
rect 10753 748 10763 752
rect 10800 749 10802 753
rect 10631 746 10728 748
rect 10751 746 10763 748
rect 10799 746 10800 748
rect 10591 745 10599 746
rect 10602 745 10737 746
rect 10748 745 10750 746
rect 10753 745 10763 746
rect 10298 741 10350 744
rect 10353 742 10354 744
rect 10292 736 10356 741
rect 10411 740 10550 745
rect 10591 744 10763 745
rect 10292 735 10358 736
rect 10213 730 10219 731
rect 10134 727 10236 730
rect 10134 724 10261 727
rect 10270 725 10277 731
rect 10298 729 10304 735
rect 10313 727 10316 732
rect 10344 729 10350 735
rect 10355 727 10358 735
rect 10317 725 10318 727
rect 10358 725 10359 727
rect 10411 726 10419 740
rect 10463 736 10550 740
rect 10465 730 10550 736
rect 10583 743 10763 744
rect 10795 743 10799 745
rect 10809 744 10827 753
rect 10931 750 10933 753
rect 10962 750 10964 753
rect 10832 744 10872 745
rect 10873 744 10884 750
rect 10583 740 10760 743
rect 10583 732 10597 740
rect 10795 735 10809 743
rect 10472 729 10473 730
rect 10473 727 10474 729
rect 8298 709 8299 712
rect 8258 707 8270 708
rect 8299 702 8300 703
rect 8258 698 8259 701
rect 8320 696 8337 714
rect 9850 713 9851 724
rect 9889 717 9890 724
rect 10134 720 10183 724
rect 10134 717 10190 720
rect 10219 719 10225 724
rect 10134 716 10142 717
rect 10134 715 10141 716
rect 8394 711 8397 713
rect 9890 711 9891 713
rect 10153 712 10155 717
rect 8387 710 8394 711
rect 10183 710 10190 717
rect 8381 708 8393 710
rect 8370 703 8393 708
rect 9849 707 9850 710
rect 10034 707 10117 710
rect 8370 696 8381 703
rect 10155 696 10158 709
rect 10190 708 10200 709
rect 10168 700 10180 708
rect 10190 700 10202 708
rect 10159 698 10164 700
rect 10166 698 10211 700
rect 10159 697 10211 698
rect 10237 697 10239 722
rect 10265 719 10271 725
rect 10318 723 10319 725
rect 10359 720 10360 722
rect 10405 720 10421 726
rect 10321 715 10323 719
rect 10360 716 10361 719
rect 10407 716 10421 720
rect 10425 716 10428 719
rect 10451 718 10453 726
rect 10463 720 10469 726
rect 10550 725 10559 730
rect 10475 723 10476 725
rect 10450 716 10453 718
rect 10457 716 10465 720
rect 10323 709 10327 715
rect 10361 710 10363 715
rect 10407 714 10417 716
rect 10407 713 10416 714
rect 10419 713 10440 716
rect 10450 713 10452 716
rect 10455 713 10465 716
rect 10416 710 10417 713
rect 10428 710 10431 713
rect 10444 712 10448 713
rect 10448 711 10453 712
rect 10455 711 10457 713
rect 10440 710 10455 711
rect 10476 710 10483 722
rect 10559 713 10564 724
rect 10591 722 10597 732
rect 10720 723 10726 729
rect 10736 727 10742 732
rect 10731 723 10736 727
rect 10766 723 10772 729
rect 10792 727 10795 735
rect 10796 727 10809 735
rect 10792 725 10796 727
rect 10817 726 10825 744
rect 10832 740 10884 744
rect 10830 735 10866 740
rect 10872 737 10884 740
rect 10933 747 10936 750
rect 10872 735 10889 737
rect 10830 731 10832 735
rect 10873 734 10889 735
rect 10933 734 10938 747
rect 10883 731 10889 734
rect 10884 730 10889 731
rect 10887 729 10891 730
rect 10936 729 10938 734
rect 10889 726 10893 729
rect 10583 719 10597 722
rect 10583 716 10599 719
rect 10651 716 10652 719
rect 10714 717 10720 723
rect 10772 717 10778 723
rect 10788 722 10792 724
rect 10793 723 10796 725
rect 10819 724 10820 726
rect 10891 725 10893 726
rect 10937 725 10938 729
rect 10825 724 10826 725
rect 10328 698 10334 708
rect 10364 698 10366 708
rect 10419 701 10431 710
rect 10432 698 10438 708
rect 10441 701 10453 710
rect 10455 709 10520 710
rect 10462 707 10520 709
rect 10469 706 10520 707
rect 10477 703 10520 706
rect 10483 700 10489 703
rect 10491 702 10520 703
rect 10492 701 10520 702
rect 10483 698 10497 700
rect 10334 697 10338 698
rect 10159 696 10338 697
rect 8300 695 8301 696
rect 8314 694 8332 696
rect 8082 690 8093 691
rect 8082 688 8091 690
rect 8082 687 8092 688
rect 8095 687 8096 690
rect 8098 688 8107 691
rect 8128 690 8130 691
rect 8235 688 8255 694
rect 8259 691 8260 692
rect 8291 690 8332 694
rect 9848 692 9849 696
rect 10155 695 10164 696
rect 10156 694 10164 695
rect 10168 694 10338 696
rect 10366 694 10370 698
rect 9853 690 9854 692
rect 8260 688 8262 690
rect 8291 688 8314 690
rect 8228 687 8322 688
rect 8079 685 8092 687
rect 8076 683 8079 685
rect 8065 677 8076 683
rect 8082 679 8090 685
rect 7981 667 7983 671
rect 7930 663 7937 667
rect 7885 661 7937 663
rect 7886 660 7945 661
rect 7869 644 7877 645
rect 7844 642 7851 643
rect 7815 637 7817 641
rect 7841 637 7851 642
rect 7860 642 7877 644
rect 7885 642 7886 659
rect 7887 649 7945 660
rect 7978 655 7981 667
rect 7977 652 7978 654
rect 8014 652 8021 672
rect 8061 668 8065 676
rect 8082 663 8090 669
rect 8094 663 8096 687
rect 8260 676 8262 687
rect 8301 682 8303 687
rect 8344 676 8354 680
rect 9851 676 9854 690
rect 8164 672 8184 673
rect 8148 664 8164 672
rect 8184 664 8236 672
rect 8144 663 8148 664
rect 8082 662 8148 663
rect 8236 663 8250 664
rect 8262 663 8264 676
rect 8338 674 8344 676
rect 8307 664 8338 674
rect 9848 670 9851 676
rect 8298 663 8307 664
rect 8236 662 8307 663
rect 7895 648 7937 649
rect 7895 645 7935 648
rect 7841 635 7848 637
rect 7860 635 7886 642
rect 7899 637 7911 645
rect 7921 644 7933 645
rect 7934 644 7935 645
rect 7921 642 7935 644
rect 7974 643 7976 647
rect 8012 645 8014 651
rect 8011 643 8012 645
rect 8059 642 8061 659
rect 8082 657 8143 662
rect 8250 661 8307 662
rect 9841 663 9851 670
rect 9853 663 9854 676
rect 9886 690 9887 692
rect 9888 690 9898 692
rect 9886 687 9913 690
rect 10153 688 10159 694
rect 9886 673 9917 687
rect 10156 684 10159 688
rect 10168 692 10264 694
rect 10168 690 10296 692
rect 10334 691 10393 694
rect 10334 690 10338 691
rect 10366 690 10370 691
rect 10393 690 10397 691
rect 10438 690 10439 696
rect 10489 695 10497 698
rect 10499 697 10520 701
rect 10561 709 10565 713
rect 10583 712 10601 716
rect 10626 712 10629 713
rect 10583 711 10599 712
rect 10583 710 10597 711
rect 10591 709 10599 710
rect 10601 709 10603 711
rect 10604 710 10629 712
rect 10644 710 10646 712
rect 10651 710 10657 715
rect 10705 710 10720 716
rect 10787 715 10792 722
rect 10780 711 10786 714
rect 10788 711 10792 715
rect 10814 716 10831 724
rect 10610 709 10712 710
rect 10561 707 10566 709
rect 10591 707 10597 709
rect 10632 707 10712 709
rect 10561 706 10567 707
rect 10594 706 10632 707
rect 10561 702 10568 706
rect 10561 701 10569 702
rect 10532 698 10542 699
rect 10561 698 10571 701
rect 10594 698 10607 706
rect 10645 703 10651 707
rect 10656 706 10712 707
rect 10780 709 10788 711
rect 10780 706 10786 709
rect 10814 708 10836 716
rect 10828 706 10836 708
rect 10847 706 10853 712
rect 10656 705 10725 706
rect 10772 705 10780 706
rect 10656 703 10780 705
rect 10656 700 10693 703
rect 10525 697 10529 698
rect 10507 695 10525 697
rect 10483 694 10525 695
rect 10543 696 10571 698
rect 10489 692 10520 694
rect 10489 691 10508 692
rect 10486 690 10494 691
rect 10168 688 10217 690
rect 10168 683 10202 688
rect 10168 682 10176 683
rect 10168 681 10175 682
rect 10068 673 10102 676
rect 9886 663 9887 673
rect 9892 663 9899 670
rect 8262 660 8264 661
rect 9841 658 9899 663
rect 9916 660 9917 673
rect 8090 656 8143 657
rect 9847 657 9892 658
rect 8090 655 8132 656
rect 8092 653 8130 655
rect 9847 653 9848 657
rect 9851 654 9889 657
rect 8094 645 8106 653
rect 8116 645 8128 653
rect 9853 646 9865 654
rect 9875 646 9887 654
rect 7921 641 7934 642
rect 7918 639 7934 641
rect 7921 637 7934 639
rect 7923 636 7934 637
rect 7913 635 7919 636
rect 7925 635 7934 636
rect 7478 626 7496 630
rect 7509 626 7546 634
rect 7581 626 7590 635
rect 7628 626 7637 635
rect 7818 630 7825 634
rect 7817 626 7825 630
rect 7478 625 7484 626
rect 7361 621 7376 625
rect 7473 621 7478 625
rect 7361 618 7383 621
rect 7469 618 7473 621
rect 7361 615 7384 618
rect 7465 615 7469 618
rect 7496 615 7533 626
rect 7818 615 7825 626
rect 7841 629 7851 635
rect 7869 630 7886 635
rect 7343 614 7384 615
rect 4291 607 4421 609
rect 4291 606 4311 607
rect 4431 606 4450 609
rect 4778 607 4901 609
rect 3772 557 3822 606
rect 3852 557 3918 606
rect 3948 557 4014 606
rect 4044 557 4110 606
rect 4140 557 4206 606
rect 4236 594 4311 606
rect 4236 557 4302 594
rect 4311 588 4318 594
rect 4318 586 4327 588
rect 4332 585 4398 606
rect 4428 594 4478 606
rect 4425 589 4478 594
rect 4421 586 4424 588
rect 4327 584 4398 585
rect 4419 584 4421 585
rect 4332 557 4398 584
rect 4412 581 4418 584
rect 4428 557 4478 589
rect 4540 557 4590 606
rect 4620 557 4686 606
rect 4716 557 4766 606
rect 4778 594 4794 607
rect 4904 598 4922 610
rect 7343 609 7398 614
rect 7459 610 7464 614
rect 7496 610 7512 615
rect 7514 610 7530 615
rect 7825 610 7829 615
rect 7841 614 7865 629
rect 7869 626 7885 630
rect 7916 626 7925 635
rect 7930 626 7931 635
rect 7935 626 7936 642
rect 7971 641 7973 642
rect 7966 637 7971 641
rect 7946 635 7966 637
rect 8008 635 8011 642
rect 7946 632 7963 635
rect 7934 624 7936 626
rect 7941 627 7963 632
rect 8003 628 8008 635
rect 8056 630 8061 642
rect 8001 627 8003 628
rect 7941 625 7953 627
rect 7916 622 7934 624
rect 7885 620 7920 622
rect 7940 620 7953 625
rect 7841 612 7869 614
rect 7841 611 7883 612
rect 7886 611 7902 620
rect 7903 618 7920 620
rect 7904 614 7920 618
rect 7922 615 7953 620
rect 7984 616 8001 627
rect 8056 626 8059 630
rect 8130 626 8131 630
rect 8248 626 8264 642
rect 8303 630 8314 642
rect 9847 630 9856 644
rect 9926 642 9927 671
rect 10209 663 10211 688
rect 10237 663 10239 690
rect 10300 688 10303 690
rect 10339 687 10340 690
rect 10397 688 10401 690
rect 10479 688 10486 690
rect 10340 678 10346 687
rect 10373 678 10380 687
rect 10389 685 10412 688
rect 10470 687 10479 688
rect 10389 684 10414 685
rect 10389 683 10435 684
rect 10439 683 10441 687
rect 10465 685 10470 687
rect 10462 684 10465 685
rect 10460 683 10462 684
rect 10389 682 10460 683
rect 10497 682 10506 691
rect 10513 690 10520 692
rect 10543 692 10573 696
rect 10543 691 10574 692
rect 10592 691 10594 698
rect 10656 691 10689 700
rect 10772 695 10780 703
rect 10814 693 10836 706
rect 10841 700 10847 706
rect 10887 700 10889 725
rect 10891 713 10901 725
rect 10937 719 10943 725
rect 10964 719 10979 750
rect 10985 749 10986 753
rect 11021 751 11108 758
rect 11136 753 11142 760
rect 11186 758 11206 760
rect 11268 758 11284 774
rect 11286 770 11302 774
rect 11304 771 11311 774
rect 11315 773 11320 774
rect 11304 770 11310 771
rect 11313 770 11315 773
rect 11350 770 11356 774
rect 11286 764 11304 770
rect 11356 764 11362 770
rect 11286 758 11302 764
rect 11364 760 11378 774
rect 11431 761 11439 774
rect 12905 771 12906 781
rect 12934 773 12935 782
rect 13056 774 13122 782
rect 13146 774 13218 783
rect 13225 777 13229 812
rect 13253 803 13262 812
rect 13282 808 13298 823
rect 13300 803 13309 812
rect 13360 808 13376 824
rect 13378 808 13394 824
rect 13425 808 13429 828
rect 13482 825 13492 828
rect 13515 825 13523 846
rect 13572 843 13585 846
rect 13589 842 13591 843
rect 13593 842 13635 851
rect 13591 839 13635 842
rect 13593 835 13635 839
rect 13651 846 13705 851
rect 13710 853 13922 856
rect 13932 855 13936 863
rect 13960 859 14002 864
rect 14031 863 14037 869
rect 14089 863 14095 869
rect 14103 868 14131 870
rect 14231 868 14232 870
rect 14123 867 14141 868
rect 14123 865 14144 867
rect 14204 865 14206 868
rect 14245 865 14251 877
rect 14132 863 14141 865
rect 13931 854 13932 855
rect 13924 853 13937 854
rect 13710 846 13937 853
rect 13651 835 13681 846
rect 13705 845 13937 846
rect 13705 843 13717 845
rect 13732 843 13750 845
rect 13593 830 13681 835
rect 13693 831 13705 843
rect 13839 842 13840 845
rect 13875 840 13881 845
rect 13593 825 13635 830
rect 13645 828 13669 830
rect 13689 828 13693 831
rect 13841 830 13844 838
rect 13882 830 13885 838
rect 13888 830 13894 845
rect 13915 839 13937 845
rect 13976 840 13981 858
rect 14037 857 14043 863
rect 14037 841 14042 857
rect 14079 841 14081 863
rect 14083 857 14089 863
rect 14131 862 14141 863
rect 14132 861 14141 862
rect 14132 859 14147 861
rect 14204 859 14210 865
rect 14251 864 14252 865
rect 14135 856 14160 859
rect 14135 853 14150 856
rect 14152 853 14158 856
rect 14188 854 14197 859
rect 14198 854 14204 859
rect 14234 857 14235 861
rect 14252 859 14254 864
rect 14254 856 14256 859
rect 14141 850 14150 853
rect 14188 850 14207 854
rect 14196 846 14207 850
rect 14207 842 14208 846
rect 14235 842 14238 854
rect 14256 850 14259 856
rect 14331 851 14347 877
rect 14384 868 14386 895
rect 14384 864 14387 868
rect 14416 864 14418 896
rect 14422 889 14430 898
rect 14422 879 14449 889
rect 14496 881 14499 885
rect 14489 879 14496 881
rect 14422 870 14489 879
rect 14424 865 14489 870
rect 14420 864 14424 865
rect 14380 856 14381 861
rect 14379 854 14381 856
rect 14259 845 14263 850
rect 14263 843 14265 845
rect 14347 844 14352 850
rect 14265 842 14266 843
rect 14266 841 14268 842
rect 14037 839 14070 841
rect 13844 828 13845 830
rect 13645 825 13654 828
rect 13480 824 13487 825
rect 13480 814 13490 824
rect 13480 812 13484 814
rect 13487 812 13490 814
rect 13512 813 13514 824
rect 13552 814 13568 824
rect 13545 813 13568 814
rect 13570 813 13593 824
rect 13637 820 13645 825
rect 13649 824 13654 825
rect 13313 803 13314 808
rect 13244 794 13257 803
rect 13309 794 13318 803
rect 13253 787 13257 794
rect 13313 792 13314 794
rect 13344 792 13360 808
rect 13395 807 13410 808
rect 13479 807 13480 811
rect 13488 808 13490 812
rect 13394 802 13410 807
rect 13396 799 13410 802
rect 13429 800 13430 807
rect 13478 804 13479 807
rect 13477 800 13478 803
rect 13490 800 13506 808
rect 13511 807 13512 812
rect 13545 808 13586 813
rect 13536 806 13557 808
rect 13568 807 13574 808
rect 13510 800 13511 806
rect 13536 802 13552 806
rect 13562 802 13568 807
rect 13533 801 13579 802
rect 13533 800 13574 801
rect 13350 790 13356 792
rect 13359 791 13360 792
rect 13387 792 13410 799
rect 13430 797 13432 800
rect 13387 791 13402 792
rect 13358 790 13360 791
rect 13344 787 13360 790
rect 13361 789 13363 790
rect 13396 789 13402 791
rect 13361 787 13402 789
rect 13432 787 13442 797
rect 13474 787 13477 797
rect 13490 792 13510 800
rect 13505 790 13510 792
rect 13533 792 13552 800
rect 13586 792 13602 808
rect 13614 807 13620 813
rect 13627 812 13637 820
rect 13648 813 13654 824
rect 13669 823 13695 828
rect 13659 822 13702 823
rect 13659 821 13700 822
rect 13689 813 13693 821
rect 13702 818 13709 822
rect 13709 816 13710 818
rect 13621 807 13627 812
rect 13648 809 13649 813
rect 13710 812 13713 816
rect 13744 813 13760 824
rect 13762 813 13778 824
rect 13813 816 13822 825
rect 13845 824 13846 828
rect 13802 815 13813 816
rect 13735 812 13737 813
rect 13775 812 13779 813
rect 13688 809 13689 812
rect 13735 810 13779 812
rect 13735 808 13769 810
rect 13620 801 13626 807
rect 13632 792 13648 808
rect 13533 790 13543 792
rect 13545 790 13552 792
rect 13344 785 13399 787
rect 13255 777 13256 785
rect 13317 777 13323 783
rect 13344 781 13367 785
rect 12935 768 12936 771
rect 13072 767 13088 774
rect 13090 767 13106 774
rect 13146 771 13154 774
rect 13158 771 13204 774
rect 13154 767 13157 769
rect 13168 767 13184 771
rect 13186 767 13202 771
rect 11364 758 11381 760
rect 11186 753 11195 758
rect 11203 755 11204 757
rect 11375 753 11381 758
rect 11411 753 11423 761
rect 11431 756 11445 761
rect 11433 753 11445 756
rect 11021 749 11106 751
rect 11131 750 11144 753
rect 10986 746 10987 748
rect 11021 745 11112 749
rect 11124 748 11144 750
rect 11180 748 11186 753
rect 11124 746 11142 748
rect 11179 746 11180 748
rect 11128 745 11142 746
rect 10987 735 10989 744
rect 11040 743 11142 745
rect 11040 740 11072 743
rect 11088 740 11142 743
rect 10989 732 10990 735
rect 10990 730 10991 731
rect 10991 726 10992 730
rect 11040 729 11142 740
rect 11165 732 11167 743
rect 11174 740 11179 746
rect 11204 742 11207 753
rect 11171 736 11174 740
rect 11170 735 11171 736
rect 11168 732 11170 735
rect 11163 730 11168 732
rect 11051 727 11055 729
rect 11092 728 11096 729
rect 11050 725 11055 727
rect 11091 725 11092 727
rect 11153 725 11163 730
rect 10983 719 10989 725
rect 10992 721 10996 724
rect 11049 722 11055 725
rect 11111 724 11163 725
rect 11048 721 11055 722
rect 11089 721 11090 722
rect 11111 721 11153 724
rect 10931 713 10937 719
rect 10989 713 10995 719
rect 10996 717 11095 721
rect 11111 717 11146 721
rect 11165 720 11167 730
rect 11207 724 11208 742
rect 11310 740 11336 753
rect 11339 748 11344 753
rect 11381 748 11384 753
rect 11407 750 11408 752
rect 11439 749 11445 753
rect 11339 747 11345 748
rect 11339 740 11344 747
rect 11384 746 11386 748
rect 11399 746 11407 749
rect 11411 747 11445 749
rect 11442 746 11445 747
rect 11345 740 11346 746
rect 11386 740 11391 746
rect 11392 740 11405 746
rect 11208 719 11211 724
rect 11164 717 11165 719
rect 11298 718 11304 731
rect 11309 724 11310 730
rect 11346 726 11348 740
rect 11310 722 11312 724
rect 11310 721 11314 722
rect 11342 721 11344 724
rect 11310 719 11344 721
rect 11348 719 11350 726
rect 11368 725 11369 727
rect 11391 726 11405 740
rect 11356 722 11362 724
rect 11356 719 11366 722
rect 11392 720 11409 726
rect 11336 718 11366 719
rect 10891 712 10893 713
rect 10891 707 10899 712
rect 10996 707 11137 717
rect 11138 712 11146 717
rect 11304 716 11310 718
rect 11346 717 11356 718
rect 11346 716 11348 717
rect 11217 715 11219 716
rect 11304 715 11348 716
rect 11160 712 11162 715
rect 10893 706 10899 707
rect 10893 700 10905 706
rect 10516 687 10520 690
rect 10518 685 10520 687
rect 10519 683 10520 685
rect 10561 690 10574 691
rect 10561 687 10575 690
rect 10561 683 10583 687
rect 10439 678 10441 682
rect 10303 673 10304 676
rect 10301 668 10304 673
rect 10346 671 10350 678
rect 10380 671 10385 678
rect 10519 677 10523 683
rect 10561 679 10580 683
rect 10583 682 10585 683
rect 10588 682 10592 690
rect 10659 686 10679 691
rect 10653 683 10679 686
rect 10652 682 10679 683
rect 10689 682 10698 691
rect 10814 690 10831 693
rect 10836 691 10837 693
rect 10838 689 10842 690
rect 10893 689 10899 700
rect 10921 698 10930 700
rect 10921 691 10934 698
rect 10830 687 10842 689
rect 10891 688 10899 689
rect 10887 687 10891 688
rect 10830 685 10845 687
rect 10876 685 10887 687
rect 10830 683 10865 685
rect 10869 683 10876 685
rect 10585 681 10592 682
rect 10639 681 10679 682
rect 10585 680 10621 681
rect 10639 680 10651 681
rect 10588 679 10609 680
rect 10630 679 10662 680
rect 10561 678 10658 679
rect 10561 677 10580 678
rect 10452 675 10462 676
rect 10523 675 10524 676
rect 10580 675 10582 676
rect 10465 674 10473 675
rect 10470 671 10484 674
rect 10350 668 10352 671
rect 10294 667 10304 668
rect 10322 667 10333 668
rect 10277 664 10294 667
rect 10266 663 10277 664
rect 10159 662 10277 663
rect 10301 662 10304 667
rect 10333 666 10354 667
rect 10333 664 10356 666
rect 10353 663 10368 664
rect 10388 663 10393 668
rect 10484 667 10486 671
rect 10500 664 10511 667
rect 10495 663 10500 664
rect 10353 662 10500 663
rect 10159 659 10266 662
rect 10159 657 10245 659
rect 10300 657 10301 659
rect 10159 656 10233 657
rect 10159 655 10229 656
rect 10159 654 10222 655
rect 10159 653 10217 654
rect 10159 648 10211 653
rect 10153 642 10217 648
rect 8301 626 8314 630
rect 8129 624 8130 625
rect 8124 619 8129 624
rect 7934 614 7953 615
rect 7903 612 7953 614
rect 7904 611 7953 612
rect 7438 609 7459 610
rect 7841 609 7953 611
rect 7975 610 7984 616
rect 8059 615 8066 619
rect 8122 616 8124 619
rect 8119 615 8122 616
rect 8066 614 8119 615
rect 8072 610 8088 614
rect 8264 610 8280 626
rect 8282 610 8298 626
rect 9017 623 9044 629
rect 9856 626 9860 630
rect 9916 626 9932 642
rect 10159 636 10165 642
rect 10175 638 10181 642
rect 10181 634 10186 638
rect 10205 636 10211 642
rect 10237 634 10239 657
rect 10296 642 10300 657
rect 10356 655 10360 660
rect 10368 659 10495 662
rect 10524 660 10531 675
rect 10581 671 10584 675
rect 10588 674 10592 678
rect 10714 675 10720 677
rect 10692 674 10720 675
rect 10587 672 10588 674
rect 10685 672 10693 674
rect 10714 671 10722 674
rect 10772 671 10778 677
rect 10830 674 10846 683
rect 10570 668 10587 671
rect 10538 664 10552 667
rect 10552 663 10558 664
rect 10565 663 10585 668
rect 10720 665 10726 671
rect 10766 665 10772 671
rect 10674 663 10677 664
rect 10893 663 10899 688
rect 10912 682 10927 691
rect 11040 689 11046 707
rect 11073 706 11088 707
rect 11073 705 11102 706
rect 10552 662 10677 663
rect 10558 660 10674 662
rect 10847 660 10899 663
rect 10565 659 10674 660
rect 10394 657 10483 659
rect 10394 654 10398 657
rect 10411 656 10476 657
rect 10415 655 10473 656
rect 10425 654 10467 655
rect 10360 652 10361 654
rect 10398 652 10399 654
rect 10431 653 10467 654
rect 10361 649 10363 652
rect 10364 642 10369 648
rect 10399 642 10408 652
rect 10441 644 10442 646
rect 10432 642 10447 644
rect 10296 634 10310 642
rect 10408 639 10410 642
rect 10432 639 10448 642
rect 10410 637 10411 639
rect 10432 637 10459 639
rect 10186 632 10253 634
rect 9860 624 9916 626
rect 9045 623 9072 624
rect 9900 610 9916 624
rect 10237 614 10239 632
rect 10244 630 10256 632
rect 10295 630 10310 634
rect 10412 633 10415 637
rect 10432 635 10441 637
rect 10445 635 10490 637
rect 10497 635 10506 644
rect 10244 626 10260 630
rect 10294 626 10310 630
rect 10260 610 10276 626
rect 10278 610 10294 626
rect 10378 615 10395 633
rect 10413 625 10435 633
rect 10441 626 10450 635
rect 10488 626 10497 635
rect 10531 630 10546 659
rect 10568 657 10666 659
rect 10568 655 10574 657
rect 10579 656 10661 657
rect 10581 655 10661 656
rect 10583 652 10655 655
rect 10841 654 10905 660
rect 10562 650 10565 652
rect 10583 651 10642 652
rect 10583 650 10598 651
rect 10608 650 10614 651
rect 10555 645 10561 649
rect 10583 645 10606 650
rect 10617 645 10636 650
rect 10847 648 10853 654
rect 10862 652 10863 654
rect 10863 650 10864 652
rect 10583 644 10603 645
rect 10583 642 10585 644
rect 10587 642 10603 644
rect 10627 642 10636 645
rect 10864 644 10866 649
rect 10893 648 10899 654
rect 10548 639 10552 642
rect 10583 641 10603 642
rect 10583 634 10598 641
rect 10624 635 10636 642
rect 10689 635 10698 644
rect 10893 642 10894 648
rect 10921 645 10927 682
rect 10947 677 10950 683
rect 10983 676 10985 683
rect 10931 667 10937 673
rect 10938 667 10947 676
rect 10937 663 10947 667
rect 10951 663 10953 673
rect 10983 671 10986 676
rect 11035 674 11040 689
rect 10982 667 10986 671
rect 10989 667 10995 673
rect 11073 672 11088 705
rect 11119 704 11123 705
rect 11143 694 11153 705
rect 11219 694 11287 715
rect 11304 712 11322 715
rect 11309 708 11322 712
rect 11350 712 11356 717
rect 11389 715 11391 718
rect 11402 716 11409 720
rect 11409 715 11411 716
rect 11443 715 11445 746
rect 11449 737 11457 749
rect 12904 743 12905 767
rect 12936 742 12939 767
rect 13072 759 13106 767
rect 13158 759 13202 767
rect 13072 758 13088 759
rect 13090 758 13109 759
rect 13168 758 13184 759
rect 13186 758 13202 759
rect 13225 763 13228 777
rect 13230 763 13236 771
rect 13094 753 13109 758
rect 13225 757 13236 763
rect 13165 753 13174 756
rect 13219 754 13236 757
rect 13253 756 13256 777
rect 13201 753 13236 754
rect 13038 740 13236 753
rect 13244 747 13256 756
rect 13322 771 13329 777
rect 13344 774 13365 781
rect 13109 738 13118 740
rect 13124 737 13230 740
rect 13253 738 13262 747
rect 13264 741 13271 747
rect 12939 733 12940 737
rect 11449 715 11457 727
rect 12940 724 12941 731
rect 13202 730 13204 737
rect 13225 730 13231 737
rect 13322 731 13323 771
rect 13350 753 13365 774
rect 13397 778 13398 785
rect 13402 778 13411 787
rect 13397 756 13399 778
rect 13403 775 13411 778
rect 13440 782 13455 787
rect 13472 782 13474 787
rect 13490 782 13510 790
rect 13440 778 13510 782
rect 13536 780 13552 790
rect 13440 774 13515 778
rect 13456 772 13472 774
rect 13474 772 13490 774
rect 13505 772 13515 774
rect 13533 774 13552 780
rect 13586 774 13602 790
rect 13632 780 13648 790
rect 13683 789 13688 808
rect 13718 803 13720 806
rect 13728 805 13744 808
rect 13779 807 13794 808
rect 13804 807 13813 815
rect 13840 810 13856 824
rect 13858 810 13874 824
rect 13885 823 13888 830
rect 13885 818 13890 823
rect 13884 816 13885 818
rect 13888 816 13890 818
rect 13915 816 13931 839
rect 13938 830 13945 838
rect 13981 830 13984 839
rect 14032 835 14043 839
rect 14032 831 14037 835
rect 13945 824 13948 830
rect 13984 828 13985 830
rect 13936 816 13952 824
rect 13880 813 13883 815
rect 13832 808 13875 810
rect 13890 808 13894 816
rect 13913 812 13915 816
rect 13936 812 13957 816
rect 13985 813 13990 828
rect 14023 817 14032 831
rect 14041 828 14043 835
rect 14036 818 14037 828
rect 14023 816 14036 817
rect 14020 815 14023 816
rect 14005 814 14017 815
rect 14003 813 14005 814
rect 13981 812 13995 813
rect 13824 807 13835 808
rect 13849 807 13851 808
rect 13875 807 13894 808
rect 13728 799 13750 805
rect 13728 798 13744 799
rect 13724 792 13744 798
rect 13750 793 13756 799
rect 13724 789 13731 792
rect 13735 789 13744 792
rect 13778 792 13794 807
rect 13802 799 13808 805
rect 13796 793 13802 799
rect 13778 790 13779 792
rect 13683 780 13698 789
rect 13728 788 13744 789
rect 13632 774 13698 780
rect 13723 778 13744 788
rect 13773 787 13775 790
rect 13778 787 13794 790
rect 13767 778 13769 787
rect 13723 776 13769 778
rect 13773 776 13794 787
rect 13811 785 13832 807
rect 13852 803 13853 805
rect 13865 799 13871 804
rect 13854 795 13855 797
rect 13875 795 13890 807
rect 13910 806 13913 812
rect 13936 810 13981 812
rect 13936 808 13957 810
rect 13985 808 13990 812
rect 13894 801 13896 805
rect 13901 795 13910 806
rect 13845 787 13861 795
rect 13875 792 13901 795
rect 13920 792 13936 808
rect 13952 806 13957 808
rect 14029 806 14036 816
rect 14041 809 14042 828
rect 14041 806 14044 809
rect 14073 807 14075 839
rect 14208 836 14210 841
rect 14238 836 14239 841
rect 14268 839 14292 841
rect 14029 805 14037 806
rect 14065 805 14075 807
rect 14079 805 14087 817
rect 14128 815 14144 824
rect 14146 815 14162 824
rect 14128 814 14162 815
rect 14210 814 14212 836
rect 14239 824 14245 836
rect 14270 830 14284 839
rect 14352 836 14354 842
rect 14377 841 14381 854
rect 14376 836 14381 841
rect 14369 834 14381 836
rect 14393 860 14421 861
rect 14393 855 14420 860
rect 14284 825 14288 830
rect 14128 813 14163 814
rect 14126 811 14128 813
rect 14161 812 14162 813
rect 14126 808 14162 811
rect 14224 809 14258 824
rect 14288 815 14292 825
rect 14292 809 14294 814
rect 14354 809 14355 825
rect 14221 808 14258 809
rect 14294 808 14295 809
rect 13957 801 13959 805
rect 13990 800 13992 805
rect 14037 802 14041 805
rect 14041 801 14065 802
rect 14073 801 14075 805
rect 14112 801 14138 808
rect 14148 801 14160 808
rect 13992 797 13993 800
rect 13961 795 13962 797
rect 13889 790 13901 792
rect 13962 791 13965 795
rect 13728 774 13739 776
rect 13774 774 13794 776
rect 13456 766 13521 772
rect 13533 768 13543 774
rect 13545 771 13579 774
rect 13582 771 13586 774
rect 13545 768 13586 771
rect 13456 758 13515 766
rect 13541 764 13543 768
rect 13552 764 13568 768
rect 13396 753 13399 756
rect 13402 753 13405 754
rect 13350 744 13405 753
rect 13463 749 13515 758
rect 13545 758 13568 764
rect 13570 758 13586 768
rect 13648 761 13664 774
rect 13545 756 13557 758
rect 13562 755 13568 758
rect 13620 755 13626 761
rect 13645 758 13664 761
rect 13666 758 13682 774
rect 13744 772 13760 774
rect 13762 772 13778 774
rect 13697 761 13703 767
rect 13735 764 13778 772
rect 13808 768 13812 785
rect 13845 780 13862 787
rect 13832 768 13838 773
rect 13858 772 13862 780
rect 13875 780 13905 790
rect 13875 774 13890 780
rect 13901 779 13905 780
rect 13884 773 13889 774
rect 13862 771 13863 772
rect 13645 755 13651 758
rect 13703 755 13709 761
rect 13744 758 13760 764
rect 13762 758 13778 764
rect 13568 749 13574 755
rect 13614 749 13620 755
rect 13647 754 13651 755
rect 13806 754 13812 768
rect 13854 767 13875 771
rect 13879 767 13884 773
rect 13820 757 13822 758
rect 13819 755 13820 757
rect 13644 750 13648 754
rect 13815 752 13819 755
rect 13854 753 13879 767
rect 13905 763 13916 779
rect 13920 774 13936 790
rect 13965 779 13970 790
rect 13970 776 13978 779
rect 13993 778 14009 797
rect 14041 793 14053 801
rect 14063 793 14075 801
rect 14106 797 14128 801
rect 14152 797 14158 801
rect 14106 795 14160 797
rect 14162 795 14178 808
rect 14208 795 14221 808
rect 14239 806 14245 808
rect 14245 802 14246 806
rect 14071 778 14075 793
rect 14100 789 14128 795
rect 13993 776 14031 778
rect 13970 775 14009 776
rect 13970 774 13986 775
rect 13916 754 13922 763
rect 13936 758 13952 774
rect 13954 763 13978 774
rect 13993 764 14009 775
rect 14016 775 14031 776
rect 14016 774 14032 775
rect 14032 763 14034 774
rect 14071 763 14073 778
rect 13954 758 13970 763
rect 13978 753 13983 763
rect 14009 754 14014 763
rect 14032 758 14037 763
rect 14072 761 14073 763
rect 14106 774 14128 789
rect 14158 792 14178 795
rect 14158 790 14172 792
rect 14158 789 14178 790
rect 14158 781 14160 789
rect 14159 774 14160 781
rect 14162 774 14178 789
rect 14201 784 14211 795
rect 14213 787 14214 795
rect 14246 786 14249 800
rect 14258 792 14274 808
rect 14199 780 14201 784
rect 14214 782 14215 786
rect 14249 781 14250 786
rect 14197 774 14199 780
rect 14250 778 14251 781
rect 14251 774 14253 778
rect 14258 774 14274 790
rect 14295 786 14303 808
rect 14369 806 14376 834
rect 14393 826 14414 855
rect 14368 802 14369 806
rect 14381 803 14390 812
rect 14393 808 14404 826
rect 14430 824 14440 847
rect 14416 818 14450 824
rect 14912 819 14913 1015
rect 15102 819 15103 1015
rect 15188 819 15189 1015
rect 15461 819 15462 1015
rect 15658 819 15659 1015
rect 16256 1012 16257 1015
rect 16315 1013 16316 1016
rect 16312 1012 16316 1013
rect 16556 1014 16572 1016
rect 16600 1015 16612 1016
rect 16574 1014 16596 1015
rect 16608 1014 16612 1015
rect 16556 1012 16617 1014
rect 16648 1012 16868 1021
rect 17039 1017 17050 1021
rect 17039 1014 17057 1017
rect 17060 1014 17125 1030
rect 17039 1012 17125 1014
rect 16246 1005 16252 1011
rect 16255 1008 16256 1012
rect 16254 1005 16255 1008
rect 16292 1005 16298 1011
rect 16240 999 16246 1005
rect 16298 999 16304 1005
rect 16266 990 16267 997
rect 16305 995 16306 1012
rect 16311 1001 16318 1012
rect 16556 1011 16614 1012
rect 16547 1008 16553 1011
rect 16554 1009 16556 1011
rect 16558 1010 16563 1011
rect 16557 1009 16563 1010
rect 16617 1009 16618 1011
rect 16639 1010 16647 1012
rect 17045 1011 17054 1012
rect 17039 1010 17052 1011
rect 17060 1010 17125 1012
rect 16554 1008 16561 1009
rect 16619 1008 16639 1010
rect 16547 1006 16555 1008
rect 16540 1005 16555 1006
rect 16557 1005 16561 1008
rect 16537 1001 16555 1005
rect 16609 1001 16612 1008
rect 16311 998 16312 1001
rect 16310 997 16311 998
rect 16304 990 16306 994
rect 16307 990 16311 997
rect 16519 994 16537 1001
rect 16540 997 16555 1001
rect 16266 989 16283 990
rect 16267 988 16283 989
rect 16252 978 16283 988
rect 16287 978 16318 990
rect 16497 986 16519 994
rect 16540 990 16556 997
rect 16610 996 16611 1000
rect 16615 998 16639 1008
rect 17039 1009 17051 1010
rect 17052 1009 17125 1010
rect 17141 1009 17222 1030
rect 17953 1015 17954 1026
rect 18143 1015 18144 1026
rect 18229 1015 18230 1026
rect 18502 1015 18503 1026
rect 18699 1015 18700 1026
rect 17039 1005 17060 1009
rect 16615 996 16624 998
rect 16610 995 16612 996
rect 16615 995 16619 996
rect 16555 988 16556 990
rect 16478 979 16497 986
rect 16252 972 16318 978
rect 16464 974 16478 979
rect 16213 967 16219 968
rect 15974 965 15976 967
rect 16029 964 16030 967
rect 16206 964 16210 967
rect 16219 964 16226 967
rect 16030 962 16032 964
rect 16193 956 16206 964
rect 16226 963 16231 964
rect 16231 959 16242 963
rect 16268 961 16284 972
rect 16286 966 16306 972
rect 16456 971 16462 973
rect 16540 972 16556 988
rect 16600 992 16615 995
rect 16621 993 16623 996
rect 16600 986 16616 992
rect 16622 988 16623 993
rect 16619 986 16622 988
rect 16765 986 16786 1002
rect 17032 1001 17039 1005
rect 17045 1001 17060 1005
rect 17018 994 17032 1001
rect 17052 998 17060 1001
rect 17078 1005 17088 1009
rect 17222 1005 17239 1009
rect 17078 1003 17091 1005
rect 17060 995 17061 998
rect 16600 985 16624 986
rect 16979 985 16985 991
rect 17003 986 17018 994
rect 17001 985 17003 986
rect 17025 985 17031 991
rect 17061 985 17068 995
rect 16599 983 16600 985
rect 16604 974 16624 985
rect 16799 974 16811 982
rect 16821 974 16833 982
rect 16973 979 16979 985
rect 17031 979 17037 985
rect 17063 980 17071 985
rect 17063 979 17072 980
rect 17063 978 17073 979
rect 17063 975 17075 978
rect 16604 971 16616 974
rect 17063 973 17077 975
rect 17078 973 17079 1003
rect 17084 993 17105 1003
rect 17239 999 17261 1005
rect 17261 997 17263 999
rect 17088 983 17105 993
rect 17263 992 17269 997
rect 17269 986 17273 992
rect 17063 971 17079 973
rect 17084 972 17105 983
rect 17273 982 17276 986
rect 17276 975 17280 982
rect 17084 971 17206 972
rect 17280 971 17282 975
rect 16451 970 16456 971
rect 16448 969 16451 970
rect 16556 968 16574 971
rect 16600 970 16616 971
rect 16793 970 16795 971
rect 16835 970 16872 971
rect 16600 969 16613 970
rect 16348 967 16352 968
rect 16354 967 16359 968
rect 16286 961 16302 966
rect 16340 965 16348 967
rect 16338 964 16340 965
rect 16359 964 16362 967
rect 16440 966 16447 968
rect 16436 964 16440 966
rect 16335 963 16338 964
rect 16334 962 16335 963
rect 16362 962 16365 964
rect 16432 963 16436 964
rect 16254 959 16302 961
rect 16231 958 16246 959
rect 16254 958 16304 959
rect 16327 958 16336 962
rect 16365 959 16369 962
rect 16412 961 16432 963
rect 16234 956 16248 958
rect 16249 957 16304 958
rect 16190 954 16193 956
rect 16234 954 16251 956
rect 16254 954 16304 957
rect 16323 956 16336 958
rect 16369 956 16372 959
rect 16420 958 16426 961
rect 16319 954 16336 956
rect 16372 954 16375 956
rect 16409 954 16417 957
rect 16541 956 16547 959
rect 16556 956 16572 968
rect 16574 967 16581 968
rect 16581 965 16592 967
rect 16600 966 16612 969
rect 16599 965 16612 966
rect 16592 964 16612 965
rect 16632 964 16638 970
rect 16678 966 16684 970
rect 16787 969 16793 970
rect 16668 964 16684 966
rect 16600 962 16612 964
rect 16519 954 16547 956
rect 16030 946 16031 949
rect 16029 945 16068 946
rect 16027 944 16029 945
rect 16012 934 16027 944
rect 16010 933 16012 934
rect 16002 928 16010 933
rect 15993 923 16002 928
rect 15988 920 15993 923
rect 15985 918 15988 920
rect 15981 915 15985 918
rect 15978 913 15981 915
rect 16030 913 16031 945
rect 16068 944 16095 945
rect 16172 944 16190 954
rect 16234 953 16304 954
rect 16234 951 16256 953
rect 16285 951 16286 953
rect 16292 951 16298 953
rect 16312 951 16336 954
rect 16234 948 16336 951
rect 16234 947 16289 948
rect 16292 947 16298 948
rect 16234 946 16268 947
rect 16270 946 16289 947
rect 16301 946 16336 948
rect 16234 944 16289 946
rect 16299 945 16336 946
rect 16298 944 16336 945
rect 16375 952 16398 954
rect 16406 953 16409 954
rect 16403 952 16406 953
rect 16375 948 16403 952
rect 16375 944 16398 948
rect 16095 938 16336 944
rect 16365 938 16380 944
rect 16388 939 16398 944
rect 16394 938 16398 939
rect 16447 938 16537 954
rect 16541 953 16567 954
rect 16599 953 16605 959
rect 16626 958 16690 964
rect 16737 963 16743 969
rect 16783 968 16789 969
rect 16778 966 16789 968
rect 16772 964 16777 966
rect 16768 963 16772 964
rect 16783 963 16789 966
rect 16799 968 16833 970
rect 16837 969 16845 970
rect 16632 954 16684 958
rect 16731 957 16737 963
rect 16789 957 16795 963
rect 16547 947 16553 953
rect 16593 947 16599 953
rect 16632 938 16646 954
rect 16156 922 16172 938
rect 16218 937 16241 938
rect 16218 934 16246 937
rect 16218 933 16254 934
rect 16256 933 16264 935
rect 16285 934 16286 938
rect 16360 937 16365 938
rect 16351 935 16359 936
rect 16287 934 16334 935
rect 16346 934 16351 935
rect 16271 933 16334 934
rect 16398 933 16414 938
rect 16441 936 16447 938
rect 16632 936 16647 938
rect 16437 935 16440 936
rect 16432 933 16436 934
rect 16218 925 16326 933
rect 16285 924 16286 925
rect 16224 922 16241 924
rect 16156 916 16172 920
rect 16207 917 16222 922
rect 16245 920 16270 922
rect 16058 913 16099 916
rect 16103 913 16172 916
rect 15975 911 15978 913
rect 16030 911 16058 913
rect 16156 911 16200 913
rect 16206 911 16222 917
rect 16243 917 16270 920
rect 16289 918 16348 922
rect 16396 920 16432 933
rect 16630 931 16647 936
rect 16626 928 16630 931
rect 16619 924 16626 928
rect 16611 920 16619 924
rect 16632 920 16647 931
rect 16678 920 16680 954
rect 16684 950 16697 954
rect 16799 953 16820 968
rect 16830 967 16833 968
rect 16838 963 16845 969
rect 16873 966 16880 970
rect 17063 969 17077 971
rect 17078 970 17206 971
rect 17088 969 17105 970
rect 17109 969 17206 970
rect 16841 960 16843 963
rect 17059 960 17062 961
rect 16846 954 16853 957
rect 16798 952 16820 953
rect 16798 950 16799 952
rect 16684 942 16692 950
rect 16797 938 16798 949
rect 16853 940 16876 954
rect 16978 953 16979 957
rect 17037 954 17059 960
rect 17063 957 17082 969
rect 17037 952 17064 954
rect 16684 920 16692 932
rect 16391 918 16396 920
rect 16271 917 16348 918
rect 16243 915 16255 917
rect 16315 916 16326 917
rect 16263 914 16275 916
rect 16314 915 16316 916
rect 15971 909 15975 911
rect 16029 910 16031 911
rect 16026 904 16027 906
rect 16030 904 16031 910
rect 16156 904 16172 911
rect 16200 910 16225 911
rect 16191 908 16222 910
rect 16225 909 16236 910
rect 16236 908 16243 909
rect 16181 906 16222 908
rect 16243 907 16256 908
rect 16264 906 16271 907
rect 16191 905 16222 906
rect 16206 904 16222 905
rect 15974 903 15975 904
rect 15965 894 15966 899
rect 16019 896 16020 904
rect 16024 895 16026 903
rect 16018 876 16020 895
rect 16172 888 16188 904
rect 16190 888 16206 904
rect 16283 888 16285 911
rect 16348 909 16364 917
rect 16380 913 16391 918
rect 16375 911 16379 913
rect 16369 909 16375 911
rect 16398 909 16414 920
rect 16598 912 16611 920
rect 16630 918 16684 920
rect 16695 918 16697 926
rect 16734 920 16737 937
rect 16876 935 16885 940
rect 16972 939 16978 952
rect 16982 946 17003 949
rect 17019 946 17020 949
rect 17031 948 17037 952
rect 17048 946 17064 952
rect 16972 936 16979 939
rect 16980 938 16982 946
rect 17003 939 17064 946
rect 17077 942 17082 957
rect 17105 968 17206 969
rect 17283 968 17284 970
rect 17011 938 17064 939
rect 17030 937 17080 938
rect 16797 925 16800 929
rect 16885 928 16896 935
rect 16972 933 16980 936
rect 17030 933 17037 937
rect 16626 912 16696 918
rect 16731 917 16733 919
rect 16800 918 16815 925
rect 16896 923 16900 928
rect 16900 920 16901 923
rect 16815 917 16838 918
rect 16731 916 16737 917
rect 16729 912 16737 916
rect 16596 911 16598 912
rect 16630 911 16645 912
rect 16646 911 16647 912
rect 16348 908 16414 909
rect 16334 907 16414 908
rect 16590 907 16596 911
rect 16630 907 16651 911
rect 16668 908 16684 912
rect 16292 906 16315 907
rect 16348 904 16414 907
rect 16382 888 16398 904
rect 16576 900 16590 907
rect 16630 904 16645 907
rect 16646 904 16647 907
rect 16678 906 16684 908
rect 16687 904 16696 912
rect 16731 911 16737 912
rect 16789 916 16838 917
rect 16789 911 16795 916
rect 16806 914 16838 916
rect 16815 913 16839 914
rect 16815 911 16838 913
rect 16841 911 16866 913
rect 16880 911 16894 920
rect 16901 918 16902 920
rect 16967 918 16972 933
rect 16978 927 16985 933
rect 16978 925 16980 927
rect 16902 911 16905 918
rect 16965 911 16967 915
rect 16726 907 16728 911
rect 16631 900 16644 904
rect 16685 900 16687 904
rect 16722 900 16726 907
rect 16737 905 16743 911
rect 16556 888 16579 900
rect 16626 897 16631 900
rect 16610 888 16626 897
rect 16643 896 16646 899
rect 16680 896 16685 899
rect 16720 897 16722 900
rect 16646 888 16662 896
rect 16664 888 16680 896
rect 16714 888 16720 897
rect 16024 875 16032 888
rect 16220 880 16350 888
rect 16553 883 16556 888
rect 16602 883 16610 888
rect 16711 883 16714 888
rect 16468 880 16516 883
rect 16198 875 16240 880
rect 16018 873 16024 875
rect 16187 873 16240 875
rect 15975 870 15979 873
rect 16008 871 16018 873
rect 16021 872 16024 873
rect 16008 870 16020 871
rect 16168 870 16240 873
rect 16283 870 16285 880
rect 16327 879 16468 880
rect 16330 875 16468 879
rect 16516 875 16517 880
rect 16549 875 16553 883
rect 16588 876 16602 883
rect 16706 876 16711 883
rect 16582 875 16588 876
rect 16749 875 16773 910
rect 16783 905 16789 911
rect 16815 909 16894 911
rect 16905 909 16906 911
rect 16828 904 16894 909
rect 16906 904 16908 908
rect 16844 888 16860 904
rect 16862 893 16878 904
rect 16908 899 16910 903
rect 16910 893 16912 899
rect 16953 898 16965 910
rect 16974 909 16978 925
rect 17011 916 17019 933
rect 17025 927 17031 933
rect 16973 904 16974 909
rect 16991 905 17011 915
rect 16978 903 16990 905
rect 16991 903 17012 905
rect 17030 904 17031 927
rect 17064 922 17080 937
rect 17082 936 17083 941
rect 17105 938 17126 968
rect 17146 965 17206 968
rect 17284 967 17285 968
rect 17285 965 17288 967
rect 17175 963 17206 965
rect 17288 963 17290 965
rect 17184 961 17206 963
rect 17290 961 17294 963
rect 17138 938 17154 954
rect 17156 938 17172 954
rect 17196 949 17224 961
rect 17294 954 17303 961
rect 17182 938 17183 949
rect 17224 947 17228 949
rect 17303 947 17311 954
rect 17228 946 17229 947
rect 17229 944 17230 946
rect 17311 944 17313 947
rect 17499 944 17500 949
rect 17528 944 17544 954
rect 17230 939 17236 944
rect 17313 940 17318 944
rect 17482 940 17549 944
rect 17318 939 17320 940
rect 17459 939 17482 940
rect 17105 936 17138 938
rect 17143 936 17188 938
rect 17236 936 17238 938
rect 17320 936 17323 939
rect 17456 936 17459 939
rect 17499 938 17500 940
rect 17549 938 17550 939
rect 17083 916 17088 933
rect 17105 922 17137 936
rect 17174 934 17188 936
rect 17238 934 17240 936
rect 17323 934 17327 936
rect 17453 934 17456 936
rect 17168 932 17188 934
rect 17240 932 17241 934
rect 17327 932 17329 934
rect 17452 932 17453 934
rect 17089 915 17095 921
rect 17105 919 17126 922
rect 17130 921 17137 922
rect 17126 915 17129 919
rect 17130 915 17141 921
rect 17083 909 17089 915
rect 17088 908 17089 909
rect 17130 906 17137 915
rect 17141 909 17147 915
rect 17179 904 17215 932
rect 17241 925 17248 932
rect 17329 925 17340 932
rect 17449 925 17452 932
rect 17248 924 17262 925
rect 17240 915 17262 924
rect 17340 919 17349 925
rect 17446 919 17449 925
rect 17349 916 17352 919
rect 17445 916 17446 919
rect 17248 907 17262 915
rect 17352 912 17357 916
rect 17443 912 17445 916
rect 17357 907 17361 912
rect 17440 910 17443 912
rect 17256 905 17265 907
rect 17262 904 17265 905
rect 17361 904 17363 907
rect 16975 901 17015 903
rect 16972 900 16973 901
rect 16971 899 16972 900
rect 16975 899 17011 901
rect 16970 898 16975 899
rect 16953 896 16975 898
rect 16913 893 16965 896
rect 16970 893 16975 896
rect 16862 888 16881 893
rect 16912 888 16965 893
rect 16809 877 16818 881
rect 16856 877 16865 881
rect 16875 879 16881 888
rect 16907 886 16921 888
rect 16902 883 16907 886
rect 16912 883 16921 886
rect 16901 882 16921 883
rect 16893 880 16921 882
rect 16890 879 16921 880
rect 16875 877 16921 879
rect 16801 875 16921 877
rect 16330 870 16432 875
rect 16470 874 16624 875
rect 16470 872 16617 874
rect 16443 871 16470 872
rect 16435 870 16443 871
rect 15979 869 16008 870
rect 16016 867 16020 870
rect 16164 869 16168 870
rect 16430 869 16435 870
rect 16015 866 16020 867
rect 16151 866 16164 869
rect 16421 868 16430 869
rect 16413 866 16421 868
rect 16517 867 16520 872
rect 16549 871 16553 872
rect 16582 871 16588 872
rect 16624 871 16638 874
rect 16704 871 16706 875
rect 16720 872 16801 875
rect 16809 872 16921 875
rect 16953 872 16965 888
rect 16966 881 16971 893
rect 16970 880 16971 881
rect 16638 870 16642 871
rect 15963 859 15964 866
rect 16013 864 16020 866
rect 16129 865 16163 866
rect 16408 865 16413 866
rect 16013 859 16015 864
rect 16129 862 16151 865
rect 16128 859 16151 862
rect 16163 859 16170 865
rect 16375 859 16408 865
rect 16012 855 16013 859
rect 16124 855 16129 859
rect 16132 854 16151 859
rect 16170 857 16173 859
rect 16369 858 16375 859
rect 16362 857 16369 858
rect 16346 854 16361 857
rect 16520 854 16525 866
rect 16547 863 16549 870
rect 16579 863 16582 870
rect 16642 868 16654 870
rect 16546 860 16547 863
rect 16578 860 16579 863
rect 16654 859 16692 868
rect 16697 863 16702 870
rect 16720 868 16809 872
rect 16810 870 16921 872
rect 16991 871 17011 899
rect 17015 893 17019 901
rect 17019 873 17024 893
rect 17127 887 17130 904
rect 17187 903 17190 904
rect 17183 902 17187 903
rect 17182 899 17183 901
rect 17215 899 17222 904
rect 17175 887 17182 899
rect 17187 897 17188 899
rect 17221 893 17222 899
rect 17257 893 17264 898
rect 17265 893 17280 904
rect 17130 877 17155 887
rect 17181 877 17182 887
rect 17264 885 17276 893
rect 17280 887 17289 893
rect 17363 887 17376 904
rect 17436 902 17448 910
rect 17458 902 17470 910
rect 17510 904 17511 938
rect 17549 934 17560 938
rect 17550 922 17560 934
rect 17550 903 17551 922
rect 17436 898 17439 902
rect 17472 899 17474 902
rect 17424 886 17432 898
rect 17436 896 17470 898
rect 17436 895 17439 896
rect 17155 870 17182 877
rect 17276 876 17283 885
rect 17289 879 17295 886
rect 17376 879 17381 886
rect 17295 877 17297 879
rect 17381 877 17383 879
rect 17187 870 17188 872
rect 16718 866 16720 868
rect 16715 864 16718 866
rect 16745 864 16748 868
rect 16695 860 16697 863
rect 16011 851 16012 854
rect 16122 851 16124 854
rect 16131 850 16132 854
rect 15962 838 15963 845
rect 16007 838 16011 850
rect 16115 838 16122 850
rect 14416 812 14432 818
rect 14434 812 14450 818
rect 15961 816 15962 837
rect 16000 816 16007 838
rect 16115 835 16121 838
rect 16109 829 16115 835
rect 16123 828 16128 842
rect 16161 835 16167 841
rect 16173 839 16174 854
rect 16250 850 16346 854
rect 16525 850 16526 854
rect 16544 853 16546 859
rect 16575 853 16578 859
rect 16687 858 16697 859
rect 16687 853 16694 858
rect 16697 857 16703 858
rect 16712 857 16715 864
rect 16800 863 16809 868
rect 16865 863 16874 870
rect 16883 868 16884 870
rect 16921 868 16922 870
rect 16743 860 16745 863
rect 16884 861 16886 868
rect 16922 860 16925 868
rect 16951 864 16952 866
rect 16950 861 16951 863
rect 16966 859 16972 870
rect 16988 864 16991 870
rect 17024 866 17026 870
rect 17063 868 17064 869
rect 17061 865 17063 868
rect 17054 864 17061 865
rect 16978 859 16980 861
rect 16703 855 16726 857
rect 16741 856 16743 859
rect 16802 856 16808 857
rect 16848 856 16854 857
rect 16887 856 16888 857
rect 16926 856 16927 857
rect 16948 856 16949 859
rect 16974 856 16982 859
rect 16703 854 16716 855
rect 16736 854 16741 856
rect 16687 852 16690 853
rect 16687 851 16689 852
rect 16711 851 16712 854
rect 16716 851 16757 854
rect 16190 843 16251 850
rect 16189 841 16190 842
rect 16167 832 16173 835
rect 16174 832 16175 838
rect 16167 829 16175 832
rect 16183 829 16189 841
rect 16193 840 16204 842
rect 16250 840 16251 843
rect 16261 843 16451 850
rect 16526 846 16529 850
rect 16536 846 16544 851
rect 16567 847 16575 851
rect 16562 846 16623 847
rect 16473 843 16555 846
rect 16261 839 16346 843
rect 16439 842 16457 843
rect 16526 842 16529 843
rect 16421 839 16439 842
rect 16457 841 16469 842
rect 16472 839 16475 841
rect 16259 838 16261 839
rect 16254 835 16258 838
rect 16248 830 16254 835
rect 16281 831 16283 839
rect 16413 838 16421 839
rect 16397 835 16413 838
rect 16171 828 16175 829
rect 16247 828 16248 830
rect 14416 809 14450 812
rect 15960 811 15961 816
rect 15999 811 16000 816
rect 16028 811 16044 824
rect 16122 813 16123 828
rect 16167 826 16169 827
rect 16171 826 16183 828
rect 16169 816 16191 826
rect 16220 817 16236 824
rect 16167 812 16191 816
rect 16210 812 16236 817
rect 16167 811 16169 812
rect 14416 808 14462 809
rect 14365 790 14368 800
rect 14372 794 14381 803
rect 14393 792 14416 808
rect 14428 803 14437 808
rect 14462 805 14467 808
rect 15997 807 15999 810
rect 16173 808 16183 812
rect 14437 794 14446 803
rect 14355 787 14370 790
rect 14303 779 14309 786
rect 14328 780 14370 787
rect 14376 786 14380 792
rect 14393 790 14403 792
rect 14393 787 14416 790
rect 14372 780 14374 784
rect 14393 781 14430 787
rect 14304 774 14320 779
rect 14328 774 14372 780
rect 14400 774 14430 781
rect 14467 774 14483 805
rect 15959 800 15960 805
rect 15994 800 15996 805
rect 15993 798 15994 800
rect 15989 790 15993 798
rect 16012 792 16023 808
rect 16172 806 16173 808
rect 16191 807 16200 812
rect 16208 809 16236 812
rect 16206 808 16217 809
rect 16220 808 16236 809
rect 16238 808 16254 824
rect 16277 818 16283 831
rect 16363 830 16397 835
rect 16321 823 16363 830
rect 16475 829 16477 839
rect 16529 829 16534 842
rect 16536 828 16544 843
rect 16313 822 16321 823
rect 16288 818 16313 822
rect 16277 816 16288 818
rect 16273 812 16283 816
rect 16204 807 16220 808
rect 16200 806 16220 807
rect 16200 805 16217 806
rect 16254 805 16270 808
rect 16122 790 16123 805
rect 15987 786 15989 790
rect 16108 787 16123 790
rect 16161 789 16172 805
rect 16198 803 16231 805
rect 16198 794 16226 803
rect 16248 797 16270 805
rect 16198 793 16220 794
rect 16204 792 16220 793
rect 16210 790 16220 792
rect 16244 792 16270 797
rect 16244 791 16254 792
rect 16161 787 16173 789
rect 15958 782 15959 786
rect 16108 783 16173 787
rect 16204 787 16220 790
rect 16237 790 16254 791
rect 16237 787 16270 790
rect 16204 783 16270 787
rect 16108 782 16172 783
rect 14106 761 14162 774
rect 14164 763 14172 774
rect 14194 763 14197 774
rect 14215 764 14216 770
rect 14034 753 14037 758
rect 14073 758 14162 761
rect 14193 760 14196 763
rect 14247 760 14258 774
rect 13463 745 13522 749
rect 13644 746 13651 750
rect 13805 748 13815 752
rect 13852 749 13854 753
rect 13683 746 13780 748
rect 13803 746 13815 748
rect 13851 746 13852 748
rect 13643 745 13651 746
rect 13654 745 13789 746
rect 13800 745 13802 746
rect 13805 745 13815 746
rect 13350 741 13402 744
rect 13405 742 13406 744
rect 13344 736 13408 741
rect 13463 740 13602 745
rect 13643 744 13815 745
rect 13344 735 13410 736
rect 13265 730 13271 731
rect 13186 727 13288 730
rect 13186 724 13313 727
rect 13322 725 13329 731
rect 13350 729 13356 735
rect 13365 727 13368 732
rect 13396 729 13402 735
rect 13407 727 13410 735
rect 13369 725 13370 727
rect 13410 725 13411 727
rect 13463 726 13471 740
rect 13515 736 13602 740
rect 13517 730 13602 736
rect 13635 743 13815 744
rect 13847 743 13851 745
rect 13861 744 13879 753
rect 13983 750 13985 753
rect 14014 750 14016 753
rect 13884 744 13924 745
rect 13925 744 13936 750
rect 13635 740 13812 743
rect 13635 732 13649 740
rect 13847 735 13861 743
rect 13524 729 13525 730
rect 13525 727 13526 729
rect 11350 709 11351 712
rect 11310 707 11322 708
rect 11351 702 11352 703
rect 11310 698 11311 701
rect 11372 696 11389 714
rect 12902 713 12903 724
rect 12941 717 12942 724
rect 13186 720 13235 724
rect 13186 717 13242 720
rect 13271 719 13277 724
rect 13186 716 13194 717
rect 13186 715 13193 716
rect 11446 711 11449 713
rect 12942 711 12943 713
rect 13205 712 13207 717
rect 11439 710 11446 711
rect 13235 710 13242 717
rect 11433 708 11445 710
rect 11422 703 11445 708
rect 12901 707 12902 710
rect 13086 707 13169 710
rect 11422 696 11433 703
rect 13207 696 13210 709
rect 13242 708 13252 709
rect 13220 700 13232 708
rect 13242 700 13254 708
rect 13211 698 13216 700
rect 13218 698 13263 700
rect 13211 697 13263 698
rect 13289 697 13291 722
rect 13317 719 13323 725
rect 13370 723 13371 725
rect 13411 720 13412 722
rect 13457 720 13473 726
rect 13373 715 13375 719
rect 13412 716 13413 719
rect 13459 716 13473 720
rect 13477 716 13480 719
rect 13503 718 13505 726
rect 13515 720 13521 726
rect 13602 725 13611 730
rect 13527 723 13528 725
rect 13502 716 13505 718
rect 13509 716 13517 720
rect 13375 709 13379 715
rect 13413 710 13415 715
rect 13459 714 13469 716
rect 13459 713 13468 714
rect 13471 713 13492 716
rect 13502 713 13504 716
rect 13507 713 13517 716
rect 13468 710 13469 713
rect 13480 710 13483 713
rect 13496 712 13500 713
rect 13500 711 13505 712
rect 13507 711 13509 713
rect 13492 710 13507 711
rect 13528 710 13535 722
rect 13611 713 13616 724
rect 13643 722 13649 732
rect 13772 723 13778 729
rect 13788 727 13794 732
rect 13783 723 13788 727
rect 13818 723 13824 729
rect 13844 727 13847 735
rect 13848 727 13861 735
rect 13844 725 13848 727
rect 13869 726 13877 744
rect 13884 740 13936 744
rect 13882 735 13918 740
rect 13924 737 13936 740
rect 13985 747 13988 750
rect 13924 735 13941 737
rect 13882 731 13884 735
rect 13925 734 13941 735
rect 13985 734 13990 747
rect 13935 731 13941 734
rect 13936 730 13941 731
rect 13939 729 13943 730
rect 13988 729 13990 734
rect 13941 726 13945 729
rect 13635 719 13649 722
rect 13635 716 13651 719
rect 13703 716 13704 719
rect 13766 717 13772 723
rect 13824 717 13830 723
rect 13840 722 13844 724
rect 13845 723 13848 725
rect 13871 724 13872 726
rect 13943 725 13945 726
rect 13989 725 13990 729
rect 13877 724 13878 725
rect 13380 698 13386 708
rect 13416 698 13418 708
rect 13471 701 13483 710
rect 13484 698 13490 708
rect 13493 701 13505 710
rect 13507 709 13572 710
rect 13514 707 13572 709
rect 13521 706 13572 707
rect 13529 703 13572 706
rect 13535 700 13541 703
rect 13543 702 13572 703
rect 13544 701 13572 702
rect 13535 698 13549 700
rect 13386 697 13390 698
rect 13211 696 13390 697
rect 11352 695 11353 696
rect 11366 694 11384 696
rect 11134 690 11145 691
rect 11134 688 11143 690
rect 11134 687 11144 688
rect 11147 687 11148 690
rect 11150 688 11159 691
rect 11180 690 11182 691
rect 11287 688 11307 694
rect 11311 691 11312 692
rect 11343 690 11384 694
rect 12900 692 12901 696
rect 13207 695 13216 696
rect 13208 694 13216 695
rect 13220 694 13390 696
rect 13418 694 13422 698
rect 12905 690 12906 692
rect 11312 688 11314 690
rect 11343 688 11366 690
rect 11280 687 11374 688
rect 11131 685 11144 687
rect 11128 683 11131 685
rect 11117 677 11128 683
rect 11134 679 11142 685
rect 11033 667 11035 671
rect 10982 663 10989 667
rect 10937 661 10989 663
rect 10938 660 10997 661
rect 10921 644 10929 645
rect 10896 642 10903 643
rect 10867 637 10869 641
rect 10893 637 10903 642
rect 10912 642 10929 644
rect 10937 642 10938 659
rect 10939 649 10997 660
rect 11030 655 11033 667
rect 11029 652 11030 654
rect 11066 652 11073 672
rect 11113 668 11117 676
rect 11134 663 11142 669
rect 11146 663 11148 687
rect 11312 676 11314 687
rect 11353 682 11355 687
rect 11396 676 11406 680
rect 12903 676 12906 690
rect 11216 672 11236 673
rect 11200 664 11216 672
rect 11236 664 11288 672
rect 11196 663 11200 664
rect 11134 662 11200 663
rect 11288 663 11302 664
rect 11314 663 11316 676
rect 11390 674 11396 676
rect 11359 664 11390 674
rect 12900 670 12903 676
rect 11350 663 11359 664
rect 11288 662 11359 663
rect 10947 648 10989 649
rect 10947 645 10987 648
rect 10893 635 10900 637
rect 10912 635 10938 642
rect 10951 637 10963 645
rect 10973 644 10985 645
rect 10986 644 10987 645
rect 10973 642 10987 644
rect 11026 643 11028 647
rect 11064 645 11066 651
rect 11063 643 11064 645
rect 11111 642 11113 659
rect 11134 657 11195 662
rect 11302 661 11359 662
rect 12893 663 12903 670
rect 12905 663 12906 676
rect 12938 687 12939 692
rect 12940 687 12965 692
rect 13205 688 13211 694
rect 12938 673 12969 687
rect 13208 684 13211 688
rect 13220 692 13316 694
rect 13220 690 13348 692
rect 13386 691 13445 694
rect 13386 690 13390 691
rect 13418 690 13422 691
rect 13445 690 13449 691
rect 13490 690 13491 696
rect 13541 695 13549 698
rect 13551 697 13572 701
rect 13613 709 13617 713
rect 13635 712 13653 716
rect 13678 712 13681 713
rect 13635 711 13651 712
rect 13635 710 13649 711
rect 13656 710 13681 712
rect 13696 710 13698 712
rect 13703 710 13709 715
rect 13757 710 13772 716
rect 13839 715 13844 722
rect 13832 711 13838 714
rect 13840 711 13844 715
rect 13866 716 13883 724
rect 13643 709 13651 710
rect 13654 709 13657 710
rect 13662 709 13764 710
rect 13613 706 13619 709
rect 13643 707 13649 709
rect 13684 707 13764 709
rect 13646 706 13764 707
rect 13832 709 13840 711
rect 13832 706 13838 709
rect 13866 708 13888 716
rect 13880 706 13888 708
rect 13899 706 13905 712
rect 13613 702 13620 706
rect 13613 701 13621 702
rect 13584 698 13594 699
rect 13613 698 13623 701
rect 13646 698 13659 706
rect 13697 703 13703 706
rect 13708 705 13777 706
rect 13824 705 13832 706
rect 13708 703 13832 705
rect 13708 700 13745 703
rect 13577 697 13581 698
rect 13595 697 13623 698
rect 13559 695 13577 697
rect 13535 694 13577 695
rect 13541 692 13572 694
rect 13541 691 13560 692
rect 13538 690 13546 691
rect 13220 688 13269 690
rect 13220 683 13254 688
rect 13220 682 13228 683
rect 13220 681 13227 682
rect 13120 673 13154 676
rect 12938 663 12939 673
rect 12944 663 12951 670
rect 11314 660 11316 661
rect 12893 658 12951 663
rect 12968 660 12969 673
rect 11142 656 11195 657
rect 12899 657 12944 658
rect 11142 655 11184 656
rect 11144 653 11182 655
rect 12899 653 12900 657
rect 12903 654 12941 657
rect 11146 645 11158 653
rect 11168 645 11180 653
rect 12905 646 12917 654
rect 12927 646 12939 654
rect 10973 641 10986 642
rect 10970 639 10986 641
rect 10973 637 10986 639
rect 10975 636 10986 637
rect 10965 635 10971 636
rect 10977 635 10986 636
rect 10530 626 10548 630
rect 10561 626 10598 634
rect 10633 626 10642 635
rect 10680 626 10689 635
rect 10870 630 10877 634
rect 10869 626 10877 630
rect 10530 625 10536 626
rect 10413 621 10428 625
rect 10525 621 10530 625
rect 10413 618 10435 621
rect 10521 618 10525 621
rect 10413 615 10436 618
rect 10517 615 10521 618
rect 10548 615 10585 626
rect 10870 615 10877 626
rect 10893 629 10903 635
rect 10921 630 10938 635
rect 10395 614 10436 615
rect 7343 607 7473 609
rect 7343 606 7363 607
rect 7483 606 7502 609
rect 7830 607 7953 609
rect 4789 593 4792 594
rect 4794 589 4800 594
rect 4800 586 4803 588
rect 4883 586 4904 598
rect 4905 596 4916 598
rect 4803 585 4807 586
rect 4807 584 4854 585
rect 4874 584 4879 585
rect 4924 557 4974 606
rect 5004 557 5070 606
rect 5100 557 5166 606
rect 5196 557 5262 606
rect 5292 557 5342 606
rect 6824 557 6874 606
rect 6904 557 6970 606
rect 7000 557 7066 606
rect 7096 557 7162 606
rect 7192 557 7258 606
rect 7288 594 7363 606
rect 7288 557 7354 594
rect 7363 588 7370 594
rect 7370 586 7379 588
rect 7384 585 7450 606
rect 7480 594 7530 606
rect 7477 589 7530 594
rect 7473 586 7476 588
rect 7379 584 7450 585
rect 7471 584 7473 585
rect 7384 557 7450 584
rect 7464 581 7470 584
rect 7480 557 7530 589
rect 7592 557 7642 606
rect 7672 557 7738 606
rect 7768 557 7818 606
rect 7830 594 7846 607
rect 7956 598 7974 610
rect 10395 609 10450 614
rect 10511 610 10516 614
rect 10548 610 10564 615
rect 10566 610 10582 615
rect 10877 610 10881 615
rect 10893 614 10917 629
rect 10921 626 10937 630
rect 10968 626 10977 635
rect 10982 626 10983 635
rect 10987 626 10988 642
rect 11023 641 11025 642
rect 11018 637 11023 641
rect 10998 635 11018 637
rect 11060 635 11063 642
rect 10998 632 11015 635
rect 10986 624 10988 626
rect 10993 627 11015 632
rect 11055 628 11060 635
rect 11108 630 11113 642
rect 11053 627 11055 628
rect 10993 625 11005 627
rect 10968 622 10986 624
rect 10937 620 10972 622
rect 10992 620 11005 625
rect 10893 612 10921 614
rect 10893 611 10935 612
rect 10938 611 10954 620
rect 10955 618 10972 620
rect 10956 614 10972 618
rect 10974 615 11005 620
rect 11036 616 11053 627
rect 11108 626 11111 630
rect 11182 626 11183 630
rect 11300 626 11316 642
rect 11355 630 11366 642
rect 12899 630 12908 644
rect 12978 642 12979 671
rect 13261 663 13263 688
rect 13289 663 13291 690
rect 13352 688 13355 690
rect 13391 687 13392 690
rect 13449 688 13453 690
rect 13531 688 13538 690
rect 13392 678 13398 687
rect 13425 678 13432 687
rect 13441 685 13464 688
rect 13522 687 13531 688
rect 13441 684 13466 685
rect 13441 683 13487 684
rect 13491 683 13493 687
rect 13517 685 13522 687
rect 13514 684 13517 685
rect 13512 683 13514 684
rect 13441 682 13512 683
rect 13549 682 13558 691
rect 13565 690 13572 692
rect 13595 691 13626 697
rect 13644 691 13646 698
rect 13708 691 13741 700
rect 13824 695 13832 703
rect 13866 693 13888 706
rect 13893 700 13899 706
rect 13939 700 13941 725
rect 13943 713 13953 725
rect 13989 719 13995 725
rect 14016 719 14031 750
rect 14037 749 14038 753
rect 14073 751 14160 758
rect 14188 753 14194 760
rect 14238 758 14258 760
rect 14320 758 14336 774
rect 14338 770 14354 774
rect 14356 771 14363 774
rect 14367 773 14372 774
rect 14356 770 14362 771
rect 14365 770 14367 773
rect 14402 770 14408 774
rect 14338 764 14356 770
rect 14408 764 14414 770
rect 14338 758 14354 764
rect 14416 760 14430 774
rect 14483 761 14491 774
rect 15957 771 15958 777
rect 15986 773 15987 782
rect 16108 774 16174 782
rect 16198 774 16270 783
rect 16277 777 16281 812
rect 16305 803 16314 812
rect 16334 808 16350 823
rect 16352 803 16361 812
rect 16412 808 16428 824
rect 16430 808 16446 824
rect 16477 808 16481 828
rect 16534 825 16544 828
rect 16567 825 16575 846
rect 16624 843 16637 846
rect 16641 842 16643 843
rect 16645 842 16687 851
rect 16643 839 16687 842
rect 16645 835 16687 839
rect 16703 846 16757 851
rect 16762 853 16974 856
rect 16984 855 16988 863
rect 17012 859 17054 864
rect 17083 863 17089 869
rect 17141 863 17147 869
rect 17155 868 17183 870
rect 17283 868 17284 870
rect 17175 867 17193 868
rect 17175 865 17196 867
rect 17256 865 17258 868
rect 17297 865 17303 877
rect 17184 863 17193 865
rect 16983 854 16984 855
rect 16976 853 16989 854
rect 16762 846 16989 853
rect 16703 835 16733 846
rect 16757 845 16989 846
rect 16757 843 16769 845
rect 16784 843 16802 845
rect 16645 830 16733 835
rect 16745 831 16757 843
rect 16891 842 16892 845
rect 16927 840 16933 845
rect 16645 825 16687 830
rect 16697 828 16721 830
rect 16741 828 16745 831
rect 16893 830 16896 838
rect 16934 830 16937 838
rect 16940 830 16946 845
rect 16967 839 16989 845
rect 17028 840 17033 858
rect 17089 857 17095 863
rect 17089 841 17094 857
rect 17131 841 17133 863
rect 17135 857 17141 863
rect 17183 862 17193 863
rect 17184 861 17193 862
rect 17184 859 17199 861
rect 17256 859 17262 865
rect 17303 864 17304 865
rect 17187 856 17212 859
rect 17187 853 17202 856
rect 17204 853 17210 856
rect 17240 854 17249 859
rect 17250 854 17256 859
rect 17286 857 17287 861
rect 17304 859 17306 864
rect 17306 856 17308 859
rect 17193 850 17202 853
rect 17240 850 17259 854
rect 17248 846 17259 850
rect 17259 842 17260 846
rect 17287 842 17290 854
rect 17308 850 17311 856
rect 17383 851 17399 877
rect 17436 868 17438 895
rect 17436 864 17439 868
rect 17468 864 17470 896
rect 17474 889 17482 898
rect 17474 879 17501 889
rect 17548 881 17551 885
rect 17541 879 17548 881
rect 17474 870 17541 879
rect 17476 865 17541 870
rect 17472 864 17476 865
rect 17432 856 17433 861
rect 17431 854 17433 856
rect 17311 845 17315 850
rect 17315 843 17317 845
rect 17399 844 17404 850
rect 17317 842 17318 843
rect 17318 841 17320 842
rect 17089 839 17122 841
rect 16896 828 16897 830
rect 16697 825 16706 828
rect 16532 824 16539 825
rect 16532 814 16542 824
rect 16532 812 16536 814
rect 16539 812 16542 814
rect 16564 813 16566 824
rect 16604 814 16620 824
rect 16597 813 16620 814
rect 16622 813 16645 824
rect 16689 820 16697 825
rect 16701 824 16706 825
rect 16365 803 16366 808
rect 16296 794 16309 803
rect 16361 794 16370 803
rect 16305 787 16309 794
rect 16365 792 16366 794
rect 16396 792 16412 808
rect 16447 807 16462 808
rect 16531 807 16532 811
rect 16540 808 16542 812
rect 16446 802 16462 807
rect 16448 799 16462 802
rect 16481 800 16482 807
rect 16530 804 16531 807
rect 16529 800 16530 803
rect 16542 800 16558 808
rect 16563 807 16564 812
rect 16597 808 16638 813
rect 16588 806 16609 808
rect 16620 807 16626 808
rect 16562 800 16563 806
rect 16588 802 16604 806
rect 16614 802 16620 807
rect 16585 801 16631 802
rect 16585 800 16626 801
rect 16402 790 16408 792
rect 16411 791 16412 792
rect 16439 792 16462 799
rect 16482 797 16484 800
rect 16439 791 16454 792
rect 16410 790 16412 791
rect 16396 787 16412 790
rect 16413 789 16415 790
rect 16448 789 16454 791
rect 16413 787 16454 789
rect 16484 787 16494 797
rect 16526 787 16529 797
rect 16542 792 16562 800
rect 16557 790 16562 792
rect 16585 792 16604 800
rect 16638 792 16654 808
rect 16666 807 16672 813
rect 16679 812 16689 820
rect 16700 813 16706 824
rect 16721 823 16747 828
rect 16711 822 16754 823
rect 16711 821 16752 822
rect 16741 813 16745 821
rect 16754 818 16761 822
rect 16761 816 16762 818
rect 16673 807 16679 812
rect 16700 809 16701 813
rect 16762 812 16765 816
rect 16796 813 16812 824
rect 16814 813 16830 824
rect 16865 816 16874 825
rect 16897 824 16898 828
rect 16854 815 16865 816
rect 16787 812 16789 813
rect 16827 812 16831 813
rect 16740 809 16741 812
rect 16787 810 16831 812
rect 16787 808 16821 810
rect 16672 801 16678 807
rect 16684 792 16700 808
rect 16585 790 16595 792
rect 16597 790 16604 792
rect 16396 785 16451 787
rect 16307 777 16308 785
rect 16369 777 16375 783
rect 16396 781 16419 785
rect 15987 768 15988 771
rect 16124 767 16140 774
rect 16142 767 16158 774
rect 16198 771 16206 774
rect 16210 771 16256 774
rect 16206 767 16209 769
rect 16220 767 16236 771
rect 16238 767 16254 771
rect 14416 758 14433 760
rect 14238 753 14247 758
rect 14255 755 14256 757
rect 14427 753 14433 758
rect 14463 753 14475 761
rect 14483 756 14497 761
rect 14485 753 14497 756
rect 14073 749 14158 751
rect 14183 750 14196 753
rect 14038 746 14039 748
rect 14073 745 14164 749
rect 14176 748 14196 750
rect 14232 748 14238 753
rect 14176 746 14194 748
rect 14231 746 14232 748
rect 14180 745 14194 746
rect 14039 735 14041 744
rect 14092 743 14194 745
rect 14092 740 14124 743
rect 14140 740 14194 743
rect 14041 732 14042 735
rect 14042 730 14043 731
rect 14043 726 14044 730
rect 14092 729 14194 740
rect 14217 732 14219 743
rect 14226 740 14231 746
rect 14256 742 14259 753
rect 14223 736 14226 740
rect 14222 735 14223 736
rect 14220 732 14222 735
rect 14215 730 14220 732
rect 14103 727 14107 729
rect 14144 728 14148 729
rect 14102 725 14107 727
rect 14143 725 14144 727
rect 14205 725 14215 730
rect 14035 719 14041 725
rect 14044 721 14048 724
rect 14101 722 14107 725
rect 14163 724 14215 725
rect 14100 721 14107 722
rect 14141 721 14142 722
rect 14163 721 14205 724
rect 13983 713 13989 719
rect 14041 713 14047 719
rect 14048 717 14147 721
rect 14163 717 14198 721
rect 14217 720 14219 730
rect 14259 724 14260 742
rect 14362 740 14388 753
rect 14391 748 14396 753
rect 14433 748 14436 753
rect 14459 750 14460 752
rect 14491 749 14497 753
rect 14391 747 14397 748
rect 14391 740 14396 747
rect 14436 746 14438 748
rect 14451 746 14459 749
rect 14463 747 14497 749
rect 14494 746 14497 747
rect 14397 740 14398 746
rect 14438 740 14443 746
rect 14444 740 14457 746
rect 14260 719 14263 724
rect 14216 717 14217 719
rect 14350 718 14356 731
rect 14361 724 14362 730
rect 14398 726 14400 740
rect 14362 722 14364 724
rect 14362 721 14366 722
rect 14394 721 14396 724
rect 14362 719 14396 721
rect 14400 719 14402 726
rect 14420 725 14421 727
rect 14443 726 14457 740
rect 14408 722 14414 724
rect 14408 719 14418 722
rect 14444 720 14461 726
rect 14388 718 14418 719
rect 13943 712 13945 713
rect 13943 707 13951 712
rect 14048 707 14189 717
rect 14190 712 14198 717
rect 14356 716 14362 718
rect 14398 717 14408 718
rect 14398 716 14400 717
rect 14269 715 14271 716
rect 14356 715 14400 716
rect 14212 712 14214 715
rect 13945 706 13951 707
rect 13945 700 13957 706
rect 13568 687 13572 690
rect 13570 685 13572 687
rect 13571 683 13572 685
rect 13613 690 13626 691
rect 13613 687 13627 690
rect 13613 683 13635 687
rect 13491 678 13493 682
rect 13355 673 13356 676
rect 13353 668 13356 673
rect 13398 671 13402 678
rect 13432 671 13437 678
rect 13571 677 13575 683
rect 13613 679 13632 683
rect 13635 682 13637 683
rect 13640 682 13644 690
rect 13711 686 13731 691
rect 13705 683 13731 686
rect 13704 682 13731 683
rect 13741 682 13750 691
rect 13866 690 13883 693
rect 13888 691 13889 693
rect 13890 689 13894 690
rect 13945 689 13951 700
rect 13973 698 13982 700
rect 13973 691 13986 698
rect 13882 687 13894 689
rect 13943 688 13951 689
rect 13939 687 13943 688
rect 13882 685 13897 687
rect 13928 685 13939 687
rect 13882 683 13917 685
rect 13921 683 13928 685
rect 13637 681 13644 682
rect 13691 681 13731 682
rect 13637 680 13673 681
rect 13691 680 13703 681
rect 13640 679 13661 680
rect 13682 679 13714 680
rect 13613 678 13710 679
rect 13613 677 13632 678
rect 13504 675 13514 676
rect 13575 675 13576 676
rect 13632 675 13634 676
rect 13517 674 13525 675
rect 13522 671 13536 674
rect 13402 668 13404 671
rect 13346 667 13356 668
rect 13374 667 13385 668
rect 13329 664 13346 667
rect 13318 663 13329 664
rect 13211 662 13329 663
rect 13353 662 13356 667
rect 13385 666 13406 667
rect 13385 664 13408 666
rect 13405 663 13420 664
rect 13440 663 13445 668
rect 13536 667 13538 671
rect 13552 664 13563 667
rect 13547 663 13552 664
rect 13405 662 13552 663
rect 13211 659 13318 662
rect 13211 657 13297 659
rect 13352 657 13353 660
rect 13211 656 13285 657
rect 13211 655 13281 656
rect 13211 654 13274 655
rect 13211 653 13269 654
rect 13211 648 13263 653
rect 13205 642 13269 648
rect 11353 626 11366 630
rect 11181 624 11182 625
rect 11176 619 11181 624
rect 10986 614 11005 615
rect 10955 612 11005 614
rect 10956 611 11005 612
rect 10490 609 10511 610
rect 10893 609 11005 611
rect 11027 610 11036 616
rect 11111 615 11118 619
rect 11174 616 11176 619
rect 11171 615 11174 616
rect 11118 614 11171 615
rect 11124 610 11140 614
rect 11316 610 11332 626
rect 11334 610 11350 626
rect 12069 623 12096 629
rect 12908 626 12912 630
rect 12968 626 12984 642
rect 13211 636 13217 642
rect 13227 638 13233 642
rect 13233 634 13238 638
rect 13257 636 13263 642
rect 13289 634 13291 657
rect 13348 642 13352 657
rect 13408 655 13412 660
rect 13420 659 13547 662
rect 13576 660 13583 675
rect 13633 671 13636 675
rect 13640 674 13644 678
rect 13766 675 13772 677
rect 13744 674 13772 675
rect 13639 672 13640 674
rect 13737 672 13745 674
rect 13766 671 13774 674
rect 13824 671 13830 677
rect 13882 674 13898 683
rect 13622 668 13639 671
rect 13590 664 13604 667
rect 13604 663 13610 664
rect 13617 663 13637 668
rect 13772 665 13778 671
rect 13818 665 13824 671
rect 13726 663 13729 664
rect 13945 663 13951 688
rect 13964 682 13979 691
rect 14092 689 14098 707
rect 14125 706 14140 707
rect 14125 705 14154 706
rect 13604 662 13729 663
rect 13610 660 13726 662
rect 13899 660 13951 663
rect 13446 657 13535 659
rect 13446 654 13450 657
rect 13463 656 13528 657
rect 13467 655 13525 656
rect 13477 654 13519 655
rect 13412 652 13413 654
rect 13450 652 13451 654
rect 13483 653 13519 654
rect 13413 649 13415 652
rect 13416 642 13421 648
rect 13451 642 13460 652
rect 13493 644 13494 646
rect 13484 642 13499 644
rect 13348 634 13362 642
rect 13460 639 13462 642
rect 13484 639 13500 642
rect 13462 637 13463 639
rect 13484 637 13511 639
rect 13238 632 13305 634
rect 12912 624 12968 626
rect 12097 623 12124 624
rect 12952 610 12968 624
rect 13289 614 13291 632
rect 13296 630 13308 632
rect 13347 630 13362 634
rect 13464 633 13467 637
rect 13484 635 13493 637
rect 13497 635 13542 637
rect 13549 635 13558 644
rect 13583 642 13600 660
rect 13617 659 13726 660
rect 13620 657 13718 659
rect 13620 655 13626 657
rect 13631 656 13713 657
rect 13633 655 13713 656
rect 13635 652 13707 655
rect 13893 654 13957 660
rect 13614 650 13617 652
rect 13635 651 13694 652
rect 13635 650 13650 651
rect 13660 650 13666 651
rect 13607 645 13613 649
rect 13635 645 13658 650
rect 13669 645 13688 650
rect 13899 648 13905 654
rect 13914 652 13915 654
rect 13915 650 13916 652
rect 13635 644 13655 645
rect 13635 642 13637 644
rect 13639 642 13655 644
rect 13679 642 13688 645
rect 13916 644 13918 649
rect 13945 648 13951 654
rect 13583 639 13604 642
rect 13296 626 13312 630
rect 13346 626 13362 630
rect 13312 610 13328 626
rect 13330 610 13346 626
rect 13430 615 13447 633
rect 13465 625 13487 633
rect 13493 626 13502 635
rect 13540 626 13549 635
rect 13583 630 13600 639
rect 13635 634 13650 642
rect 13676 635 13688 642
rect 13741 635 13750 644
rect 13945 643 13948 648
rect 13973 645 13979 682
rect 13999 677 14002 683
rect 14035 676 14037 683
rect 13983 667 13989 673
rect 13990 667 13999 676
rect 13989 663 13999 667
rect 14003 663 14005 673
rect 14035 671 14038 676
rect 14087 674 14092 689
rect 14034 667 14038 671
rect 14041 667 14047 673
rect 14125 672 14140 705
rect 14171 704 14175 705
rect 14195 694 14205 705
rect 14271 694 14339 715
rect 14356 712 14374 715
rect 14361 708 14374 712
rect 14362 707 14374 708
rect 14402 712 14408 717
rect 14441 715 14443 718
rect 14454 716 14461 720
rect 14461 715 14463 716
rect 14495 715 14497 746
rect 14501 737 14509 749
rect 15956 743 15957 767
rect 15988 742 15991 767
rect 16124 759 16158 767
rect 16210 759 16254 767
rect 16124 758 16140 759
rect 16142 758 16161 759
rect 16220 758 16236 759
rect 16238 758 16254 759
rect 16277 763 16280 777
rect 16282 763 16288 771
rect 16146 753 16161 758
rect 16277 757 16288 763
rect 16217 753 16226 756
rect 16271 754 16288 757
rect 16305 756 16308 777
rect 16253 753 16288 754
rect 16090 740 16288 753
rect 16296 747 16308 756
rect 16374 771 16381 777
rect 16396 774 16417 781
rect 16161 738 16170 740
rect 16176 737 16282 740
rect 16305 738 16314 747
rect 16316 741 16323 747
rect 15991 733 15992 737
rect 14501 715 14509 727
rect 15992 724 15993 731
rect 16254 730 16256 737
rect 16277 730 16283 737
rect 16374 731 16375 771
rect 16402 753 16417 774
rect 16449 778 16450 785
rect 16454 778 16463 787
rect 16449 756 16451 778
rect 16455 775 16463 778
rect 16492 782 16507 787
rect 16524 782 16526 787
rect 16542 782 16562 790
rect 16492 778 16562 782
rect 16588 780 16604 790
rect 16492 774 16567 778
rect 16508 772 16524 774
rect 16526 772 16542 774
rect 16557 772 16567 774
rect 16585 774 16604 780
rect 16638 774 16654 790
rect 16684 780 16700 790
rect 16735 789 16740 808
rect 16770 803 16772 806
rect 16780 805 16796 808
rect 16831 807 16846 808
rect 16856 807 16865 815
rect 16892 810 16908 824
rect 16910 810 16926 824
rect 16937 823 16940 830
rect 16937 818 16942 823
rect 16936 816 16937 818
rect 16940 816 16942 818
rect 16967 816 16983 839
rect 16990 830 16997 838
rect 17033 830 17036 839
rect 17084 835 17095 839
rect 17084 831 17089 835
rect 16997 824 17000 830
rect 17036 828 17037 830
rect 16988 816 17004 824
rect 16932 813 16935 815
rect 16884 808 16927 810
rect 16942 808 16946 816
rect 16965 812 16967 816
rect 16988 812 17009 816
rect 17037 813 17042 828
rect 17075 817 17084 831
rect 17093 828 17095 835
rect 17088 818 17089 828
rect 17075 816 17088 817
rect 17072 815 17075 816
rect 17057 814 17069 815
rect 17055 813 17057 814
rect 17033 812 17047 813
rect 16876 807 16887 808
rect 16901 807 16903 808
rect 16927 807 16946 808
rect 16780 799 16802 805
rect 16780 798 16796 799
rect 16776 792 16796 798
rect 16802 793 16808 799
rect 16776 789 16783 792
rect 16787 789 16796 792
rect 16830 792 16846 807
rect 16854 799 16860 805
rect 16848 793 16854 799
rect 16830 790 16831 792
rect 16735 780 16750 789
rect 16780 788 16796 789
rect 16684 774 16750 780
rect 16775 778 16796 788
rect 16825 787 16827 790
rect 16830 787 16846 790
rect 16819 778 16821 787
rect 16775 776 16821 778
rect 16825 776 16846 787
rect 16863 785 16884 807
rect 16904 803 16905 805
rect 16917 799 16923 804
rect 16906 795 16907 797
rect 16927 795 16942 807
rect 16962 806 16965 812
rect 16988 810 17033 812
rect 16988 808 17009 810
rect 17037 808 17042 812
rect 16946 801 16948 805
rect 16953 795 16962 806
rect 16897 787 16913 795
rect 16927 792 16953 795
rect 16972 792 16988 808
rect 17004 806 17009 808
rect 17081 806 17088 816
rect 17093 809 17094 828
rect 17093 806 17096 809
rect 17125 807 17127 839
rect 17260 836 17262 841
rect 17290 836 17291 841
rect 17320 839 17344 841
rect 17081 805 17089 806
rect 17117 805 17127 807
rect 17131 805 17139 817
rect 17180 815 17196 824
rect 17198 815 17214 824
rect 17180 814 17214 815
rect 17262 814 17264 836
rect 17291 824 17297 836
rect 17322 830 17336 839
rect 17404 836 17406 842
rect 17429 841 17433 854
rect 17428 836 17433 841
rect 17421 834 17433 836
rect 17445 860 17473 861
rect 17445 855 17472 860
rect 17336 825 17340 830
rect 17180 813 17215 814
rect 17178 811 17180 813
rect 17213 812 17214 813
rect 17178 808 17214 811
rect 17276 809 17310 824
rect 17340 815 17344 825
rect 17344 809 17346 814
rect 17406 809 17407 825
rect 17273 808 17310 809
rect 17346 808 17347 809
rect 17009 801 17011 805
rect 17042 800 17044 805
rect 17089 802 17093 805
rect 17093 801 17117 802
rect 17125 801 17127 805
rect 17164 801 17190 808
rect 17200 801 17212 808
rect 17044 797 17045 800
rect 17013 795 17014 797
rect 16941 790 16953 792
rect 17014 791 17017 795
rect 16780 774 16791 776
rect 16826 774 16846 776
rect 16508 766 16573 772
rect 16585 768 16595 774
rect 16597 771 16631 774
rect 16634 771 16638 774
rect 16597 768 16638 771
rect 16508 758 16567 766
rect 16593 764 16595 768
rect 16604 764 16620 768
rect 16448 753 16451 756
rect 16454 753 16457 754
rect 16402 744 16457 753
rect 16515 749 16567 758
rect 16597 758 16620 764
rect 16622 758 16638 768
rect 16700 761 16716 774
rect 16597 756 16609 758
rect 16614 755 16620 758
rect 16672 755 16678 761
rect 16697 758 16716 761
rect 16718 758 16734 774
rect 16796 772 16812 774
rect 16814 772 16830 774
rect 16749 761 16755 767
rect 16787 764 16830 772
rect 16860 768 16864 785
rect 16897 780 16914 787
rect 16884 768 16890 773
rect 16910 772 16914 780
rect 16927 780 16957 790
rect 16927 774 16942 780
rect 16953 779 16957 780
rect 16936 773 16941 774
rect 16914 771 16915 772
rect 16697 755 16703 758
rect 16755 755 16761 761
rect 16796 758 16812 764
rect 16814 758 16830 764
rect 16620 749 16626 755
rect 16666 749 16672 755
rect 16699 754 16703 755
rect 16858 754 16864 768
rect 16906 767 16927 771
rect 16931 767 16936 773
rect 16872 757 16874 758
rect 16871 755 16872 757
rect 16696 750 16700 754
rect 16867 752 16871 755
rect 16906 753 16931 767
rect 16957 763 16968 779
rect 16972 774 16988 790
rect 17017 779 17022 790
rect 17022 776 17030 779
rect 17045 778 17061 797
rect 17093 793 17105 801
rect 17115 793 17127 801
rect 17158 797 17180 801
rect 17204 797 17210 801
rect 17158 795 17212 797
rect 17214 795 17230 808
rect 17260 795 17273 808
rect 17291 806 17297 808
rect 17297 802 17298 806
rect 17123 778 17127 793
rect 17152 789 17180 795
rect 17045 776 17083 778
rect 17022 775 17061 776
rect 17022 774 17038 775
rect 16968 754 16974 763
rect 16988 758 17004 774
rect 17006 763 17030 774
rect 17045 764 17061 775
rect 17068 775 17083 776
rect 17068 774 17084 775
rect 17084 763 17086 774
rect 17123 763 17125 778
rect 17006 758 17022 763
rect 17030 753 17035 763
rect 17061 754 17066 763
rect 17084 758 17089 763
rect 17124 761 17125 763
rect 17158 774 17180 789
rect 17210 792 17230 795
rect 17210 790 17224 792
rect 17210 789 17230 790
rect 17210 781 17212 789
rect 17211 774 17212 781
rect 17214 774 17230 789
rect 17253 784 17263 795
rect 17265 787 17266 795
rect 17298 786 17301 800
rect 17310 792 17326 808
rect 17251 780 17253 784
rect 17266 782 17267 786
rect 17301 781 17302 786
rect 17249 774 17251 780
rect 17302 778 17303 781
rect 17303 774 17305 778
rect 17310 774 17326 790
rect 17347 786 17355 808
rect 17421 806 17428 834
rect 17445 826 17466 855
rect 17420 802 17421 806
rect 17433 803 17442 812
rect 17445 808 17456 826
rect 17482 824 17492 847
rect 17468 818 17502 824
rect 17964 819 17965 1015
rect 18154 819 18155 1015
rect 18240 819 18241 1015
rect 18513 819 18514 1015
rect 18710 819 18711 1015
rect 17468 812 17484 818
rect 17486 812 17502 818
rect 17468 809 17502 812
rect 17468 808 17514 809
rect 17417 790 17420 800
rect 17424 794 17433 803
rect 17445 792 17468 808
rect 17480 803 17489 808
rect 17514 805 17519 808
rect 17489 794 17498 803
rect 17407 787 17422 790
rect 17355 779 17361 786
rect 17380 780 17422 787
rect 17428 786 17432 792
rect 17445 790 17455 792
rect 17445 787 17468 790
rect 17424 780 17426 784
rect 17445 781 17482 787
rect 17356 774 17372 779
rect 17380 774 17424 780
rect 17452 774 17482 781
rect 17519 774 17535 805
rect 17158 761 17214 774
rect 17216 763 17224 774
rect 17246 763 17249 774
rect 17267 764 17268 770
rect 17086 753 17089 758
rect 17125 758 17214 761
rect 17245 760 17248 763
rect 17299 760 17310 774
rect 16515 745 16574 749
rect 16696 746 16703 750
rect 16857 748 16867 752
rect 16904 749 16906 753
rect 16735 746 16832 748
rect 16855 746 16867 748
rect 16903 746 16904 748
rect 16695 745 16703 746
rect 16706 745 16841 746
rect 16852 745 16854 746
rect 16857 745 16867 746
rect 16402 741 16454 744
rect 16457 742 16458 744
rect 16396 736 16460 741
rect 16515 740 16654 745
rect 16695 744 16867 745
rect 16396 735 16462 736
rect 16317 730 16323 731
rect 16238 727 16340 730
rect 16238 724 16365 727
rect 16374 725 16381 731
rect 16402 729 16408 735
rect 16417 727 16420 732
rect 16448 729 16454 735
rect 16459 727 16462 735
rect 16421 725 16422 727
rect 16462 725 16463 727
rect 16515 726 16523 740
rect 16567 736 16654 740
rect 16569 730 16654 736
rect 16687 743 16867 744
rect 16899 743 16903 745
rect 16913 744 16931 753
rect 17035 750 17037 753
rect 17066 750 17068 753
rect 16936 744 16976 745
rect 16977 744 16988 750
rect 16687 740 16864 743
rect 16687 732 16701 740
rect 16899 735 16913 743
rect 16576 729 16577 730
rect 16577 727 16578 729
rect 14186 689 14197 691
rect 14186 688 14195 689
rect 14186 687 14196 688
rect 14199 687 14200 690
rect 14202 688 14211 691
rect 14232 690 14234 691
rect 14339 688 14359 694
rect 14362 691 14364 706
rect 14402 694 14407 712
rect 14424 696 14441 714
rect 15954 713 15955 724
rect 15993 717 15994 724
rect 16238 720 16287 724
rect 16238 717 16294 720
rect 16323 719 16329 724
rect 16238 716 16246 717
rect 16238 715 16245 716
rect 14498 711 14501 713
rect 15994 711 15995 713
rect 16257 712 16259 717
rect 14491 710 14498 711
rect 16287 710 16294 717
rect 14485 708 14497 710
rect 14474 703 14497 708
rect 15953 707 15954 710
rect 16138 707 16221 710
rect 14474 696 14485 703
rect 16259 696 16262 709
rect 16294 708 16304 709
rect 16272 700 16284 708
rect 16294 700 16306 708
rect 16263 698 16268 700
rect 16270 698 16315 700
rect 16263 697 16315 698
rect 16341 697 16343 722
rect 16369 719 16375 725
rect 16422 723 16423 725
rect 16463 720 16464 722
rect 16509 720 16525 726
rect 16425 715 16427 719
rect 16464 716 16465 719
rect 16511 716 16525 720
rect 16529 716 16532 719
rect 16555 718 16557 726
rect 16567 720 16573 726
rect 16654 725 16663 730
rect 16579 723 16580 725
rect 16554 716 16557 718
rect 16561 716 16569 720
rect 16427 709 16431 715
rect 16465 710 16467 715
rect 16511 714 16521 716
rect 16511 713 16520 714
rect 16523 713 16544 716
rect 16554 713 16556 716
rect 16559 713 16569 716
rect 16520 710 16521 713
rect 16532 710 16535 713
rect 16548 712 16552 713
rect 16552 711 16557 712
rect 16559 711 16561 713
rect 16544 710 16559 711
rect 16580 710 16587 722
rect 16663 713 16668 724
rect 16695 722 16701 732
rect 16824 723 16830 729
rect 16840 727 16846 732
rect 16835 723 16840 727
rect 16870 723 16876 729
rect 16896 727 16899 735
rect 16900 727 16913 735
rect 16896 725 16900 727
rect 16921 726 16929 744
rect 16936 740 16988 744
rect 16934 735 16970 740
rect 16976 737 16988 740
rect 17037 747 17040 750
rect 16976 735 16993 737
rect 16934 731 16936 735
rect 16977 734 16993 735
rect 17037 734 17042 747
rect 16987 731 16993 734
rect 16988 730 16993 731
rect 16991 729 16995 730
rect 17040 729 17042 734
rect 16993 726 16997 729
rect 16687 719 16701 722
rect 16687 716 16703 719
rect 16755 716 16756 719
rect 16818 717 16824 723
rect 16876 717 16882 723
rect 16892 722 16896 724
rect 16897 723 16900 725
rect 16923 724 16924 726
rect 16995 725 16997 726
rect 17041 725 17042 729
rect 16929 724 16930 725
rect 16432 698 16438 708
rect 16468 698 16470 708
rect 16523 701 16535 710
rect 16536 698 16542 708
rect 16545 701 16557 710
rect 16559 709 16624 710
rect 16566 707 16624 709
rect 16573 706 16624 707
rect 16581 703 16624 706
rect 16587 700 16593 703
rect 16595 702 16624 703
rect 16596 701 16624 702
rect 16587 698 16601 700
rect 16438 697 16442 698
rect 16263 696 16442 697
rect 14418 694 14436 696
rect 14364 688 14366 691
rect 14395 690 14436 694
rect 15952 692 15953 696
rect 16259 695 16268 696
rect 16260 694 16268 695
rect 16272 694 16442 696
rect 16470 694 16474 698
rect 15957 690 15958 692
rect 14395 688 14418 690
rect 14332 687 14426 688
rect 14183 685 14196 687
rect 14180 683 14183 685
rect 14169 677 14180 683
rect 14186 679 14194 685
rect 14085 667 14087 671
rect 14034 663 14041 667
rect 13989 661 14041 663
rect 13990 660 14049 661
rect 13973 644 13981 645
rect 13919 637 13921 641
rect 13945 637 13955 643
rect 13964 642 13981 644
rect 13989 642 13990 659
rect 13991 649 14049 660
rect 14082 655 14085 667
rect 14081 652 14082 654
rect 14118 652 14125 672
rect 14165 668 14169 676
rect 14186 663 14194 669
rect 14198 663 14200 687
rect 14364 676 14366 687
rect 14402 682 14407 687
rect 14448 676 14458 680
rect 15955 676 15958 690
rect 14268 672 14288 673
rect 14252 664 14268 672
rect 14288 664 14340 672
rect 14248 663 14252 664
rect 14186 662 14252 663
rect 14340 663 14354 664
rect 14366 663 14368 676
rect 14442 674 14448 676
rect 14411 664 14442 674
rect 15952 670 15955 676
rect 14402 663 14411 664
rect 14340 662 14411 663
rect 13999 648 14041 649
rect 13999 645 14040 648
rect 13945 635 13952 637
rect 13964 635 13990 642
rect 14003 637 14015 645
rect 14025 644 14037 645
rect 14038 644 14040 645
rect 14025 641 14040 644
rect 14078 643 14080 647
rect 14116 645 14118 651
rect 14115 643 14116 645
rect 14075 641 14078 643
rect 14022 639 14040 641
rect 14025 637 14040 639
rect 14070 637 14075 641
rect 14027 636 14040 637
rect 14017 635 14023 636
rect 14029 635 14040 636
rect 13582 626 13600 630
rect 13613 626 13650 634
rect 13685 626 13694 635
rect 13732 626 13741 635
rect 13582 625 13588 626
rect 13465 621 13480 625
rect 13577 621 13582 625
rect 13465 618 13487 621
rect 13573 618 13577 621
rect 13465 615 13488 618
rect 13569 615 13573 618
rect 13613 615 13637 626
rect 13922 615 13929 634
rect 13945 629 13955 635
rect 13447 614 13488 615
rect 10395 607 10525 609
rect 10395 606 10415 607
rect 10535 606 10554 609
rect 10882 607 11005 609
rect 7841 593 7844 594
rect 7846 589 7852 594
rect 7852 586 7855 588
rect 7935 586 7956 598
rect 7957 596 7968 598
rect 7855 585 7859 586
rect 7859 584 7906 585
rect 7926 584 7931 585
rect 7976 557 8026 606
rect 8056 557 8122 606
rect 8152 557 8218 606
rect 8248 557 8314 606
rect 8344 557 8394 606
rect 9876 557 9926 606
rect 9956 557 10022 606
rect 10052 557 10118 606
rect 10148 557 10214 606
rect 10244 557 10310 606
rect 10340 594 10415 606
rect 10340 557 10406 594
rect 10415 588 10422 594
rect 10422 586 10431 588
rect 10436 585 10502 606
rect 10532 594 10582 606
rect 10529 589 10582 594
rect 10525 586 10528 588
rect 10431 584 10502 585
rect 10523 584 10525 585
rect 10436 557 10502 584
rect 10516 581 10522 584
rect 10532 557 10582 589
rect 10644 557 10694 606
rect 10724 557 10790 606
rect 10820 557 10870 606
rect 10882 594 10898 607
rect 11008 598 11026 610
rect 13447 609 13502 614
rect 13563 610 13568 614
rect 13607 610 13613 615
rect 13618 610 13634 615
rect 13929 610 13933 615
rect 13945 614 13969 629
rect 13973 626 13990 635
rect 14020 626 14029 635
rect 14034 626 14035 635
rect 14038 624 14040 635
rect 14050 635 14070 637
rect 14112 635 14115 643
rect 14163 642 14165 660
rect 14186 657 14247 662
rect 14354 661 14411 662
rect 15945 663 15955 670
rect 15957 663 15958 676
rect 15990 687 15991 692
rect 15992 687 16017 692
rect 16257 688 16263 694
rect 15990 673 16021 687
rect 16260 684 16263 688
rect 16272 692 16368 694
rect 16272 690 16400 692
rect 16438 691 16497 694
rect 16438 690 16442 691
rect 16470 690 16474 691
rect 16497 690 16501 691
rect 16542 690 16543 696
rect 16593 695 16601 698
rect 16603 697 16624 701
rect 16665 709 16669 713
rect 16687 712 16705 716
rect 16730 712 16733 713
rect 16687 711 16703 712
rect 16687 710 16701 711
rect 16708 710 16733 712
rect 16748 710 16750 712
rect 16755 710 16761 715
rect 16809 710 16824 716
rect 16891 715 16896 722
rect 16884 711 16890 714
rect 16892 711 16896 715
rect 16918 716 16935 724
rect 16695 709 16703 710
rect 16706 709 16709 710
rect 16714 709 16816 710
rect 16665 706 16671 709
rect 16695 707 16701 709
rect 16736 707 16816 709
rect 16698 706 16816 707
rect 16884 709 16892 711
rect 16884 706 16890 709
rect 16918 708 16940 716
rect 16932 706 16940 708
rect 16951 706 16957 712
rect 16665 702 16672 706
rect 16665 701 16673 702
rect 16636 698 16646 699
rect 16665 698 16675 701
rect 16698 698 16711 706
rect 16749 703 16755 706
rect 16760 705 16829 706
rect 16876 705 16884 706
rect 16760 703 16884 705
rect 16760 700 16797 703
rect 16629 697 16633 698
rect 16647 697 16675 698
rect 16611 695 16629 697
rect 16587 694 16629 695
rect 16593 692 16624 694
rect 16593 691 16612 692
rect 16590 690 16598 691
rect 16272 688 16321 690
rect 16272 683 16306 688
rect 16272 682 16280 683
rect 16272 681 16279 682
rect 16172 673 16206 676
rect 15990 663 15991 673
rect 15996 663 16003 670
rect 14366 660 14368 661
rect 15945 658 16003 663
rect 16020 660 16021 673
rect 14194 656 14247 657
rect 15951 657 15996 658
rect 14194 655 14236 656
rect 14196 653 14234 655
rect 15951 653 15952 657
rect 15955 654 15993 657
rect 14198 645 14210 653
rect 14220 645 14232 653
rect 15957 646 15969 654
rect 15979 646 15991 654
rect 15951 642 15952 644
rect 16030 642 16031 671
rect 16313 663 16315 688
rect 16341 663 16343 690
rect 16404 688 16407 690
rect 16443 687 16444 690
rect 16501 688 16505 690
rect 16583 688 16590 690
rect 16444 678 16450 687
rect 16477 678 16484 687
rect 16493 685 16516 688
rect 16574 687 16583 688
rect 16493 684 16518 685
rect 16493 683 16539 684
rect 16543 683 16545 687
rect 16569 685 16574 687
rect 16566 684 16569 685
rect 16564 683 16566 684
rect 16493 682 16564 683
rect 16601 682 16610 691
rect 16617 690 16624 692
rect 16647 691 16678 697
rect 16696 691 16698 698
rect 16760 691 16793 700
rect 16876 695 16884 703
rect 16918 693 16940 706
rect 16945 700 16951 706
rect 16991 700 16993 725
rect 16995 713 17005 725
rect 17041 719 17047 725
rect 17068 719 17083 750
rect 17089 749 17090 753
rect 17125 751 17212 758
rect 17240 753 17246 760
rect 17290 758 17310 760
rect 17372 758 17388 774
rect 17390 770 17406 774
rect 17408 771 17415 774
rect 17419 773 17424 774
rect 17408 770 17414 771
rect 17417 770 17419 773
rect 17454 770 17460 774
rect 17390 764 17408 770
rect 17460 764 17466 770
rect 17390 758 17406 764
rect 17468 760 17482 774
rect 17535 761 17543 774
rect 17468 758 17485 760
rect 17290 753 17299 758
rect 17307 755 17308 757
rect 17479 753 17485 758
rect 17515 753 17527 761
rect 17535 756 17549 761
rect 17537 753 17549 756
rect 17125 749 17210 751
rect 17235 750 17248 753
rect 17090 746 17091 748
rect 17125 745 17216 749
rect 17228 748 17248 750
rect 17284 748 17290 753
rect 17228 746 17246 748
rect 17283 746 17284 748
rect 17232 745 17246 746
rect 17091 735 17093 744
rect 17144 743 17246 745
rect 17144 740 17176 743
rect 17192 740 17246 743
rect 17093 732 17094 735
rect 17094 730 17095 731
rect 17095 726 17096 730
rect 17144 729 17246 740
rect 17269 732 17271 743
rect 17278 740 17283 746
rect 17308 742 17311 753
rect 17275 736 17278 740
rect 17274 735 17275 736
rect 17272 732 17274 735
rect 17267 730 17272 732
rect 17155 727 17159 729
rect 17196 728 17200 729
rect 17154 725 17159 727
rect 17195 725 17196 727
rect 17257 725 17267 730
rect 17087 719 17093 725
rect 17096 721 17100 724
rect 17153 722 17159 725
rect 17215 724 17267 725
rect 17152 721 17159 722
rect 17193 721 17194 722
rect 17215 721 17257 724
rect 17035 713 17041 719
rect 17093 713 17099 719
rect 17100 717 17199 721
rect 17215 717 17250 721
rect 17269 720 17271 730
rect 17311 724 17312 742
rect 17414 740 17440 753
rect 17443 748 17448 753
rect 17485 748 17488 753
rect 17511 750 17512 752
rect 17543 749 17549 753
rect 17443 747 17449 748
rect 17443 740 17448 747
rect 17488 746 17490 748
rect 17503 746 17511 749
rect 17515 747 17549 749
rect 17546 746 17549 747
rect 17449 740 17450 746
rect 17490 740 17495 746
rect 17496 740 17509 746
rect 17312 719 17315 724
rect 17268 717 17269 719
rect 17402 718 17408 731
rect 17413 724 17414 730
rect 17450 726 17452 740
rect 17414 722 17416 724
rect 17414 721 17418 722
rect 17446 721 17448 724
rect 17414 719 17448 721
rect 17452 719 17454 726
rect 17472 725 17473 727
rect 17495 726 17509 740
rect 17460 722 17466 724
rect 17460 719 17470 722
rect 17496 720 17513 726
rect 17440 718 17470 719
rect 16995 712 16997 713
rect 16995 707 17003 712
rect 17100 707 17241 717
rect 17242 712 17250 717
rect 17408 716 17414 718
rect 17450 717 17460 718
rect 17450 716 17452 717
rect 17321 715 17323 716
rect 17408 715 17452 716
rect 17264 712 17266 715
rect 16997 706 17003 707
rect 16997 700 17009 706
rect 16620 687 16624 690
rect 16622 685 16624 687
rect 16623 683 16624 685
rect 16665 690 16678 691
rect 16665 687 16679 690
rect 16665 683 16687 687
rect 16543 678 16545 682
rect 16407 673 16408 676
rect 16405 668 16408 673
rect 16450 671 16454 678
rect 16484 671 16489 678
rect 16623 677 16627 683
rect 16665 679 16684 683
rect 16687 682 16689 683
rect 16692 682 16696 690
rect 16763 686 16783 691
rect 16757 683 16783 686
rect 16756 682 16783 683
rect 16793 682 16802 691
rect 16918 690 16935 693
rect 16940 691 16941 693
rect 16942 689 16946 690
rect 16997 689 17003 700
rect 17025 698 17034 700
rect 17025 691 17038 698
rect 16934 687 16946 689
rect 16995 688 17003 689
rect 16991 687 16995 688
rect 16934 685 16949 687
rect 16980 685 16991 687
rect 16934 683 16969 685
rect 16973 683 16980 685
rect 16689 681 16696 682
rect 16743 681 16783 682
rect 16689 680 16725 681
rect 16743 680 16755 681
rect 16692 679 16713 680
rect 16734 679 16766 680
rect 16665 678 16762 679
rect 16665 677 16684 678
rect 16556 675 16566 676
rect 16627 675 16628 676
rect 16684 675 16686 676
rect 16569 674 16577 675
rect 16574 671 16588 674
rect 16454 668 16456 671
rect 16398 667 16408 668
rect 16426 667 16437 668
rect 16381 664 16398 667
rect 16370 663 16381 664
rect 16263 662 16381 663
rect 16405 662 16408 667
rect 16437 666 16458 667
rect 16437 664 16460 666
rect 16457 663 16472 664
rect 16492 663 16497 668
rect 16588 667 16590 671
rect 16604 664 16615 667
rect 16599 663 16604 664
rect 16457 662 16604 663
rect 16263 659 16370 662
rect 16263 657 16349 659
rect 16404 657 16405 660
rect 16263 656 16337 657
rect 16263 655 16333 656
rect 16263 654 16326 655
rect 16263 653 16321 654
rect 16263 648 16315 653
rect 16257 642 16321 648
rect 14050 632 14067 635
rect 14045 627 14067 632
rect 14107 628 14112 635
rect 14105 627 14107 628
rect 14045 625 14057 627
rect 14020 622 14038 624
rect 13989 620 14024 622
rect 14044 620 14057 625
rect 13945 612 13973 614
rect 13945 611 13987 612
rect 13990 611 14006 620
rect 14008 614 14024 620
rect 14026 615 14057 620
rect 14088 616 14105 627
rect 14160 626 14165 642
rect 14234 626 14235 631
rect 14352 626 14368 642
rect 14407 630 14418 642
rect 15952 630 15960 641
rect 14405 626 14418 630
rect 14228 619 14234 625
rect 14038 614 14057 615
rect 14007 612 14057 614
rect 14008 611 14057 612
rect 13542 609 13563 610
rect 13945 609 14057 611
rect 14079 610 14088 616
rect 14163 615 14170 619
rect 14226 616 14228 619
rect 14223 615 14226 616
rect 14170 614 14223 615
rect 14176 610 14192 614
rect 14368 610 14384 626
rect 14386 610 14402 626
rect 15121 623 15148 629
rect 15960 626 15964 630
rect 16020 626 16036 642
rect 16263 636 16269 642
rect 16279 638 16285 642
rect 16285 634 16290 638
rect 16309 636 16315 642
rect 16341 634 16343 657
rect 16400 642 16404 657
rect 16460 655 16464 660
rect 16472 659 16599 662
rect 16628 660 16635 675
rect 16685 671 16688 675
rect 16692 674 16696 678
rect 16818 675 16824 677
rect 16796 674 16824 675
rect 16691 672 16692 674
rect 16789 672 16797 674
rect 16818 671 16826 674
rect 16876 671 16882 677
rect 16934 674 16950 683
rect 16674 668 16691 671
rect 16642 664 16656 667
rect 16656 663 16662 664
rect 16669 663 16689 668
rect 16824 665 16830 671
rect 16870 665 16876 671
rect 16778 663 16781 664
rect 16997 663 17003 688
rect 17016 682 17031 691
rect 17144 689 17150 707
rect 17177 706 17192 707
rect 17177 705 17206 706
rect 16656 662 16781 663
rect 16662 660 16778 662
rect 16951 660 17003 663
rect 16498 657 16587 659
rect 16498 654 16502 657
rect 16515 656 16580 657
rect 16519 655 16577 656
rect 16529 654 16571 655
rect 16464 652 16465 654
rect 16502 652 16503 654
rect 16535 653 16571 654
rect 16465 649 16467 652
rect 16468 642 16473 648
rect 16503 642 16512 652
rect 16545 644 16546 646
rect 16536 642 16551 644
rect 16400 634 16414 642
rect 16512 639 16514 642
rect 16536 639 16552 642
rect 16514 637 16515 639
rect 16536 637 16563 639
rect 16290 632 16357 634
rect 15964 624 16020 626
rect 15149 623 15176 624
rect 16004 610 16020 624
rect 16341 614 16343 632
rect 16348 630 16360 632
rect 16399 630 16414 634
rect 16516 633 16519 637
rect 16536 635 16545 637
rect 16549 635 16594 637
rect 16601 635 16610 644
rect 16635 642 16652 660
rect 16669 659 16778 660
rect 16672 657 16770 659
rect 16672 655 16678 657
rect 16683 656 16765 657
rect 16685 655 16765 656
rect 16687 652 16759 655
rect 16945 654 17009 660
rect 16666 650 16669 652
rect 16687 651 16746 652
rect 16687 650 16702 651
rect 16712 650 16718 651
rect 16659 645 16665 649
rect 16687 645 16710 650
rect 16721 645 16740 650
rect 16951 648 16957 654
rect 16966 652 16967 654
rect 16967 650 16968 652
rect 16687 644 16707 645
rect 16687 642 16689 644
rect 16691 642 16707 644
rect 16731 642 16740 645
rect 16968 644 16970 649
rect 16997 648 17003 654
rect 16635 639 16656 642
rect 16348 626 16364 630
rect 16398 626 16414 630
rect 16364 610 16380 626
rect 16382 610 16398 626
rect 16482 615 16499 633
rect 16517 625 16539 633
rect 16545 626 16554 635
rect 16592 626 16601 635
rect 16635 630 16652 639
rect 16687 634 16702 642
rect 16728 635 16740 642
rect 16793 635 16802 644
rect 16997 643 17000 648
rect 17025 645 17031 682
rect 17051 677 17054 683
rect 17087 676 17089 683
rect 17035 667 17041 673
rect 17042 667 17051 676
rect 17041 663 17051 667
rect 17055 663 17057 673
rect 17087 671 17090 676
rect 17139 674 17144 689
rect 17086 667 17090 671
rect 17093 667 17099 673
rect 17177 672 17192 705
rect 17223 704 17227 705
rect 17247 694 17257 705
rect 17323 694 17391 715
rect 17408 712 17426 715
rect 17413 708 17426 712
rect 17414 707 17426 708
rect 17454 712 17460 717
rect 17493 715 17495 718
rect 17506 716 17513 720
rect 17513 715 17515 716
rect 17547 715 17549 746
rect 17553 737 17561 749
rect 17553 715 17561 727
rect 17238 689 17249 691
rect 17238 688 17247 689
rect 17238 687 17248 688
rect 17251 687 17252 690
rect 17254 688 17263 691
rect 17284 690 17286 691
rect 17391 688 17411 694
rect 17414 691 17416 706
rect 17454 694 17459 712
rect 17476 696 17493 714
rect 17550 711 17553 713
rect 17543 710 17550 711
rect 17537 708 17549 710
rect 17526 703 17549 708
rect 17526 696 17537 703
rect 17470 694 17488 696
rect 17416 688 17418 691
rect 17447 690 17488 694
rect 17447 688 17470 690
rect 17384 687 17478 688
rect 17235 685 17248 687
rect 17232 683 17235 685
rect 17221 677 17232 683
rect 17238 679 17246 685
rect 17137 667 17139 671
rect 17086 663 17093 667
rect 17041 661 17093 663
rect 17042 660 17101 661
rect 17025 644 17033 645
rect 16971 637 16973 641
rect 16997 637 17007 643
rect 17016 642 17033 644
rect 17041 642 17042 659
rect 17043 649 17101 660
rect 17134 655 17137 667
rect 17133 652 17134 654
rect 17170 652 17177 672
rect 17217 668 17221 676
rect 17238 663 17246 669
rect 17250 663 17252 687
rect 17416 676 17418 687
rect 17454 682 17459 687
rect 17500 676 17510 680
rect 17320 672 17340 673
rect 17304 664 17320 672
rect 17340 664 17392 672
rect 17300 663 17304 664
rect 17238 662 17304 663
rect 17392 663 17406 664
rect 17418 663 17420 676
rect 17494 674 17500 676
rect 17463 664 17494 674
rect 17454 663 17463 664
rect 17392 662 17463 663
rect 17051 648 17093 649
rect 17051 645 17092 648
rect 16997 635 17004 637
rect 17016 635 17042 642
rect 17055 637 17067 645
rect 17077 644 17089 645
rect 17090 644 17092 645
rect 17077 641 17092 644
rect 17130 643 17132 647
rect 17168 645 17170 651
rect 17167 643 17168 645
rect 17127 641 17130 643
rect 17074 639 17092 641
rect 17077 637 17092 639
rect 17122 637 17127 641
rect 17079 636 17092 637
rect 17069 635 17075 636
rect 17081 635 17092 636
rect 16634 626 16652 630
rect 16665 626 16702 634
rect 16737 626 16746 635
rect 16784 626 16793 635
rect 16634 625 16640 626
rect 16517 621 16532 625
rect 16629 621 16634 625
rect 16517 618 16539 621
rect 16625 618 16629 621
rect 16517 615 16540 618
rect 16621 615 16625 618
rect 16665 615 16689 626
rect 16974 615 16981 634
rect 16997 629 17007 635
rect 16499 614 16540 615
rect 13447 607 13577 609
rect 13447 606 13467 607
rect 13587 606 13606 609
rect 13934 607 14057 609
rect 10893 593 10896 594
rect 10898 589 10904 594
rect 10904 586 10907 588
rect 10987 586 11008 598
rect 11009 596 11020 598
rect 10907 585 10911 586
rect 10911 584 10958 585
rect 10978 584 10983 585
rect 11028 557 11078 606
rect 11108 557 11174 606
rect 11204 557 11270 606
rect 11300 557 11366 606
rect 11396 557 11446 606
rect 12928 557 12978 606
rect 13008 557 13074 606
rect 13104 557 13170 606
rect 13200 557 13266 606
rect 13296 557 13362 606
rect 13392 594 13467 606
rect 13392 557 13458 594
rect 13467 588 13474 594
rect 13474 586 13483 588
rect 13488 585 13554 606
rect 13584 594 13634 606
rect 13581 589 13634 594
rect 13577 586 13580 588
rect 13483 584 13554 585
rect 13575 584 13577 585
rect 13488 557 13554 584
rect 13568 581 13574 584
rect 13584 557 13634 589
rect 13696 557 13746 606
rect 13776 557 13842 606
rect 13872 557 13922 606
rect 13934 594 13950 607
rect 14060 598 14078 610
rect 16499 609 16554 614
rect 16615 610 16620 614
rect 16659 610 16665 615
rect 16670 610 16686 615
rect 16981 610 16985 615
rect 16997 614 17021 629
rect 17025 626 17042 635
rect 17072 626 17081 635
rect 17086 626 17087 635
rect 17090 624 17092 635
rect 17102 635 17122 637
rect 17164 635 17167 643
rect 17215 642 17217 660
rect 17238 657 17299 662
rect 17406 661 17463 662
rect 17418 660 17420 661
rect 17246 656 17299 657
rect 17246 655 17288 656
rect 17248 653 17286 655
rect 17250 645 17262 653
rect 17272 645 17284 653
rect 17102 632 17119 635
rect 17097 627 17119 632
rect 17159 628 17164 635
rect 17157 627 17159 628
rect 17097 625 17109 627
rect 17072 622 17090 624
rect 17041 620 17076 622
rect 17096 620 17109 625
rect 16997 612 17025 614
rect 16997 611 17039 612
rect 17042 611 17058 620
rect 17060 614 17076 620
rect 17078 615 17109 620
rect 17140 616 17157 627
rect 17212 626 17217 642
rect 17286 626 17287 631
rect 17404 626 17420 642
rect 17459 630 17470 642
rect 17457 626 17470 630
rect 17280 619 17286 625
rect 17090 614 17109 615
rect 17059 612 17109 614
rect 17060 611 17109 612
rect 16594 609 16615 610
rect 16997 609 17109 611
rect 17131 610 17140 616
rect 17215 615 17222 619
rect 17278 616 17280 619
rect 17275 615 17278 616
rect 17222 614 17275 615
rect 17228 610 17244 614
rect 17420 610 17436 626
rect 17438 610 17454 626
rect 18173 623 18200 629
rect 18201 623 18228 624
rect 16499 607 16629 609
rect 16499 606 16519 607
rect 16639 606 16658 609
rect 16986 607 17109 609
rect 13945 593 13948 594
rect 13950 589 13956 594
rect 13956 586 13959 588
rect 14039 586 14060 598
rect 14061 596 14072 598
rect 13959 585 13963 586
rect 13963 584 14010 585
rect 14030 584 14035 585
rect 14080 557 14130 606
rect 14160 557 14226 606
rect 14256 557 14322 606
rect 14352 557 14418 606
rect 14448 557 14498 606
rect 15980 557 16030 606
rect 16060 557 16126 606
rect 16156 557 16222 606
rect 16252 557 16318 606
rect 16348 557 16414 606
rect 16444 594 16519 606
rect 16444 557 16510 594
rect 16519 588 16526 594
rect 16526 586 16535 588
rect 16540 585 16606 606
rect 16636 594 16686 606
rect 16633 589 16686 594
rect 16629 586 16632 588
rect 16535 584 16606 585
rect 16627 584 16629 585
rect 16540 557 16606 584
rect 16620 581 16626 584
rect 16636 557 16686 589
rect 16748 557 16798 606
rect 16828 557 16894 606
rect 16924 557 16974 606
rect 16986 594 17002 607
rect 17112 598 17130 610
rect 16997 593 17000 594
rect 17002 589 17008 594
rect 17008 586 17011 588
rect 17091 586 17112 598
rect 17113 596 17124 598
rect 17011 585 17015 586
rect 17015 584 17062 585
rect 17082 584 17087 585
rect 17132 557 17182 606
rect 17212 557 17278 606
rect 17308 557 17374 606
rect 17404 557 17470 606
rect 17500 557 17550 606
rect 6536 481 6537 487
rect 9588 481 9589 487
rect 12640 481 12641 487
rect 15692 481 15693 487
rect 18744 481 18745 487
rect 6502 441 6537 475
rect 6548 463 6549 475
rect 6548 441 6549 453
rect 9554 441 9589 475
rect 9600 463 9601 475
rect 9600 441 9601 453
rect 12606 441 12641 475
rect 12652 463 12653 475
rect 12652 441 12653 453
rect 15658 441 15693 475
rect 15704 463 15705 475
rect 15704 441 15705 453
rect 18710 441 18745 475
rect 18756 463 18757 475
rect 18756 441 18757 453
rect 5745 429 5746 440
rect 5935 429 5936 440
rect 6021 429 6022 440
rect 6294 429 6295 440
rect 6491 429 6492 440
rect 6525 429 6537 435
rect 8797 429 8798 440
rect 8987 429 8988 440
rect 9073 429 9074 440
rect 9346 429 9347 440
rect 9543 429 9544 440
rect 9577 429 9589 435
rect 11849 429 11850 440
rect 12039 429 12040 440
rect 12125 429 12126 440
rect 12398 429 12399 440
rect 12595 429 12596 440
rect 12629 429 12641 435
rect 14901 429 14902 440
rect 15091 429 15092 440
rect 15177 429 15178 440
rect 15450 429 15451 440
rect 15647 429 15648 440
rect 15681 429 15693 435
rect 17953 429 17954 440
rect 18143 429 18144 440
rect 18229 429 18230 440
rect 18502 429 18503 440
rect 18699 429 18700 440
rect 18733 429 18745 435
rect 5756 389 5757 429
rect 5946 389 5947 429
rect 6032 389 6033 429
rect 6305 389 6306 429
rect 6502 389 6503 429
rect 8808 389 8809 429
rect 8998 389 8999 429
rect 9084 389 9085 429
rect 9357 389 9358 429
rect 9554 389 9555 429
rect 11860 389 11861 429
rect 12050 389 12051 429
rect 12136 389 12137 429
rect 12409 389 12410 429
rect 12606 389 12607 429
rect 14912 389 14913 429
rect 15102 389 15103 429
rect 15188 389 15189 429
rect 15461 389 15462 429
rect 15658 389 15659 429
rect 17964 389 17965 429
rect 18154 389 18155 429
rect 18240 389 18241 429
rect 18513 389 18514 429
rect 18710 389 18711 429
<< nwell >>
rect 2995 1407 5844 1749
rect 7598 1647 7632 1681
rect 10650 1647 10684 1681
rect 13702 1647 13736 1681
rect 16754 1647 16788 1681
rect 2995 1275 18820 1407
rect 2995 1272 13735 1275
rect 2995 1221 13711 1272
rect 2995 1199 13735 1221
rect 13815 1199 18820 1275
rect 2995 1087 18820 1199
rect 2995 820 5844 1087
<< ndiff >>
rect 6503 441 6537 475
rect 9555 441 9589 475
rect 12607 441 12641 475
rect 15659 441 15693 475
rect 18711 441 18745 475
<< pdiff >>
rect 4546 1647 4580 1681
rect 7598 1647 7632 1681
rect 10650 1647 10684 1681
rect 13702 1647 13736 1681
rect 16754 1647 16788 1681
<< locali >>
rect 2 2173 18820 2493
rect 3407 1407 3441 1476
rect 0 1275 18820 1407
rect 0 1272 13735 1275
rect 0 1221 13711 1272
rect 0 1199 13735 1221
rect 13815 1199 18820 1275
rect 0 1087 18820 1199
rect 1 0 18820 320
<< metal1 >>
rect 2 2173 18820 2493
rect 18735 1983 18746 2014
rect 18706 1977 18776 1983
rect 3303 1863 3309 1921
rect 3367 1863 3373 1921
rect 18706 1919 18712 1977
rect 18770 1919 18776 1977
rect 18706 1913 18776 1919
rect 6502 1854 6572 1860
rect 4934 1843 5004 1849
rect 4934 1785 4940 1843
rect 4998 1785 5004 1843
rect 6502 1796 6508 1854
rect 6566 1796 6572 1854
rect 9553 1854 9624 1861
rect 6502 1790 6572 1796
rect 7986 1845 8056 1851
rect 4934 1779 5004 1785
rect 7986 1787 7992 1845
rect 8050 1787 8056 1845
rect 9553 1796 9560 1854
rect 9618 1796 9624 1854
rect 12597 1854 12667 1860
rect 9553 1790 9624 1796
rect 11038 1845 11108 1851
rect 7986 1781 8056 1787
rect 11038 1787 11044 1845
rect 11102 1787 11108 1845
rect 12597 1796 12603 1854
rect 12661 1796 12667 1854
rect 15649 1854 15719 1860
rect 12597 1790 12667 1796
rect 14090 1845 14160 1851
rect 11038 1781 11108 1787
rect 14090 1787 14096 1845
rect 14154 1787 14160 1845
rect 15649 1796 15655 1854
rect 15713 1796 15719 1854
rect 15649 1790 15719 1796
rect 17142 1845 17212 1851
rect 14090 1781 14160 1787
rect 17142 1787 17148 1845
rect 17206 1787 17212 1845
rect 17142 1781 17212 1787
rect 3228 1715 3234 1773
rect 3292 1715 3298 1773
rect 3035 1641 3093 1687
rect 4546 1647 4580 1681
rect 7598 1647 7632 1681
rect 10650 1647 10684 1681
rect 13702 1647 13736 1681
rect 16754 1647 16788 1681
rect 0 1275 18820 1407
rect 0 1272 13735 1275
rect 0 1221 13711 1272
rect 0 1199 13735 1221
rect 13815 1199 18820 1275
rect 0 1087 18820 1199
rect 6503 441 6537 475
rect 9555 441 9589 475
rect 12607 441 12641 475
rect 15659 441 15693 475
rect 18711 441 18745 475
rect 1 0 18820 320
<< via1 >>
rect 3309 1863 3367 1921
rect 18712 1919 18770 1977
rect 4940 1785 4998 1843
rect 6508 1796 6566 1854
rect 7992 1787 8050 1845
rect 9560 1796 9618 1854
rect 11044 1787 11102 1845
rect 12603 1796 12661 1854
rect 14096 1787 14154 1845
rect 15655 1796 15713 1854
rect 17148 1787 17206 1845
rect 3234 1715 3292 1773
<< metal2 >>
rect 3247 2138 18746 2172
rect 3247 1779 3281 2138
rect 18712 1983 18746 2138
rect 18706 1977 18776 1983
rect 3309 1921 3367 1927
rect 18706 1919 18712 1977
rect 18770 1919 18776 1977
rect 18706 1913 18776 1919
rect 3367 1869 3575 1903
rect 3309 1857 3367 1863
rect 3541 1829 3575 1869
rect 6502 1854 6572 1860
rect 4934 1843 5004 1849
rect 4934 1829 4940 1843
rect 3541 1795 4940 1829
rect 4934 1785 4940 1795
rect 4998 1785 5004 1843
rect 6502 1796 6508 1854
rect 6566 1836 6572 1854
rect 9554 1854 9624 1860
rect 7986 1845 8056 1851
rect 7986 1836 7992 1845
rect 6566 1796 7992 1836
rect 6502 1790 6572 1796
rect 4934 1779 5004 1785
rect 7986 1787 7992 1796
rect 8050 1787 8056 1845
rect 9554 1796 9560 1854
rect 9618 1836 9624 1854
rect 12597 1854 12667 1860
rect 11038 1845 11108 1851
rect 11038 1836 11044 1845
rect 9618 1796 11044 1836
rect 9554 1790 9624 1796
rect 7986 1781 8056 1787
rect 11038 1787 11044 1796
rect 11102 1787 11108 1845
rect 12597 1796 12603 1854
rect 12661 1836 12667 1854
rect 15649 1854 15719 1860
rect 14090 1845 14160 1851
rect 14090 1836 14096 1845
rect 12661 1796 14096 1836
rect 12597 1790 12667 1796
rect 11038 1781 11108 1787
rect 14090 1787 14096 1796
rect 14154 1787 14160 1845
rect 15649 1796 15655 1854
rect 15713 1836 15719 1854
rect 17142 1845 17212 1851
rect 17142 1836 17148 1845
rect 15713 1796 17148 1836
rect 15649 1790 15719 1796
rect 14090 1781 14160 1787
rect 17142 1787 17148 1796
rect 17206 1787 17212 1845
rect 17142 1781 17212 1787
rect 3234 1773 3292 1779
rect 3234 1709 3292 1715
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1698882961
transform 1 0 3010 0 -1 2234
box -8 0 552 902
use sky130_osu_single_mpr2ya_8_b0r1  sky130_osu_single_mpr2ya_8_b0r1_0
timestamp 1708003747
transform 1 0 15768 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2ya_8_b0r1  sky130_osu_single_mpr2ya_8_b0r1_1
timestamp 1708003747
transform 1 0 3560 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2ya_8_b0r1  sky130_osu_single_mpr2ya_8_b0r1_2
timestamp 1708003747
transform 1 0 6612 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2ya_8_b0r1  sky130_osu_single_mpr2ya_8_b0r1_3
timestamp 1708003747
transform 1 0 9664 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2ya_8_b0r1  sky130_osu_single_mpr2ya_8_b0r1_4
timestamp 1708003747
transform 1 0 12716 0 1 0
box 0 0 3052 2493
<< labels >>
flabel metal1 s 3035 1641 3093 1687 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 4546 1647 4580 1681 0 FreeSans 100 0 0 0 s1
port 1 nsew signal input
flabel metal1 s 7598 1647 7632 1681 0 FreeSans 100 0 0 0 s2
port 2 nsew signal input
flabel metal1 s 10650 1647 10684 1681 0 FreeSans 100 0 0 0 s3
port 3 nsew signal input
flabel metal1 s 13702 1647 13736 1681 0 FreeSans 100 0 0 0 s4
port 4 nsew signal input
flabel metal1 s 16754 1647 16788 1681 0 FreeSans 100 0 0 0 s5
port 5 nsew signal input
flabel metal1 s 6503 441 6537 475 0 FreeSans 100 0 0 0 X1_Y1
port 6 nsew signal output
flabel metal1 s 9555 441 9589 475 0 FreeSans 100 0 0 0 X2_Y1
port 7 nsew signal output
flabel metal1 s 12607 441 12641 475 0 FreeSans 100 0 0 0 X3_Y1
port 8 nsew signal output
flabel metal1 s 15659 441 15693 475 0 FreeSans 100 0 0 0 X4_Y1
port 9 nsew signal output
flabel metal1 s 18711 441 18745 475 0 FreeSans 100 0 0 0 X5_Y1
port 10 nsew signal output
flabel metal1 s 3000 1087 18820 1407 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 2 2173 18820 2493 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 0 1087 13711 1407 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 1 0 18820 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
<< end >>
