magic
tech sky130A
magscale 1 2
timestamp 1696006315
<< error_p >>
rect 1080 495 1089 496
rect 1000 490 1080 495
rect 1089 491 1125 495
rect 1125 490 1127 491
rect 732 482 1000 490
rect 1127 482 1144 490
rect 721 481 732 482
rect 701 479 732 481
rect 1145 479 1149 482
rect 683 468 721 479
rect 1151 471 1157 477
rect 350 466 389 467
rect 350 465 387 466
rect 389 465 390 466
rect 348 463 350 465
rect 376 457 388 465
rect 390 463 391 465
rect 650 463 683 468
rect 1055 466 1111 468
rect 391 457 397 463
rect 638 461 683 463
rect 950 462 1055 466
rect 1111 462 1121 466
rect 638 457 694 461
rect 339 456 391 457
rect 338 453 339 456
rect 397 454 398 457
rect 394 453 398 454
rect 638 455 654 457
rect 682 456 694 457
rect 656 455 678 456
rect 690 455 694 456
rect 638 453 699 455
rect 730 453 950 462
rect 1121 458 1132 462
rect 1121 455 1139 458
rect 1142 455 1207 471
rect 1121 453 1207 455
rect 328 446 334 452
rect 337 449 338 453
rect 336 446 337 449
rect 322 440 328 446
rect 348 431 349 447
rect 374 446 380 452
rect 380 440 386 446
rect 387 436 388 453
rect 393 442 400 453
rect 638 452 696 453
rect 629 449 635 452
rect 636 450 638 452
rect 640 451 645 452
rect 639 450 645 451
rect 699 450 700 452
rect 721 451 729 453
rect 1127 452 1136 453
rect 1121 451 1134 452
rect 1142 451 1207 453
rect 636 449 643 450
rect 701 449 721 451
rect 629 447 637 449
rect 622 446 638 447
rect 639 446 643 449
rect 619 442 638 446
rect 691 442 694 449
rect 386 431 388 435
rect 389 431 394 442
rect 601 435 619 442
rect 348 430 365 431
rect 349 429 365 430
rect 334 419 365 429
rect 369 419 400 431
rect 560 420 601 435
rect 622 431 638 442
rect 692 437 693 441
rect 697 439 721 449
rect 1121 450 1133 451
rect 1134 450 1207 451
rect 1223 450 1304 471
rect 1121 446 1142 450
rect 697 437 706 439
rect 692 436 694 437
rect 697 436 705 437
rect 636 429 638 431
rect 334 413 400 419
rect 546 415 560 420
rect 295 408 301 409
rect 56 406 58 408
rect 111 405 112 408
rect 288 405 292 408
rect 301 405 308 408
rect 112 403 114 405
rect 275 397 288 405
rect 308 404 313 405
rect 313 400 324 404
rect 350 402 366 413
rect 368 407 388 413
rect 538 412 544 414
rect 622 413 638 429
rect 682 433 697 436
rect 700 434 705 436
rect 682 427 698 433
rect 704 429 705 434
rect 701 427 704 429
rect 847 427 868 443
rect 1114 442 1121 446
rect 1127 442 1142 446
rect 1100 435 1114 442
rect 1134 439 1142 442
rect 1160 446 1170 450
rect 1304 446 1321 450
rect 1160 444 1173 446
rect 1142 436 1143 439
rect 682 426 706 427
rect 1061 426 1067 432
rect 1083 426 1100 435
rect 1107 426 1113 432
rect 1143 426 1150 436
rect 681 424 682 426
rect 686 415 706 426
rect 881 415 893 423
rect 903 415 915 423
rect 1055 420 1061 426
rect 1113 420 1119 426
rect 1145 421 1153 426
rect 1145 420 1154 421
rect 1145 419 1155 420
rect 1145 416 1157 419
rect 686 412 698 415
rect 1145 414 1159 416
rect 1160 414 1161 444
rect 1166 434 1187 444
rect 1321 440 1343 446
rect 1170 424 1187 434
rect 1343 433 1351 440
rect 1351 427 1355 433
rect 1145 412 1161 414
rect 1166 413 1187 424
rect 1355 423 1358 427
rect 1358 416 1362 423
rect 1166 412 1288 413
rect 1362 412 1364 416
rect 533 411 538 412
rect 530 410 533 411
rect 638 409 656 412
rect 682 411 698 412
rect 875 411 877 412
rect 917 411 954 412
rect 682 410 695 411
rect 368 402 384 407
rect 422 406 434 409
rect 436 408 441 409
rect 420 405 422 406
rect 441 405 444 408
rect 522 407 529 409
rect 518 405 522 407
rect 417 404 420 405
rect 416 403 417 404
rect 444 403 447 405
rect 514 404 518 405
rect 336 400 384 402
rect 313 399 328 400
rect 336 399 386 400
rect 409 399 418 403
rect 447 400 451 403
rect 494 402 514 404
rect 316 397 330 399
rect 331 398 386 399
rect 272 395 275 397
rect 316 395 333 397
rect 336 395 386 398
rect 405 397 418 399
rect 451 397 454 400
rect 502 399 508 402
rect 401 395 418 397
rect 454 395 457 397
rect 491 395 499 398
rect 623 397 629 400
rect 638 397 654 409
rect 656 408 663 409
rect 663 406 674 408
rect 682 407 694 410
rect 681 406 694 407
rect 674 405 694 406
rect 714 405 720 411
rect 760 407 766 411
rect 869 410 875 411
rect 750 405 766 407
rect 682 403 694 405
rect 601 395 629 397
rect 112 387 113 390
rect 111 386 150 387
rect 109 385 111 386
rect 94 375 109 385
rect 70 361 94 375
rect 67 359 70 361
rect 60 354 67 359
rect 112 354 113 386
rect 150 385 177 386
rect 254 385 272 395
rect 316 394 386 395
rect 316 392 338 394
rect 367 392 368 394
rect 374 392 380 394
rect 394 392 418 395
rect 316 389 418 392
rect 316 388 371 389
rect 374 388 380 389
rect 316 387 350 388
rect 352 387 371 388
rect 383 387 418 389
rect 316 385 371 387
rect 381 386 418 387
rect 380 385 418 386
rect 457 387 491 395
rect 457 385 480 387
rect 177 379 418 385
rect 447 379 462 385
rect 470 380 480 385
rect 476 379 480 380
rect 529 379 619 395
rect 623 394 649 395
rect 681 394 687 400
rect 708 399 772 405
rect 819 404 825 410
rect 865 409 871 410
rect 860 407 871 409
rect 854 405 859 407
rect 850 404 854 405
rect 865 404 871 407
rect 881 409 915 411
rect 919 410 927 411
rect 714 395 766 399
rect 813 398 819 404
rect 871 398 877 404
rect 629 388 635 394
rect 675 388 681 394
rect 714 379 728 395
rect 238 363 254 379
rect 300 378 323 379
rect 300 375 328 378
rect 300 374 336 375
rect 338 374 346 376
rect 367 375 368 379
rect 442 378 447 379
rect 433 376 441 377
rect 369 375 416 376
rect 428 375 433 376
rect 353 374 416 375
rect 480 374 496 379
rect 523 377 529 379
rect 714 377 729 379
rect 519 376 522 377
rect 514 374 518 375
rect 300 366 408 374
rect 367 365 368 366
rect 306 363 323 365
rect 238 357 254 361
rect 289 358 304 363
rect 327 361 352 363
rect 140 354 181 357
rect 185 354 254 357
rect 57 352 60 354
rect 112 352 140 354
rect 238 352 282 354
rect 288 352 304 358
rect 325 358 352 361
rect 371 359 430 363
rect 478 361 514 374
rect 712 372 729 377
rect 708 369 712 372
rect 701 365 708 369
rect 693 361 701 365
rect 714 361 729 372
rect 760 361 762 395
rect 766 391 779 395
rect 881 394 902 409
rect 912 408 915 409
rect 920 404 927 410
rect 955 407 962 411
rect 1145 410 1159 412
rect 1160 411 1288 412
rect 1170 410 1187 411
rect 1191 410 1288 411
rect 923 401 925 404
rect 1141 401 1144 402
rect 928 395 935 398
rect 880 393 902 394
rect 880 391 881 393
rect 766 383 774 391
rect 879 379 880 390
rect 935 381 958 395
rect 1060 394 1061 398
rect 1119 395 1141 401
rect 1145 398 1164 410
rect 1119 393 1146 395
rect 766 361 774 373
rect 473 359 478 361
rect 353 358 430 359
rect 325 356 337 358
rect 397 357 408 358
rect 345 355 357 357
rect 396 356 398 357
rect 53 350 57 352
rect 111 351 113 352
rect 109 347 114 351
rect 56 344 57 345
rect 47 335 48 340
rect 101 337 102 345
rect 108 344 114 347
rect 238 345 254 352
rect 282 351 307 352
rect 273 349 304 351
rect 307 350 318 351
rect 318 349 325 350
rect 263 347 304 349
rect 325 348 338 349
rect 346 347 353 348
rect 273 346 304 347
rect 288 345 304 346
rect 106 340 114 344
rect 106 336 108 340
rect 100 317 102 336
rect 254 329 270 345
rect 272 329 288 345
rect 365 329 367 352
rect 430 350 446 358
rect 462 354 473 359
rect 457 352 461 354
rect 451 350 457 352
rect 480 350 496 361
rect 680 353 693 361
rect 712 359 766 361
rect 777 359 779 367
rect 816 361 819 378
rect 958 376 967 381
rect 1054 380 1060 393
rect 1064 387 1085 390
rect 1101 387 1102 390
rect 1113 389 1119 393
rect 1130 387 1146 393
rect 1054 377 1061 380
rect 1062 379 1064 387
rect 1085 380 1146 387
rect 1159 383 1164 398
rect 1187 409 1288 410
rect 1365 409 1366 411
rect 1093 379 1146 380
rect 1112 378 1162 379
rect 879 366 882 370
rect 967 369 978 376
rect 1054 374 1062 377
rect 1112 374 1119 378
rect 708 353 778 359
rect 813 358 815 360
rect 882 359 897 366
rect 978 364 982 369
rect 982 361 983 364
rect 897 358 920 359
rect 813 357 819 358
rect 811 353 819 357
rect 678 352 680 353
rect 712 352 727 353
rect 728 352 729 353
rect 430 349 496 350
rect 416 348 496 349
rect 672 348 678 352
rect 712 348 733 352
rect 750 349 766 353
rect 374 347 397 348
rect 430 345 496 348
rect 464 329 480 345
rect 658 341 672 348
rect 712 345 727 348
rect 728 345 729 348
rect 760 347 766 349
rect 769 345 778 353
rect 813 352 819 353
rect 871 357 920 358
rect 871 352 877 357
rect 888 355 920 357
rect 897 354 921 355
rect 897 352 920 354
rect 923 352 948 354
rect 962 352 976 361
rect 983 359 984 361
rect 1049 359 1054 374
rect 1060 368 1067 374
rect 1060 366 1062 368
rect 984 352 987 359
rect 1047 352 1049 356
rect 808 348 810 352
rect 713 341 726 345
rect 767 341 769 345
rect 804 341 808 348
rect 819 346 825 352
rect 638 329 661 341
rect 708 338 713 341
rect 692 329 708 338
rect 725 337 728 340
rect 762 337 767 340
rect 728 329 744 337
rect 746 329 762 337
rect 796 329 804 341
rect 106 316 114 329
rect 302 321 432 329
rect 635 324 638 329
rect 684 324 692 329
rect 793 324 796 329
rect 550 321 598 324
rect 280 316 322 321
rect 100 314 106 316
rect 269 314 322 316
rect 57 311 61 314
rect 90 312 100 314
rect 103 313 106 314
rect 90 311 102 312
rect 250 311 322 314
rect 61 310 90 311
rect 98 308 102 311
rect 246 310 250 311
rect 97 307 102 308
rect 233 307 246 310
rect 45 300 46 307
rect 95 305 102 307
rect 211 306 245 307
rect 95 300 97 305
rect 211 303 233 306
rect 210 300 233 303
rect 245 300 252 306
rect 365 304 367 321
rect 409 320 550 321
rect 412 316 550 320
rect 598 316 599 321
rect 631 316 635 324
rect 670 317 684 324
rect 788 317 793 324
rect 664 316 670 317
rect 831 316 855 351
rect 865 346 871 352
rect 897 350 976 352
rect 987 350 988 352
rect 910 345 976 350
rect 988 345 990 349
rect 926 329 942 345
rect 944 334 960 345
rect 990 340 992 344
rect 992 334 994 340
rect 1035 339 1047 351
rect 1056 350 1060 366
rect 1093 357 1101 374
rect 1107 368 1113 374
rect 1055 345 1056 350
rect 1070 346 1093 356
rect 1060 344 1094 346
rect 1112 345 1113 368
rect 1146 363 1162 378
rect 1164 377 1165 382
rect 1187 379 1208 409
rect 1228 406 1288 409
rect 1366 408 1367 409
rect 1367 406 1370 408
rect 1257 404 1288 406
rect 1370 404 1372 406
rect 1266 402 1288 404
rect 1372 402 1376 404
rect 1220 379 1236 395
rect 1238 379 1254 395
rect 1278 390 1306 402
rect 1376 395 1385 402
rect 1264 379 1265 390
rect 1306 388 1310 390
rect 1385 388 1393 395
rect 1310 387 1311 388
rect 1311 385 1312 387
rect 1393 385 1395 388
rect 1581 385 1582 390
rect 1610 385 1626 395
rect 1312 380 1318 385
rect 1395 381 1400 385
rect 1564 381 1631 385
rect 1400 380 1402 381
rect 1541 380 1564 381
rect 1187 377 1220 379
rect 1225 377 1270 379
rect 1165 357 1170 374
rect 1187 363 1219 377
rect 1256 375 1270 377
rect 1318 375 1322 379
rect 1402 377 1405 380
rect 1538 377 1541 380
rect 1581 379 1582 381
rect 1631 379 1632 380
rect 1405 375 1409 377
rect 1535 375 1538 377
rect 1250 373 1270 375
rect 1322 373 1323 375
rect 1409 373 1411 375
rect 1534 373 1535 375
rect 1171 356 1177 362
rect 1187 360 1208 363
rect 1212 362 1219 363
rect 1208 356 1211 360
rect 1212 356 1223 362
rect 1165 350 1171 356
rect 1170 349 1171 350
rect 1212 347 1219 356
rect 1223 350 1229 356
rect 1261 345 1297 373
rect 1323 366 1330 373
rect 1411 366 1422 373
rect 1531 366 1534 373
rect 1330 365 1344 366
rect 1322 356 1344 365
rect 1422 360 1431 366
rect 1528 360 1531 366
rect 1431 357 1434 360
rect 1527 357 1528 360
rect 1330 348 1344 356
rect 1434 353 1439 357
rect 1525 353 1527 357
rect 1439 348 1443 353
rect 1522 351 1525 353
rect 1338 346 1347 348
rect 1344 345 1347 346
rect 1443 345 1445 348
rect 1057 342 1097 344
rect 1053 340 1055 342
rect 1057 340 1093 342
rect 1052 339 1057 340
rect 1035 337 1057 339
rect 995 334 1047 337
rect 1052 334 1057 337
rect 944 329 963 334
rect 994 329 1047 334
rect 891 318 900 322
rect 938 318 947 322
rect 957 320 963 329
rect 989 327 1004 329
rect 984 324 989 327
rect 994 324 1004 327
rect 983 323 1004 324
rect 975 321 1004 323
rect 972 320 1004 321
rect 957 318 1004 320
rect 883 316 1004 318
rect 412 311 514 316
rect 552 315 706 316
rect 552 313 699 315
rect 525 312 552 313
rect 517 311 525 312
rect 512 310 517 311
rect 503 309 512 310
rect 495 307 503 309
rect 599 308 602 313
rect 631 312 635 313
rect 664 312 670 313
rect 706 312 720 315
rect 786 312 788 316
rect 802 313 883 316
rect 891 313 1004 316
rect 490 306 495 307
rect 457 300 490 306
rect 94 296 95 300
rect 206 296 211 300
rect 214 295 233 300
rect 252 298 255 300
rect 451 299 457 300
rect 444 298 451 299
rect 428 295 443 298
rect 602 295 607 307
rect 629 304 631 312
rect 661 304 664 312
rect 720 311 724 312
rect 724 309 736 311
rect 628 301 629 304
rect 660 301 661 304
rect 736 300 774 309
rect 779 304 785 312
rect 802 309 891 313
rect 892 311 1004 313
rect 1035 312 1047 329
rect 1048 322 1054 334
rect 800 307 802 309
rect 797 305 800 307
rect 827 305 831 309
rect 777 301 779 304
rect 93 292 94 295
rect 204 292 206 295
rect 213 291 214 295
rect 44 279 45 291
rect 89 279 93 291
rect 197 279 204 291
rect 43 257 44 278
rect 82 257 89 279
rect 197 276 203 279
rect 191 270 197 276
rect 205 269 210 283
rect 243 276 249 282
rect 255 280 256 295
rect 332 291 428 295
rect 607 291 608 295
rect 626 293 628 300
rect 657 293 660 300
rect 769 299 779 300
rect 769 293 776 299
rect 779 298 785 299
rect 794 298 797 305
rect 882 304 891 309
rect 947 304 956 311
rect 965 309 966 311
rect 994 309 1004 311
rect 1034 310 1035 312
rect 1052 309 1054 322
rect 825 301 827 304
rect 966 302 968 309
rect 1004 301 1007 309
rect 1033 305 1034 307
rect 1032 302 1033 304
rect 1048 300 1054 309
rect 1070 305 1093 340
rect 1097 334 1101 342
rect 1101 307 1108 334
rect 1209 328 1212 345
rect 1269 344 1272 345
rect 1265 343 1269 344
rect 1264 340 1265 342
rect 1297 340 1304 345
rect 1257 328 1264 340
rect 1269 338 1270 340
rect 1303 334 1304 340
rect 1339 334 1346 339
rect 1347 334 1362 345
rect 1212 318 1237 328
rect 1263 318 1264 328
rect 1346 326 1358 334
rect 1362 328 1371 334
rect 1445 328 1458 345
rect 1518 343 1530 351
rect 1540 343 1552 351
rect 1592 345 1593 379
rect 1631 375 1642 379
rect 1632 363 1642 375
rect 1632 344 1633 363
rect 1518 339 1521 343
rect 1554 340 1556 343
rect 1506 327 1514 339
rect 1518 337 1552 339
rect 1518 336 1521 337
rect 1237 314 1269 318
rect 1358 317 1365 326
rect 1371 320 1377 327
rect 1458 320 1463 327
rect 1377 318 1379 320
rect 1463 318 1465 320
rect 1237 310 1270 314
rect 1145 309 1146 310
rect 1143 306 1145 309
rect 1136 305 1143 306
rect 1060 300 1062 303
rect 785 296 808 298
rect 823 297 825 300
rect 884 297 890 298
rect 930 297 936 298
rect 969 297 970 298
rect 1008 297 1009 298
rect 1030 297 1031 300
rect 1056 297 1064 300
rect 785 295 798 296
rect 816 295 823 297
rect 844 296 1056 297
rect 1066 296 1070 304
rect 1094 300 1136 305
rect 1165 304 1171 310
rect 1223 304 1229 310
rect 1237 309 1269 310
rect 1365 309 1366 317
rect 1237 308 1275 309
rect 1237 306 1278 308
rect 1338 306 1340 309
rect 1379 306 1385 318
rect 1266 304 1275 306
rect 844 295 1066 296
rect 769 292 771 293
rect 793 292 794 295
rect 798 292 839 295
rect 272 284 333 291
rect 271 282 272 283
rect 249 273 255 276
rect 256 273 257 279
rect 249 270 257 273
rect 265 270 271 282
rect 275 281 286 283
rect 332 281 333 284
rect 343 284 533 291
rect 608 287 611 291
rect 618 287 626 292
rect 649 288 657 292
rect 644 287 705 288
rect 555 284 637 287
rect 343 280 428 284
rect 521 283 539 284
rect 608 283 611 284
rect 503 280 521 283
rect 539 282 551 283
rect 554 280 557 282
rect 341 279 343 280
rect 336 276 340 279
rect 330 271 336 276
rect 363 272 365 280
rect 495 279 503 280
rect 479 276 495 279
rect 253 269 257 270
rect 329 269 330 271
rect 42 251 43 257
rect 81 252 82 257
rect 110 251 126 265
rect 128 251 144 265
rect 204 254 205 269
rect 249 267 251 268
rect 253 267 265 269
rect 251 257 282 267
rect 302 258 318 265
rect 249 252 282 257
rect 292 253 318 258
rect 78 246 81 251
rect 108 249 110 251
rect 148 249 153 251
rect 94 247 108 249
rect 94 246 105 247
rect 148 246 160 249
rect 251 248 282 252
rect 290 250 318 253
rect 288 249 299 250
rect 302 249 318 250
rect 320 249 336 265
rect 359 259 365 272
rect 445 271 479 276
rect 403 265 445 271
rect 557 270 559 280
rect 611 270 616 283
rect 618 269 626 284
rect 398 264 445 265
rect 395 263 414 264
rect 370 259 395 263
rect 359 257 370 259
rect 355 253 365 257
rect 286 248 302 249
rect 254 247 265 248
rect 282 247 302 248
rect 282 246 299 247
rect 336 246 352 249
rect 41 239 42 246
rect 75 239 78 246
rect 71 231 75 239
rect 94 233 107 246
rect 39 212 41 231
rect 69 226 71 231
rect 68 214 69 226
rect 105 216 107 233
rect 153 215 161 246
rect 204 231 206 246
rect 190 223 206 231
rect 241 231 254 246
rect 280 244 313 246
rect 280 235 308 244
rect 280 234 302 235
rect 286 233 302 234
rect 292 231 302 233
rect 335 233 352 246
rect 359 248 365 253
rect 387 249 396 253
rect 398 249 414 263
rect 416 249 432 264
rect 434 249 443 253
rect 494 249 510 265
rect 512 249 528 265
rect 559 249 563 269
rect 616 266 626 269
rect 649 266 657 287
rect 706 284 719 287
rect 723 283 725 284
rect 727 283 769 292
rect 725 280 769 283
rect 727 276 769 280
rect 785 287 839 292
rect 844 287 1071 295
rect 785 276 815 287
rect 839 286 1071 287
rect 839 284 851 286
rect 866 284 884 286
rect 727 271 815 276
rect 827 272 839 284
rect 973 283 974 286
rect 1009 281 1015 286
rect 727 266 769 271
rect 779 269 803 271
rect 823 269 827 272
rect 975 271 978 279
rect 1016 271 1019 279
rect 1022 271 1028 286
rect 1049 280 1071 286
rect 1110 281 1115 299
rect 1171 298 1177 304
rect 1171 282 1176 298
rect 1213 282 1215 304
rect 1217 298 1223 304
rect 1265 303 1275 304
rect 1266 302 1275 303
rect 1266 300 1281 302
rect 1338 300 1344 306
rect 1385 305 1386 306
rect 1269 297 1294 300
rect 1269 294 1284 297
rect 1286 294 1292 297
rect 1322 295 1331 300
rect 1332 295 1338 300
rect 1368 298 1369 302
rect 1386 300 1388 305
rect 1388 297 1390 300
rect 1275 291 1284 294
rect 1322 291 1341 295
rect 1330 287 1341 291
rect 1341 283 1342 287
rect 1369 283 1372 295
rect 1390 291 1393 297
rect 1465 292 1481 318
rect 1518 309 1520 336
rect 1518 305 1521 309
rect 1550 305 1552 337
rect 1556 327 1564 339
rect 1630 322 1633 326
rect 1623 320 1630 322
rect 1558 317 1623 320
rect 1556 306 1623 317
rect 1554 305 1564 306
rect 1514 297 1515 302
rect 1513 295 1515 297
rect 1548 296 1554 301
rect 1393 286 1397 291
rect 1397 283 1400 286
rect 1481 285 1486 291
rect 1400 282 1402 283
rect 1171 280 1204 282
rect 978 269 979 271
rect 779 266 788 269
rect 613 265 621 266
rect 613 255 624 265
rect 382 248 397 249
rect 335 231 336 233
rect 210 223 214 224
rect 190 219 230 223
rect 241 219 256 231
rect 286 224 302 231
rect 333 229 334 231
rect 190 215 256 219
rect 280 219 302 224
rect 280 215 314 219
rect 324 217 326 226
rect 335 224 352 231
rect 330 220 352 224
rect 328 217 352 220
rect 324 215 352 217
rect 359 218 363 248
rect 382 247 396 248
rect 377 244 396 247
rect 432 244 448 249
rect 377 227 394 244
rect 432 235 452 244
rect 432 233 448 235
rect 478 233 494 249
rect 529 248 544 249
rect 613 248 618 255
rect 621 253 624 255
rect 622 249 624 253
rect 528 243 544 248
rect 530 240 544 243
rect 563 241 564 248
rect 611 241 613 248
rect 624 241 640 249
rect 645 248 648 265
rect 686 255 702 265
rect 679 254 702 255
rect 704 254 727 265
rect 771 261 779 266
rect 783 265 788 266
rect 679 249 727 254
rect 670 247 691 249
rect 702 248 708 249
rect 644 241 645 247
rect 670 243 686 247
rect 696 243 702 248
rect 667 242 713 243
rect 667 241 708 242
rect 484 231 490 233
rect 493 232 494 233
rect 521 233 544 240
rect 564 238 566 241
rect 521 232 536 233
rect 492 231 494 232
rect 395 227 407 229
rect 478 228 494 231
rect 495 230 497 231
rect 530 230 536 232
rect 495 228 536 230
rect 566 228 576 238
rect 608 228 611 238
rect 624 233 644 241
rect 639 231 644 233
rect 667 233 686 241
rect 720 233 736 249
rect 748 248 754 254
rect 755 249 771 261
rect 782 254 788 265
rect 803 264 829 269
rect 793 263 836 264
rect 793 262 834 263
rect 823 254 827 262
rect 836 259 843 263
rect 843 257 844 259
rect 782 250 783 254
rect 844 253 847 257
rect 878 254 894 265
rect 896 254 912 265
rect 947 257 956 266
rect 979 265 980 269
rect 936 256 947 257
rect 869 253 871 254
rect 909 253 913 254
rect 822 250 823 253
rect 869 251 913 253
rect 869 249 903 251
rect 755 248 782 249
rect 754 242 760 248
rect 766 233 782 248
rect 667 231 677 233
rect 679 231 686 233
rect 377 226 436 227
rect 377 223 394 226
rect 436 223 440 226
rect 443 223 447 228
rect 478 226 533 228
rect 161 212 162 215
rect 69 209 70 212
rect 162 211 163 212
rect 38 184 39 208
rect 70 183 73 208
rect 107 207 108 211
rect 163 207 164 211
rect 164 204 165 207
rect 108 194 112 204
rect 165 200 166 204
rect 206 200 240 215
rect 280 212 288 215
rect 292 212 338 215
rect 288 208 291 210
rect 302 208 318 212
rect 320 208 336 212
rect 292 200 336 208
rect 166 195 171 200
rect 206 199 222 200
rect 224 199 243 200
rect 302 199 318 200
rect 320 199 336 200
rect 359 204 362 218
rect 373 216 377 223
rect 384 219 392 223
rect 440 219 447 223
rect 389 218 390 219
rect 443 218 447 219
rect 451 218 457 224
rect 478 222 501 226
rect 372 215 373 216
rect 370 212 372 215
rect 369 211 370 212
rect 366 207 370 211
rect 383 208 384 217
rect 364 204 370 207
rect 171 194 176 195
rect 112 190 114 194
rect 176 190 192 194
rect 228 193 243 199
rect 359 198 370 204
rect 114 189 115 190
rect 172 189 195 190
rect 234 189 243 193
rect 73 174 74 178
rect 36 154 37 172
rect 74 158 76 172
rect 115 165 125 189
rect 172 188 243 189
rect 299 188 308 197
rect 355 195 370 198
rect 383 197 384 206
rect 387 197 390 218
rect 354 194 370 195
rect 311 188 320 189
rect 322 188 370 194
rect 378 192 390 197
rect 456 212 463 218
rect 478 215 499 222
rect 378 188 392 192
rect 172 185 241 188
rect 243 185 252 188
rect 277 187 370 188
rect 277 185 312 187
rect 314 185 370 187
rect 172 181 370 185
rect 383 184 384 188
rect 383 183 385 184
rect 243 179 252 181
rect 258 178 365 181
rect 387 179 396 188
rect 398 182 405 188
rect 392 178 397 179
rect 335 171 338 178
rect 359 171 365 178
rect 395 177 405 178
rect 429 177 432 180
rect 391 171 429 177
rect 320 169 429 171
rect 456 172 457 212
rect 484 194 499 215
rect 531 219 532 226
rect 536 219 545 228
rect 531 197 533 219
rect 537 216 545 219
rect 574 223 589 228
rect 606 223 608 228
rect 624 223 644 231
rect 574 219 644 223
rect 670 221 686 231
rect 574 215 649 219
rect 590 213 606 215
rect 608 213 624 215
rect 639 213 649 215
rect 667 215 686 221
rect 720 215 736 231
rect 766 221 782 231
rect 817 230 822 249
rect 852 244 854 247
rect 862 246 878 249
rect 913 248 928 249
rect 938 248 947 256
rect 974 251 990 265
rect 992 251 1008 265
rect 1019 264 1022 271
rect 1019 259 1024 264
rect 1018 257 1019 259
rect 1022 257 1024 259
rect 1049 257 1066 280
rect 1072 271 1079 279
rect 1115 271 1118 280
rect 1166 276 1177 280
rect 1166 272 1171 276
rect 1079 265 1082 271
rect 1118 269 1119 271
rect 1070 257 1086 265
rect 1014 254 1017 256
rect 966 249 1009 251
rect 1024 249 1028 257
rect 958 248 969 249
rect 983 248 985 249
rect 1009 248 1028 249
rect 862 240 884 246
rect 862 239 878 240
rect 858 233 878 239
rect 884 234 890 240
rect 858 230 865 233
rect 869 230 878 233
rect 912 233 928 248
rect 936 240 942 246
rect 930 234 936 240
rect 912 231 913 233
rect 817 221 832 230
rect 862 229 878 230
rect 766 215 832 221
rect 857 219 878 229
rect 907 228 909 231
rect 912 228 928 231
rect 901 219 903 228
rect 857 217 903 219
rect 907 217 928 228
rect 945 226 966 248
rect 986 244 987 246
rect 999 240 1005 245
rect 988 236 989 238
rect 1009 236 1024 248
rect 1044 247 1049 257
rect 1070 253 1091 257
rect 1119 254 1124 269
rect 1157 258 1166 272
rect 1175 269 1177 276
rect 1170 259 1171 269
rect 1157 257 1170 258
rect 1154 256 1157 257
rect 1139 255 1151 256
rect 1137 254 1139 255
rect 1115 253 1129 254
rect 1070 251 1115 253
rect 1070 249 1091 251
rect 1119 249 1124 253
rect 1028 239 1032 246
rect 1035 236 1044 247
rect 979 228 995 236
rect 1009 233 1035 236
rect 1054 233 1070 249
rect 1086 247 1091 249
rect 1163 247 1170 257
rect 1175 250 1176 269
rect 1175 247 1178 250
rect 1207 248 1209 280
rect 1342 277 1344 282
rect 1372 277 1373 282
rect 1402 280 1426 282
rect 1163 246 1171 247
rect 1199 246 1209 248
rect 1213 246 1221 258
rect 1262 256 1278 265
rect 1280 256 1296 265
rect 1262 255 1296 256
rect 1262 254 1297 255
rect 1260 252 1262 254
rect 1295 253 1296 254
rect 1260 249 1296 252
rect 1344 249 1347 277
rect 1373 265 1380 277
rect 1404 271 1418 280
rect 1486 277 1488 283
rect 1511 282 1515 295
rect 1510 277 1515 282
rect 1502 275 1515 277
rect 1538 293 1552 296
rect 1418 266 1422 271
rect 1358 250 1392 265
rect 1422 256 1426 266
rect 1426 250 1428 255
rect 1488 250 1489 266
rect 1355 249 1392 250
rect 1428 249 1429 250
rect 1091 239 1095 246
rect 1124 241 1126 246
rect 1171 243 1175 246
rect 1175 242 1199 243
rect 1207 242 1209 246
rect 1246 242 1272 249
rect 1282 242 1294 249
rect 1126 238 1127 241
rect 1095 236 1096 238
rect 1023 231 1035 233
rect 1096 232 1099 236
rect 862 215 873 217
rect 908 215 928 217
rect 590 207 655 213
rect 667 209 677 215
rect 679 212 713 215
rect 716 212 720 215
rect 679 209 720 212
rect 590 199 649 207
rect 675 205 677 209
rect 686 205 702 209
rect 530 194 533 197
rect 536 194 539 195
rect 484 185 539 194
rect 597 190 649 199
rect 679 199 702 205
rect 704 199 720 209
rect 782 202 798 215
rect 679 197 691 199
rect 696 196 702 199
rect 754 196 760 202
rect 779 199 798 202
rect 800 199 816 215
rect 878 213 894 215
rect 896 213 912 215
rect 831 202 837 208
rect 869 205 912 213
rect 942 209 946 226
rect 979 221 996 228
rect 992 214 996 221
rect 1009 221 1039 231
rect 1009 215 1024 221
rect 1035 220 1039 221
rect 1018 214 1023 215
rect 966 209 972 214
rect 992 213 1018 214
rect 995 212 1018 213
rect 779 196 785 199
rect 837 196 843 202
rect 878 199 894 205
rect 896 199 912 205
rect 702 190 708 196
rect 748 190 754 196
rect 781 195 785 196
rect 940 195 946 209
rect 954 198 956 199
rect 953 196 954 198
rect 778 191 782 195
rect 949 193 953 196
rect 988 194 1018 212
rect 1039 204 1050 220
rect 1054 215 1070 231
rect 1099 220 1104 231
rect 1104 217 1117 220
rect 1127 219 1143 238
rect 1175 234 1187 242
rect 1197 234 1209 242
rect 1240 238 1262 242
rect 1286 238 1292 242
rect 1240 236 1294 238
rect 1296 236 1312 249
rect 1342 236 1355 249
rect 1373 243 1380 249
rect 1205 219 1209 234
rect 1234 234 1263 236
rect 1234 230 1262 234
rect 1127 217 1165 219
rect 1104 216 1143 217
rect 1104 215 1120 216
rect 1050 195 1056 204
rect 1070 199 1086 215
rect 1088 199 1117 215
rect 1127 205 1143 216
rect 1150 216 1165 217
rect 1150 215 1166 216
rect 1166 204 1168 215
rect 1205 204 1207 219
rect 1104 194 1117 199
rect 1143 195 1148 204
rect 1166 199 1171 204
rect 1206 202 1207 204
rect 1240 215 1262 230
rect 1292 233 1312 236
rect 1292 231 1306 233
rect 1292 230 1312 231
rect 1292 222 1294 230
rect 1293 215 1294 222
rect 1296 215 1312 230
rect 1335 225 1345 236
rect 1347 228 1348 236
rect 1380 227 1383 241
rect 1392 233 1408 249
rect 1333 221 1335 225
rect 1348 223 1349 227
rect 1383 222 1384 227
rect 1331 215 1333 221
rect 1384 219 1385 222
rect 1385 215 1387 219
rect 1392 215 1408 231
rect 1429 227 1437 249
rect 1502 244 1510 275
rect 1538 267 1548 293
rect 1515 244 1524 253
rect 1536 249 1538 267
rect 1550 253 1566 265
rect 1568 253 1584 265
rect 1550 250 1584 253
rect 1550 249 1596 250
rect 1502 243 1515 244
rect 1499 231 1502 241
rect 1506 235 1515 243
rect 1534 233 1550 249
rect 1562 244 1571 249
rect 1596 246 1601 249
rect 1571 235 1580 244
rect 1489 228 1504 231
rect 1437 220 1443 227
rect 1462 221 1504 228
rect 1510 227 1514 233
rect 1536 231 1538 233
rect 1534 228 1550 231
rect 1506 221 1508 225
rect 1438 215 1454 220
rect 1462 215 1506 221
rect 1534 215 1564 228
rect 1601 215 1617 246
rect 1240 202 1296 215
rect 1298 204 1306 215
rect 1328 204 1331 215
rect 1349 205 1350 211
rect 1168 194 1171 199
rect 1207 199 1296 202
rect 1327 201 1330 204
rect 1381 201 1392 215
rect 597 186 656 190
rect 778 187 785 191
rect 939 190 949 193
rect 986 190 988 194
rect 817 187 914 189
rect 937 187 949 190
rect 985 187 986 189
rect 777 186 785 187
rect 788 186 923 187
rect 934 186 936 187
rect 939 186 949 187
rect 995 186 1018 194
rect 1117 191 1119 194
rect 1148 191 1150 194
rect 484 182 536 185
rect 539 183 540 185
rect 478 177 542 182
rect 597 181 736 186
rect 777 185 949 186
rect 478 176 544 177
rect 320 165 391 169
rect 399 166 405 169
rect 456 166 463 172
rect 484 170 490 176
rect 499 168 502 173
rect 530 170 536 176
rect 541 168 544 176
rect 125 156 129 165
rect 327 161 369 165
rect 370 164 375 165
rect 327 158 368 161
rect 318 156 327 158
rect 129 154 130 156
rect 312 154 318 156
rect 76 152 77 154
rect 130 152 133 154
rect 303 152 311 154
rect 339 153 341 158
rect 35 148 36 151
rect 133 150 141 152
rect 300 151 303 152
rect 369 151 376 161
rect 405 160 411 166
rect 451 160 457 166
rect 503 162 506 168
rect 544 166 545 168
rect 597 167 605 181
rect 649 177 736 181
rect 651 171 736 177
rect 769 184 949 185
rect 981 184 985 186
rect 995 185 1058 186
rect 1059 185 1070 191
rect 769 181 946 184
rect 769 173 783 181
rect 979 176 995 184
rect 658 170 659 171
rect 659 168 660 170
rect 545 161 546 164
rect 591 161 607 167
rect 507 156 509 160
rect 546 157 547 160
rect 593 158 607 161
rect 593 157 608 158
rect 611 157 614 160
rect 637 159 639 167
rect 649 161 655 167
rect 736 166 745 171
rect 636 157 639 159
rect 643 157 651 161
rect 220 150 300 151
rect 509 150 513 156
rect 547 151 549 156
rect 593 154 603 157
rect 605 154 626 157
rect 636 154 638 157
rect 641 154 651 157
rect 601 151 603 154
rect 614 151 617 154
rect 630 152 639 154
rect 641 152 643 154
rect 626 151 641 152
rect 661 151 669 166
rect 745 154 750 165
rect 777 163 783 173
rect 906 164 912 170
rect 922 168 928 173
rect 917 164 922 168
rect 952 164 958 170
rect 978 166 995 176
rect 1003 167 1011 185
rect 1018 181 1070 185
rect 1016 176 1052 181
rect 1058 178 1070 181
rect 1119 188 1122 191
rect 1058 176 1075 178
rect 1016 172 1018 176
rect 1059 175 1075 176
rect 1119 175 1124 188
rect 1069 172 1075 175
rect 1070 171 1075 172
rect 1073 170 1077 171
rect 1122 170 1124 175
rect 1075 167 1079 170
rect 974 164 978 165
rect 979 164 995 166
rect 1005 165 1006 167
rect 1077 166 1079 167
rect 1123 166 1124 170
rect 1011 165 1013 166
rect 769 160 783 163
rect 769 157 785 160
rect 837 157 838 160
rect 900 158 906 164
rect 958 158 964 164
rect 141 148 295 150
rect 341 137 344 150
rect 376 149 386 150
rect 354 141 366 149
rect 376 141 388 149
rect 345 137 350 141
rect 376 137 386 141
rect 389 139 397 141
rect 514 139 520 149
rect 550 139 552 149
rect 605 142 617 151
rect 618 139 624 149
rect 627 142 639 151
rect 641 150 706 151
rect 648 148 706 150
rect 655 147 706 148
rect 663 144 706 147
rect 669 141 675 144
rect 677 143 706 144
rect 678 142 706 143
rect 669 139 683 141
rect 391 138 397 139
rect 520 138 524 139
rect 391 137 524 138
rect 34 133 35 137
rect 341 136 350 137
rect 342 135 350 136
rect 354 135 524 137
rect 552 135 556 139
rect 39 131 40 133
rect 37 117 40 131
rect 34 111 37 117
rect 27 101 37 111
rect 39 102 40 117
rect 72 102 73 133
rect 74 128 99 133
rect 339 129 345 135
rect 354 129 373 135
rect 386 133 450 135
rect 386 129 388 133
rect 397 129 403 133
rect 450 131 482 133
rect 520 132 579 135
rect 520 131 524 132
rect 552 131 556 132
rect 579 131 583 132
rect 624 131 625 137
rect 675 136 683 139
rect 685 138 706 142
rect 747 150 751 154
rect 769 153 787 157
rect 812 153 815 154
rect 769 152 785 153
rect 769 151 783 152
rect 790 151 815 153
rect 826 151 832 153
rect 837 151 843 156
rect 891 151 906 157
rect 973 156 979 164
rect 1000 157 1017 165
rect 966 152 972 155
rect 974 152 978 156
rect 777 150 785 151
rect 788 150 791 151
rect 796 150 898 151
rect 747 147 753 150
rect 777 148 783 150
rect 818 148 898 150
rect 780 147 898 148
rect 966 150 974 152
rect 966 147 972 150
rect 1000 149 1022 157
rect 1014 147 1022 149
rect 1033 147 1039 153
rect 747 143 754 147
rect 747 142 755 143
rect 718 139 728 140
rect 747 139 757 142
rect 780 139 793 147
rect 831 144 837 147
rect 842 146 911 147
rect 958 146 966 147
rect 842 144 966 146
rect 842 141 879 144
rect 711 138 715 139
rect 729 138 757 139
rect 693 136 711 138
rect 669 135 711 136
rect 675 132 706 135
rect 729 132 760 138
rect 778 132 780 139
rect 842 132 875 141
rect 958 136 966 144
rect 1000 134 1022 147
rect 1027 141 1033 147
rect 1073 141 1075 166
rect 1077 154 1087 166
rect 1123 160 1129 166
rect 1150 160 1165 191
rect 1171 190 1172 194
rect 1207 192 1294 199
rect 1322 194 1328 201
rect 1372 199 1392 201
rect 1454 199 1470 215
rect 1472 211 1488 215
rect 1490 212 1497 215
rect 1501 214 1506 215
rect 1490 211 1496 212
rect 1499 211 1501 214
rect 1536 211 1542 215
rect 1472 205 1490 211
rect 1542 205 1548 211
rect 1472 199 1488 205
rect 1550 201 1564 215
rect 1617 202 1625 215
rect 1550 199 1567 201
rect 1372 194 1381 199
rect 1389 196 1390 198
rect 1561 194 1567 199
rect 1207 190 1292 192
rect 1317 191 1330 194
rect 1172 187 1173 189
rect 1207 186 1298 190
rect 1310 189 1330 191
rect 1310 187 1328 189
rect 1314 186 1328 187
rect 1173 176 1175 185
rect 1226 184 1328 186
rect 1226 181 1258 184
rect 1274 181 1328 184
rect 1175 173 1176 176
rect 1176 171 1177 172
rect 1177 167 1178 171
rect 1226 170 1328 181
rect 1351 173 1353 191
rect 1366 189 1372 194
rect 1365 187 1366 189
rect 1360 181 1365 187
rect 1390 183 1393 194
rect 1357 177 1360 181
rect 1356 176 1357 177
rect 1354 173 1356 176
rect 1349 171 1354 173
rect 1236 166 1241 170
rect 1277 166 1282 170
rect 1339 166 1349 171
rect 1169 160 1175 166
rect 1178 162 1182 165
rect 1235 163 1241 166
rect 1297 165 1349 166
rect 1234 162 1241 163
rect 1275 162 1276 164
rect 1297 162 1339 165
rect 1117 154 1123 160
rect 1175 154 1181 160
rect 1182 158 1281 162
rect 1297 158 1332 162
rect 1351 161 1353 171
rect 1393 165 1394 183
rect 1496 181 1522 194
rect 1525 189 1530 194
rect 1567 189 1570 194
rect 1571 189 1580 197
rect 1597 194 1609 202
rect 1617 197 1631 202
rect 1619 194 1631 197
rect 1593 191 1594 193
rect 1625 190 1631 194
rect 1525 188 1531 189
rect 1570 188 1580 189
rect 1525 181 1530 188
rect 1555 187 1572 188
rect 1585 187 1593 190
rect 1597 188 1631 190
rect 1628 187 1631 188
rect 1531 181 1532 187
rect 1394 160 1397 165
rect 1350 158 1351 160
rect 1484 159 1490 172
rect 1495 165 1496 171
rect 1532 167 1534 181
rect 1555 179 1571 187
rect 1572 181 1577 187
rect 1578 181 1591 187
rect 1555 168 1566 179
rect 1496 163 1498 165
rect 1496 162 1500 163
rect 1528 162 1530 165
rect 1496 160 1530 162
rect 1534 160 1536 167
rect 1554 166 1555 168
rect 1577 167 1591 181
rect 1542 163 1548 165
rect 1542 160 1552 163
rect 1578 161 1595 167
rect 1522 159 1552 160
rect 1077 153 1079 154
rect 1077 148 1085 153
rect 1182 148 1323 158
rect 1324 153 1332 158
rect 1490 157 1496 159
rect 1532 158 1542 159
rect 1532 157 1534 158
rect 1403 156 1405 157
rect 1490 156 1534 157
rect 1346 153 1348 156
rect 1079 147 1085 148
rect 1079 141 1091 147
rect 672 131 680 132
rect 486 129 489 131
rect 99 120 103 128
rect 342 125 345 129
rect 525 128 526 131
rect 583 129 587 131
rect 665 129 672 131
rect 526 119 532 128
rect 559 119 566 128
rect 575 126 598 129
rect 656 128 665 129
rect 575 125 600 126
rect 575 124 621 125
rect 625 124 627 128
rect 651 126 656 128
rect 648 125 651 126
rect 646 124 648 125
rect 575 123 646 124
rect 683 123 692 132
rect 693 131 706 132
rect 702 128 706 131
rect 704 126 706 128
rect 705 124 706 126
rect 747 131 760 132
rect 747 128 761 131
rect 747 124 769 128
rect 625 119 627 123
rect 39 101 41 102
rect 71 101 73 102
rect 27 99 34 101
rect 39 99 73 101
rect 78 99 85 111
rect 102 101 103 117
rect 489 114 490 117
rect 33 94 34 99
rect 39 87 51 95
rect 61 87 73 95
rect 33 71 42 85
rect 112 83 113 112
rect 487 109 490 114
rect 532 112 536 119
rect 566 112 571 119
rect 705 118 709 124
rect 747 120 766 124
rect 769 123 771 124
rect 774 123 778 131
rect 845 127 865 132
rect 839 124 865 127
rect 838 123 865 124
rect 875 123 884 132
rect 1000 131 1017 134
rect 1022 132 1023 134
rect 1024 130 1028 131
rect 1079 130 1085 141
rect 1107 139 1116 141
rect 1107 132 1120 139
rect 1016 128 1028 130
rect 1077 129 1085 130
rect 1073 128 1077 129
rect 1016 126 1031 128
rect 1062 126 1073 128
rect 1016 124 1051 126
rect 1055 124 1062 126
rect 771 122 778 123
rect 825 122 865 123
rect 771 121 807 122
rect 825 121 837 122
rect 774 120 795 121
rect 816 120 848 121
rect 747 119 844 120
rect 747 118 766 119
rect 638 116 648 117
rect 709 116 710 117
rect 766 116 768 117
rect 651 115 659 116
rect 656 112 670 115
rect 536 109 538 112
rect 480 108 490 109
rect 508 108 519 109
rect 452 103 480 108
rect 487 103 490 108
rect 519 103 554 108
rect 574 103 579 109
rect 670 108 672 112
rect 686 105 697 108
rect 681 103 686 105
rect 354 101 359 103
rect 359 98 361 101
rect 431 100 452 103
rect 554 101 581 103
rect 419 98 431 100
rect 486 98 487 101
rect 339 83 345 89
rect 42 67 46 71
rect 102 67 118 83
rect 345 77 351 83
rect 361 79 367 98
rect 415 97 419 98
rect 408 96 415 97
rect 403 95 408 96
rect 397 94 403 95
rect 397 83 403 89
rect 482 83 486 98
rect 542 96 546 101
rect 554 100 584 101
rect 669 100 681 103
rect 710 101 717 116
rect 767 112 770 116
rect 774 115 778 119
rect 900 116 906 118
rect 878 115 906 116
rect 773 113 774 115
rect 871 113 879 115
rect 900 112 908 115
rect 958 112 964 118
rect 1016 115 1032 124
rect 756 109 773 112
rect 724 105 738 108
rect 738 103 744 105
rect 751 103 771 109
rect 906 106 912 112
rect 952 106 958 112
rect 860 103 863 105
rect 744 102 771 103
rect 744 101 763 102
rect 580 98 597 100
rect 662 98 669 100
rect 580 95 584 98
rect 597 97 601 98
rect 659 97 662 98
rect 601 96 611 97
rect 653 96 659 97
rect 611 95 617 96
rect 642 95 653 96
rect 546 93 547 95
rect 547 90 549 93
rect 550 83 555 89
rect 584 83 594 95
rect 617 94 653 95
rect 627 85 628 87
rect 618 83 633 85
rect 367 75 372 79
rect 391 77 397 83
rect 482 75 496 83
rect 594 80 596 83
rect 618 80 634 83
rect 596 78 597 80
rect 618 78 645 80
rect 372 73 439 75
rect 430 71 442 73
rect 481 71 496 75
rect 598 74 601 78
rect 618 76 627 78
rect 631 76 676 78
rect 683 76 692 85
rect 717 83 734 101
rect 751 100 762 101
rect 754 98 765 100
rect 754 96 760 98
rect 765 97 767 98
rect 769 97 784 101
rect 852 100 860 103
rect 1079 101 1085 129
rect 1098 123 1113 132
rect 1226 130 1232 148
rect 1259 147 1274 148
rect 1259 146 1288 147
rect 847 98 852 100
rect 767 96 784 97
rect 841 96 847 98
rect 769 93 784 96
rect 829 93 841 96
rect 1027 95 1033 101
rect 1079 95 1091 101
rect 748 91 751 93
rect 769 92 785 93
rect 818 92 828 93
rect 769 91 784 92
rect 794 91 800 92
rect 741 86 747 90
rect 769 86 792 91
rect 803 86 822 91
rect 1033 89 1039 95
rect 1048 91 1050 95
rect 769 85 789 86
rect 769 83 771 85
rect 773 83 789 85
rect 813 83 822 86
rect 1050 85 1052 90
rect 1079 89 1085 95
rect 717 80 738 83
rect 430 67 446 71
rect 480 67 496 71
rect 46 65 102 67
rect 86 51 102 65
rect 446 51 462 67
rect 464 51 480 67
rect 564 56 581 74
rect 599 66 621 74
rect 627 67 636 76
rect 674 67 683 76
rect 717 71 734 80
rect 769 75 784 83
rect 810 76 822 83
rect 875 76 884 85
rect 1079 84 1082 89
rect 1107 86 1113 123
rect 1133 118 1136 124
rect 1169 117 1171 124
rect 1117 108 1123 114
rect 1124 108 1133 117
rect 1123 102 1133 108
rect 1124 101 1133 102
rect 1107 85 1115 86
rect 1053 78 1055 82
rect 1079 78 1089 84
rect 1098 83 1115 85
rect 1123 83 1124 100
rect 1125 90 1133 101
rect 1137 92 1139 114
rect 1169 112 1172 117
rect 1221 115 1226 130
rect 1168 108 1172 112
rect 1175 108 1181 114
rect 1259 113 1274 146
rect 1305 145 1309 146
rect 1329 135 1339 146
rect 1405 135 1473 156
rect 1490 153 1508 156
rect 1495 149 1508 153
rect 1496 148 1508 149
rect 1536 153 1542 158
rect 1575 156 1577 159
rect 1588 157 1595 161
rect 1595 156 1597 157
rect 1629 156 1631 187
rect 1635 178 1643 190
rect 1635 156 1643 168
rect 1320 130 1331 132
rect 1320 129 1329 130
rect 1320 128 1330 129
rect 1333 128 1334 131
rect 1336 129 1345 132
rect 1366 131 1368 132
rect 1473 129 1493 135
rect 1496 129 1500 147
rect 1536 135 1541 153
rect 1558 137 1575 155
rect 1632 152 1635 154
rect 1625 151 1632 152
rect 1619 149 1631 151
rect 1608 144 1631 149
rect 1608 137 1619 144
rect 1552 135 1570 137
rect 1529 131 1570 135
rect 1529 129 1552 131
rect 1466 128 1560 129
rect 1314 124 1330 128
rect 1303 118 1314 124
rect 1320 120 1328 124
rect 1219 108 1221 112
rect 1168 102 1175 108
rect 1168 92 1171 102
rect 1137 90 1171 92
rect 1133 86 1135 89
rect 1168 86 1169 90
rect 716 67 734 71
rect 747 67 784 75
rect 819 67 828 76
rect 866 67 875 76
rect 1055 75 1056 78
rect 1079 76 1086 78
rect 1098 76 1124 83
rect 1137 78 1149 86
rect 1159 85 1171 86
rect 1172 85 1174 100
rect 1175 90 1183 102
rect 1216 96 1219 108
rect 1215 93 1216 95
rect 1159 82 1174 85
rect 1212 84 1214 88
rect 1250 86 1259 113
rect 1299 109 1303 117
rect 1249 84 1250 86
rect 1209 82 1212 84
rect 1156 80 1174 82
rect 1159 78 1174 80
rect 1204 78 1209 82
rect 1161 77 1174 78
rect 1151 76 1157 77
rect 1163 76 1174 77
rect 1191 76 1204 78
rect 1246 76 1249 84
rect 1297 83 1299 101
rect 1320 98 1328 110
rect 1332 100 1334 128
rect 1496 117 1500 128
rect 1536 123 1541 128
rect 1582 117 1592 121
rect 1402 113 1422 114
rect 1382 103 1402 113
rect 1422 103 1488 113
rect 1500 103 1502 117
rect 1576 115 1582 117
rect 1536 103 1576 115
rect 1364 100 1366 103
rect 1488 102 1576 103
rect 1332 98 1366 100
rect 1371 97 1381 102
rect 1500 101 1502 102
rect 1332 86 1344 94
rect 1354 86 1366 94
rect 716 66 722 67
rect 599 62 614 66
rect 711 62 716 66
rect 599 59 621 62
rect 599 56 622 59
rect 703 56 711 62
rect 747 56 771 67
rect 1056 56 1063 75
rect 1079 70 1089 76
rect 581 55 622 56
rect 581 50 636 55
rect 697 51 702 55
rect 741 51 747 56
rect 752 51 768 56
rect 1063 51 1067 56
rect 1079 55 1103 70
rect 1107 67 1124 76
rect 1154 67 1163 76
rect 1168 67 1169 76
rect 1172 65 1174 76
rect 1184 73 1204 76
rect 1179 68 1204 73
rect 1241 69 1246 76
rect 1239 68 1241 69
rect 1179 66 1191 68
rect 1154 63 1172 65
rect 1123 61 1158 63
rect 1178 61 1191 66
rect 1079 53 1107 55
rect 1079 52 1121 53
rect 1124 52 1140 61
rect 1142 55 1158 61
rect 1160 57 1191 61
rect 1222 57 1239 68
rect 1294 67 1299 83
rect 1368 67 1369 72
rect 1486 67 1502 83
rect 1541 71 1552 83
rect 1539 67 1552 71
rect 1362 60 1368 66
rect 1172 55 1191 57
rect 1141 53 1191 55
rect 1142 52 1191 53
rect 676 50 697 51
rect 1079 50 1191 52
rect 1213 51 1222 57
rect 1297 56 1304 60
rect 1360 57 1362 60
rect 1357 56 1360 57
rect 1304 55 1357 56
rect 1310 51 1326 55
rect 1502 51 1518 67
rect 1520 51 1536 67
rect 581 48 711 50
rect 581 47 601 48
rect 721 47 740 50
rect 1068 48 1191 50
rect 62 -2 112 47
rect 142 -2 208 47
rect 238 -2 304 47
rect 334 -2 400 47
rect 430 -2 496 47
rect 526 35 601 47
rect 526 -2 592 35
rect 601 29 608 35
rect 608 27 617 29
rect 622 26 688 47
rect 718 35 768 47
rect 715 30 768 35
rect 711 27 714 29
rect 617 25 688 26
rect 709 25 711 26
rect 622 -2 688 25
rect 702 22 708 25
rect 718 -2 768 30
rect 830 -2 880 47
rect 910 -2 976 47
rect 1006 -2 1056 47
rect 1068 35 1084 48
rect 1194 47 1221 51
rect 1194 46 1264 47
rect 1194 39 1212 46
rect 1079 34 1082 35
rect 1084 30 1090 35
rect 1090 27 1093 29
rect 1173 27 1194 39
rect 1195 37 1206 39
rect 1093 26 1097 27
rect 1097 25 1144 26
rect 1164 25 1169 26
rect 1214 -2 1264 46
rect 1294 -2 1360 47
rect 1390 -2 1456 47
rect 1486 -2 1552 47
rect 1582 -2 1632 47
<< nwell >>
rect -48 261 1796 582
<< pwell >>
rect 77 -17 111 17
<< nmos >>
rect 112 48 142 177
rect 208 48 238 177
rect 304 48 334 177
rect 400 48 430 177
rect 496 48 526 177
rect 592 48 622 177
rect 688 48 718 177
rect 784 47 814 177
rect 880 48 910 177
rect 976 48 1006 177
rect 1168 47 1198 177
rect 1264 48 1294 177
rect 1360 48 1390 177
rect 1456 48 1486 177
rect 1552 48 1582 177
<< scnmos >>
rect 112 47 142 48
rect 208 47 238 48
rect 304 47 334 48
rect 400 47 430 48
rect 496 47 526 48
rect 592 47 622 48
rect 688 47 718 48
rect 880 47 910 48
rect 976 47 1006 48
rect 1264 47 1294 48
rect 1360 47 1390 48
rect 1456 47 1486 48
rect 1552 47 1582 48
<< pmos >>
rect 112 297 142 497
rect 208 297 238 497
rect 304 297 334 497
rect 400 297 430 497
rect 496 297 526 497
rect 592 297 622 497
rect 688 297 718 497
rect 880 297 910 497
rect 976 297 1006 497
rect 1072 297 1102 497
rect 1264 297 1294 497
rect 1360 297 1390 497
rect 1456 297 1486 497
rect 1552 297 1582 497
<< ndiff >>
rect 58 101 112 177
rect 58 67 68 101
rect 102 67 112 101
rect 58 47 112 67
rect 142 47 208 177
rect 238 101 304 177
rect 238 67 254 101
rect 288 67 304 101
rect 238 47 304 67
rect 334 47 400 177
rect 430 101 496 177
rect 430 67 446 101
rect 480 67 496 101
rect 430 47 496 67
rect 526 47 592 177
rect 622 101 688 177
rect 622 67 638 101
rect 672 67 688 101
rect 622 47 688 67
rect 718 101 784 177
rect 718 67 734 101
rect 768 67 784 101
rect 718 47 784 67
rect 814 101 880 177
rect 814 67 830 101
rect 864 67 880 101
rect 814 47 880 67
rect 910 47 976 177
rect 1006 165 1060 177
rect 1006 131 1016 165
rect 1050 131 1060 165
rect 1006 47 1060 131
rect 1114 101 1168 177
rect 1114 67 1124 101
rect 1158 67 1168 101
rect 1114 47 1168 67
rect 1198 101 1264 177
rect 1198 67 1214 101
rect 1248 67 1264 101
rect 1198 47 1264 67
rect 1294 101 1360 177
rect 1294 67 1310 101
rect 1344 67 1360 101
rect 1294 47 1360 67
rect 1390 101 1456 177
rect 1390 67 1406 101
rect 1440 67 1456 101
rect 1390 47 1456 67
rect 1486 101 1552 177
rect 1486 67 1502 101
rect 1536 67 1552 101
rect 1486 47 1552 67
rect 1582 101 1636 177
rect 1582 67 1594 101
rect 1628 67 1636 101
rect 1582 47 1636 67
<< pdiff >>
rect 58 379 112 497
rect 58 345 68 379
rect 102 345 112 379
rect 58 297 112 345
rect 142 477 208 497
rect 142 443 158 477
rect 192 443 208 477
rect 142 297 208 443
rect 238 379 304 497
rect 238 345 254 379
rect 288 345 304 379
rect 238 297 304 345
rect 334 447 400 497
rect 334 413 350 447
rect 384 413 400 447
rect 334 297 400 413
rect 430 379 496 497
rect 430 345 446 379
rect 480 345 496 379
rect 430 297 496 345
rect 526 477 592 497
rect 526 443 542 477
rect 576 443 592 477
rect 526 297 592 443
rect 622 447 688 497
rect 622 413 638 447
rect 672 413 688 447
rect 622 297 688 413
rect 718 379 772 497
rect 718 345 728 379
rect 762 345 772 379
rect 718 297 772 345
rect 826 477 880 497
rect 826 443 834 477
rect 868 443 880 477
rect 826 297 880 443
rect 910 379 976 497
rect 910 345 926 379
rect 960 345 976 379
rect 910 297 976 345
rect 1006 477 1072 497
rect 1006 443 1022 477
rect 1056 443 1072 477
rect 1006 297 1072 443
rect 1102 379 1156 497
rect 1102 345 1112 379
rect 1146 345 1156 379
rect 1102 297 1156 345
rect 1210 379 1264 497
rect 1210 345 1220 379
rect 1254 345 1264 379
rect 1210 297 1264 345
rect 1294 297 1360 497
rect 1390 477 1456 497
rect 1390 443 1406 477
rect 1440 443 1456 477
rect 1390 297 1456 443
rect 1486 297 1552 497
rect 1582 379 1636 497
rect 1582 345 1592 379
rect 1626 345 1636 379
rect 1582 297 1636 345
<< ndiffc >>
rect 68 67 102 101
rect 254 67 288 101
rect 446 67 480 101
rect 638 67 672 101
rect 734 67 768 101
rect 830 67 864 101
rect 1016 131 1050 165
rect 1124 67 1158 101
rect 1214 67 1248 101
rect 1310 67 1344 101
rect 1406 67 1440 101
rect 1502 67 1536 101
rect 1594 67 1628 101
<< pdiffc >>
rect 68 345 102 379
rect 158 443 192 477
rect 254 345 288 379
rect 350 413 384 447
rect 446 345 480 379
rect 542 443 576 477
rect 638 413 672 447
rect 728 345 762 379
rect 834 443 868 477
rect 926 345 960 379
rect 1022 443 1056 477
rect 1112 345 1146 379
rect 1220 345 1254 379
rect 1406 443 1440 477
rect 1592 345 1626 379
<< poly >>
rect 112 497 142 523
rect 208 497 238 523
rect 304 497 334 523
rect 400 497 430 523
rect 496 497 526 523
rect 592 497 622 523
rect 688 497 718 523
rect 880 497 910 523
rect 976 497 1006 523
rect 1072 497 1102 523
rect 1264 497 1294 523
rect 1360 497 1390 523
rect 1456 497 1486 523
rect 1552 497 1582 523
rect 112 265 142 297
rect 208 265 238 297
rect 304 265 334 297
rect 400 265 430 297
rect 496 265 526 297
rect 592 265 622 297
rect 688 265 718 297
rect 880 265 910 297
rect 976 265 1006 297
rect 1072 265 1102 297
rect 1264 265 1294 297
rect 1360 265 1390 297
rect 1456 265 1486 297
rect 1552 265 1582 297
rect 100 249 154 265
rect 100 215 110 249
rect 144 215 154 249
rect 100 199 154 215
rect 196 249 250 265
rect 196 215 206 249
rect 240 215 250 249
rect 196 199 250 215
rect 292 249 346 265
rect 292 215 302 249
rect 336 215 346 249
rect 292 199 346 215
rect 388 249 442 265
rect 388 215 398 249
rect 432 215 442 249
rect 388 199 442 215
rect 484 249 538 265
rect 484 215 494 249
rect 528 215 538 249
rect 484 199 538 215
rect 580 249 634 265
rect 580 215 590 249
rect 624 215 634 249
rect 580 199 634 215
rect 676 249 730 265
rect 676 215 686 249
rect 720 215 730 249
rect 676 199 730 215
rect 772 249 826 265
rect 772 215 782 249
rect 816 215 826 249
rect 772 199 826 215
rect 868 249 922 265
rect 868 215 878 249
rect 912 215 922 249
rect 868 199 922 215
rect 964 249 1018 265
rect 964 215 974 249
rect 1008 215 1018 249
rect 964 199 1018 215
rect 1060 249 1114 265
rect 1060 215 1070 249
rect 1104 215 1114 249
rect 1060 199 1114 215
rect 1156 249 1210 265
rect 1156 215 1166 249
rect 1200 215 1210 249
rect 1156 199 1210 215
rect 1252 249 1306 265
rect 1252 215 1262 249
rect 1296 215 1306 249
rect 1252 199 1306 215
rect 1348 249 1402 265
rect 1348 215 1358 249
rect 1392 215 1402 249
rect 1348 199 1402 215
rect 1444 249 1498 265
rect 1444 215 1454 249
rect 1488 215 1498 249
rect 1444 199 1498 215
rect 1540 249 1594 265
rect 1540 215 1550 249
rect 1584 215 1594 249
rect 1540 199 1594 215
rect 112 177 142 199
rect 208 177 238 199
rect 304 177 334 199
rect 400 177 430 199
rect 496 177 526 199
rect 592 177 622 199
rect 688 177 718 199
rect 784 177 814 199
rect 880 177 910 199
rect 976 177 1006 199
rect 1168 177 1198 199
rect 1264 177 1294 199
rect 1360 177 1390 199
rect 1456 177 1486 199
rect 1552 177 1582 199
rect 112 21 142 47
rect 208 21 238 47
rect 304 21 334 47
rect 400 21 430 47
rect 496 21 526 47
rect 592 21 622 47
rect 688 21 718 47
rect 784 21 814 47
rect 880 21 910 47
rect 976 21 1006 47
rect 1168 21 1198 47
rect 1264 21 1294 47
rect 1360 21 1390 47
rect 1456 21 1486 47
rect 1552 21 1582 47
<< polycont >>
rect 110 215 144 249
rect 206 215 240 249
rect 302 215 336 249
rect 398 215 432 249
rect 494 215 528 249
rect 590 215 624 249
rect 686 215 720 249
rect 782 215 816 249
rect 878 215 912 249
rect 974 215 1008 249
rect 1070 215 1104 249
rect 1166 215 1200 249
rect 1262 215 1296 249
rect 1358 215 1392 249
rect 1454 215 1488 249
rect 1550 215 1584 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 158 477 192 527
rect 542 477 576 527
tri 350 465 387 467 se
tri 387 466 389 467 sw
rect 387 465 389 466
tri 389 465 390 466 sw
rect 158 427 192 443
tri 348 463 350 465 se
rect 350 463 390 465
tri 390 463 391 465 sw
rect 348 457 391 463
tri 391 457 397 463 sw
rect 348 454 397 457
tri 397 454 398 457 sw
rect 348 453 394 454
rect 348 447 354 453
tri 348 430 349 447 ne
rect 349 423 350 447
tri 349 413 350 423 ne
rect 388 442 394 453
tri 394 443 398 454 nw
rect 834 477 868 527
tri 638 452 696 455 se
tri 696 453 699 455 sw
rect 696 452 699 453
rect 388 423 389 442
tri 389 428 394 442 nw
rect 542 427 576 443
tri 636 449 638 452 se
rect 638 450 699 452
tri 699 450 700 452 sw
rect 638 449 700 450
rect 636 447 660 449
tri 636 429 638 447 ne
tri 388 419 389 423 nw
tri 384 413 388 419 nw
rect 694 434 700 449
tri 700 434 705 449 sw
rect 694 429 704 434
tri 704 429 705 434 nw
rect 694 423 701 429
tri 701 423 704 429 nw
rect 834 427 868 443
rect 1022 477 1056 527
rect 1406 477 1440 527
tri 1142 450 1207 471 se
rect 1207 450 1223 471
tri 1223 450 1304 471 sw
rect 1022 427 1056 443
tri 1127 446 1142 450 se
rect 1142 446 1304 450
tri 1304 446 1321 450 sw
rect 694 416 698 423
tri 698 416 701 423 nw
rect 694 415 697 416
tri 697 415 698 416 nw
rect 672 413 693 415
rect 638 412 693 413
tri 693 412 697 415 nw
rect 1161 440 1321 446
tri 1321 440 1343 446 sw
rect 1161 433 1343 440
tri 1343 433 1351 440 sw
rect 1161 427 1351 433
tri 1351 427 1355 433 sw
rect 1406 427 1440 443
rect 1161 423 1355 427
tri 1355 423 1358 427 sw
rect 1161 416 1358 423
tri 1358 416 1362 423 sw
rect 1161 412 1362 416
tri 1362 412 1364 416 sw
tri 638 409 656 412 ne
rect 656 409 682 412
tri 295 408 298 409 se
tri 298 408 301 409 sw
tri 56 406 58 408 se
rect 58 406 111 408
rect 56 405 111 406
tri 111 405 112 408 sw
tri 288 405 292 408 se
rect 292 405 301 408
tri 301 405 308 408 sw
tri 422 406 434 409 se
rect 434 408 436 409
tri 436 408 441 409 sw
tri 656 408 663 409 ne
rect 663 408 682 409
rect 434 406 441 408
tri 420 405 422 406 se
rect 422 405 441 406
tri 441 405 444 408 sw
tri 663 406 674 408 ne
rect 674 406 682 408
tri 682 406 693 412 nw
tri 917 411 953 412 se
tri 953 411 954 412 sw
tri 1160 411 1172 412 ne
rect 1172 411 1365 412
tri 674 405 678 406 ne
tri 678 405 682 406 nw
rect 56 403 112 405
tri 112 403 114 405 sw
rect 56 379 114 403
tri 275 397 288 405 se
rect 288 404 308 405
tri 308 404 313 405 sw
tri 417 404 420 405 se
rect 420 404 444 405
rect 288 399 313 404
tri 313 399 324 404 sw
tri 416 403 417 404 se
rect 417 403 444 404
tri 444 403 447 405 sw
tri 409 400 416 403 se
rect 416 400 447 403
tri 447 400 451 403 sw
rect 288 397 324 399
tri 324 397 330 399 sw
tri 405 397 409 399 se
rect 409 397 451 400
tri 451 397 454 400 sw
tri 272 395 275 397 se
rect 275 395 331 397
tri 331 395 333 397 sw
tri 401 395 403 397 se
rect 403 395 454 397
tri 454 395 457 397 sw
tri 727 395 729 397 se
tri 729 395 766 397 sw
tri 257 385 272 395 se
rect 272 392 333 395
tri 333 392 338 395 sw
tri 394 392 401 395 se
rect 401 392 457 395
rect 272 387 338 392
tri 338 387 350 392 sw
tri 383 387 394 392 se
rect 394 387 457 392
rect 272 385 350 387
tri 350 385 362 387 sw
tri 381 386 383 387 se
rect 383 386 457 387
tri 380 385 381 386 se
rect 381 385 457 386
tri 457 385 469 395 sw
rect 56 345 68 379
tri 56 344 57 345 ne
rect 57 317 68 345
rect 102 327 114 379
tri 254 379 257 385 se
rect 257 380 470 385
tri 470 380 476 385 sw
rect 257 379 476 380
tri 476 379 480 380 sw
rect 288 365 446 379
rect 288 363 306 365
tri 306 363 314 365 nw
tri 314 363 323 365 ne
rect 323 363 446 365
rect 288 358 300 363
tri 300 358 304 363 nw
tri 327 358 352 363 ne
rect 352 358 371 363
tri 371 358 424 363 nw
tri 424 358 430 363 ne
rect 430 358 446 363
tri 288 345 299 358 nw
tri 430 345 446 358 ne
tri 725 345 727 379 se
rect 727 345 728 395
rect 762 391 774 395
tri 774 391 779 395 sw
rect 762 367 779 391
tri 880 391 881 394 se
rect 762 359 777 367
tri 777 359 779 367 nw
tri 879 379 880 390 se
rect 880 379 881 391
rect 879 377 881 379
rect 915 407 955 411
tri 955 407 962 411 sw
tri 1191 409 1228 411 ne
rect 1228 409 1365 411
tri 1365 409 1366 411 sw
rect 915 379 962 407
tri 1228 406 1257 409 ne
rect 1257 408 1366 409
tri 1366 408 1367 409 sw
rect 1257 406 1367 408
tri 1367 406 1370 408 sw
tri 1257 404 1266 406 ne
rect 1266 404 1370 406
tri 1370 404 1372 406 sw
tri 1266 402 1278 404 ne
rect 1278 402 1372 404
tri 1372 402 1376 404 sw
tri 1278 390 1306 402 ne
rect 1306 395 1376 402
tri 1376 395 1385 402 sw
rect 1306 390 1385 395
tri 1064 387 1067 390 se
tri 1067 387 1085 390 sw
tri 1306 388 1310 390 ne
rect 1310 388 1385 390
tri 1385 388 1393 395 sw
tri 1310 387 1311 388 ne
rect 1311 387 1393 388
rect 915 377 926 379
rect 879 370 926 377
tri 879 366 882 370 ne
rect 882 366 926 370
tri 882 359 897 366 ne
rect 897 359 926 366
rect 762 345 769 359
tri 769 345 777 359 nw
tri 897 350 920 359 ne
rect 920 350 926 359
tri 920 345 926 350 ne
rect 960 352 962 379
tri 1062 379 1064 387 se
rect 1064 380 1085 387
tri 1085 380 1145 387 sw
tri 1311 385 1312 387 ne
rect 1312 385 1393 387
tri 1393 385 1395 388 sw
tri 1312 380 1318 385 ne
rect 1318 381 1395 385
tri 1395 381 1400 385 sw
tri 1564 381 1626 385 se
tri 1626 381 1631 385 sw
rect 1318 380 1400 381
tri 1400 380 1402 381 sw
tri 1541 380 1564 381 se
rect 1564 380 1631 381
rect 1064 379 1145 380
rect 1318 379 1402 380
tri 1060 366 1062 377 se
rect 1062 366 1112 379
rect 960 350 961 352
tri 961 350 962 352 nw
tri 1056 350 1060 366 se
rect 1060 350 1112 366
tri 960 345 961 350 nw
tri 1055 345 1056 350 se
rect 1056 345 1112 350
tri 1219 377 1220 379 se
tri 1212 347 1219 377 se
rect 1219 347 1220 377
rect 1212 345 1220 347
tri 1254 377 1256 379 sw
rect 1254 373 1256 377
tri 1256 373 1261 377 sw
tri 1318 375 1322 379 ne
rect 1322 377 1402 379
tri 1402 377 1405 380 sw
tri 1538 377 1541 380 se
rect 1541 379 1631 380
rect 1541 377 1592 379
rect 1322 375 1405 377
tri 1405 375 1409 377 sw
tri 1535 375 1538 377 se
rect 1538 375 1592 377
tri 1322 373 1323 375 ne
rect 1323 373 1409 375
tri 1409 373 1411 375 sw
tri 1534 373 1535 375 se
rect 1535 373 1592 375
rect 1254 345 1261 373
tri 1261 345 1297 373 sw
tri 1323 366 1330 373 ne
rect 1330 366 1411 373
tri 1411 366 1422 373 sw
tri 1531 366 1534 373 se
rect 1534 366 1592 373
tri 1330 348 1344 366 ne
rect 1344 360 1422 366
tri 1422 360 1431 366 sw
tri 1528 360 1531 366 se
rect 1531 360 1592 366
rect 1344 357 1431 360
tri 1431 357 1434 360 sw
tri 1527 357 1528 360 se
rect 1528 357 1592 360
rect 1344 353 1434 357
tri 1434 353 1439 357 sw
tri 1525 353 1527 357 se
rect 1527 353 1592 357
rect 1344 348 1439 353
tri 1439 348 1443 353 sw
tri 1522 348 1525 353 se
rect 1525 348 1592 353
tri 1344 345 1347 348 ne
rect 1347 345 1443 348
tri 1443 345 1445 348 sw
tri 1521 345 1522 347 se
rect 1522 345 1592 348
rect 1626 375 1631 379
tri 1631 375 1632 380 sw
rect 1626 345 1632 375
rect 725 340 767 345
tri 767 341 769 345 nw
tri 725 337 728 340 ne
rect 728 337 762 340
tri 762 337 767 340 nw
tri 1053 340 1055 342 se
rect 1055 340 1146 345
tri 1043 337 1053 339 se
rect 1053 337 1146 340
tri 995 329 1038 337 se
rect 1038 334 1146 337
rect 1038 329 1060 334
rect 102 317 106 327
rect 57 316 106 317
tri 106 316 114 327 nw
tri 302 321 350 329 se
tri 350 321 432 329 sw
tri 989 327 995 329 se
rect 995 327 1060 329
tri 984 324 989 327 se
rect 989 324 1060 327
tri 550 321 593 324 se
tri 593 321 598 324 sw
tri 983 323 984 324 se
rect 984 323 1060 324
tri 975 321 983 323 se
rect 983 321 1060 323
tri 280 316 302 321 se
rect 302 316 432 321
tri 432 316 481 321 sw
tri 481 316 550 321 se
rect 550 316 598 321
tri 598 316 599 321 sw
tri 972 320 975 321 se
rect 975 320 1060 321
tri 962 318 972 320 se
rect 972 318 1060 320
tri 883 316 910 318 se
rect 910 316 1060 318
rect 57 314 100 316
tri 100 314 106 316 nw
tri 269 314 280 316 se
rect 280 314 599 316
tri 57 311 61 314 ne
rect 61 311 90 314
tri 90 311 100 314 nw
tri 250 311 269 314 se
rect 269 311 599 314
tri 61 310 88 311 ne
tri 88 310 90 311 nw
tri 246 310 250 311 se
rect 250 310 599 311
tri 233 307 246 310 se
rect 246 308 599 310
tri 599 308 602 316 sw
tri 802 309 883 316 se
rect 883 309 1060 316
rect 246 307 602 308
tri 800 307 802 309 se
rect 802 307 1060 309
tri 214 295 233 307 se
rect 233 295 602 307
tri 602 295 607 307 sw
tri 797 305 800 307 se
rect 800 305 1060 307
tri 794 295 797 305 se
rect 797 300 1060 305
rect 1094 310 1146 334
tri 1209 334 1212 345 se
rect 1212 340 1297 345
tri 1297 340 1304 345 sw
tri 1209 328 1212 334 ne
rect 1212 328 1269 340
tri 1212 318 1237 328 ne
rect 1237 318 1269 328
rect 1094 309 1145 310
tri 1145 309 1146 310 nw
rect 1094 306 1143 309
tri 1143 306 1145 309 nw
tri 1237 306 1269 318 ne
tri 1303 334 1304 340 nw
tri 1347 334 1362 345 ne
rect 1362 334 1445 345
tri 1362 328 1371 334 ne
rect 1371 328 1445 334
tri 1445 328 1458 345 sw
rect 1371 327 1458 328
tri 1518 339 1521 345 se
rect 1521 344 1632 345
tri 1632 344 1633 375 sw
rect 1521 339 1633 344
tri 1371 320 1377 327 ne
rect 1377 320 1458 327
tri 1458 320 1463 327 sw
tri 1377 318 1379 320 ne
rect 1379 318 1463 320
tri 1463 318 1465 320 sw
tri 1379 306 1385 318 ne
rect 1385 306 1465 318
rect 1094 305 1136 306
tri 1136 305 1143 306 nw
tri 1385 305 1386 306 ne
rect 1386 305 1465 306
tri 1094 300 1136 305 nw
tri 1386 300 1388 305 ne
rect 1388 300 1465 305
rect 797 297 1056 300
tri 1056 297 1064 300 nw
tri 1388 297 1390 300 ne
rect 1390 297 1465 300
rect 797 295 844 297
tri 213 291 214 295 se
rect 214 291 332 295
tri 332 291 367 295 nw
tri 367 291 428 295 ne
rect 428 291 607 295
tri 607 291 608 295 sw
tri 793 291 794 295 se
rect 794 291 844 295
tri 205 269 210 283 se
tri 204 254 205 269 se
rect 205 257 210 269
rect 244 283 272 291
tri 272 284 332 291 nw
tri 428 284 533 291 ne
rect 533 284 608 291
tri 533 283 539 284 ne
rect 539 283 608 284
tri 608 283 611 291 sw
tri 791 283 793 291 se
rect 793 286 844 291
tri 844 286 1056 297 nw
tri 1390 291 1393 297 ne
rect 1393 292 1465 297
tri 1465 292 1481 318 sw
rect 1552 326 1633 339
rect 1552 322 1630 326
tri 1630 322 1633 326 nw
rect 1552 320 1623 322
tri 1623 320 1630 322 nw
rect 1552 306 1558 320
tri 1558 306 1623 320 nw
rect 1552 305 1554 306
tri 1554 305 1558 306 nw
rect 1393 291 1481 292
tri 1393 286 1397 291 ne
rect 1397 286 1481 291
rect 793 284 839 286
tri 839 284 844 286 nw
rect 793 283 827 284
rect 244 282 271 283
tri 271 282 272 283 nw
tri 539 282 551 283 ne
rect 551 282 611 283
rect 244 269 265 282
tri 265 270 271 282 nw
tri 554 280 557 282 ne
rect 557 280 611 282
tri 557 270 559 280 ne
rect 559 270 611 280
tri 611 270 616 283 sw
rect 244 257 254 269
rect 205 254 254 257
tri 108 249 110 251 se
rect 110 249 148 251
tri 105 247 108 249 se
rect 108 247 110 249
rect 105 246 110 247
tri 105 216 107 246 ne
rect 107 215 110 246
rect 144 246 148 249
tri 148 246 153 251 sw
rect 204 249 254 254
rect 204 246 206 249
rect 144 215 153 246
tri 153 215 161 246 sw
tri 204 216 206 246 ne
rect 240 246 254 249
tri 254 247 265 269 nw
rect 559 269 616 270
tri 788 270 791 283 se
rect 791 272 827 283
tri 827 272 839 284 nw
tri 1397 283 1400 286 ne
rect 1400 285 1481 286
tri 1481 285 1486 291 sw
rect 1400 283 1486 285
tri 1400 282 1402 283 ne
rect 1402 282 1486 283
tri 1171 280 1173 282 se
tri 1173 280 1204 282 sw
tri 1402 280 1404 282 ne
rect 1404 280 1486 282
tri 1166 272 1171 280 se
rect 1171 272 1175 280
rect 791 270 823 272
tri 559 249 563 269 ne
rect 563 255 616 269
tri 616 255 621 269 sw
rect 563 253 621 255
tri 783 254 788 269 se
rect 788 254 823 270
tri 823 254 827 272 nw
tri 1157 257 1166 272 se
rect 1166 257 1175 272
tri 1154 256 1157 257 se
rect 1157 256 1175 257
tri 1139 255 1151 256 se
rect 1151 255 1175 256
tri 1137 254 1139 255 se
rect 1139 254 1175 255
tri 621 253 622 254 sw
rect 783 253 823 254
rect 563 249 622 253
tri 622 249 623 253 sw
tri 782 250 783 253 se
rect 783 250 822 253
tri 822 250 823 253 nw
tri 869 253 871 254 se
rect 871 253 909 254
rect 869 252 909 253
tri 909 252 913 254 sw
tri 1115 253 1129 254 se
rect 1129 253 1175 254
rect 869 251 913 252
tri 1090 251 1115 253 se
rect 1115 251 1175 253
tri 689 249 720 250 se
tri 295 247 302 249 se
tri 293 246 295 247 se
rect 295 246 302 247
tri 395 248 397 249 se
rect 397 248 398 249
tri 394 247 395 248 se
rect 395 247 398 248
rect 240 219 241 246
tri 241 219 254 246 nw
tri 377 223 394 247 se
rect 394 223 398 247
tri 373 216 377 223 se
rect 377 217 398 223
tri 493 233 494 248 se
rect 377 216 395 217
tri 372 215 373 216 se
rect 373 215 395 216
rect 107 212 161 215
tri 161 212 162 215 sw
tri 370 212 372 215 se
rect 372 212 395 215
rect 107 211 162 212
tri 162 211 163 212 sw
tri 107 207 108 211 ne
rect 108 207 163 211
tri 163 207 164 211 sw
tri 366 207 369 211 se
rect 369 207 395 212
rect 108 204 164 207
tri 164 204 165 207 sw
tri 364 205 366 207 se
rect 366 205 395 207
tri 108 194 112 204 ne
rect 112 200 165 204
tri 165 200 166 204 sw
tri 361 200 364 204 se
rect 364 200 395 205
rect 112 195 166 200
tri 166 195 171 200 sw
tri 359 198 361 200 se
rect 361 198 395 200
tri 355 195 359 198 se
rect 359 195 395 198
rect 112 194 171 195
tri 171 194 176 195 sw
tri 354 194 355 195 se
rect 355 194 395 195
tri 112 190 114 194 ne
rect 114 190 176 194
tri 176 190 192 194 sw
tri 349 190 354 194 se
rect 354 190 395 194
tri 114 189 115 190 ne
rect 115 189 192 190
tri 192 189 195 190 sw
tri 115 165 125 189 ne
rect 125 183 196 189
tri 196 183 241 189 sw
tri 343 188 349 190 se
rect 349 188 395 190
tri 314 185 343 188 se
rect 343 185 395 188
tri 241 183 292 185 se
rect 292 183 395 185
rect 429 183 432 215
tri 492 217 493 232 se
rect 493 217 494 233
rect 528 248 529 249
tri 529 248 530 249 sw
rect 563 248 590 249
rect 528 228 530 248
tri 530 228 533 248 sw
tri 563 241 564 248 ne
rect 564 241 590 248
tri 564 238 566 241 ne
rect 566 238 590 241
tri 566 228 576 238 ne
rect 576 228 590 238
rect 492 215 494 217
tri 576 216 589 228 ne
rect 589 216 590 228
tri 679 243 686 249 se
rect 782 249 822 250
rect 816 215 817 249
tri 817 230 822 249 nw
rect 903 249 913 251
rect 912 248 913 249
tri 966 248 969 251 se
tri 969 249 1009 251 sw
tri 1071 249 1090 251 se
rect 1090 249 1175 251
tri 1404 271 1418 280 ne
rect 1418 277 1486 280
tri 1486 277 1488 283 sw
rect 1418 271 1488 277
tri 1418 266 1422 271 ne
rect 1422 266 1488 271
tri 1422 256 1426 266 ne
tri 1263 255 1294 256 se
tri 1294 255 1295 256 sw
rect 1426 255 1488 266
rect 1263 254 1295 255
rect 969 248 974 249
tri 912 226 913 248 nw
tri 945 226 966 248 se
rect 966 226 974 248
tri 869 216 870 217 ne
rect 870 216 878 217
tri 870 215 872 216 ne
rect 872 215 878 216
tri 942 220 945 226 se
rect 945 220 974 226
rect 942 215 974 220
rect 1008 215 1009 249
rect 1104 219 1166 249
rect 1104 217 1129 219
tri 1129 217 1162 219 nw
tri 1162 217 1165 219 ne
tri 1104 216 1129 217 nw
rect 1165 216 1166 219
tri 1165 215 1166 216 ne
rect 1200 215 1207 246
tri 1207 219 1209 246 nw
tri 1260 252 1262 254 se
rect 1262 253 1295 254
tri 1295 253 1296 255 sw
rect 1262 252 1296 253
rect 1260 249 1296 252
tri 1426 250 1428 255 ne
rect 1428 250 1488 255
tri 1488 250 1489 266 sw
tri 1355 249 1356 250 se
tri 1356 249 1390 250 sw
tri 1428 249 1429 250 ne
rect 1429 249 1489 250
rect 1260 238 1262 249
rect 492 212 499 215
tri 492 207 493 212 ne
rect 493 207 499 212
tri 493 194 499 207 ne
rect 713 212 716 215
tri 716 212 720 215 nw
rect 942 212 1009 215
tri 713 209 716 212 nw
tri 940 195 942 209 se
rect 942 195 988 212
rect 940 194 988 195
tri 988 194 1009 212 nw
tri 1166 204 1168 215 ne
rect 1168 204 1205 215
tri 1205 204 1207 215 nw
tri 1345 236 1355 249 se
rect 1355 236 1358 249
tri 1335 225 1345 236 se
rect 1345 225 1358 236
tri 1333 221 1335 225 se
rect 1335 221 1358 225
tri 1331 215 1333 221 se
rect 1333 215 1358 221
tri 1429 227 1437 249 ne
rect 1437 227 1454 249
tri 1437 220 1443 227 ne
rect 1443 220 1454 227
tri 1443 215 1454 220 ne
rect 1488 220 1489 249
tri 1488 215 1489 220 nw
tri 1550 249 1595 250 se
tri 1595 249 1596 250 sw
rect 1584 246 1596 249
tri 1596 246 1601 249 sw
rect 1584 215 1601 246
tri 1601 215 1617 246 sw
tri 1328 204 1331 215 se
rect 1331 204 1381 215
tri 1168 194 1171 204 ne
rect 1171 202 1206 204
tri 1206 202 1207 204 sw
tri 1327 202 1328 204 se
rect 1328 202 1381 204
tri 1381 202 1392 215 nw
tri 1550 202 1561 215 ne
rect 1171 194 1207 202
rect 125 180 432 183
rect 125 177 429 180
tri 429 177 432 180 nw
rect 605 188 639 189
rect 125 169 391 177
tri 391 169 429 177 nw
rect 125 165 368 169
tri 368 165 391 169 nw
tri 125 156 129 165 ne
rect 129 158 327 165
tri 327 158 368 165 nw
rect 129 156 318 158
tri 318 156 327 158 nw
tri 129 154 130 156 ne
rect 130 154 312 156
tri 312 154 318 156 nw
tri 639 187 649 189 sw
tri 817 187 874 189 se
tri 874 187 914 189 sw
tri 937 187 940 190 se
rect 940 189 986 194
tri 986 190 988 194 nw
tri 1171 190 1172 194 ne
rect 940 187 985 189
tri 985 187 986 189 nw
rect 1172 189 1207 194
tri 1172 187 1173 189 ne
rect 639 186 649 187
tri 649 186 651 187 sw
tri 788 186 804 187 se
rect 804 186 914 187
tri 914 186 923 187 sw
tri 934 186 936 187 se
rect 936 186 985 187
rect 1173 186 1207 189
tri 1207 186 1244 202 sw
rect 1327 201 1381 202
tri 1322 194 1327 201 se
rect 1327 194 1372 201
tri 1372 194 1381 201 nw
rect 1561 201 1617 215
tri 1561 194 1567 201 ne
rect 1567 197 1617 201
tri 1617 197 1625 215 sw
rect 1567 194 1625 197
tri 1317 187 1322 194 se
rect 1322 189 1366 194
tri 1366 189 1372 194 nw
rect 1322 187 1365 189
tri 1365 187 1366 189 nw
tri 1314 186 1317 187 se
rect 1317 186 1360 187
rect 639 171 651 186
tri 651 171 736 186 sw
rect 781 185 981 186
rect 639 166 736 171
tri 736 166 745 171 sw
rect 639 154 745 166
tri 745 154 750 165 sw
tri 130 152 133 154 ne
rect 133 152 303 154
tri 303 152 311 154 nw
tri 630 152 639 154 ne
rect 639 152 750 154
tri 133 150 141 152 ne
rect 141 151 300 152
tri 300 151 303 152 nw
tri 639 151 641 152 ne
rect 641 151 750 152
tri 750 151 751 154 sw
rect 141 150 296 151
tri 296 150 300 151 nw
tri 641 150 646 151 ne
rect 646 150 751 151
rect 815 176 981 185
tri 981 176 985 186 nw
tri 1018 176 1052 186 se
tri 1052 185 1058 186 sw
rect 1173 185 1244 186
rect 1052 176 1058 185
tri 1058 176 1069 185 sw
tri 1173 176 1175 185 ne
rect 1175 178 1244 185
tri 1244 178 1258 186 sw
tri 1306 181 1314 186 se
rect 1314 181 1360 186
tri 1360 181 1365 187 nw
tri 1301 178 1306 181 se
rect 1306 178 1357 181
rect 1175 177 1258 178
tri 1258 177 1275 178 sw
tri 1297 177 1301 178 se
rect 1301 177 1357 178
tri 1357 177 1360 181 nw
rect 1175 176 1275 177
tri 1275 176 1290 177 sw
tri 1290 176 1297 177 se
rect 1297 176 1356 177
tri 1356 176 1357 177 nw
rect 815 165 978 176
tri 978 166 981 176 nw
tri 1016 172 1018 176 se
rect 1018 172 1069 176
tri 1069 172 1073 176 sw
tri 1175 173 1176 176 ne
rect 1176 173 1354 176
tri 1354 173 1356 176 nw
rect 1176 172 1349 173
rect 1016 171 1073 172
tri 1073 171 1075 172 sw
tri 1176 171 1177 172 ne
rect 1177 171 1349 172
tri 1349 171 1354 173 nw
rect 1016 167 1075 171
tri 1075 167 1077 171 sw
tri 1177 167 1178 171 ne
rect 1016 166 1077 167
rect 815 152 974 165
tri 974 152 978 165 nw
rect 1016 165 1041 166
rect 815 151 972 152
rect 781 150 972 151
tri 972 150 974 152 nw
tri 141 148 150 150 ne
tri 150 148 295 150 nw
tri 648 148 655 150 ne
rect 655 148 751 150
tri 655 147 663 148 ne
rect 663 147 751 148
tri 751 147 753 150 sw
tri 818 147 870 150 ne
rect 870 147 968 150
tri 968 147 972 150 nw
tri 663 144 677 147 ne
rect 677 144 753 147
tri 753 144 754 147 sw
tri 870 144 911 147 ne
rect 911 146 960 147
tri 960 146 966 147 nw
tri 911 144 960 146 nw
tri 677 143 678 144 ne
rect 678 143 754 144
tri 678 142 685 143 ne
rect 685 142 754 143
tri 754 142 755 143 sw
tri 685 138 693 142 ne
rect 693 138 755 142
tri 755 138 757 142 sw
rect 693 137 757 138
tri 37 117 39 131 se
tri 34 101 37 117 se
rect 37 101 39 117
rect 73 128 74 133
tri 74 128 99 133 sw
rect 73 120 99 128
tri 99 120 103 128 sw
rect 73 117 103 120
rect 73 101 102 117
tri 102 101 103 117 nw
rect 254 101 288 117
tri 388 133 450 137 sw
rect 388 131 450 133
tri 450 131 482 133 sw
tri 693 131 702 137 ne
rect 702 131 757 137
tri 757 131 760 138 sw
rect 1075 148 1077 166
tri 1077 148 1079 167 sw
rect 1178 165 1339 171
tri 1339 165 1349 171 nw
tri 1495 165 1496 171 se
tri 1178 162 1182 165 ne
rect 1182 162 1332 165
tri 1332 162 1339 165 nw
tri 1182 148 1281 162 ne
rect 1281 158 1323 162
tri 1323 158 1332 162 nw
rect 1495 160 1496 165
tri 1567 189 1570 194 ne
rect 1570 190 1625 194
tri 1625 190 1631 197 sw
rect 1570 189 1597 190
tri 1530 188 1531 189 sw
rect 1530 181 1531 188
tri 1570 187 1572 189 ne
rect 1572 187 1597 189
tri 1531 181 1532 187 sw
tri 1572 181 1577 187 ne
rect 1577 181 1597 187
rect 1530 167 1532 181
tri 1532 167 1534 181 sw
tri 1577 167 1588 181 ne
rect 1588 167 1597 181
rect 1530 160 1534 167
rect 1495 158 1534 160
tri 1534 158 1536 167 sw
tri 1281 148 1323 158 nw
rect 1495 157 1536 158
tri 1588 157 1595 167 ne
rect 1595 157 1597 167
tri 1495 149 1496 157 ne
rect 1075 134 1079 148
rect 1496 147 1536 157
tri 1079 134 1080 147 sw
rect 1075 132 1080 134
rect 1050 131 1080 132
rect 388 129 486 131
tri 486 129 489 131 sw
rect 388 114 489 129
tri 702 128 704 131 ne
rect 704 128 760 131
tri 760 128 761 131 sw
rect 1016 130 1079 131
tri 1079 130 1080 131 nw
tri 1326 130 1331 132 se
rect 1331 130 1332 132
tri 1016 128 1024 130 ne
rect 1024 129 1077 130
tri 1077 129 1079 130 nw
tri 1322 129 1326 130 se
rect 1326 129 1332 130
rect 1024 128 1073 129
tri 1073 128 1077 129 nw
tri 1320 128 1322 129 se
rect 1322 128 1332 129
tri 704 126 705 128 ne
rect 705 124 761 128
tri 705 118 709 124 ne
rect 709 118 761 124
tri 761 118 766 128 sw
tri 1024 126 1031 128 ne
rect 1031 126 1062 128
tri 1062 126 1073 128 nw
tri 1031 124 1051 126 ne
rect 1051 124 1055 126
tri 1055 124 1062 126 nw
tri 1314 124 1320 128 se
rect 1320 124 1332 128
rect 709 117 766 118
tri 1133 118 1136 124 se
rect 1136 118 1137 124
tri 489 114 490 117 sw
rect 388 103 487 114
tri 487 103 490 114 nw
tri 354 101 359 103 ne
rect 359 101 487 103
tri 33 94 34 100 se
rect 34 99 39 101
rect 34 94 68 99
rect 33 85 68 94
tri 33 71 42 85 ne
rect 42 71 68 85
tri 42 67 46 71 ne
rect 46 67 68 71
tri 359 98 361 101 ne
rect 361 98 446 101
tri 361 79 367 98 ne
rect 367 79 446 98
tri 367 75 372 79 ne
rect 372 75 446 79
tri 372 73 439 75 ne
rect 439 73 446 75
tri 439 71 442 73 ne
rect 442 71 446 73
tri 442 67 446 71 ne
rect 480 98 486 101
tri 486 98 487 101 nw
rect 638 101 672 117
tri 709 116 710 117 ne
rect 710 116 766 117
tri 766 116 767 117 sw
tri 710 101 717 116 ne
rect 717 109 767 116
tri 767 109 770 116 sw
rect 717 102 770 109
tri 770 102 771 109 sw
rect 717 101 771 102
rect 480 75 482 98
tri 482 79 486 98 nw
rect 480 71 481 75
tri 481 73 482 75 nw
tri 480 67 481 71 nw
tri 717 67 734 101 ne
rect 768 70 769 101
tri 769 70 771 101 nw
rect 830 101 864 117
tri 768 68 769 70 nw
tri 1124 101 1133 117 se
rect 1133 101 1137 118
tri 1303 118 1314 124 se
rect 1314 118 1332 124
tri 1171 104 1172 117 sw
tri 46 65 49 67 ne
tri 49 65 101 67 nw
rect 254 17 288 67
rect 638 17 672 67
rect 830 17 864 67
tri 1123 67 1124 100 se
rect 1171 90 1172 104
rect 1214 101 1248 117
tri 1299 109 1303 117 se
rect 1303 109 1332 118
rect 1299 101 1332 109
tri 1366 131 1368 132 sw
rect 1366 117 1368 131
tri 1496 117 1500 147 ne
rect 1500 123 1536 147
tri 1536 123 1541 157 sw
tri 1595 156 1597 157 ne
rect 1500 117 1541 123
rect 1158 67 1172 90
tri 1172 67 1174 100 sw
rect 1123 65 1172 67
tri 1172 65 1174 67 nw
rect 1123 63 1154 65
tri 1154 63 1172 65 nw
tri 1123 61 1127 63 ne
tri 1127 61 1154 63 nw
rect 1214 17 1248 67
tri 1297 67 1299 101 se
rect 1299 67 1310 101
rect 1366 98 1369 117
rect 1344 72 1369 98
rect 1344 67 1368 72
tri 1368 67 1369 72 nw
rect 1406 101 1440 117
tri 1500 101 1502 117 ne
rect 1502 101 1541 117
rect 1536 71 1541 101
rect 1536 67 1539 71
tri 1539 67 1541 71 nw
rect 1594 101 1628 117
rect 1297 66 1368 67
rect 1297 60 1362 66
tri 1362 60 1368 66 nw
tri 1297 56 1304 60 ne
rect 1304 57 1360 60
tri 1360 57 1362 60 nw
rect 1304 56 1357 57
tri 1357 56 1360 57 nw
tri 1304 55 1355 56 ne
tri 1355 55 1357 56 nw
rect 1406 17 1440 67
rect 1594 17 1628 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 354 447 388 453
rect 354 419 384 447
rect 384 419 388 447
rect 660 447 694 449
rect 660 415 672 447
rect 672 415 694 447
rect 1127 412 1161 446
rect 68 345 102 351
rect 68 317 102 345
rect 728 379 762 395
rect 728 361 762 379
rect 881 377 915 411
rect 1060 300 1094 334
rect 1269 306 1303 340
rect 210 257 244 291
rect 1518 305 1552 339
rect 292 215 302 246
rect 302 215 326 246
rect 395 215 398 217
rect 398 215 429 217
rect 292 212 326 215
rect 395 183 429 215
rect 499 215 528 228
rect 528 215 533 228
rect 679 215 686 243
rect 686 215 713 243
rect 869 249 903 251
rect 869 217 878 249
rect 878 217 903 249
rect 1175 249 1209 280
rect 1175 246 1200 249
rect 1200 246 1209 249
rect 499 194 533 215
rect 679 209 713 215
rect 1260 215 1262 238
rect 1262 215 1294 238
rect 1260 204 1294 215
rect 605 154 639 188
rect 781 151 815 185
rect 1041 165 1075 166
rect 39 101 73 133
rect 354 103 388 137
rect 1041 132 1050 165
rect 1050 132 1075 165
rect 1496 160 1530 194
rect 39 99 68 101
rect 68 99 73 101
rect 1137 101 1171 124
rect 1137 90 1158 101
rect 1158 90 1171 101
rect 1332 101 1366 132
rect 1597 156 1631 190
rect 1332 98 1344 101
rect 1344 98 1366 101
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
tri 339 456 391 457 se
tri 338 453 339 456 se
rect 339 455 391 456
tri 391 455 393 457 sw
tri 656 455 678 456 se
rect 678 455 690 456
tri 690 455 691 456 sw
tri 1146 455 1148 456 se
rect 1148 455 1150 456
rect 339 453 393 455
tri 650 453 656 455 se
rect 656 454 691 455
tri 691 454 696 455 sw
rect 656 453 696 454
tri 1136 453 1146 455 se
rect 1146 454 1150 455
tri 1150 454 1160 456 sw
rect 1146 453 1160 454
tri 1160 453 1161 454 sw
tri 337 449 338 453 se
rect 338 449 354 453
tri 336 446 337 449 se
rect 337 446 354 449
rect 388 439 393 453
tri 645 452 650 453 se
rect 650 452 696 453
tri 1133 452 1136 453 se
rect 1136 452 1161 453
tri 640 450 645 452 se
rect 645 451 696 452
tri 696 451 697 452 sw
rect 645 450 697 451
tri 637 449 640 450 se
rect 640 449 697 450
tri 632 447 637 449 se
rect 637 447 660 449
tri 629 446 632 447 se
rect 632 446 660 447
tri 619 442 629 446 se
rect 388 419 392 439
tri 392 435 393 439 nw
tri 601 435 619 442 se
rect 619 435 629 442
tri 560 420 601 435 se
rect 601 420 629 435
rect 380 418 392 419
rect 380 415 390 418
tri 390 415 392 418 nw
tri 546 415 560 420 se
rect 560 415 629 420
rect 694 437 697 449
tri 1121 446 1133 452 se
rect 1133 450 1161 452
tri 1161 450 1166 453 sw
rect 1133 446 1166 450
tri 1114 442 1121 446 se
rect 1121 442 1127 446
tri 697 437 698 442 sw
rect 694 415 698 437
tri 1100 435 1114 442 se
rect 1114 435 1127 442
tri 1083 426 1100 435 se
rect 1100 426 1127 435
tri 380 414 390 415 nw
tri 538 412 544 414 se
rect 544 412 629 415
tri 533 411 538 412 se
rect 538 411 629 412
tri 530 410 533 411 se
rect 533 410 629 411
tri 529 409 530 410 se
rect 530 409 629 410
tri 522 407 529 409 se
rect 529 407 629 409
tri 518 405 522 407 se
rect 522 405 629 407
tri 514 404 518 405 se
rect 518 404 629 405
tri 511 402 514 404 se
rect 514 402 629 404
tri 502 399 508 402 se
rect 508 399 629 402
tri 500 398 501 399 se
rect 501 398 629 399
tri 491 395 499 398 se
rect 499 397 629 398
rect 499 395 621 397
tri 621 395 629 397 nw
tri 468 387 491 395 se
rect 491 387 529 395
tri 111 386 118 387 se
tri 118 386 150 387 sw
tri 464 386 468 387 se
rect 468 386 529 387
tri 109 385 111 386 se
rect 111 385 150 386
tri 150 385 177 386 sw
tri 462 385 464 386 se
rect 464 385 529 386
tri 94 375 109 385 se
rect 109 379 177 385
tri 177 379 317 385 sw
tri 447 379 462 385 se
rect 462 379 529 385
tri 529 379 619 395 nw
rect 681 413 698 415
rect 681 411 696 413
tri 696 411 698 413 nw
tri 877 412 879 414 se
rect 879 412 916 415
tri 916 412 919 415 sw
tri 875 411 877 412 se
rect 877 411 919 412
rect 681 410 692 411
tri 692 410 695 411 nw
tri 871 410 875 411 se
rect 875 410 881 411
rect 681 409 691 410
tri 691 409 692 410 nw
tri 869 409 871 410 se
rect 871 409 881 410
rect 681 407 687 409
tri 687 407 691 409 nw
tri 860 407 869 409 se
rect 869 407 881 409
tri 681 405 687 407 nw
tri 854 405 859 407 se
rect 859 405 881 407
tri 850 404 854 405 se
rect 854 404 881 405
rect 109 378 317 379
tri 317 378 323 379 sw
tri 442 378 447 379 se
rect 447 378 523 379
rect 109 375 323 378
tri 323 375 328 378 sw
tri 441 377 442 378 se
rect 442 377 523 378
tri 523 377 529 379 nw
tri 433 376 441 377 se
rect 441 376 519 377
tri 519 376 522 377 nw
tri 428 375 433 376 se
rect 433 375 518 376
tri 518 375 519 376 nw
tri 70 361 94 375 se
rect 94 374 328 375
tri 328 374 336 375 sw
tri 399 374 416 375 se
rect 416 374 514 375
tri 514 374 518 375 nw
rect 94 361 478 374
tri 478 361 514 374 nw
tri 67 359 70 361 se
rect 70 359 473 361
tri 473 359 478 361 nw
tri 60 354 67 359 se
rect 67 357 462 359
rect 67 354 140 357
tri 140 354 181 357 nw
tri 185 354 244 357 ne
rect 244 354 462 357
tri 462 354 473 359 nw
tri 57 352 60 354 se
rect 60 352 113 354
tri 113 352 140 354 nw
tri 244 352 282 354 ne
rect 282 352 457 354
tri 457 352 461 354 nw
rect 871 377 881 404
rect 915 410 919 411
tri 919 410 920 411 sw
rect 915 404 920 410
tri 920 404 923 410 sw
rect 915 401 923 404
tri 923 401 925 404 sw
rect 915 398 925 401
tri 925 398 928 401 sw
rect 915 395 928 398
tri 928 395 935 398 sw
rect 915 381 935 395
tri 935 381 958 395 sw
rect 915 377 958 381
rect 871 376 958 377
tri 958 376 967 381 sw
rect 871 369 967 376
tri 967 369 978 376 sw
rect 1113 412 1127 426
rect 1161 412 1166 446
rect 1113 410 1166 412
rect 1113 407 1163 410
tri 1163 407 1166 410 nw
rect 1113 405 1152 407
tri 1152 405 1163 407 nw
rect 1113 404 1149 405
tri 1149 404 1152 405 nw
rect 1113 402 1146 404
tri 1146 402 1149 404 nw
rect 1113 401 1141 402
tri 1141 401 1144 402 nw
rect 1113 393 1119 401
tri 1119 393 1141 401 nw
tri 1113 389 1119 393 nw
rect 871 364 978 369
tri 978 364 982 369 sw
rect 871 361 982 364
tri 982 361 983 364 sw
rect 871 359 983 361
tri 983 359 984 361 sw
rect 871 358 984 359
tri 871 357 888 358 ne
rect 888 357 984 358
tri 888 355 904 357 ne
rect 904 355 984 357
tri 910 354 921 355 ne
rect 921 354 984 355
tri 923 352 948 354 ne
rect 948 352 984 354
tri 984 352 987 359 sw
tri 53 350 57 352 se
rect 57 351 111 352
tri 111 351 113 352 nw
tri 282 351 307 352 ne
rect 307 351 451 352
rect 57 350 68 351
tri 48 345 53 350 se
rect 53 345 68 350
tri 47 335 48 340 se
rect 48 335 68 345
rect 47 317 68 335
rect 102 347 109 351
tri 109 349 111 351 nw
tri 307 350 318 351 ne
rect 318 350 451 351
tri 451 350 457 352 nw
tri 948 350 952 352 ne
rect 952 350 987 352
tri 987 350 988 352 sw
tri 318 349 325 350 ne
rect 325 349 450 350
tri 450 349 451 350 nw
rect 952 349 988 350
tri 325 348 338 349 ne
rect 338 348 416 349
tri 416 348 443 349 nw
tri 346 347 353 348 ne
rect 353 347 374 348
tri 374 347 397 348 nw
rect 953 347 988 349
rect 102 344 108 347
tri 108 345 109 347 nw
tri 953 345 954 347 ne
rect 954 345 988 347
tri 988 345 990 349 sw
rect 102 317 106 344
tri 106 336 108 344 nw
rect 954 344 990 345
tri 954 340 956 344 ne
rect 956 340 990 344
tri 990 340 992 344 sw
tri 1057 340 1093 344 se
tri 1093 342 1097 344 sw
rect 1093 340 1097 342
tri 956 336 957 340 ne
rect 47 316 106 317
rect 957 334 992 340
tri 992 334 994 340 sw
tri 1052 334 1057 340 se
rect 1057 334 1097 340
tri 1097 334 1101 342 sw
tri 957 316 963 334 ne
rect 963 316 994 334
rect 46 315 106 316
rect 46 313 103 315
tri 103 313 106 315 nw
tri 552 313 699 316 se
tri 699 315 706 316 sw
rect 964 315 994 316
rect 699 313 706 315
rect 46 312 102 313
tri 102 312 103 313 nw
tri 525 312 552 313 se
rect 552 312 706 313
tri 706 312 720 315 sw
tri 964 312 965 315 ne
rect 46 308 98 312
tri 98 310 102 312 nw
tri 517 311 525 312 se
rect 525 311 720 312
tri 720 311 724 312 sw
rect 965 311 994 315
tri 512 310 517 311 se
rect 517 310 724 311
tri 503 309 512 310 se
rect 512 309 724 310
tri 724 309 736 311 sw
tri 965 309 966 311 ne
rect 966 309 994 311
tri 994 309 1004 334 sw
tri 1052 309 1054 334 ne
rect 46 307 97 308
tri 97 307 98 308 nw
tri 495 307 503 309 se
rect 503 307 736 309
tri 45 300 46 307 se
rect 46 300 95 307
tri 95 300 97 307 nw
tri 211 300 220 307 se
tri 220 306 245 307 sw
tri 490 306 495 307 se
rect 495 306 736 307
rect 220 300 245 306
tri 245 300 252 306 sw
tri 457 300 490 306 se
rect 490 300 736 306
tri 736 300 774 309 sw
tri 966 302 968 309 ne
rect 968 301 1004 309
tri 1004 301 1007 309 sw
rect 968 300 1007 301
rect 1054 300 1060 334
rect 1094 307 1101 334
tri 1101 307 1108 334 sw
rect 1094 300 1108 307
tri 1108 300 1110 305 sw
tri 1269 344 1272 346 se
rect 1272 344 1286 346
tri 1265 343 1269 344 se
rect 1269 343 1286 344
tri 1264 340 1265 342 se
rect 1265 340 1286 343
tri 1514 340 1517 343 se
rect 1517 340 1554 343
tri 1554 340 1556 343 sw
tri 1263 334 1264 339 se
tri 1263 313 1264 334 ne
rect 1264 313 1269 340
tri 1264 309 1265 313 ne
rect 1265 306 1269 313
tri 1338 339 1339 340 sw
rect 1514 339 1556 340
rect 1338 334 1339 339
tri 1339 334 1346 339 sw
rect 1338 326 1346 334
tri 1346 326 1358 334 sw
rect 1338 317 1358 326
tri 1358 317 1365 326 sw
rect 1338 309 1365 317
tri 1365 309 1366 317 sw
rect 1338 308 1366 309
tri 1366 308 1367 309 sw
rect 1265 304 1286 306
rect 45 295 94 300
tri 94 296 95 300 nw
tri 206 296 211 300 se
rect 211 298 252 300
tri 252 298 255 300 sw
tri 451 299 457 300 se
rect 457 299 774 300
tri 774 299 779 300 sw
tri 968 299 969 300 ne
rect 969 299 1007 300
tri 1007 299 1008 300 sw
tri 444 298 451 299 se
rect 451 298 779 299
tri 779 298 785 299 sw
rect 969 298 1008 299
rect 1054 299 1110 300
tri 1175 299 1176 304 se
rect 1176 299 1213 304
rect 211 296 255 298
rect 45 291 93 295
tri 93 292 94 295 nw
tri 204 292 206 295 se
rect 206 292 255 296
tri 428 295 443 298 se
rect 443 295 785 298
tri 785 295 798 298 sw
tri 969 296 970 298 ne
rect 970 295 1008 298
tri 1008 295 1009 298 sw
tri 1054 295 1058 299 ne
rect 1058 295 1110 299
rect 204 291 255 292
tri 44 279 45 291 se
rect 45 279 89 291
tri 89 279 93 291 nw
tri 197 279 204 291 se
rect 204 279 210 291
tri 43 257 44 278 se
rect 44 257 82 279
tri 82 257 89 279 nw
rect 197 276 210 279
rect 244 280 255 291
tri 255 280 256 295 sw
tri 343 280 428 295 se
rect 428 288 798 295
rect 428 287 644 288
tri 644 287 699 288 nw
tri 699 287 705 288 ne
rect 705 287 798 288
tri 798 287 839 295 sw
rect 428 284 555 287
tri 555 284 637 287 nw
tri 706 284 719 287 ne
rect 719 284 839 287
tri 839 284 851 287 sw
tri 866 284 884 286 se
rect 428 283 521 284
tri 521 283 535 284 nw
tri 723 283 725 284 ne
rect 725 283 884 284
rect 428 280 503 283
tri 503 280 521 283 nw
tri 725 280 741 283 ne
rect 741 280 884 283
rect 244 276 256 280
tri 341 279 343 280 se
rect 343 279 495 280
tri 495 279 503 280 nw
tri 741 279 747 280 ne
rect 747 279 884 280
rect 249 273 256 276
tri 256 273 257 279 sw
tri 336 276 340 279 se
rect 340 276 479 279
tri 479 276 495 279 nw
tri 747 276 761 279 ne
rect 761 276 884 279
rect 249 264 253 273
tri 253 264 257 273 nw
tri 330 271 336 276 se
rect 336 271 445 276
tri 445 271 479 276 nw
tri 761 271 792 276 ne
rect 792 271 884 276
tri 329 269 330 271 se
rect 330 269 403 271
tri 324 264 329 269 se
rect 329 264 403 269
tri 403 264 445 271 nw
tri 792 269 803 271 ne
rect 803 269 884 271
tri 803 264 829 269 ne
rect 829 264 884 269
rect 249 257 251 264
tri 251 257 253 264 nw
tri 42 251 43 257 se
rect 43 251 81 257
tri 81 252 82 257 nw
rect 42 246 78 251
tri 78 246 81 251 nw
tri 41 239 42 246 se
rect 42 239 75 246
tri 75 239 78 246 nw
rect 41 231 71 239
tri 71 231 75 239 nw
tri 39 212 41 231 se
rect 41 226 69 231
tri 69 226 71 231 nw
rect 41 214 68 226
tri 68 220 69 226 nw
tri 249 252 251 257 nw
tri 313 253 324 264 se
rect 324 263 395 264
tri 395 263 403 264 nw
tri 829 263 836 264 ne
rect 836 263 884 264
rect 324 259 370 263
tri 370 259 395 263 nw
tri 836 259 843 263 ne
rect 843 259 884 263
rect 324 257 362 259
tri 362 257 370 259 nw
tri 843 257 844 259 ne
rect 844 257 884 259
rect 324 253 355 257
tri 355 253 362 257 nw
tri 844 253 847 257 ne
rect 847 253 884 257
tri 307 250 313 253 se
rect 313 252 353 253
tri 847 252 848 253 ne
rect 313 250 349 252
tri 288 248 291 250 se
rect 291 248 349 250
tri 349 248 353 252 nw
rect 848 251 884 253
tri 970 288 973 295 ne
rect 973 286 1009 295
tri 973 283 974 286 ne
rect 974 281 1009 286
tri 1009 281 1015 295 sw
rect 974 280 1015 281
tri 1058 280 1071 295 ne
rect 1071 281 1110 295
tri 1110 281 1115 299 sw
rect 1071 280 1115 281
tri 1171 282 1175 299 se
rect 1175 282 1213 299
tri 1213 282 1215 304 nw
tri 1265 303 1267 304 ne
rect 1267 302 1286 304
tri 1272 300 1281 302 ne
rect 1281 300 1286 302
rect 1338 303 1367 308
rect 1514 305 1518 339
rect 1552 305 1556 339
tri 1367 303 1368 304 sw
rect 1514 303 1556 305
rect 1338 300 1368 303
tri 1281 297 1294 300 ne
rect 1294 298 1368 300
tri 1368 298 1369 302 sw
rect 1294 297 1369 298
tri 1514 297 1515 302 se
rect 1515 301 1554 303
tri 1554 301 1556 303 nw
rect 1515 297 1548 301
tri 1324 295 1330 297 ne
rect 1330 295 1369 297
tri 1513 295 1514 297 se
rect 1514 296 1548 297
tri 1548 296 1554 301 nw
rect 1514 295 1538 296
tri 1330 287 1341 295 ne
rect 1341 287 1369 295
tri 1341 283 1342 287 ne
rect 1342 283 1369 287
tri 1369 283 1372 295 sw
rect 1342 282 1372 283
tri 1511 287 1513 295 se
rect 1513 287 1538 295
rect 1171 280 1213 282
tri 974 279 975 280 ne
rect 975 279 1015 280
tri 1015 279 1016 280 sw
tri 1071 279 1072 280 ne
rect 1072 279 1115 280
tri 975 271 978 279 ne
rect 978 271 1016 279
tri 1016 271 1019 279 sw
tri 1072 271 1079 279 ne
rect 1079 271 1115 279
tri 1115 271 1118 280 sw
tri 978 269 979 271 ne
rect 979 269 1019 271
tri 979 265 980 269 ne
rect 980 265 1019 269
tri 1019 265 1022 271 sw
tri 1079 265 1082 271 ne
rect 1082 269 1118 271
tri 1118 269 1119 271 sw
rect 980 264 1022 265
rect 1082 264 1119 269
tri 980 258 982 264 ne
rect 982 257 1022 264
tri 1022 257 1024 264 sw
tri 1082 257 1086 264 ne
rect 1086 257 1119 264
tri 982 254 983 257 ne
rect 288 247 349 248
rect 288 246 340 247
tri 68 214 69 220 sw
rect 41 212 69 214
rect 288 212 292 246
rect 326 238 340 246
tri 340 238 349 247 nw
tri 675 245 677 247 se
rect 677 245 702 247
rect 675 243 702 245
tri 848 247 852 251 ne
rect 852 247 869 251
tri 852 244 854 247 ne
rect 854 244 869 247
rect 326 236 339 238
tri 339 236 340 238 nw
rect 326 231 335 236
tri 335 232 339 236 nw
tri 497 231 498 232 se
rect 498 231 533 232
rect 326 229 333 231
tri 333 229 334 231 nw
tri 495 230 497 231 se
rect 497 230 533 231
tri 533 230 536 232 sw
rect 326 212 330 229
tri 330 226 333 229 nw
rect 495 228 536 230
tri 392 226 393 227 se
tri 393 226 436 227 sw
rect 39 209 69 212
tri 69 209 70 212 sw
tri 38 184 39 208 se
rect 39 184 70 209
rect 288 210 330 212
tri 288 208 291 210 ne
rect 291 208 328 210
tri 328 208 330 210 nw
tri 384 219 392 226 se
rect 392 223 436 226
tri 436 223 440 226 sw
rect 392 219 440 223
tri 440 219 443 223 sw
rect 384 218 443 219
tri 443 218 444 219 sw
rect 384 217 405 218
rect 38 183 70 184
tri 70 183 73 208 sw
tri 383 184 384 206 se
rect 384 184 395 217
tri 383 183 385 184 ne
rect 385 183 395 184
tri 37 179 38 180 se
rect 38 179 73 183
tri 385 180 388 183 ne
rect 388 180 405 183
tri 388 179 392 180 ne
rect 392 179 405 180
rect 37 174 73 179
tri 392 178 397 179 ne
rect 397 178 405 179
tri 73 174 74 178 sw
tri 397 176 405 178 ne
tri 36 154 37 172 se
rect 37 158 74 174
tri 74 158 76 172 sw
tri 536 219 537 228 sw
rect 536 191 537 219
rect 675 209 679 243
tri 854 242 856 244 ne
rect 856 241 869 244
tri 856 239 858 241 ne
rect 858 239 869 241
rect 983 251 1024 257
tri 983 248 985 251 ne
rect 985 248 1024 251
tri 1024 248 1028 257 sw
rect 985 247 1028 248
tri 1086 247 1091 257 ne
rect 1091 249 1119 257
tri 1119 249 1124 269 sw
rect 986 246 1028 247
rect 1091 246 1124 249
tri 1170 259 1171 269 se
rect 1171 259 1175 280
rect 1170 247 1175 259
tri 1170 246 1171 247 ne
rect 1171 246 1175 247
rect 1209 246 1213 280
tri 1342 277 1344 282 ne
rect 1344 277 1372 282
tri 1372 277 1373 282 sw
tri 1510 278 1511 282 se
rect 1511 278 1538 287
tri 986 244 987 246 ne
rect 987 242 1028 246
tri 987 241 988 242 ne
tri 858 230 865 239 ne
rect 865 217 869 239
rect 903 231 909 240
tri 909 231 918 240 nw
rect 988 239 1028 242
tri 1028 239 1032 246 sw
tri 1091 239 1095 246 ne
rect 1095 241 1124 246
tri 1124 241 1126 246 sw
tri 1171 243 1175 246 ne
rect 1175 245 1213 246
rect 1175 243 1211 245
tri 1211 243 1213 245 nw
tri 1344 244 1347 277 ne
rect 1347 243 1373 277
tri 1373 243 1380 277 sw
tri 1175 242 1199 243 ne
rect 1199 242 1211 243
rect 988 238 1032 239
rect 1095 238 1126 241
tri 1126 238 1127 241 sw
tri 1255 238 1259 242 se
rect 1259 239 1296 242
tri 1296 239 1298 242 sw
rect 1259 238 1298 239
tri 988 236 989 238 ne
rect 989 237 1032 238
tri 1032 237 1033 238 sw
rect 989 236 1033 237
tri 1095 236 1096 238 ne
rect 1096 236 1127 238
tri 989 232 990 236 ne
rect 990 232 1033 236
tri 1033 232 1034 236 sw
tri 1096 232 1099 236 ne
tri 990 231 991 232 ne
rect 991 231 1034 232
tri 1034 231 1035 232 sw
rect 1099 231 1127 236
rect 903 217 907 231
tri 907 228 909 231 nw
tri 991 228 992 231 ne
rect 992 228 1035 231
rect 865 215 907 217
tri 865 213 867 215 ne
rect 867 213 904 215
tri 904 213 907 215 nw
tri 992 213 996 228 ne
rect 996 220 1035 228
tri 1035 220 1039 231 sw
tri 1099 220 1104 231 ne
rect 1104 220 1127 231
rect 996 213 1039 220
tri 996 210 997 213 ne
rect 675 207 702 209
tri 675 205 677 207 ne
rect 677 205 702 207
rect 997 209 1039 213
tri 997 207 998 209 ne
rect 998 205 1039 209
tri 998 203 1000 205 ne
rect 1000 204 1039 205
tri 1039 204 1050 220 sw
rect 1000 202 1050 204
tri 778 191 782 195 se
rect 782 191 785 195
tri 777 186 778 187 se
rect 778 186 785 191
rect 777 185 785 186
tri 1000 196 1002 202 ne
rect 1002 195 1050 202
tri 1050 195 1056 204 sw
rect 1002 194 1056 195
tri 1104 194 1117 220 ne
rect 1117 205 1127 220
tri 1127 205 1143 238 sw
tri 1254 236 1255 238 se
rect 1255 236 1260 238
rect 1117 195 1143 205
rect 1294 204 1298 238
rect 1347 241 1380 243
tri 1502 243 1510 277 se
rect 1510 267 1538 278
tri 1538 267 1548 296 nw
rect 1510 243 1536 267
tri 1347 228 1348 241 ne
rect 1348 227 1380 241
tri 1380 227 1383 241 sw
tri 1499 227 1502 241 se
rect 1502 227 1536 243
tri 1348 223 1349 227 ne
rect 1349 222 1383 227
tri 1383 222 1384 227 sw
tri 1498 222 1499 227 se
rect 1499 222 1536 227
tri 1298 215 1299 222 sw
tri 1298 211 1299 215 nw
rect 1349 219 1384 222
tri 1384 219 1385 222 sw
tri 1497 219 1498 222 se
rect 1498 219 1536 222
tri 1536 219 1538 267 nw
rect 1349 212 1385 219
tri 1385 212 1387 219 sw
rect 1349 211 1387 212
tri 1496 212 1497 219 se
rect 1497 212 1536 219
rect 1496 211 1536 212
tri 1349 205 1350 211 ne
tri 1143 195 1148 204 sw
rect 1117 194 1148 195
tri 1002 192 1003 194 ne
rect 37 154 76 158
rect 601 157 605 161
rect 36 152 76 154
tri 76 152 77 154 sw
tri 35 148 36 151 se
rect 36 148 77 152
tri 601 151 603 157 ne
rect 603 154 605 157
rect 639 157 643 161
rect 639 154 641 157
rect 603 152 641 154
tri 641 152 643 157 nw
rect 603 151 626 152
tri 626 151 641 152 nw
rect 777 151 781 185
rect 1003 191 1056 194
tri 1056 191 1059 194 sw
tri 1117 191 1119 194 ne
rect 1119 191 1148 194
tri 1148 191 1150 194 sw
tri 1003 167 1011 191 ne
rect 1011 175 1059 191
tri 1059 175 1070 191 sw
tri 1119 175 1122 191 ne
rect 1011 171 1070 175
tri 1070 171 1073 175 sw
rect 1122 171 1150 191
rect 1011 170 1073 171
tri 1073 170 1077 171 sw
tri 1122 170 1123 171 ne
rect 1123 170 1150 171
rect 1011 167 1077 170
tri 1077 167 1079 170 sw
rect 1011 166 1079 167
tri 891 151 906 157 se
rect 777 150 785 151
tri 888 150 891 151 se
rect 891 150 906 151
tri 777 148 781 150 ne
rect 781 148 820 150
tri 820 148 821 150 nw
tri 884 148 888 150 se
rect 888 148 906 150
rect 35 146 77 148
tri 781 147 790 148 ne
rect 790 147 816 148
tri 816 147 818 148 nw
tri 880 147 882 148 se
rect 882 147 906 148
tri 77 146 78 147 sw
tri 34 133 35 137 se
rect 35 133 78 146
tri 863 141 879 147 se
rect 879 141 906 147
tri 350 139 352 141 se
rect 352 139 389 141
tri 389 139 392 141 sw
tri 859 140 863 141 se
rect 863 140 906 141
tri 718 139 728 140 se
tri 728 139 729 140 sw
rect 350 137 392 139
tri 711 138 715 139 se
rect 715 138 729 139
rect 350 135 354 137
rect 388 135 392 137
tri 392 135 458 138 se
tri 458 135 522 138 sw
tri 694 135 711 138 se
rect 711 135 729 138
rect 34 99 39 133
rect 73 99 78 133
rect 34 98 78 99
tri 34 95 37 98 ne
rect 37 95 75 98
tri 75 95 78 98 nw
rect 397 132 522 135
tri 522 132 579 135 sw
tri 680 132 694 135 se
rect 694 132 729 135
tri 729 132 748 139 sw
tri 851 134 859 139 se
rect 859 134 906 140
rect 397 131 579 132
tri 579 131 583 132 sw
tri 672 131 680 132 se
rect 680 131 748 132
rect 397 129 583 131
tri 583 129 587 131 sw
tri 665 129 672 131 se
rect 672 129 748 131
rect 397 126 587 129
tri 587 126 598 129 sw
tri 656 128 665 129 se
rect 665 128 748 129
tri 748 128 760 132 sw
tri 845 128 851 134 se
rect 851 128 906 134
tri 651 126 656 128 se
rect 656 126 760 128
rect 397 125 598 126
tri 598 125 600 126 sw
tri 648 125 651 126 se
rect 651 125 760 126
rect 397 124 600 125
tri 600 124 621 125 sw
tri 646 124 648 125 se
rect 648 124 760 125
tri 760 124 769 128 sw
tri 839 124 845 127 se
rect 845 124 906 128
rect 397 123 621 124
tri 621 123 633 124 sw
tri 633 123 646 124 se
rect 646 123 769 124
tri 769 123 771 124 sw
tri 838 123 839 124 se
rect 839 123 906 124
rect 397 121 771 123
tri 771 121 777 123 sw
tri 825 121 837 123 se
rect 837 121 906 123
rect 397 120 777 121
tri 777 120 795 121 sw
tri 816 120 825 121 se
rect 825 120 906 121
rect 397 119 795 120
tri 795 119 804 120 sw
tri 804 119 811 120 se
rect 811 119 906 120
rect 397 116 906 119
rect 397 115 880 116
tri 880 115 906 116 nw
rect 397 113 871 115
tri 871 113 879 115 nw
rect 397 109 863 113
rect 397 108 480 109
tri 480 108 488 109 nw
tri 508 108 519 109 ne
rect 519 108 863 109
rect 397 103 452 108
tri 452 103 480 108 nw
tri 519 103 554 108 ne
rect 554 105 686 108
tri 686 105 697 108 nw
tri 724 105 738 108 ne
rect 738 105 863 108
tri 863 105 871 113 nw
tri 1011 162 1013 166 ne
rect 1013 161 1041 166
tri 1013 159 1014 161 ne
rect 1014 157 1041 161
tri 1014 134 1022 157 ne
rect 1022 147 1041 157
rect 1075 147 1079 166
tri 1123 164 1124 170 ne
rect 1124 160 1150 170
tri 1150 160 1165 191 sw
rect 1292 202 1298 204
rect 1292 200 1296 202
tri 1296 200 1298 202 nw
rect 1350 203 1387 211
tri 1387 203 1388 211 sw
rect 1350 202 1388 203
tri 1388 202 1389 203 sw
tri 1292 199 1296 200 nw
rect 1350 198 1389 202
tri 1350 197 1351 198 ne
rect 1351 196 1389 198
tri 1389 196 1390 198 sw
rect 1351 191 1390 196
tri 1351 168 1353 191 ne
rect 1353 183 1390 191
tri 1390 183 1393 194 sw
tri 1351 161 1353 168 se
rect 1353 165 1393 183
tri 1393 165 1394 183 sw
rect 1353 161 1394 165
rect 1351 160 1394 161
tri 1394 160 1397 165 sw
tri 1594 193 1595 194 se
rect 1595 193 1632 194
tri 1593 191 1594 193 se
rect 1594 191 1632 193
tri 1632 191 1635 194 sw
rect 1593 190 1635 191
tri 1591 187 1593 190 se
rect 1593 187 1597 190
tri 1578 161 1591 187 se
rect 1591 161 1597 187
rect 1022 134 1033 147
tri 1022 132 1023 134 ne
rect 1023 132 1033 134
tri 1023 131 1024 132 ne
rect 1024 131 1033 132
tri 1024 124 1028 131 ne
rect 1028 124 1033 131
tri 1028 120 1032 124 ne
rect 1032 119 1033 124
tri 1032 118 1033 119 ne
rect 554 103 681 105
tri 681 103 686 105 nw
tri 738 103 744 105 ne
rect 744 103 860 105
tri 860 103 863 105 nw
rect 397 100 431 103
tri 431 100 452 103 nw
tri 554 100 581 103 ne
rect 581 100 669 103
tri 669 100 681 103 nw
tri 744 101 755 103 ne
rect 755 101 852 103
tri 755 100 758 101 ne
rect 758 100 852 101
tri 852 100 860 103 nw
rect 397 98 419 100
tri 419 98 431 100 nw
tri 581 98 597 100 ne
rect 597 98 662 100
tri 662 98 669 100 nw
tri 758 98 765 100 ne
rect 765 98 847 100
tri 847 98 852 100 nw
rect 397 97 415 98
tri 415 97 419 98 nw
tri 597 97 601 98 ne
rect 601 97 659 98
tri 659 97 662 98 nw
tri 765 97 767 98 ne
rect 767 97 841 98
rect 397 96 408 97
tri 408 96 415 97 nw
tri 601 96 611 97 ne
rect 611 96 653 97
tri 653 96 659 97 nw
tri 767 96 771 97 ne
rect 771 96 841 97
tri 841 96 847 98 nw
rect 397 95 403 96
tri 403 95 408 96 nw
tri 611 95 617 96 ne
rect 617 95 642 96
tri 397 94 403 95 nw
tri 617 94 642 95 ne
tri 642 94 653 96 nw
tri 771 94 777 96 ne
rect 777 94 829 96
rect 779 93 829 94
tri 829 93 841 96 nw
tri 1350 158 1351 160 se
rect 1351 158 1397 160
tri 1348 156 1350 158 se
rect 1350 157 1397 158
tri 1397 157 1400 160 sw
tri 1577 159 1578 160 se
rect 1578 159 1597 161
tri 1492 158 1493 159 ne
rect 1493 157 1532 159
rect 1350 156 1403 157
tri 1403 156 1405 157 sw
rect 1494 156 1532 157
tri 1532 156 1534 159 nw
tri 1575 156 1577 159 se
rect 1577 156 1597 159
rect 1631 156 1635 190
tri 1346 153 1348 156 se
rect 1348 153 1405 156
tri 1339 146 1346 153 se
rect 1346 146 1405 153
tri 1329 135 1339 146 se
rect 1339 135 1405 146
tri 1405 135 1473 156 sw
tri 1558 137 1575 155 se
rect 1575 154 1635 156
rect 1575 152 1632 154
tri 1632 152 1635 154 nw
rect 1575 151 1625 152
tri 1625 151 1632 152 nw
rect 1575 149 1619 151
tri 1619 149 1625 151 nw
rect 1575 137 1608 149
tri 1608 137 1619 149 nw
tri 1552 135 1558 137 se
rect 1558 135 1592 137
rect 1329 132 1473 135
tri 782 92 785 93 ne
rect 785 92 818 93
tri 818 92 828 93 nw
rect 1133 90 1137 108
rect 1171 90 1175 108
tri 1328 128 1329 132 se
rect 1329 128 1332 132
rect 1328 98 1332 128
rect 1366 129 1473 132
tri 1473 129 1493 135 sw
tri 1529 129 1552 135 se
rect 1552 129 1592 135
rect 1366 121 1592 129
tri 1592 121 1608 137 nw
rect 1366 117 1582 121
tri 1582 117 1592 121 nw
rect 1366 115 1576 117
tri 1576 115 1582 117 nw
rect 1366 114 1536 115
rect 1366 113 1402 114
tri 1402 113 1415 114 nw
tri 1415 113 1422 114 ne
rect 1422 113 1536 114
rect 1366 103 1382 113
tri 1382 103 1402 113 nw
tri 1422 103 1488 113 ne
rect 1488 103 1536 113
rect 1366 102 1381 103
tri 1381 102 1382 103 nw
tri 1488 102 1536 103 ne
tri 1536 102 1576 115 nw
rect 1366 98 1371 102
rect 1328 97 1371 98
tri 1371 97 1381 102 nw
rect 1328 96 1370 97
tri 1328 94 1330 96 ne
rect 1330 94 1368 96
tri 1368 94 1370 96 nw
rect 1133 89 1175 90
tri 1133 86 1135 89 ne
rect 1135 86 1172 89
tri 1172 86 1175 89 nw
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< via1 >>
rect 328 419 354 446
rect 354 419 380 446
rect 328 394 380 419
rect 629 415 660 446
rect 660 415 681 446
rect 629 394 681 415
rect 714 395 766 405
rect 714 361 728 395
rect 728 361 762 395
rect 762 361 766 395
rect 714 353 766 361
rect 819 352 871 404
rect 1061 374 1113 426
rect 1171 304 1223 356
rect 1286 340 1338 352
rect 1286 306 1303 340
rect 1303 306 1338 340
rect 197 257 210 276
rect 210 257 244 276
rect 244 257 249 276
rect 197 224 249 257
rect 884 251 936 292
rect 1286 300 1338 306
rect 702 243 754 248
rect 405 217 457 218
rect 405 183 429 217
rect 429 183 457 217
rect 405 166 457 183
rect 484 194 499 228
rect 499 194 533 228
rect 533 194 536 228
rect 484 176 536 194
rect 597 188 649 213
rect 702 209 713 243
rect 713 209 754 243
rect 884 240 903 251
rect 903 240 936 251
rect 702 196 754 209
rect 597 161 605 188
rect 605 161 639 188
rect 639 161 649 188
rect 785 185 837 202
rect 1240 204 1260 236
rect 1260 204 1292 236
rect 785 151 815 185
rect 815 151 837 185
rect 785 150 837 151
rect 345 103 354 135
rect 354 103 388 135
rect 388 103 397 135
rect 906 112 958 164
rect 1240 184 1292 204
rect 1490 194 1542 211
rect 1490 160 1496 194
rect 1496 160 1530 194
rect 1530 160 1542 194
rect 1033 132 1041 147
rect 1041 132 1075 147
rect 1075 132 1085 147
rect 345 83 397 103
rect 1033 95 1085 132
rect 1123 124 1175 160
rect 1490 159 1542 160
rect 1123 108 1137 124
rect 1137 108 1171 124
rect 1171 108 1175 124
<< metal2 >>
tri 1080 495 1086 496 se
tri 1086 495 1089 496 sw
tri 1000 490 1080 495 se
rect 1080 491 1089 495
tri 1089 491 1125 495 sw
rect 1080 490 1125 491
tri 1125 490 1127 491 sw
tri 732 482 1000 490 se
rect 1000 482 1127 490
tri 1127 482 1144 490 sw
tri 721 479 732 482 se
rect 732 479 1145 482
tri 1145 479 1149 482 sw
tri 683 468 721 479 se
rect 721 477 1149 479
tri 1149 477 1151 479 sw
rect 721 468 1151 477
tri 1151 468 1157 477 sw
tri 650 457 683 468 se
rect 683 466 1055 468
tri 1055 466 1102 468 nw
tri 1102 466 1111 468 ne
rect 1111 466 1157 468
rect 683 462 950 466
tri 950 462 1055 466 nw
tri 1111 462 1121 466 ne
rect 1121 462 1157 466
tri 1157 462 1160 468 sw
rect 683 457 730 462
tri 645 454 650 457 se
rect 650 454 730 457
tri 644 453 645 454 se
rect 645 453 730 454
tri 730 453 950 462 nw
tri 1121 453 1132 462 ne
rect 1132 453 1160 462
tri 643 451 644 453 se
rect 644 451 721 453
tri 721 451 729 453 nw
tri 1133 451 1134 453 ne
rect 1134 451 1160 453
tri 639 446 643 451 se
rect 643 446 701 451
rect 681 439 701 446
tri 701 439 721 451 nw
tri 1134 439 1142 451 ne
rect 1142 444 1160 451
tri 1160 444 1170 462 sw
rect 1142 439 1170 444
rect 681 436 697 439
tri 697 436 701 439 nw
tri 1142 436 1143 439 ne
rect 1143 436 1170 439
rect 681 426 682 436
tri 682 426 697 436 nw
tri 1143 426 1150 436 ne
rect 1150 426 1170 436
tri 681 424 682 426 nw
rect 332 352 367 394
tri 367 365 368 394 nw
tri 712 372 714 377 se
tri 708 369 712 372 se
rect 712 369 714 372
tri 701 365 708 369 se
rect 708 365 714 369
tri 693 361 701 365 se
rect 701 361 714 365
tri 680 353 693 361 se
rect 693 353 714 361
tri 816 361 819 378 se
tri 815 360 816 361 se
rect 816 360 819 361
tri 813 357 815 360 se
rect 815 357 819 360
tri 811 353 813 357 se
rect 813 353 819 357
tri 678 352 680 353 se
rect 680 352 733 353
tri 733 352 734 353 nw
tri 810 352 811 353 se
rect 811 352 819 353
tri 1060 394 1061 398 se
tri 1054 374 1060 393 se
rect 1060 374 1061 394
tri 1150 421 1153 426 ne
rect 1153 421 1170 426
rect 1154 420 1170 421
tri 1154 419 1155 420 ne
rect 1155 419 1170 420
tri 1155 416 1157 419 ne
rect 1157 416 1170 419
tri 1157 410 1159 416 ne
rect 1159 410 1170 416
tri 1170 410 1187 444 sw
tri 1159 383 1164 410 ne
rect 1164 382 1187 410
tri 1164 377 1165 382 ne
rect 1165 374 1187 382
tri 1049 359 1054 374 se
rect 1054 359 1093 374
rect 1049 356 1093 359
tri 1093 357 1101 374 nw
tri 1165 357 1170 374 ne
rect 1170 360 1187 374
tri 1187 360 1208 410 sw
tri 1047 352 1049 356 se
rect 1049 352 1070 356
rect 332 292 365 352
tri 365 304 367 352 nw
tri 672 348 678 352 se
rect 678 348 726 352
tri 726 348 733 352 nw
tri 808 348 810 352 se
rect 810 351 855 352
rect 810 348 831 351
tri 661 341 672 348 se
rect 672 341 713 348
tri 713 341 726 348 nw
tri 804 341 808 348 se
rect 808 341 831 348
tri 638 329 661 341 se
rect 661 338 708 341
tri 708 338 713 341 nw
rect 661 329 692 338
tri 692 329 708 338 nw
tri 796 329 804 341 se
rect 804 329 831 341
tri 635 324 638 329 se
rect 638 324 684 329
tri 684 324 692 329 nw
tri 793 324 796 329 se
rect 796 324 831 329
tri 631 312 635 324 se
rect 635 317 670 324
tri 670 317 684 324 nw
tri 788 317 793 324 se
rect 793 317 831 324
rect 635 312 664 317
tri 664 312 670 317 nw
tri 786 312 788 316 se
rect 788 312 831 317
tri 831 312 855 351 nw
tri 629 304 631 312 se
rect 631 304 661 312
tri 661 304 664 312 nw
tri 779 304 785 312 se
rect 785 304 827 312
tri 827 305 831 312 nw
tri 628 301 629 304 se
rect 629 301 660 304
tri 660 301 661 304 nw
tri 777 301 779 304 se
rect 779 301 825 304
tri 825 301 827 304 nw
rect 628 300 660 301
tri 776 300 777 301 se
rect 777 300 825 301
tri 626 293 628 300 se
rect 628 293 657 300
tri 657 293 660 300 nw
tri 771 293 776 300 se
rect 776 297 823 300
tri 823 297 825 300 nw
rect 776 293 816 297
tri 816 293 823 297 nw
rect 626 292 657 293
tri 769 292 771 293 se
rect 771 292 815 293
tri 815 292 816 293 nw
tri 1035 312 1047 351 se
rect 1047 312 1070 352
tri 1034 310 1035 312 se
rect 1035 310 1070 312
tri 1033 305 1034 307 se
rect 1034 305 1070 310
tri 1070 305 1093 356 nw
rect 1170 356 1208 360
tri 1208 356 1211 360 sw
rect 1170 354 1171 356
tri 1170 349 1171 354 ne
rect 1033 304 1070 305
tri 1032 302 1033 304 se
rect 1033 302 1066 304
tri 1031 300 1032 301 se
rect 1032 300 1066 302
tri 1030 297 1031 300 se
rect 1031 297 1066 300
tri 1029 294 1030 297 se
rect 1030 296 1066 297
tri 1066 296 1070 304 nw
rect 1030 294 1049 296
tri 332 281 333 292 ne
tri 249 267 251 268 sw
rect 249 248 251 267
tri 251 248 282 267 sw
rect 249 244 282 248
tri 282 244 289 248 sw
tri 210 218 214 224 ne
rect 214 218 243 224
tri 214 200 228 218 ne
rect 228 200 243 218
tri 228 193 243 200 ne
rect 333 228 363 292
tri 363 248 365 292 nw
tri 618 266 626 292 se
rect 626 266 649 292
tri 649 266 657 292 nw
tri 727 266 769 292 se
rect 769 271 785 292
tri 785 271 815 292 nw
rect 769 266 779 271
tri 779 266 785 271 nw
tri 613 248 618 266 se
rect 618 265 648 266
tri 648 265 649 266 nw
rect 618 248 645 265
tri 645 248 648 265 nw
tri 716 249 727 265 se
rect 727 261 771 266
tri 771 261 779 266 nw
rect 727 249 755 261
rect 716 248 755 249
tri 755 248 771 261 nw
tri 1028 292 1029 293 se
rect 1029 292 1049 294
tri 1022 271 1028 291 se
rect 1028 271 1049 292
tri 1019 259 1022 270 se
rect 1022 259 1049 271
tri 1018 257 1019 259 se
rect 1019 257 1049 259
tri 1049 257 1066 296 nw
rect 333 193 362 228
tri 362 218 363 228 nw
tri 611 241 613 248 se
rect 613 247 645 248
rect 613 241 644 247
tri 644 241 645 247 nw
rect 611 238 644 241
tri 608 228 611 238 se
rect 611 228 639 238
tri 443 218 447 228 sw
tri 333 192 334 193 ne
rect 334 190 362 193
tri 334 189 335 190 ne
rect 335 189 362 190
tri 335 171 338 189 ne
rect 338 168 362 189
tri 362 168 365 188 sw
tri 398 182 405 188 ne
rect 338 166 365 168
tri 365 166 366 168 sw
tri 606 221 608 228 se
rect 608 221 639 228
tri 605 219 606 221 se
rect 606 219 639 221
tri 604 214 605 218 se
rect 605 214 639 219
rect 604 213 639 214
tri 639 213 644 238 nw
tri 536 185 539 195 sw
rect 536 183 539 185
tri 539 183 540 185 sw
rect 536 177 540 183
tri 540 177 541 182 sw
rect 536 176 541 177
tri 497 174 499 176 ne
rect 499 173 541 176
tri 499 168 502 173 ne
rect 502 168 541 173
tri 541 168 544 177 sw
tri 338 165 339 166 ne
rect 339 161 366 166
tri 366 161 369 166 sw
tri 503 162 506 168 ne
rect 506 166 544 168
tri 544 166 545 168 sw
rect 506 161 545 166
tri 545 161 546 164 sw
tri 754 247 755 248 nw
tri 936 256 938 257 nw
tri 1017 256 1018 257 se
rect 1018 256 1044 257
tri 1014 254 1017 256 se
rect 1017 254 1044 256
tri 1005 245 1014 254 se
rect 1014 247 1044 254
tri 1044 247 1049 257 nw
rect 1014 245 1035 247
tri 999 240 1005 245 se
rect 1005 240 1035 245
tri 995 236 999 240 se
rect 999 236 1035 240
tri 1035 236 1044 247 nw
tri 979 221 995 236 se
rect 995 221 1023 236
tri 1023 221 1035 236 nw
tri 972 214 979 221 se
rect 979 214 1018 221
tri 1018 214 1023 221 nw
tri 966 209 972 214 se
rect 972 209 995 214
tri 960 203 966 209 se
rect 966 203 995 209
tri 649 177 656 190 sw
rect 649 174 656 177
tri 656 174 658 177 sw
rect 649 170 658 174
tri 658 170 659 173 sw
rect 649 168 659 170
tri 659 168 660 170 sw
rect 649 161 661 168
tri 339 153 341 161 ne
rect 341 151 369 161
tri 369 151 376 161 sw
tri 506 160 507 161 ne
rect 507 160 546 161
tri 610 160 611 161 ne
rect 611 160 661 161
tri 507 156 509 160 ne
rect 509 157 546 160
tri 546 157 547 160 sw
rect 509 156 547 157
tri 611 156 614 160 ne
rect 614 156 661 160
rect 341 150 376 151
tri 509 150 513 156 ne
rect 513 151 547 156
tri 547 151 549 156 sw
rect 513 150 549 151
tri 614 150 617 156 ne
rect 617 150 661 156
tri 661 150 669 166 sw
tri 783 152 785 160 se
rect 783 150 785 152
tri 956 199 959 202 se
rect 959 199 995 203
tri 954 198 956 199 se
rect 956 198 995 199
tri 953 196 954 198 se
rect 954 196 995 198
tri 949 193 953 196 se
rect 953 193 995 196
tri 939 184 949 193 se
rect 949 184 995 193
tri 995 185 1018 214 nw
tri 1514 234 1515 235 se
tri 1510 227 1514 233 se
rect 1514 227 1515 234
tri 1508 225 1510 227 se
rect 1510 225 1515 227
tri 1506 221 1508 225 se
rect 1508 221 1515 225
tri 1501 214 1506 221 se
rect 1506 214 1515 221
tri 1499 211 1501 214 se
rect 1501 211 1515 214
tri 928 173 939 184 se
rect 939 173 979 184
tri 922 168 928 173 se
rect 928 168 979 173
tri 917 164 922 168 se
rect 922 164 979 168
tri 979 164 995 184 nw
tri 1236 166 1241 184 se
rect 1241 182 1282 184
rect 1241 166 1277 182
tri 1277 166 1282 182 nw
tri 1235 165 1236 166 se
rect 1236 165 1276 166
tri 1276 165 1277 166 nw
rect 1235 164 1276 165
tri 837 157 838 160 sw
rect 837 153 838 157
tri 838 153 839 156 sw
rect 837 150 839 153
tri 341 136 344 150 ne
rect 344 135 376 150
tri 376 135 386 150 sw
tri 513 149 514 150 ne
rect 514 149 549 150
tri 549 149 550 150 sw
tri 617 149 618 150 ne
rect 618 149 669 150
tri 514 139 520 149 ne
rect 520 139 550 149
tri 550 139 552 149 sw
tri 618 139 624 149 ne
rect 624 139 669 149
tri 669 139 675 150 sw
tri 780 139 783 150 se
rect 783 148 839 150
tri 839 148 842 153 sw
rect 783 139 842 148
tri 344 130 345 135 ne
tri 520 131 524 139 ne
rect 524 131 552 139
tri 552 131 556 139 sw
rect 624 137 675 139
tri 624 131 625 137 ne
rect 625 132 675 137
tri 675 132 678 139 sw
tri 778 132 780 139 se
rect 780 132 842 139
tri 842 132 866 148 sw
tri 525 128 526 131 ne
rect 526 128 556 131
tri 556 128 559 131 sw
rect 625 128 627 132
tri 526 119 532 128 ne
rect 532 119 559 128
tri 559 119 566 128 sw
tri 625 119 627 128 ne
tri 532 112 536 119 ne
rect 536 112 566 119
tri 566 112 571 119 sw
tri 536 109 538 112 ne
rect 538 109 571 112
tri 571 109 574 112 sw
tri 538 108 539 109 ne
rect 539 107 574 109
tri 539 103 542 107 ne
rect 542 102 574 107
tri 574 102 579 109 sw
rect 542 101 579 102
tri 579 101 580 102 sw
tri 542 96 546 101 ne
rect 546 95 580 101
tri 580 95 584 101 sw
tri 546 93 547 95 ne
rect 547 93 584 95
tri 547 90 549 93 ne
rect 549 90 584 93
tri 549 89 550 90 ne
rect 550 89 584 90
tri 550 83 555 89 ne
rect 555 83 584 89
tri 584 83 594 95 sw
tri 555 74 564 83 ne
rect 564 80 594 83
tri 594 80 596 83 sw
rect 564 78 596 80
tri 596 78 597 80 sw
rect 564 74 598 78
tri 598 74 601 78 sw
tri 774 115 778 131 se
rect 778 115 819 132
tri 773 113 774 115 se
rect 774 113 819 115
tri 771 109 773 112 se
rect 773 109 819 113
tri 763 102 771 109 se
rect 771 102 819 109
tri 762 101 763 102 se
rect 763 101 819 102
tri 760 100 762 101 se
rect 762 100 819 101
tri 754 96 760 100 se
rect 760 96 819 100
tri 751 93 754 96 se
rect 754 93 819 96
tri 748 91 751 93 se
rect 751 92 819 93
rect 751 91 794 92
tri 794 91 800 92 nw
tri 800 91 801 92 ne
rect 801 91 819 92
tri 747 90 748 91 se
rect 748 90 785 91
tri 741 86 747 90 se
rect 747 86 785 90
tri 785 86 792 91 nw
tri 803 86 812 91 ne
rect 812 86 819 91
tri 738 83 741 86 se
rect 741 83 780 86
tri 734 80 738 83 se
rect 738 82 780 83
tri 780 82 784 86 nw
tri 813 83 819 86 ne
rect 738 80 775 82
tri 732 78 734 80 se
rect 734 78 775 80
tri 775 78 779 82 nw
tri 726 74 732 78 se
rect 732 75 771 78
tri 771 75 775 78 nw
rect 958 156 973 164
tri 973 156 979 164 nw
tri 1234 160 1235 163 se
rect 1235 160 1275 164
tri 1275 160 1276 164 nw
rect 958 155 972 156
tri 972 155 973 156 nw
rect 958 147 966 155
tri 966 147 972 155 nw
tri 958 136 966 147 nw
tri 1120 139 1123 142 se
tri 1114 132 1120 139 se
rect 1120 132 1123 139
rect 1234 159 1274 160
tri 1274 159 1275 160 nw
rect 1542 168 1555 188
tri 1555 168 1566 188 nw
rect 1542 166 1554 168
tri 1554 166 1555 168 nw
rect 1542 164 1553 166
tri 1553 165 1554 166 nw
rect 1542 163 1552 164
tri 1552 163 1553 164 nw
rect 1542 159 1546 163
tri 1546 159 1552 163 nw
tri 1233 156 1234 159 se
rect 1234 156 1259 159
tri 1232 152 1233 155 se
rect 1233 152 1259 156
tri 1226 130 1232 152 se
rect 1232 130 1259 152
tri 1221 115 1226 130 se
rect 1226 115 1259 130
rect 1221 113 1259 115
tri 1259 113 1274 159 nw
tri 1219 108 1221 112 se
rect 1221 108 1250 113
tri 1048 91 1050 95 ne
rect 1050 90 1079 95
tri 1050 85 1052 90 ne
rect 1052 83 1079 90
tri 1052 82 1053 83 ne
rect 1053 82 1079 83
tri 1053 78 1055 82 ne
rect 1055 79 1079 82
tri 1079 79 1082 89 sw
rect 1055 78 1082 79
tri 1055 75 1056 78 ne
rect 1056 75 1082 78
rect 732 74 747 75
tri 564 56 581 74 ne
rect 581 71 601 74
tri 601 71 603 74 sw
tri 722 71 726 74 se
rect 726 71 747 74
rect 581 66 603 71
tri 603 66 607 71 sw
tri 716 66 722 71 se
rect 722 66 747 71
rect 581 59 607 66
tri 607 59 614 66 sw
tri 711 62 716 66 se
rect 716 62 747 66
rect 581 56 614 59
tri 581 35 601 56 ne
rect 601 55 614 56
tri 614 55 622 59 sw
tri 703 56 711 62 se
rect 711 56 747 62
tri 747 56 771 75 nw
tri 1056 56 1063 75 ne
rect 1063 66 1082 75
tri 1082 66 1086 78 sw
tri 1216 96 1219 108 se
rect 1219 96 1250 108
tri 1215 93 1216 95 se
rect 1216 93 1250 96
tri 1214 89 1215 90 se
rect 1215 89 1250 93
tri 1212 84 1214 88 se
rect 1214 86 1250 89
tri 1250 86 1259 113 nw
rect 1214 84 1249 86
tri 1249 84 1250 86 nw
tri 1209 82 1212 84 se
rect 1212 82 1246 84
tri 1204 78 1209 82 se
rect 1209 78 1246 82
tri 1191 68 1204 78 se
rect 1204 76 1246 78
tri 1246 76 1249 84 nw
rect 1204 69 1241 76
tri 1241 69 1246 76 nw
rect 1204 68 1239 69
tri 1239 68 1241 69 nw
tri 1189 66 1191 68 se
rect 1191 66 1222 68
rect 1063 56 1086 66
tri 1086 56 1098 66 sw
tri 1178 57 1189 66 se
rect 1189 57 1222 66
tri 1222 57 1239 68 nw
tri 702 55 703 56 se
rect 703 55 741 56
rect 601 50 622 55
tri 622 50 636 55 sw
tri 697 51 702 55 se
rect 702 51 741 55
tri 741 51 747 56 nw
tri 1063 51 1067 56 ne
rect 1067 53 1098 56
tri 1098 53 1101 56 sw
tri 1172 55 1178 57 se
rect 1178 55 1213 57
tri 1161 53 1172 55 se
rect 1172 53 1213 55
rect 1067 52 1101 53
tri 1101 52 1121 53 sw
tri 1155 52 1161 53 se
rect 1161 52 1213 53
rect 1067 51 1121 52
tri 1121 51 1153 52 sw
tri 1153 51 1155 52 se
rect 1155 51 1213 52
tri 1213 51 1222 57 nw
tri 676 50 697 51 se
rect 697 50 740 51
tri 740 50 741 51 nw
tri 1067 50 1068 51 ne
rect 1068 50 1194 51
rect 601 35 721 50
tri 721 35 740 50 nw
tri 1068 35 1084 50 ne
rect 1084 39 1194 50
tri 1194 39 1212 51 nw
rect 1084 35 1173 39
tri 601 29 608 35 ne
rect 608 30 715 35
tri 715 30 721 35 nw
tri 1084 30 1090 35 ne
rect 608 29 714 30
tri 714 29 715 30 nw
rect 1090 29 1173 35
tri 608 27 617 29 ne
rect 617 26 711 29
tri 711 27 714 29 nw
tri 1090 27 1093 29 ne
rect 1093 27 1173 29
tri 1173 27 1194 39 nw
tri 1093 26 1097 27 ne
rect 1097 26 1169 27
tri 617 25 622 26 ne
rect 622 25 709 26
tri 709 25 711 26 nw
tri 1097 25 1144 26 ne
rect 1144 25 1164 26
tri 1164 25 1169 26 nw
tri 622 22 630 25 ne
rect 630 22 702 25
tri 702 22 708 25 nw
<< via2 >>
rect 891 292 947 313
rect 1275 352 1331 356
rect 1275 300 1286 352
rect 1286 300 1331 352
rect 243 224 249 244
rect 249 224 299 244
rect 243 188 299 224
rect 891 257 936 292
rect 936 257 947 292
rect 387 218 443 244
rect 387 188 405 218
rect 405 188 443 218
rect 1515 211 1571 244
rect 1515 188 1542 211
rect 1542 188 1571 211
rect 627 76 683 132
rect 819 76 875 132
rect 1107 108 1123 132
rect 1123 108 1163 132
rect 1107 76 1163 108
<< metal3 >>
rect 886 313 952 398
rect 886 257 891 313
rect 947 257 952 313
rect 1270 356 1336 422
rect 1270 300 1275 356
rect 1331 300 1336 356
rect 1270 276 1336 300
rect 886 252 952 257
rect 238 244 304 249
rect 238 188 243 244
rect 299 188 304 244
rect 238 103 304 188
rect 382 244 448 249
rect 382 188 387 244
rect 443 188 448 244
rect 1510 244 1576 249
rect 382 103 448 188
rect 622 132 688 217
rect 1510 188 1515 244
rect 1571 188 1576 244
rect 622 76 627 132
rect 683 76 688 132
rect 622 71 688 76
rect 814 132 960 137
rect 814 76 819 132
rect 875 76 960 132
rect 814 71 960 76
rect 1102 132 1248 137
rect 1102 76 1107 132
rect 1163 76 1248 132
rect 1510 103 1576 188
rect 1102 71 1248 76
<< labels >>
flabel nwell s 77 527 111 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel pwell s 77 -17 111 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel comment s 0 0 0 0 0 FreeSans 100 0 0 0 scs130hd_mpr2ya_8
flabel metal3 s 238 103 304 249 0 FreeSans 100 0 0 0 A0
port 3 nsew
flabel metal3 s 382 103 448 249 0 FreeSans 100 0 0 0 B0
port 4 nsew
flabel metal3 s 814 71 960 137 0 FreeSans 100 0 0 0 B1
port 5 nsew
flabel metal3 s 1270 276 1336 422 0 FreeSans 100 0 0 0 R3
port 6 nsew
flabel metal3 s 622 71 688 216 0 FreeSans 100 0 0 0 R2
port 7 nsew
flabel metal3 s 1510 103 1576 249 0 FreeSans 100 0 0 0 R1
port 8 nsew
flabel metal3 s 1102 71 1248 137 0 FreeSans 100 0 0 0 R0
port 9 nsew
flabel metal3 s 886 252 952 398 0 FreeSans 100 0 0 0 A1
port 10 nsew
flabel metal1 s 31 -17 65 17 0 FreeSans 100 0 0 0 vgnd
port 11 nsew
flabel metal1 s 31 527 65 561 0 FreeSans 100 0 0 0 vpwr
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 1748 544
<< end >>
