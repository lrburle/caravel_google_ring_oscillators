magic
tech sky130A
magscale 1 2
timestamp 1716047795
<< nwell >>
rect 0 1674 1180 1748
rect 1342 1674 3267 1748
rect 0 1086 3267 1674
rect 0 921 112 1086
rect 0 819 177 921
rect 2077 804 2291 1086
rect 2078 744 2291 804
rect 3073 772 3103 807
rect 3222 744 3267 1086
<< ndiff >>
rect 3159 442 3193 476
<< locali >>
rect 2 2172 3268 2492
rect 2842 1869 2920 1885
rect 2796 1851 2920 1869
rect 2983 1721 3102 1755
rect 2994 1689 2995 1721
rect 3160 1460 3194 1494
rect 1 1086 3267 1406
rect 3159 998 3193 1032
rect 2960 725 3094 759
rect 2796 623 2924 641
rect 175 567 250 578
rect 175 550 214 567
rect 627 550 705 578
rect 1060 572 1099 578
rect 1002 550 1041 572
rect 1370 550 1409 578
rect 2842 607 2924 623
rect 1740 550 1780 573
rect 2075 572 2113 576
rect 2074 550 2113 572
rect 150 320 2113 550
rect 1 0 3267 320
<< viali >>
rect 2796 1869 2842 1915
rect 3159 1742 3193 1776
rect 2796 577 2842 623
rect 3159 442 3193 476
<< metal1 >>
rect 2 2172 3268 2492
rect 1317 1757 1352 2172
rect 1463 1933 1537 1942
rect 1463 1877 1472 1933
rect 1528 1877 1537 1933
rect 2784 1915 2854 1921
rect 2636 1908 2796 1915
rect 2648 1902 2796 1908
rect 1463 1872 1537 1877
rect 2602 1881 2796 1902
rect 1463 1868 1514 1872
rect 2602 1868 2648 1881
rect 2784 1869 2796 1881
rect 2842 1869 2854 1915
rect 2784 1863 2854 1869
rect 2681 1846 2746 1853
rect 2681 1828 2688 1846
rect 1565 1794 2688 1828
rect 2740 1794 2746 1846
rect 2681 1788 2746 1794
rect 1317 1755 1367 1757
rect 1317 1754 1381 1755
rect 1317 1741 1392 1754
rect 1317 1720 1409 1741
rect 2521 1708 2527 1766
rect 2579 1708 2585 1766
rect 1189 1680 1253 1693
rect 2311 1689 2379 1695
rect 2311 1680 2317 1689
rect 1189 1675 1257 1680
rect 2308 1675 2317 1680
rect 1189 1641 2317 1675
rect 1189 1635 1253 1641
rect 2311 1631 2317 1641
rect 2375 1631 2379 1689
rect 2311 1625 2379 1631
rect 1 1086 3267 1406
rect 1920 861 1984 870
rect 1936 848 1984 861
rect 2313 868 2381 874
rect 1936 811 2113 848
rect 1936 806 1984 811
rect 175 550 214 578
rect 627 550 705 578
rect 1060 572 1099 578
rect 1002 550 1041 572
rect 1370 550 1409 578
rect 2076 576 2113 811
rect 2313 810 2319 868
rect 2377 810 2381 868
rect 2313 803 2381 810
rect 2521 783 2585 789
rect 2521 775 2527 783
rect 2523 773 2527 775
rect 2521 772 2527 773
rect 2516 769 2527 772
rect 2515 738 2527 769
rect 2521 732 2527 738
rect 2579 731 2585 783
rect 2574 729 2585 731
rect 2676 716 2746 722
rect 2676 698 2682 716
rect 2215 664 2682 698
rect 2215 621 2249 664
rect 2676 658 2682 664
rect 2740 658 2746 716
rect 2676 652 2746 658
rect 2784 624 2854 629
rect 2602 623 2636 624
rect 2648 623 2854 624
rect 2075 572 2113 576
rect 2074 550 2113 572
rect 2197 615 2265 621
rect 2197 557 2203 615
rect 2261 557 2265 615
rect 2602 590 2796 623
rect 2784 577 2796 590
rect 2842 577 2854 623
rect 2784 571 2854 577
rect 2197 551 2265 557
rect 150 320 2113 550
rect 1 0 3267 320
<< via1 >>
rect 1472 1877 1528 1933
rect 2688 1794 2740 1846
rect 2527 1708 2579 1766
rect 2317 1631 2375 1689
rect 2319 810 2377 868
rect 2527 731 2579 783
rect 2682 658 2740 716
rect 2203 557 2261 615
<< metal2 >>
rect 1463 1933 1537 1942
rect 1463 1877 1472 1933
rect 1528 1877 1537 1933
rect 1463 1868 1537 1877
rect 2681 1846 2746 1853
rect 2681 1840 2688 1846
rect 2458 1806 2688 1840
rect 2311 1689 2379 1695
rect 2311 1631 2317 1689
rect 2375 1631 2379 1689
rect 2311 1625 2379 1631
rect 2328 874 2362 1625
rect 2313 868 2381 874
rect 2313 810 2319 868
rect 2377 810 2381 868
rect 2313 804 2381 810
rect 2458 765 2490 1806
rect 2681 1794 2688 1806
rect 2740 1794 2746 1846
rect 2681 1788 2746 1794
rect 2521 1708 2527 1766
rect 2579 1708 2585 1766
rect 2521 1701 2585 1708
rect 2527 1666 2561 1701
rect 2527 1631 2562 1666
rect 2527 1596 2722 1631
rect 2521 783 2585 789
rect 2521 765 2527 783
rect 2458 731 2527 765
rect 2579 731 2585 783
rect 2521 725 2585 731
rect 2687 722 2722 1596
rect 2676 716 2746 722
rect 2676 658 2682 716
rect 2740 658 2746 716
rect 500 547 534 657
rect 2676 652 2746 658
rect 2215 621 2249 622
rect 2197 615 2265 621
rect 2197 557 2203 615
rect 2261 557 2265 615
rect 2197 551 2265 557
rect 2197 547 2249 551
rect 500 513 2249 547
<< via2 >>
rect 1472 1877 1528 1933
<< metal3 >>
rect 1463 1935 1537 1942
rect 1463 1933 1860 1935
rect 1463 1877 1472 1933
rect 1528 1877 1860 1933
rect 1463 1875 1860 1877
rect 1463 1868 1537 1875
rect 1800 775 1860 1875
rect 1032 715 1452 775
rect 1392 713 1452 715
rect 1640 715 1860 775
rect 1640 713 1701 715
rect 1392 655 1701 713
rect 1392 652 1664 655
use scs130hd_mpr2ea_8  scs130hd_mpr2ea_8_0
timestamp 1714057206
transform 1 0 150 0 1 559
box -38 -48 1970 592
use sky130_osu_sc_12T_hs__fill_2  sky130_osu_sc_12T_hs__fill_2_0
timestamp 1714057206
transform 1 0 1728 0 -1 2233
box -7 0 161 897
use sky130_osu_sc_12T_hs__fill_8  sky130_osu_sc_12T_hs__fill_8_0
timestamp 1714057206
transform 1 0 1899 0 -1 2233
box -9 0 179 897
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1714057206
transform 1 0 2840 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1714057206
transform 1 0 3038 0 1 260
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1714057206
transform 1 0 3039 0 -1 2232
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1714057206
transform 1 0 2840 0 -1 2233
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1714057206
transform 1 0 2291 0 1 259
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1714057206
transform 1 0 1168 0 -1 2233
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1714057206
transform 1 0 2291 0 -1 2233
box -10 0 552 902
<< labels >>
rlabel metal1 76 1151 76 1151 1 vccd1
port 6 n
rlabel metal1 53 293 53 293 1 vssd1
port 5 n
rlabel metal1 1565 1794 1594 1828 1 in
port 8 n
rlabel metal1 53 2200 53 2200 1 vssd1
port 5 n
rlabel viali 3159 442 3193 476 1 Y1
port 10 n
rlabel viali 3159 1742 3193 1776 1 Y0
port 9 n
rlabel metal2 2347 841 2347 841 1 sel
port 7 n
<< end >>
