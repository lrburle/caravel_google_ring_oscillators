magic
tech sky130A
magscale 1 2
timestamp 1714057206
<< error_s >>
rect -1864 1495 -1848 1524
rect -1836 1495 -1820 1496
rect -1829 1460 -1819 1461
rect -1801 1456 -1791 1461
rect -1966 1372 -1941 1386
rect -1938 1381 -1913 1386
<< nwell >>
rect -2159 1147 -1480 1489
rect 148 1386 306 1489
rect 1014 1427 1015 1465
rect 348 1386 380 1422
rect 148 1367 311 1386
rect -1476 1147 -1431 1170
rect 109 1147 311 1367
rect 1242 1147 1287 1489
rect -2159 1146 -1431 1147
rect -2159 1139 -1480 1146
rect -1476 1139 -1431 1146
rect -2159 873 -1397 1139
rect -2159 826 -1365 873
rect 70 869 1287 1147
rect 72 838 1287 869
rect 89 827 1287 838
rect -2159 824 -1423 826
rect -2159 603 -1325 824
rect 89 796 311 827
rect -273 763 311 796
rect 89 603 311 763
rect -2159 483 -1440 603
rect 148 485 311 603
rect 1093 513 1123 548
rect 1242 485 1287 827
<< ndiff >>
rect 1177 182 1212 216
<< psubdiff >>
rect 318 1947 342 1954
rect 318 1917 348 1947
rect 318 1914 349 1917
rect 474 1915 549 1947
rect 473 1914 555 1915
<< locali >>
rect -2158 1928 1287 2233
rect -2158 1927 -659 1928
rect -2158 1913 -1343 1927
rect -1400 1446 -1343 1913
rect -1286 1446 -1229 1927
rect -1172 1446 -1115 1927
rect -1058 1446 -1001 1927
rect -944 1446 -887 1927
rect -830 1446 -773 1927
rect -716 1446 -659 1927
rect -602 1446 -545 1928
rect -488 1446 -432 1928
rect -375 1446 -318 1928
rect -261 1446 -204 1928
rect -147 1446 -90 1928
rect 24 1913 1287 1928
rect 24 1446 72 1913
rect 1012 1462 1119 1497
rect -905 1206 -871 1421
rect 346 1386 382 1434
rect 1014 1427 1015 1462
rect 1179 1202 1213 1236
rect -2158 1141 -1423 1147
rect -2158 873 -1397 1141
rect -2158 826 -1365 873
rect 70 869 1287 1147
rect 89 827 1287 869
rect 1178 738 1212 772
rect 1013 466 1117 502
rect -1401 327 -1392 359
rect 70 331 131 359
rect -1226 329 131 331
rect -1401 62 -1345 327
rect -1288 62 -1231 327
rect -1174 62 -1117 329
rect -1060 62 -1003 329
rect -946 62 -889 329
rect -832 62 -775 329
rect -718 62 -661 329
rect -604 62 -547 329
rect -490 62 -433 329
rect -376 62 -319 329
rect -262 62 -205 329
rect -148 62 -91 329
rect -34 62 23 329
rect 46 325 131 329
rect 80 62 131 325
rect -1401 61 131 62
rect -2158 -259 1287 61
<< viali >>
rect 894 1617 940 1663
rect 1178 1484 1212 1518
rect 897 330 943 376
rect 1178 182 1212 216
<< metal1 >>
rect -2158 1928 1287 2233
rect -2158 1927 -659 1928
rect -2158 1913 -1343 1927
rect -1882 1495 -1848 1913
rect -1734 1668 -1660 1677
rect -1734 1612 -1725 1668
rect -1669 1612 -1660 1668
rect -1734 1603 -1660 1612
rect -1645 1513 -1639 1569
rect -1583 1513 -1577 1569
rect -1882 1494 -1801 1495
rect -1882 1463 -1802 1494
rect -1882 1461 -1800 1463
rect -1882 1460 -1819 1461
rect -1400 1446 -1343 1913
rect -1286 1446 -1229 1927
rect -1172 1446 -1115 1927
rect -1058 1446 -1001 1927
rect -944 1446 -887 1927
rect -830 1446 -773 1927
rect -716 1446 -659 1927
rect -602 1446 -545 1928
rect -488 1446 -432 1928
rect -375 1446 -318 1928
rect -261 1446 -204 1928
rect -147 1446 -90 1928
rect 24 1913 1287 1928
rect 24 1446 72 1913
rect 894 1671 940 1675
rect 888 1663 946 1671
rect 888 1656 894 1663
rect 656 1649 894 1656
rect 668 1643 894 1649
rect 622 1622 894 1643
rect 622 1609 668 1622
rect 888 1617 894 1622
rect 940 1617 946 1663
rect 888 1609 946 1617
rect 894 1604 940 1609
rect 701 1587 766 1594
rect 701 1535 708 1587
rect 760 1535 766 1587
rect 701 1529 766 1535
rect 541 1513 605 1519
rect 541 1461 547 1513
rect 599 1461 605 1513
rect 541 1454 605 1461
rect -2009 1434 -1941 1440
rect -2009 1378 -2003 1434
rect -1947 1421 -1941 1434
rect -1947 1414 -1938 1421
rect -1545 1414 -1539 1432
rect -1947 1387 -1539 1414
rect -1947 1378 -1941 1387
rect -1938 1381 -1539 1387
rect -2009 1372 -1941 1378
rect -1545 1376 -1539 1381
rect -1483 1376 -1477 1432
rect 332 1427 397 1434
rect 332 1375 339 1427
rect 391 1375 397 1427
rect 332 1369 397 1375
rect -2158 1146 -1423 1147
rect -2158 1128 -1646 1146
rect -1585 1141 -1423 1146
rect -1585 1128 -1397 1141
rect -2158 873 -1397 1128
rect -2158 826 -1365 873
rect 70 869 1287 1147
rect 72 838 1287 869
rect 89 827 1287 838
rect 332 757 397 764
rect 332 705 339 757
rect 391 705 397 757
rect 332 699 397 705
rect 348 586 382 699
rect 541 531 605 537
rect 541 513 547 531
rect 478 479 547 513
rect 599 479 605 531
rect 541 473 605 479
rect 207 457 272 464
rect 207 405 214 457
rect 266 405 272 457
rect 207 399 272 405
rect 696 457 766 463
rect 696 399 702 457
rect 760 399 766 457
rect 696 393 766 399
rect 896 386 943 388
rect 884 376 952 386
rect 884 365 897 376
rect -1401 327 -1391 365
rect 72 359 131 365
rect 70 331 131 359
rect 622 364 656 365
rect 668 364 897 365
rect 622 331 897 364
rect -1226 329 131 331
rect -1401 62 -1345 327
rect -1288 62 -1231 327
rect -1174 62 -1117 329
rect -1060 62 -1003 329
rect -946 62 -889 329
rect -832 62 -775 329
rect -718 62 -661 329
rect -604 62 -547 329
rect -490 62 -433 329
rect -376 62 -319 329
rect -262 62 -205 329
rect -148 62 -91 329
rect -34 62 23 329
rect 46 325 131 329
rect 71 294 131 325
rect 884 330 897 331
rect 943 330 952 376
rect 884 323 952 330
rect 896 318 943 323
rect 80 62 131 294
rect -1401 61 131 62
rect -2158 -259 1287 61
<< via1 >>
rect -1725 1612 -1669 1668
rect -1639 1513 -1583 1569
rect 708 1535 760 1587
rect 547 1461 599 1513
rect -2003 1378 -1947 1434
rect -1539 1376 -1483 1432
rect 339 1375 391 1427
rect 339 705 391 757
rect 547 479 599 531
rect 214 405 266 457
rect 702 399 760 457
<< metal2 >>
rect -1734 1668 -1660 1677
rect -1734 1612 -1725 1668
rect -1669 1612 -1660 1668
rect -1734 1603 -1660 1612
rect -1629 1671 510 1705
rect -1629 1575 -1595 1671
rect -1528 1605 382 1639
rect -1639 1569 -1583 1575
rect -1639 1507 -1583 1513
rect -2013 1434 -1938 1443
rect -1528 1438 -1494 1605
rect -2013 1378 -2003 1434
rect -1947 1378 -1938 1434
rect -2013 1369 -1938 1378
rect -1539 1432 -1483 1438
rect 348 1434 382 1605
rect 478 1581 510 1671
rect 701 1587 766 1594
rect 701 1581 708 1587
rect 478 1547 708 1581
rect -1539 1370 -1483 1376
rect 332 1427 397 1434
rect 332 1375 339 1427
rect 391 1375 397 1427
rect 332 1369 397 1375
rect 346 764 380 1369
rect 332 757 397 764
rect 332 705 339 757
rect 391 705 397 757
rect 332 699 397 705
rect -496 504 -461 636
rect 478 513 510 1547
rect 701 1535 708 1547
rect 760 1535 766 1587
rect 701 1529 766 1535
rect 541 1513 605 1519
rect 541 1461 547 1513
rect 599 1461 605 1513
rect 541 1454 605 1461
rect 547 1407 581 1454
rect 547 1372 582 1407
rect 547 1337 742 1372
rect 541 531 605 537
rect 541 513 547 531
rect -496 469 148 504
rect 478 479 547 513
rect 599 479 605 531
rect 541 473 605 479
rect 113 439 148 469
rect 207 457 272 464
rect 707 463 742 1337
rect 207 439 214 457
rect 113 405 214 439
rect 266 439 272 457
rect 696 457 766 463
rect 696 439 702 457
rect 266 405 702 439
rect 207 399 272 405
rect 696 399 702 405
rect 760 399 766 457
rect 696 393 766 399
<< via2 >>
rect -1725 1612 -1669 1668
rect -2003 1378 -1947 1434
<< metal3 >>
rect -2008 1443 -1942 2230
rect -1734 1668 -1660 1677
rect -1734 1612 -1725 1668
rect -1669 1665 -1660 1668
rect -1669 1612 -304 1665
rect -1734 1605 -304 1612
rect -1734 1603 -1660 1605
rect -2013 1434 -1938 1443
rect -2013 1378 -2003 1434
rect -1947 1378 -1938 1434
rect -2013 1369 -1938 1378
rect -781 1298 -721 1605
rect -575 1227 -515 1605
rect -364 1234 -304 1605
rect -583 1157 -515 1227
rect -379 1161 -304 1234
use scs130hd_mpr2ct_8  scs130hd_mpr2ct_8_1
timestamp 1710282110
transform 1 0 -1400 0 1 342
box -43 -60 1510 1148
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_0
timestamp 1714057206
transform 1 0 1057 0 1 0
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1714057206
transform 1 0 860 0 1 0
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1714057206
transform 1 0 1058 0 -1 1974
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1714057206
transform 1 0 860 0 -1 1974
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1714057206
transform 1 0 311 0 1 0
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1714057206
transform 1 0 -2026 0 -1 1972
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1714057206
transform 1 0 311 0 -1 1974
box -10 0 552 902
<< labels >>
rlabel metal2 364 733 364 733 1 sel
port 8 n
rlabel metal1 -2106 26 -2106 26 1 vssd1
port 5 n
rlabel metal1 -2097 1088 -2097 1088 1 vccd1
port 6 n
rlabel via1 -1612 1537 -1612 1537 1 in
port 11 n
rlabel metal1 -2100 1944 -2100 1944 1 vssd1
port 5 n
rlabel viali 1178 182 1212 216 1 Y1
port 10 n
rlabel viali 1178 1484 1212 1518 1 Y0
port 9 n
<< end >>
