VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -15.990 -10.630 -8.930 3530.310 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.030 -6.670 2935.610 -3.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.030 3523.250 2935.610 3526.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2928.550 -10.630 2935.610 3530.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.720 -11.470 7.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.720 -11.470 42.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.720 -11.470 77.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.720 -11.470 112.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 145.720 -11.470 147.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.720 -11.470 182.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 215.720 -11.470 217.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.720 -11.470 252.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 285.720 -11.470 287.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.720 -11.470 322.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 355.720 -11.470 357.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 390.720 -11.470 392.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.720 -11.470 427.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 460.720 -11.470 462.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.720 -11.470 497.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 530.720 -11.470 532.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 565.720 -11.470 567.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 600.720 -11.470 602.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.720 -11.470 637.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 670.720 -11.470 672.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 705.720 -11.470 707.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 740.720 -11.470 742.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.720 -11.470 777.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 810.720 -11.470 812.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 845.720 -11.470 847.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 880.720 -11.470 882.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 915.720 -11.470 917.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 950.720 -11.470 952.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 985.720 -11.470 987.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1020.720 -11.470 1022.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.720 -11.470 1057.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1090.720 -11.470 1092.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.720 -11.470 1127.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1160.720 -11.470 1162.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1195.720 -11.470 1197.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1230.720 -11.470 1232.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1265.720 -11.470 1267.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1300.720 -11.470 1302.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1335.720 -11.470 1337.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1370.720 -11.470 1372.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1405.720 -11.470 1407.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1440.720 -11.470 1442.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 -11.470 1477.320 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 1003.200 1477.320 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 1843.200 1477.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1510.720 -11.470 1512.320 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1510.720 1003.200 1512.320 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1510.720 1843.200 1512.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1545.720 -11.470 1547.320 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1545.720 1003.200 1547.320 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1545.720 1843.200 1547.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1580.720 -11.470 1582.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1615.720 -11.470 1617.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1650.720 -11.470 1652.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1685.720 -11.470 1687.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1720.720 -11.470 1722.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1755.720 -11.470 1757.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1790.720 -11.470 1792.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.720 -11.470 1827.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1860.720 -11.470 1862.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1895.720 -11.470 1897.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1930.720 -11.470 1932.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1965.720 -11.470 1967.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.720 -11.470 2002.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2035.720 -11.470 2037.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2070.720 -11.470 2072.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2105.720 -11.470 2107.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2140.720 -11.470 2142.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.720 -11.470 2177.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2210.720 -11.470 2212.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2245.720 -11.470 2247.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2280.720 -11.470 2282.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2315.720 -11.470 2317.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2350.720 -11.470 2352.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2385.720 -11.470 2387.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2420.720 -11.470 2422.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2455.720 -11.470 2457.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2490.720 -11.470 2492.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2525.720 -11.470 2527.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2560.720 -11.470 2562.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2595.720 -11.470 2597.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.720 -11.470 2632.320 1200.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.720 1308.760 2632.320 1400.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.720 1508.760 2632.320 1600.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.720 1708.760 2632.320 1800.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.720 1908.760 2632.320 2000.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.720 2108.760 2632.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2665.720 -11.470 2667.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 -11.470 2702.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2735.720 -11.470 2737.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2770.720 -11.470 2772.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2805.720 -11.470 2807.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2840.720 -11.470 2842.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2875.720 -11.470 2877.320 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2910.720 -11.470 2912.320 3531.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 11.080 2944.370 12.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 46.080 2944.370 47.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 81.080 2944.370 82.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 116.080 2944.370 117.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 151.080 2944.370 152.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 186.080 2944.370 187.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 221.080 2944.370 222.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 256.080 2944.370 257.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 291.080 2944.370 292.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 326.080 2944.370 327.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 361.080 2944.370 362.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 396.080 2944.370 397.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 431.080 2944.370 432.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 466.080 2944.370 467.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 501.080 2944.370 502.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 536.080 2944.370 537.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 571.080 2944.370 572.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 606.080 2944.370 607.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 641.080 2944.370 642.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 676.080 2944.370 677.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 711.080 2944.370 712.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 746.080 2944.370 747.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 781.080 2944.370 782.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 816.080 2944.370 817.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 851.080 2944.370 852.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 886.080 2944.370 887.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 921.080 2944.370 922.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 956.080 2944.370 957.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 991.080 2944.370 992.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1026.080 2944.370 1027.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1061.080 2944.370 1062.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1096.080 2944.370 1097.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1131.080 2944.370 1132.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1166.080 2944.370 1167.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1201.080 2944.370 1202.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1236.080 2944.370 1237.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1271.080 2944.370 1272.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1306.080 2944.370 1307.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1341.080 2944.370 1342.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1376.080 2944.370 1377.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1411.080 2944.370 1412.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1446.080 2944.370 1447.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1481.080 2944.370 1482.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1516.080 2944.370 1517.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1551.080 2944.370 1552.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1586.080 2944.370 1587.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1621.080 2944.370 1622.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1656.080 2944.370 1657.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1691.080 2944.370 1692.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1726.080 2944.370 1727.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1761.080 2944.370 1762.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1796.080 2944.370 1797.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1831.080 2944.370 1832.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1866.080 2944.370 1867.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1901.080 2944.370 1902.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1936.080 2944.370 1937.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1971.080 2944.370 1972.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2006.080 2944.370 2007.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2041.080 2944.370 2042.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2076.080 2944.370 2077.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2111.080 2944.370 2112.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2146.080 2944.370 2147.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2181.080 2944.370 2182.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2216.080 2944.370 2217.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2251.080 2944.370 2252.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2286.080 2944.370 2287.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2321.080 2944.370 2322.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2356.080 2944.370 2357.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2391.080 2944.370 2392.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2426.080 2944.370 2427.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2461.080 2944.370 2462.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2496.080 2944.370 2497.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2531.080 2944.370 2532.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2566.080 2944.370 2567.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2601.080 2944.370 2602.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2636.080 2944.370 2637.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2671.080 2944.370 2672.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2706.080 2944.370 2707.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2741.080 2944.370 2742.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2776.080 2944.370 2777.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2811.080 2944.370 2812.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2846.080 2944.370 2847.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2881.080 2944.370 2882.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2916.080 2944.370 2917.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2951.080 2944.370 2952.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2986.080 2944.370 2987.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3021.080 2944.370 3022.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3056.080 2944.370 3057.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3091.080 2944.370 3092.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3126.080 2944.370 3127.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3161.080 2944.370 3162.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3196.080 2944.370 3197.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3231.080 2944.370 3232.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3266.080 2944.370 3267.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3301.080 2944.370 3302.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3336.080 2944.370 3337.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3371.080 2944.370 3372.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3406.080 2944.370 3407.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3441.080 2944.370 3442.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3476.080 2944.370 3477.680 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.750 -19.390 -17.690 3539.070 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.830 -11.470 2936.450 -8.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.830 3528.050 2936.450 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2937.310 -19.390 2944.370 3539.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.380 -11.470 15.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.380 -11.470 50.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.380 -11.470 85.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.380 -11.470 120.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.380 -11.470 155.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.380 -11.470 190.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.380 -11.470 225.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 259.380 -11.470 260.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.380 -11.470 295.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.380 -11.470 330.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.380 -11.470 365.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 399.380 -11.470 400.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 434.380 -11.470 435.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.380 -11.470 470.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.380 -11.470 505.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 539.380 -11.470 540.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.380 -11.470 575.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 609.380 -11.470 610.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 644.380 -11.470 645.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.380 -11.470 680.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.380 -11.470 715.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 749.380 -11.470 750.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.380 -11.470 785.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.380 -11.470 820.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.380 -11.470 855.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 889.380 -11.470 890.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 924.380 -11.470 925.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.380 -11.470 960.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 994.380 -11.470 995.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1029.380 -11.470 1030.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1064.380 -11.470 1065.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.380 -11.470 1100.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1134.380 -11.470 1135.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1169.380 -11.470 1170.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1204.380 -11.470 1205.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1239.380 -11.470 1240.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1274.380 -11.470 1275.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1309.380 -11.470 1310.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1344.380 -11.470 1345.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1379.380 -11.470 1380.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.380 -11.470 1415.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1449.380 -11.470 1450.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1484.380 -11.470 1485.980 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1484.380 1003.200 1485.980 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1484.380 1843.200 1485.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1519.380 -11.470 1520.980 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1519.380 1003.200 1520.980 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1519.380 1843.200 1520.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1554.380 -11.470 1555.980 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1554.380 1002.735 1555.980 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1554.380 1842.735 1555.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1589.380 -11.470 1590.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1624.380 -11.470 1625.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1659.380 -11.470 1660.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1694.380 -11.470 1695.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1729.380 -11.470 1730.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1764.380 -11.470 1765.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1799.380 -11.470 1800.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1834.380 -11.470 1835.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1869.380 -11.470 1870.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.380 -11.470 1905.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1939.380 -11.470 1940.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1974.380 -11.470 1975.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.380 -11.470 2010.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.380 -11.470 2045.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2079.380 -11.470 2080.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.380 -11.470 2115.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2149.380 -11.470 2150.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.380 -11.470 2185.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2219.380 -11.470 2220.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.380 -11.470 2255.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.380 -11.470 2290.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2324.380 -11.470 2325.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2359.380 -11.470 2360.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.380 -11.470 2395.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2429.380 -11.470 2430.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.380 -11.470 2465.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2499.380 -11.470 2500.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2534.380 -11.470 2535.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2569.380 -11.470 2570.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.380 -11.470 2605.980 1200.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.380 1308.760 2605.980 1400.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.380 1508.760 2605.980 1600.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.380 1708.760 2605.980 1800.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.380 1908.760 2605.980 2000.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.380 2108.760 2605.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2639.380 -11.470 2640.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.380 -11.470 2675.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.380 -11.470 2710.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2744.380 -11.470 2745.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2779.380 -11.470 2780.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2814.380 -11.470 2815.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2849.380 -11.470 2850.980 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2884.380 -11.470 2885.980 3531.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 16.415 2944.370 18.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 51.415 2944.370 53.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 86.415 2944.370 88.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 121.415 2944.370 123.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 156.415 2944.370 158.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 191.415 2944.370 193.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 226.415 2944.370 228.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 261.415 2944.370 263.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 296.415 2944.370 298.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 331.415 2944.370 333.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 366.415 2944.370 368.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 401.415 2944.370 403.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 436.415 2944.370 438.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 471.415 2944.370 473.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 506.415 2944.370 508.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 541.415 2944.370 543.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 576.415 2944.370 578.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 611.415 2944.370 613.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 646.415 2944.370 648.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 681.415 2944.370 683.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 716.415 2944.370 718.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 751.415 2944.370 753.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 786.415 2944.370 788.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 821.415 2944.370 823.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 856.415 2944.370 858.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 891.415 2944.370 893.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 926.415 2944.370 928.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 961.415 2944.370 963.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 996.415 2944.370 998.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1031.415 2944.370 1033.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1066.415 2944.370 1068.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1101.415 2944.370 1103.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1136.415 2944.370 1138.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1171.415 2944.370 1173.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1206.415 2944.370 1208.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1241.415 2944.370 1243.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1276.415 2944.370 1278.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1311.415 2944.370 1313.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1346.415 2944.370 1348.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1381.415 2944.370 1383.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1416.415 2944.370 1418.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1451.415 2944.370 1453.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1486.415 2944.370 1488.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1521.415 2944.370 1523.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1556.415 2944.370 1558.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1591.415 2944.370 1593.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1626.415 2944.370 1628.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1661.415 2944.370 1663.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1696.415 2944.370 1698.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1731.415 2944.370 1733.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1766.415 2944.370 1768.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1801.415 2944.370 1803.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1836.415 2944.370 1838.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1871.415 2944.370 1873.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1906.415 2944.370 1908.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1941.415 2944.370 1943.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 1976.415 2944.370 1978.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2011.415 2944.370 2013.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2046.415 2944.370 2048.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2081.415 2944.370 2083.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2116.415 2944.370 2118.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2151.415 2944.370 2153.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2186.415 2944.370 2188.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2221.415 2944.370 2223.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2256.415 2944.370 2258.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2291.415 2944.370 2293.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2326.415 2944.370 2328.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2361.415 2944.370 2363.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2396.415 2944.370 2398.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2431.415 2944.370 2433.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2466.415 2944.370 2468.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2501.415 2944.370 2503.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2536.415 2944.370 2538.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2571.415 2944.370 2573.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2606.415 2944.370 2608.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2641.415 2944.370 2643.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2676.415 2944.370 2678.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2711.415 2944.370 2713.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2746.415 2944.370 2748.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2781.415 2944.370 2783.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2816.415 2944.370 2818.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2851.415 2944.370 2853.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2886.415 2944.370 2888.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2921.415 2944.370 2923.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2956.415 2944.370 2958.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 2991.415 2944.370 2993.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3026.415 2944.370 3028.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3061.415 2944.370 3063.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3096.415 2944.370 3098.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3131.415 2944.370 3133.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3166.415 2944.370 3168.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3201.415 2944.370 3203.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3236.415 2944.370 3238.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3271.415 2944.370 3273.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3306.415 2944.370 3308.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3341.415 2944.370 3343.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3376.415 2944.370 3378.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3411.415 2944.370 3413.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3446.415 2944.370 3448.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.750 3481.415 2944.370 3483.015 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 1475.720 884.000 2634.160 2458.310 ;
      LAYER met1 ;
        RECT 1462.410 884.000 2901.150 2458.310 ;
      LAYER met2 ;
        RECT 1462.440 32.795 2902.050 2464.165 ;
      LAYER met3 ;
        RECT 1469.305 2424.180 2917.600 2464.145 ;
        RECT 1469.305 2422.180 2917.200 2424.180 ;
        RECT 1469.305 2358.220 2917.600 2422.180 ;
        RECT 1469.305 2356.220 2917.200 2358.220 ;
        RECT 1469.305 2291.580 2917.600 2356.220 ;
        RECT 1469.305 2289.580 2917.200 2291.580 ;
        RECT 1469.305 2224.940 2917.600 2289.580 ;
        RECT 1469.305 2222.940 2917.200 2224.940 ;
        RECT 1469.305 2158.980 2917.600 2222.940 ;
        RECT 1469.305 2156.980 2917.200 2158.980 ;
        RECT 1469.305 2092.340 2917.600 2156.980 ;
        RECT 1469.305 2090.340 2917.200 2092.340 ;
        RECT 1469.305 2025.700 2917.600 2090.340 ;
        RECT 1469.305 2023.700 2917.200 2025.700 ;
        RECT 1469.305 1959.740 2917.600 2023.700 ;
        RECT 1469.305 1957.740 2917.200 1959.740 ;
        RECT 1469.305 1893.100 2917.600 1957.740 ;
        RECT 1469.305 1891.100 2917.200 1893.100 ;
        RECT 1469.305 1826.460 2917.600 1891.100 ;
        RECT 1469.305 1824.460 2917.200 1826.460 ;
        RECT 1469.305 1760.500 2917.600 1824.460 ;
        RECT 1469.305 1758.500 2917.200 1760.500 ;
        RECT 1469.305 1693.860 2917.600 1758.500 ;
        RECT 1469.305 1691.860 2917.200 1693.860 ;
        RECT 1469.305 1627.220 2917.600 1691.860 ;
        RECT 1469.305 1625.220 2917.200 1627.220 ;
        RECT 1469.305 1561.260 2917.600 1625.220 ;
        RECT 1469.305 1559.260 2917.200 1561.260 ;
        RECT 1469.305 1494.620 2917.600 1559.260 ;
        RECT 1469.305 1492.620 2917.200 1494.620 ;
        RECT 1469.305 1427.980 2917.600 1492.620 ;
        RECT 1469.305 1425.980 2917.200 1427.980 ;
        RECT 1469.305 1362.020 2917.600 1425.980 ;
        RECT 1469.305 1360.020 2917.200 1362.020 ;
        RECT 1469.305 1295.380 2917.600 1360.020 ;
        RECT 1469.305 1293.380 2917.200 1295.380 ;
        RECT 1469.305 1228.740 2917.600 1293.380 ;
        RECT 1469.305 1226.740 2917.200 1228.740 ;
        RECT 1469.305 1162.780 2917.600 1226.740 ;
        RECT 1469.305 1160.780 2917.200 1162.780 ;
        RECT 1469.305 1096.140 2917.600 1160.780 ;
        RECT 1469.305 1094.140 2917.200 1096.140 ;
        RECT 1469.305 1029.500 2917.600 1094.140 ;
        RECT 1469.305 1027.500 2917.200 1029.500 ;
        RECT 1469.305 963.540 2917.600 1027.500 ;
        RECT 1469.305 961.540 2917.200 963.540 ;
        RECT 1469.305 896.900 2917.600 961.540 ;
        RECT 1469.305 894.900 2917.200 896.900 ;
        RECT 1469.305 830.260 2917.600 894.900 ;
        RECT 1469.305 828.260 2917.200 830.260 ;
        RECT 1469.305 764.300 2917.600 828.260 ;
        RECT 1469.305 762.300 2917.200 764.300 ;
        RECT 1469.305 697.660 2917.600 762.300 ;
        RECT 1469.305 695.660 2917.200 697.660 ;
        RECT 1469.305 631.020 2917.600 695.660 ;
        RECT 1469.305 629.020 2917.200 631.020 ;
        RECT 1469.305 565.060 2917.600 629.020 ;
        RECT 1469.305 563.060 2917.200 565.060 ;
        RECT 1469.305 498.420 2917.600 563.060 ;
        RECT 1469.305 496.420 2917.200 498.420 ;
        RECT 1469.305 431.780 2917.600 496.420 ;
        RECT 1469.305 429.780 2917.200 431.780 ;
        RECT 1469.305 365.820 2917.600 429.780 ;
        RECT 1469.305 363.820 2917.200 365.820 ;
        RECT 1469.305 299.180 2917.600 363.820 ;
        RECT 1469.305 297.180 2917.200 299.180 ;
        RECT 1469.305 232.540 2917.600 297.180 ;
        RECT 1469.305 230.540 2917.200 232.540 ;
        RECT 1469.305 166.580 2917.600 230.540 ;
        RECT 1469.305 164.580 2917.200 166.580 ;
        RECT 1469.305 99.940 2917.600 164.580 ;
        RECT 1469.305 97.940 2917.200 99.940 ;
        RECT 1469.305 33.980 2917.600 97.940 ;
        RECT 1469.305 32.815 2917.200 33.980 ;
      LAYER met4 ;
        RECT 1481.415 1842.800 1483.980 2098.160 ;
        RECT 1486.380 1842.800 1510.320 2098.160 ;
        RECT 1512.720 1842.800 1518.980 2098.160 ;
        RECT 1521.380 1842.800 1545.320 2098.160 ;
        RECT 1547.720 1842.800 1553.980 2098.160 ;
        RECT 1481.415 1842.335 1553.980 1842.800 ;
        RECT 1556.380 1842.335 1580.320 2098.160 ;
        RECT 1481.415 1821.580 1580.320 1842.335 ;
        RECT 1481.415 1002.800 1483.980 1821.580 ;
        RECT 1486.380 1002.800 1510.320 1821.580 ;
        RECT 1512.720 1002.800 1518.980 1821.580 ;
        RECT 1521.380 1002.800 1545.320 1821.580 ;
        RECT 1547.720 1002.800 1553.980 1821.580 ;
        RECT 1481.415 1002.335 1553.980 1002.800 ;
        RECT 1556.380 1002.335 1580.320 1821.580 ;
        RECT 1481.415 991.780 1580.320 1002.335 ;
        RECT 1582.720 991.780 1588.980 2098.160 ;
        RECT 1591.380 991.780 1615.320 2098.160 ;
        RECT 1617.720 991.780 1623.980 2098.160 ;
        RECT 1626.380 991.780 1650.320 2098.160 ;
        RECT 1652.720 991.780 1658.980 2098.160 ;
        RECT 1661.380 991.780 1685.320 2098.160 ;
        RECT 1687.720 991.780 1693.980 2098.160 ;
        RECT 1696.380 991.780 1720.320 2098.160 ;
        RECT 1722.720 991.780 1728.980 2098.160 ;
        RECT 1731.380 991.780 1755.320 2098.160 ;
        RECT 1757.720 991.780 1763.980 2098.160 ;
        RECT 1766.380 991.780 1790.320 2098.160 ;
        RECT 1792.720 991.780 1798.980 2098.160 ;
        RECT 1801.380 991.780 1825.320 2098.160 ;
        RECT 1827.720 991.780 1833.980 2098.160 ;
        RECT 1836.380 991.780 1860.320 2098.160 ;
        RECT 1862.720 991.780 1868.980 2098.160 ;
        RECT 1871.380 991.780 1895.320 2098.160 ;
        RECT 1897.720 991.780 1903.980 2098.160 ;
        RECT 1906.380 991.780 1930.320 2098.160 ;
        RECT 1932.720 991.780 1938.980 2098.160 ;
        RECT 1941.380 991.780 1965.320 2098.160 ;
        RECT 1967.720 991.780 1973.980 2098.160 ;
        RECT 1976.380 991.780 2000.320 2098.160 ;
        RECT 2002.720 991.780 2008.980 2098.160 ;
        RECT 2011.380 991.780 2035.320 2098.160 ;
        RECT 2037.720 991.780 2043.980 2098.160 ;
        RECT 2046.380 991.780 2070.320 2098.160 ;
        RECT 2072.720 991.780 2078.980 2098.160 ;
        RECT 2081.380 991.780 2105.320 2098.160 ;
        RECT 2107.720 991.780 2113.980 2098.160 ;
        RECT 2116.380 991.780 2140.320 2098.160 ;
        RECT 2142.720 991.780 2148.980 2098.160 ;
        RECT 2151.380 991.780 2175.320 2098.160 ;
        RECT 2177.720 991.780 2183.980 2098.160 ;
        RECT 2186.380 991.780 2210.320 2098.160 ;
        RECT 2212.720 991.780 2218.980 2098.160 ;
        RECT 2221.380 991.780 2245.320 2098.160 ;
        RECT 2247.720 991.780 2253.980 2098.160 ;
        RECT 2256.380 991.780 2280.320 2098.160 ;
        RECT 2282.720 991.780 2288.980 2098.160 ;
        RECT 2291.380 991.780 2315.320 2098.160 ;
        RECT 2317.720 991.780 2323.980 2098.160 ;
        RECT 2326.380 991.780 2350.320 2098.160 ;
        RECT 2352.720 991.780 2358.980 2098.160 ;
        RECT 2361.380 991.780 2385.320 2098.160 ;
        RECT 2387.720 991.780 2393.980 2098.160 ;
        RECT 2396.380 991.780 2420.320 2098.160 ;
        RECT 2422.720 991.780 2428.980 2098.160 ;
        RECT 2431.380 991.780 2455.320 2098.160 ;
        RECT 2457.720 991.780 2463.980 2098.160 ;
        RECT 2466.380 991.780 2490.320 2098.160 ;
        RECT 2492.720 991.780 2498.980 2098.160 ;
        RECT 2501.380 991.780 2525.320 2098.160 ;
        RECT 2527.720 991.780 2533.980 2098.160 ;
        RECT 2536.380 991.780 2560.320 2098.160 ;
        RECT 2562.720 991.780 2568.980 2098.160 ;
        RECT 2571.380 991.780 2595.320 2098.160 ;
        RECT 2597.720 2000.440 2634.960 2098.160 ;
        RECT 2597.720 1908.360 2603.980 2000.440 ;
        RECT 2606.380 1908.360 2630.320 2000.440 ;
        RECT 2632.720 1908.360 2634.960 2000.440 ;
        RECT 2597.720 1800.440 2634.960 1908.360 ;
        RECT 2597.720 1708.360 2603.980 1800.440 ;
        RECT 2606.380 1708.360 2630.320 1800.440 ;
        RECT 2632.720 1708.360 2634.960 1800.440 ;
        RECT 2597.720 1600.440 2634.960 1708.360 ;
        RECT 2597.720 1508.360 2603.980 1600.440 ;
        RECT 2606.380 1508.360 2630.320 1600.440 ;
        RECT 2632.720 1508.360 2634.960 1600.440 ;
        RECT 2597.720 1400.440 2634.960 1508.360 ;
        RECT 2597.720 1308.360 2603.980 1400.440 ;
        RECT 2606.380 1308.360 2630.320 1400.440 ;
        RECT 2632.720 1308.360 2634.960 1400.440 ;
        RECT 2597.720 1200.440 2634.960 1308.360 ;
        RECT 2597.720 991.780 2603.980 1200.440 ;
        RECT 2606.380 991.780 2630.320 1200.440 ;
        RECT 2632.720 991.780 2634.960 1200.440 ;
  END
END user_project_wrapper
END LIBRARY

