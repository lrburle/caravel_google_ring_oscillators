magic
tech sky130A
magscale 1 2
timestamp 1604095901
<< checkpaint >>
rect -1267 2461 1310 2601
rect -1760 -1129 6260 2461
rect -1267 -1260 1310 -1129
<< error_p >>
rect 0 1271 44 1332
rect 50 581 161 1341
rect 0 0 44 61
<< nwell >>
rect -7 485 50 897
<< locali >>
rect 0 827 44 888
rect 0 0 44 61
<< metal1 >>
rect 0 827 44 888
rect 0 0 44 61
<< labels >>
rlabel metal1 22 856 22 856 1 vccd1
rlabel metal1 23 28 23 28 1 vssd1
<< end >>
