VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0.005 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r1 ;
  SIZE 81.78 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 18.11 0.915 18.28 1.085 ;
        RECT 18.105 0.91 18.275 1.08 ;
        RECT 18.105 2.39 18.275 2.56 ;
      LAYER li1 ;
        RECT 18.11 0.915 18.28 1.085 ;
        RECT 18.105 0.57 18.275 1.08 ;
        RECT 18.105 2.39 18.275 3.86 ;
      LAYER met1 ;
        RECT 18.045 2.36 18.335 2.59 ;
        RECT 18.045 0.88 18.335 1.11 ;
        RECT 18.105 0.88 18.275 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 33.89 0.915 34.06 1.085 ;
        RECT 33.885 0.91 34.055 1.08 ;
        RECT 33.885 2.39 34.055 2.56 ;
      LAYER li1 ;
        RECT 33.89 0.915 34.06 1.085 ;
        RECT 33.885 0.57 34.055 1.08 ;
        RECT 33.885 2.39 34.055 3.86 ;
      LAYER met1 ;
        RECT 33.825 2.36 34.115 2.59 ;
        RECT 33.825 0.88 34.115 1.11 ;
        RECT 33.885 0.88 34.055 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 49.665 0.915 49.835 1.085 ;
        RECT 49.66 0.91 49.83 1.08 ;
        RECT 49.66 2.39 49.83 2.56 ;
      LAYER li1 ;
        RECT 49.665 0.915 49.835 1.085 ;
        RECT 49.66 0.57 49.83 1.08 ;
        RECT 49.66 2.39 49.83 3.86 ;
      LAYER met1 ;
        RECT 49.6 2.36 49.89 2.59 ;
        RECT 49.6 0.88 49.89 1.11 ;
        RECT 49.66 0.88 49.83 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 65.45 0.915 65.62 1.085 ;
        RECT 65.445 0.91 65.615 1.08 ;
        RECT 65.445 2.39 65.615 2.56 ;
      LAYER li1 ;
        RECT 65.45 0.915 65.62 1.085 ;
        RECT 65.445 0.57 65.615 1.08 ;
        RECT 65.445 2.39 65.615 3.86 ;
      LAYER met1 ;
        RECT 65.385 2.36 65.675 2.59 ;
        RECT 65.385 0.88 65.675 1.11 ;
        RECT 65.445 0.88 65.615 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 81.235 0.915 81.405 1.085 ;
        RECT 81.23 0.91 81.4 1.08 ;
        RECT 81.23 2.39 81.4 2.56 ;
      LAYER li1 ;
        RECT 81.235 0.915 81.405 1.085 ;
        RECT 81.23 0.57 81.4 1.08 ;
        RECT 81.23 2.39 81.4 3.86 ;
      LAYER met1 ;
        RECT 81.17 2.36 81.46 2.59 ;
        RECT 81.17 0.88 81.46 1.11 ;
        RECT 81.23 0.88 81.4 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 13.87 5.855 14.22 6.205 ;
        RECT 13.865 2.705 14.215 3.055 ;
        RECT 13.94 2.705 14.115 6.205 ;
      LAYER li1 ;
        RECT 13.955 1.66 14.125 2.935 ;
        RECT 13.955 5.945 14.125 7.22 ;
        RECT 9.175 5.945 9.345 7.22 ;
      LAYER met1 ;
        RECT 13.865 2.765 14.355 2.935 ;
        RECT 13.865 2.705 14.215 3.055 ;
        RECT 9.115 5.945 14.355 6.115 ;
        RECT 13.87 5.855 14.22 6.205 ;
        RECT 9.115 5.915 9.405 6.145 ;
      LAYER mcon ;
        RECT 9.175 5.945 9.345 6.115 ;
        RECT 13.955 5.945 14.125 6.115 ;
        RECT 13.955 2.765 14.125 2.935 ;
      LAYER via1 ;
        RECT 13.965 2.805 14.115 2.955 ;
        RECT 13.97 5.955 14.12 6.105 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 29.65 5.855 30 6.205 ;
        RECT 29.645 2.705 29.995 3.055 ;
        RECT 29.72 2.705 29.895 6.205 ;
      LAYER li1 ;
        RECT 29.735 1.66 29.905 2.935 ;
        RECT 29.735 5.945 29.905 7.22 ;
        RECT 24.955 5.945 25.125 7.22 ;
      LAYER met1 ;
        RECT 29.645 2.765 30.135 2.935 ;
        RECT 29.645 2.705 29.995 3.055 ;
        RECT 24.895 5.945 30.135 6.115 ;
        RECT 29.65 5.855 30 6.205 ;
        RECT 24.895 5.915 25.185 6.145 ;
      LAYER mcon ;
        RECT 24.955 5.945 25.125 6.115 ;
        RECT 29.735 5.945 29.905 6.115 ;
        RECT 29.735 2.765 29.905 2.935 ;
      LAYER via1 ;
        RECT 29.745 2.805 29.895 2.955 ;
        RECT 29.75 5.955 29.9 6.105 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 45.425 5.855 45.775 6.205 ;
        RECT 45.42 2.705 45.77 3.055 ;
        RECT 45.495 2.705 45.67 6.205 ;
      LAYER li1 ;
        RECT 45.51 1.66 45.68 2.935 ;
        RECT 45.51 5.945 45.68 7.22 ;
        RECT 40.73 5.945 40.9 7.22 ;
      LAYER met1 ;
        RECT 45.42 2.765 45.91 2.935 ;
        RECT 45.42 2.705 45.77 3.055 ;
        RECT 40.67 5.945 45.91 6.115 ;
        RECT 45.425 5.855 45.775 6.205 ;
        RECT 40.67 5.915 40.96 6.145 ;
      LAYER mcon ;
        RECT 40.73 5.945 40.9 6.115 ;
        RECT 45.51 5.945 45.68 6.115 ;
        RECT 45.51 2.765 45.68 2.935 ;
      LAYER via1 ;
        RECT 45.52 2.805 45.67 2.955 ;
        RECT 45.525 5.955 45.675 6.105 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 61.21 5.855 61.56 6.205 ;
        RECT 61.205 2.705 61.555 3.055 ;
        RECT 61.28 2.705 61.455 6.205 ;
      LAYER li1 ;
        RECT 61.295 1.66 61.465 2.935 ;
        RECT 61.295 5.945 61.465 7.22 ;
        RECT 56.515 5.945 56.685 7.22 ;
      LAYER met1 ;
        RECT 61.205 2.765 61.695 2.935 ;
        RECT 61.205 2.705 61.555 3.055 ;
        RECT 56.455 5.945 61.695 6.115 ;
        RECT 61.21 5.855 61.56 6.205 ;
        RECT 56.455 5.915 56.745 6.145 ;
      LAYER mcon ;
        RECT 56.515 5.945 56.685 6.115 ;
        RECT 61.295 5.945 61.465 6.115 ;
        RECT 61.295 2.765 61.465 2.935 ;
      LAYER via1 ;
        RECT 61.305 2.805 61.455 2.955 ;
        RECT 61.31 5.955 61.46 6.105 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 76.995 5.855 77.345 6.205 ;
        RECT 76.99 2.705 77.34 3.055 ;
        RECT 77.065 2.705 77.24 6.205 ;
      LAYER li1 ;
        RECT 77.08 1.66 77.25 2.935 ;
        RECT 77.08 5.945 77.25 7.22 ;
        RECT 72.3 5.945 72.47 7.22 ;
      LAYER met1 ;
        RECT 76.99 2.765 77.48 2.935 ;
        RECT 76.99 2.705 77.34 3.055 ;
        RECT 72.24 5.945 77.48 6.115 ;
        RECT 76.995 5.855 77.345 6.205 ;
        RECT 72.24 5.915 72.53 6.145 ;
      LAYER mcon ;
        RECT 72.3 5.945 72.47 6.115 ;
        RECT 77.08 5.945 77.25 6.115 ;
        RECT 77.08 2.765 77.25 2.935 ;
      LAYER via1 ;
        RECT 77.09 2.805 77.24 2.955 ;
        RECT 77.095 5.955 77.245 6.105 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.24 5.945 0.41 7.22 ;
      LAYER met1 ;
        RECT 0.18 5.945 0.64 6.115 ;
        RECT 0.18 5.915 0.47 6.145 ;
      LAYER mcon ;
        RECT 0.24 5.945 0.41 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 4.135 81.775 4.745 ;
        RECT 79.64 4.13 81.62 4.75 ;
        RECT 80.8 3.4 80.97 5.48 ;
        RECT 79.81 3.4 79.98 5.48 ;
        RECT 77.07 3.405 77.24 5.475 ;
        RECT 75.27 3.635 75.44 4.745 ;
        RECT 74.31 3.635 74.48 4.745 ;
        RECT 72.29 4.135 72.46 5.475 ;
        RECT 71.87 3.635 72.04 4.745 ;
        RECT 70.87 3.635 71.04 4.745 ;
        RECT 69.91 3.635 70.08 4.745 ;
        RECT 67.47 3.635 67.64 4.745 ;
        RECT 63.855 4.13 65.835 4.75 ;
        RECT 65.015 3.4 65.185 5.48 ;
        RECT 64.025 3.4 64.195 5.48 ;
        RECT 61.285 3.405 61.455 5.475 ;
        RECT 59.485 3.635 59.655 4.745 ;
        RECT 58.525 3.635 58.695 4.745 ;
        RECT 56.505 4.135 56.675 5.475 ;
        RECT 56.085 3.635 56.255 4.745 ;
        RECT 55.085 3.635 55.255 4.745 ;
        RECT 54.125 3.635 54.295 4.745 ;
        RECT 51.685 3.635 51.855 4.745 ;
        RECT 48.07 4.13 50.05 4.75 ;
        RECT 49.23 3.4 49.4 5.48 ;
        RECT 48.24 3.4 48.41 5.48 ;
        RECT 45.5 3.405 45.67 5.475 ;
        RECT 43.7 3.635 43.87 4.745 ;
        RECT 42.74 3.635 42.91 4.745 ;
        RECT 40.72 4.135 40.89 5.475 ;
        RECT 40.3 3.635 40.47 4.745 ;
        RECT 39.3 3.635 39.47 4.745 ;
        RECT 38.34 3.635 38.51 4.745 ;
        RECT 35.9 3.635 36.07 4.745 ;
        RECT 32.295 4.13 34.275 4.75 ;
        RECT 33.455 3.4 33.625 5.48 ;
        RECT 32.465 3.4 32.635 5.48 ;
        RECT 29.725 3.405 29.895 5.475 ;
        RECT 27.925 3.635 28.095 4.745 ;
        RECT 26.965 3.635 27.135 4.745 ;
        RECT 24.945 4.135 25.115 5.475 ;
        RECT 24.525 3.635 24.695 4.745 ;
        RECT 23.525 3.635 23.695 4.745 ;
        RECT 22.565 3.635 22.735 4.745 ;
        RECT 20.125 3.635 20.295 4.745 ;
        RECT 16.515 4.13 18.495 4.75 ;
        RECT 17.675 3.4 17.845 5.48 ;
        RECT 16.685 3.4 16.855 5.48 ;
        RECT 13.945 3.405 14.115 5.475 ;
        RECT 12.145 3.635 12.315 4.745 ;
        RECT 11.185 3.635 11.355 4.745 ;
        RECT 9.165 4.135 9.335 5.475 ;
        RECT 8.745 3.635 8.915 4.745 ;
        RECT 7.745 3.635 7.915 4.745 ;
        RECT 6.785 3.635 6.955 4.745 ;
        RECT 4.345 3.635 4.515 4.745 ;
        RECT 2.04 4.135 2.21 8.305 ;
        RECT 0.23 4.135 0.4 5.475 ;
      LAYER met1 ;
        RECT 0 4.135 81.775 4.745 ;
        RECT 79.64 4.13 81.62 4.75 ;
        RECT 66.18 3.98 75.84 4.745 ;
        RECT 63.855 4.13 65.835 4.75 ;
        RECT 50.395 3.98 60.055 4.745 ;
        RECT 48.07 4.13 50.05 4.75 ;
        RECT 34.61 3.98 44.27 4.745 ;
        RECT 32.295 4.13 34.275 4.75 ;
        RECT 18.835 3.98 28.495 4.745 ;
        RECT 16.515 4.13 18.495 4.75 ;
        RECT 3.055 3.98 12.715 4.745 ;
        RECT 1.98 6.655 2.27 6.885 ;
        RECT 1.81 6.685 2.27 6.855 ;
      LAYER mcon ;
        RECT 0.315 4.36 0.485 4.53 ;
        RECT 1.45 4.355 1.62 4.525 ;
        RECT 2.04 6.685 2.21 6.855 ;
        RECT 2.35 4.545 2.52 4.715 ;
        RECT 3.2 4.135 3.37 4.305 ;
        RECT 3.66 4.135 3.83 4.305 ;
        RECT 4.12 4.135 4.29 4.305 ;
        RECT 4.58 4.135 4.75 4.305 ;
        RECT 5.04 4.135 5.21 4.305 ;
        RECT 5.5 4.135 5.67 4.305 ;
        RECT 5.96 4.135 6.13 4.305 ;
        RECT 6.42 4.135 6.59 4.305 ;
        RECT 6.88 4.135 7.05 4.305 ;
        RECT 7.34 4.135 7.51 4.305 ;
        RECT 7.8 4.135 7.97 4.305 ;
        RECT 8.26 4.135 8.43 4.305 ;
        RECT 8.72 4.135 8.89 4.305 ;
        RECT 9.18 4.135 9.35 4.305 ;
        RECT 9.64 4.135 9.81 4.305 ;
        RECT 10.1 4.135 10.27 4.305 ;
        RECT 10.56 4.135 10.73 4.305 ;
        RECT 11.02 4.135 11.19 4.305 ;
        RECT 11.285 4.545 11.455 4.715 ;
        RECT 11.48 4.135 11.65 4.305 ;
        RECT 11.94 4.135 12.11 4.305 ;
        RECT 12.4 4.135 12.57 4.305 ;
        RECT 16.065 4.545 16.235 4.715 ;
        RECT 16.065 4.165 16.235 4.335 ;
        RECT 16.765 4.55 16.935 4.72 ;
        RECT 16.765 4.16 16.935 4.33 ;
        RECT 17.755 4.55 17.925 4.72 ;
        RECT 17.755 4.16 17.925 4.33 ;
        RECT 18.98 4.135 19.15 4.305 ;
        RECT 19.44 4.135 19.61 4.305 ;
        RECT 19.9 4.135 20.07 4.305 ;
        RECT 20.36 4.135 20.53 4.305 ;
        RECT 20.82 4.135 20.99 4.305 ;
        RECT 21.28 4.135 21.45 4.305 ;
        RECT 21.74 4.135 21.91 4.305 ;
        RECT 22.2 4.135 22.37 4.305 ;
        RECT 22.66 4.135 22.83 4.305 ;
        RECT 23.12 4.135 23.29 4.305 ;
        RECT 23.58 4.135 23.75 4.305 ;
        RECT 24.04 4.135 24.21 4.305 ;
        RECT 24.5 4.135 24.67 4.305 ;
        RECT 24.96 4.135 25.13 4.305 ;
        RECT 25.42 4.135 25.59 4.305 ;
        RECT 25.88 4.135 26.05 4.305 ;
        RECT 26.34 4.135 26.51 4.305 ;
        RECT 26.8 4.135 26.97 4.305 ;
        RECT 27.065 4.545 27.235 4.715 ;
        RECT 27.26 4.135 27.43 4.305 ;
        RECT 27.72 4.135 27.89 4.305 ;
        RECT 28.18 4.135 28.35 4.305 ;
        RECT 31.845 4.545 32.015 4.715 ;
        RECT 31.845 4.165 32.015 4.335 ;
        RECT 32.545 4.55 32.715 4.72 ;
        RECT 32.545 4.16 32.715 4.33 ;
        RECT 33.535 4.55 33.705 4.72 ;
        RECT 33.535 4.16 33.705 4.33 ;
        RECT 34.755 4.135 34.925 4.305 ;
        RECT 35.215 4.135 35.385 4.305 ;
        RECT 35.675 4.135 35.845 4.305 ;
        RECT 36.135 4.135 36.305 4.305 ;
        RECT 36.595 4.135 36.765 4.305 ;
        RECT 37.055 4.135 37.225 4.305 ;
        RECT 37.515 4.135 37.685 4.305 ;
        RECT 37.975 4.135 38.145 4.305 ;
        RECT 38.435 4.135 38.605 4.305 ;
        RECT 38.895 4.135 39.065 4.305 ;
        RECT 39.355 4.135 39.525 4.305 ;
        RECT 39.815 4.135 39.985 4.305 ;
        RECT 40.275 4.135 40.445 4.305 ;
        RECT 40.735 4.135 40.905 4.305 ;
        RECT 41.195 4.135 41.365 4.305 ;
        RECT 41.655 4.135 41.825 4.305 ;
        RECT 42.115 4.135 42.285 4.305 ;
        RECT 42.575 4.135 42.745 4.305 ;
        RECT 42.84 4.545 43.01 4.715 ;
        RECT 43.035 4.135 43.205 4.305 ;
        RECT 43.495 4.135 43.665 4.305 ;
        RECT 43.955 4.135 44.125 4.305 ;
        RECT 47.62 4.545 47.79 4.715 ;
        RECT 47.62 4.165 47.79 4.335 ;
        RECT 48.32 4.55 48.49 4.72 ;
        RECT 48.32 4.16 48.49 4.33 ;
        RECT 49.31 4.55 49.48 4.72 ;
        RECT 49.31 4.16 49.48 4.33 ;
        RECT 50.54 4.135 50.71 4.305 ;
        RECT 51 4.135 51.17 4.305 ;
        RECT 51.46 4.135 51.63 4.305 ;
        RECT 51.92 4.135 52.09 4.305 ;
        RECT 52.38 4.135 52.55 4.305 ;
        RECT 52.84 4.135 53.01 4.305 ;
        RECT 53.3 4.135 53.47 4.305 ;
        RECT 53.76 4.135 53.93 4.305 ;
        RECT 54.22 4.135 54.39 4.305 ;
        RECT 54.68 4.135 54.85 4.305 ;
        RECT 55.14 4.135 55.31 4.305 ;
        RECT 55.6 4.135 55.77 4.305 ;
        RECT 56.06 4.135 56.23 4.305 ;
        RECT 56.52 4.135 56.69 4.305 ;
        RECT 56.98 4.135 57.15 4.305 ;
        RECT 57.44 4.135 57.61 4.305 ;
        RECT 57.9 4.135 58.07 4.305 ;
        RECT 58.36 4.135 58.53 4.305 ;
        RECT 58.625 4.545 58.795 4.715 ;
        RECT 58.82 4.135 58.99 4.305 ;
        RECT 59.28 4.135 59.45 4.305 ;
        RECT 59.74 4.135 59.91 4.305 ;
        RECT 63.405 4.545 63.575 4.715 ;
        RECT 63.405 4.165 63.575 4.335 ;
        RECT 64.105 4.55 64.275 4.72 ;
        RECT 64.105 4.16 64.275 4.33 ;
        RECT 65.095 4.55 65.265 4.72 ;
        RECT 65.095 4.16 65.265 4.33 ;
        RECT 66.325 4.135 66.495 4.305 ;
        RECT 66.785 4.135 66.955 4.305 ;
        RECT 67.245 4.135 67.415 4.305 ;
        RECT 67.705 4.135 67.875 4.305 ;
        RECT 68.165 4.135 68.335 4.305 ;
        RECT 68.625 4.135 68.795 4.305 ;
        RECT 69.085 4.135 69.255 4.305 ;
        RECT 69.545 4.135 69.715 4.305 ;
        RECT 70.005 4.135 70.175 4.305 ;
        RECT 70.465 4.135 70.635 4.305 ;
        RECT 70.925 4.135 71.095 4.305 ;
        RECT 71.385 4.135 71.555 4.305 ;
        RECT 71.845 4.135 72.015 4.305 ;
        RECT 72.305 4.135 72.475 4.305 ;
        RECT 72.765 4.135 72.935 4.305 ;
        RECT 73.225 4.135 73.395 4.305 ;
        RECT 73.685 4.135 73.855 4.305 ;
        RECT 74.145 4.135 74.315 4.305 ;
        RECT 74.41 4.545 74.58 4.715 ;
        RECT 74.605 4.135 74.775 4.305 ;
        RECT 75.065 4.135 75.235 4.305 ;
        RECT 75.525 4.135 75.695 4.305 ;
        RECT 79.19 4.545 79.36 4.715 ;
        RECT 79.19 4.165 79.36 4.335 ;
        RECT 79.89 4.55 80.06 4.72 ;
        RECT 79.89 4.16 80.06 4.33 ;
        RECT 80.88 4.55 81.05 4.72 ;
        RECT 80.88 4.16 81.05 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -0.005 8.58 81.775 8.88 ;
        RECT 81.595 8.575 81.775 8.88 ;
        RECT 80.8 7.95 80.97 8.88 ;
        RECT 79.81 7.95 79.98 8.88 ;
        RECT 65.81 8.575 79.645 8.88 ;
        RECT 77.07 7.945 77.24 8.88 ;
        RECT 72.29 7.945 72.46 8.88 ;
        RECT 65.015 7.95 65.185 8.88 ;
        RECT 64.025 7.95 64.195 8.88 ;
        RECT 50.025 8.575 63.86 8.88 ;
        RECT 61.285 7.945 61.455 8.88 ;
        RECT 56.505 7.945 56.675 8.88 ;
        RECT 49.23 7.95 49.4 8.88 ;
        RECT 48.24 7.95 48.41 8.88 ;
        RECT 34.25 8.575 48.075 8.88 ;
        RECT 45.5 7.945 45.67 8.88 ;
        RECT 40.72 7.945 40.89 8.88 ;
        RECT 33.455 7.95 33.625 8.88 ;
        RECT 32.465 7.95 32.635 8.88 ;
        RECT 18.47 8.575 32.3 8.88 ;
        RECT 29.725 7.945 29.895 8.88 ;
        RECT 24.945 7.945 25.115 8.88 ;
        RECT 17.675 7.95 17.845 8.88 ;
        RECT 16.685 7.95 16.855 8.88 ;
        RECT -0.005 8.575 16.52 8.88 ;
        RECT 13.945 7.945 14.115 8.88 ;
        RECT 9.165 7.945 9.335 8.88 ;
        RECT 0.23 7.945 0.4 8.88 ;
        RECT 73.295 6.075 73.465 8.025 ;
        RECT 73.24 7.855 73.41 8.305 ;
        RECT 73.24 5.015 73.41 6.245 ;
        RECT 57.51 6.075 57.68 8.025 ;
        RECT 57.455 7.855 57.625 8.305 ;
        RECT 57.455 5.015 57.625 6.245 ;
        RECT 41.725 6.075 41.895 8.025 ;
        RECT 41.67 7.855 41.84 8.305 ;
        RECT 41.67 5.015 41.84 6.245 ;
        RECT 25.95 6.075 26.12 8.025 ;
        RECT 25.895 7.855 26.065 8.305 ;
        RECT 25.895 5.015 26.065 6.245 ;
        RECT 10.17 6.075 10.34 8.025 ;
        RECT 10.115 7.855 10.285 8.305 ;
        RECT 10.115 5.015 10.285 6.245 ;
      LAYER met1 ;
        RECT -0.005 8.575 81.775 8.88 ;
        RECT 73.235 6.285 73.525 6.515 ;
        RECT 72.865 6.315 73.525 6.485 ;
        RECT 72.865 6.315 73.035 8.88 ;
        RECT 57.45 6.285 57.74 6.515 ;
        RECT 57.08 6.315 57.74 6.485 ;
        RECT 57.08 6.315 57.25 8.88 ;
        RECT 41.665 6.285 41.955 6.515 ;
        RECT 41.295 6.315 41.955 6.485 ;
        RECT 41.295 6.315 41.465 8.88 ;
        RECT 25.89 6.285 26.18 6.515 ;
        RECT 25.52 6.315 26.18 6.485 ;
        RECT 25.52 6.315 25.69 8.88 ;
        RECT 10.11 6.285 10.4 6.515 ;
        RECT 9.74 6.315 10.4 6.485 ;
        RECT 9.74 6.315 9.91 8.88 ;
      LAYER mcon ;
        RECT 0.31 8.605 0.48 8.775 ;
        RECT 0.99 8.605 1.16 8.775 ;
        RECT 1.67 8.605 1.84 8.775 ;
        RECT 2.35 8.605 2.52 8.775 ;
        RECT 9.245 8.605 9.415 8.775 ;
        RECT 9.925 8.605 10.095 8.775 ;
        RECT 10.17 6.315 10.34 6.485 ;
        RECT 10.605 8.605 10.775 8.775 ;
        RECT 11.285 8.605 11.455 8.775 ;
        RECT 14.025 8.605 14.195 8.775 ;
        RECT 14.705 8.605 14.875 8.775 ;
        RECT 15.385 8.605 15.555 8.775 ;
        RECT 16.065 8.605 16.235 8.775 ;
        RECT 16.765 8.61 16.935 8.78 ;
        RECT 17.755 8.61 17.925 8.78 ;
        RECT 25.025 8.605 25.195 8.775 ;
        RECT 25.705 8.605 25.875 8.775 ;
        RECT 25.95 6.315 26.12 6.485 ;
        RECT 26.385 8.605 26.555 8.775 ;
        RECT 27.065 8.605 27.235 8.775 ;
        RECT 29.805 8.605 29.975 8.775 ;
        RECT 30.485 8.605 30.655 8.775 ;
        RECT 31.165 8.605 31.335 8.775 ;
        RECT 31.845 8.605 32.015 8.775 ;
        RECT 32.545 8.61 32.715 8.78 ;
        RECT 33.535 8.61 33.705 8.78 ;
        RECT 40.8 8.605 40.97 8.775 ;
        RECT 41.48 8.605 41.65 8.775 ;
        RECT 41.725 6.315 41.895 6.485 ;
        RECT 42.16 8.605 42.33 8.775 ;
        RECT 42.84 8.605 43.01 8.775 ;
        RECT 45.58 8.605 45.75 8.775 ;
        RECT 46.26 8.605 46.43 8.775 ;
        RECT 46.94 8.605 47.11 8.775 ;
        RECT 47.62 8.605 47.79 8.775 ;
        RECT 48.32 8.61 48.49 8.78 ;
        RECT 49.31 8.61 49.48 8.78 ;
        RECT 56.585 8.605 56.755 8.775 ;
        RECT 57.265 8.605 57.435 8.775 ;
        RECT 57.51 6.315 57.68 6.485 ;
        RECT 57.945 8.605 58.115 8.775 ;
        RECT 58.625 8.605 58.795 8.775 ;
        RECT 61.365 8.605 61.535 8.775 ;
        RECT 62.045 8.605 62.215 8.775 ;
        RECT 62.725 8.605 62.895 8.775 ;
        RECT 63.405 8.605 63.575 8.775 ;
        RECT 64.105 8.61 64.275 8.78 ;
        RECT 65.095 8.61 65.265 8.78 ;
        RECT 72.37 8.605 72.54 8.775 ;
        RECT 73.05 8.605 73.22 8.775 ;
        RECT 73.295 6.315 73.465 6.485 ;
        RECT 73.73 8.605 73.9 8.775 ;
        RECT 74.41 8.605 74.58 8.775 ;
        RECT 77.15 8.605 77.32 8.775 ;
        RECT 77.83 8.605 78 8.775 ;
        RECT 78.51 8.605 78.68 8.775 ;
        RECT 79.19 8.605 79.36 8.775 ;
        RECT 79.89 8.61 80.06 8.78 ;
        RECT 80.88 8.61 81.05 8.78 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 73.57 7.04 73.94 7.41 ;
      RECT 73.61 6.72 73.945 7.085 ;
      RECT 73.61 6.72 73.995 7.03 ;
      RECT 73.61 6.72 76.4 7.025 ;
      RECT 76.095 2.85 76.4 7.025 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 75.32 0.815 75.625 4.02 ;
      RECT 75.07 2.975 75.625 3.705 ;
      RECT 75.28 0.815 75.65 1.185 ;
      RECT 71.43 1.85 71.76 2.745 ;
      RECT 70.55 2.015 70.88 2.745 ;
      RECT 71.425 1.85 71.795 2.65 ;
      RECT 74.59 1.85 74.92 2.58 ;
      RECT 74.55 1.735 74.73 2.385 ;
      RECT 70.56 1.85 74.92 2.22 ;
      RECT 71.05 3.535 71.38 3.865 ;
      RECT 69.845 3.55 71.38 3.85 ;
      RECT 69.845 2.43 70.145 3.85 ;
      RECT 69.59 2.415 69.92 2.745 ;
      RECT 57.785 7.04 58.155 7.41 ;
      RECT 57.825 6.72 58.16 7.085 ;
      RECT 57.825 6.72 58.21 7.03 ;
      RECT 57.825 6.72 60.615 7.025 ;
      RECT 60.31 2.85 60.615 7.025 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 59.535 0.815 59.84 4.02 ;
      RECT 59.285 2.975 59.84 3.705 ;
      RECT 59.495 0.815 59.865 1.185 ;
      RECT 55.645 1.85 55.975 2.745 ;
      RECT 54.765 2.015 55.095 2.745 ;
      RECT 55.64 1.85 56.01 2.65 ;
      RECT 58.805 1.85 59.135 2.58 ;
      RECT 58.765 1.735 58.945 2.385 ;
      RECT 54.775 1.85 59.135 2.22 ;
      RECT 55.265 3.535 55.595 3.865 ;
      RECT 54.06 3.55 55.595 3.85 ;
      RECT 54.06 2.43 54.36 3.85 ;
      RECT 53.805 2.415 54.135 2.745 ;
      RECT 42 7.04 42.37 7.41 ;
      RECT 42.04 6.72 42.375 7.085 ;
      RECT 42.04 6.72 42.425 7.03 ;
      RECT 42.04 6.72 44.83 7.025 ;
      RECT 44.525 2.85 44.83 7.025 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 43.75 0.815 44.055 4.02 ;
      RECT 43.5 2.975 44.055 3.705 ;
      RECT 43.71 0.815 44.08 1.185 ;
      RECT 39.86 1.85 40.19 2.745 ;
      RECT 38.98 2.015 39.31 2.745 ;
      RECT 39.855 1.85 40.225 2.65 ;
      RECT 43.02 1.85 43.35 2.58 ;
      RECT 42.98 1.735 43.16 2.385 ;
      RECT 38.99 1.85 43.35 2.22 ;
      RECT 39.48 3.535 39.81 3.865 ;
      RECT 38.275 3.55 39.81 3.85 ;
      RECT 38.275 2.43 38.575 3.85 ;
      RECT 38.02 2.415 38.35 2.745 ;
      RECT 26.225 7.04 26.595 7.41 ;
      RECT 26.265 6.72 26.6 7.085 ;
      RECT 26.265 6.72 26.65 7.03 ;
      RECT 26.265 6.72 29.055 7.025 ;
      RECT 28.75 2.85 29.055 7.025 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 27.975 0.815 28.28 4.02 ;
      RECT 27.725 2.975 28.28 3.705 ;
      RECT 27.935 0.815 28.305 1.185 ;
      RECT 24.085 1.85 24.415 2.745 ;
      RECT 23.205 2.015 23.535 2.745 ;
      RECT 24.08 1.85 24.45 2.65 ;
      RECT 27.245 1.85 27.575 2.58 ;
      RECT 27.205 1.735 27.385 2.385 ;
      RECT 23.215 1.85 27.575 2.22 ;
      RECT 23.705 3.535 24.035 3.865 ;
      RECT 22.5 3.55 24.035 3.85 ;
      RECT 22.5 2.43 22.8 3.85 ;
      RECT 22.245 2.415 22.575 2.745 ;
      RECT 10.445 7.04 10.815 7.41 ;
      RECT 10.485 6.72 10.82 7.085 ;
      RECT 10.485 6.72 10.87 7.03 ;
      RECT 10.485 6.72 13.275 7.025 ;
      RECT 12.97 2.85 13.275 7.025 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 12.195 0.815 12.5 4.02 ;
      RECT 11.945 2.975 12.5 3.705 ;
      RECT 12.155 0.815 12.525 1.185 ;
      RECT 8.305 1.85 8.635 2.745 ;
      RECT 7.425 2.015 7.755 2.745 ;
      RECT 8.3 1.85 8.67 2.65 ;
      RECT 11.465 1.85 11.795 2.58 ;
      RECT 11.425 1.735 11.605 2.385 ;
      RECT 7.435 1.85 11.795 2.22 ;
      RECT 7.925 3.535 8.255 3.865 ;
      RECT 6.72 3.55 8.255 3.85 ;
      RECT 6.72 2.43 7.02 3.85 ;
      RECT 6.465 2.415 6.795 2.745 ;
      RECT 72.99 2.575 73.32 3.305 ;
      RECT 68.87 2.415 69.2 3.145 ;
      RECT 67.87 1.855 68.2 2.585 ;
      RECT 66.43 2.575 66.76 3.305 ;
      RECT 57.205 2.575 57.535 3.305 ;
      RECT 53.085 2.415 53.415 3.145 ;
      RECT 52.085 1.855 52.415 2.585 ;
      RECT 50.645 2.575 50.975 3.305 ;
      RECT 41.42 2.575 41.75 3.305 ;
      RECT 37.3 2.415 37.63 3.145 ;
      RECT 36.3 1.855 36.63 2.585 ;
      RECT 34.86 2.575 35.19 3.305 ;
      RECT 25.645 2.575 25.975 3.305 ;
      RECT 21.525 2.415 21.855 3.145 ;
      RECT 20.525 1.855 20.855 2.585 ;
      RECT 19.085 2.575 19.415 3.305 ;
      RECT 9.865 2.575 10.195 3.305 ;
      RECT 5.745 2.415 6.075 3.145 ;
      RECT 4.745 1.855 5.075 2.585 ;
      RECT 3.305 2.575 3.635 3.305 ;
    LAYER via2 ;
      RECT 76.145 2.935 76.345 3.135 ;
      RECT 75.365 0.9 75.565 1.1 ;
      RECT 75.135 3.04 75.335 3.24 ;
      RECT 74.655 2.315 74.855 2.515 ;
      RECT 73.655 7.125 73.855 7.325 ;
      RECT 73.055 3.04 73.255 3.24 ;
      RECT 71.495 2.48 71.695 2.68 ;
      RECT 71.115 3.6 71.315 3.8 ;
      RECT 70.615 2.48 70.815 2.68 ;
      RECT 69.655 2.48 69.855 2.68 ;
      RECT 68.935 2.48 69.135 2.68 ;
      RECT 67.935 1.92 68.135 2.12 ;
      RECT 66.495 3.04 66.695 3.24 ;
      RECT 60.36 2.935 60.56 3.135 ;
      RECT 59.58 0.9 59.78 1.1 ;
      RECT 59.35 3.04 59.55 3.24 ;
      RECT 58.87 2.315 59.07 2.515 ;
      RECT 57.87 7.125 58.07 7.325 ;
      RECT 57.27 3.04 57.47 3.24 ;
      RECT 55.71 2.48 55.91 2.68 ;
      RECT 55.33 3.6 55.53 3.8 ;
      RECT 54.83 2.48 55.03 2.68 ;
      RECT 53.87 2.48 54.07 2.68 ;
      RECT 53.15 2.48 53.35 2.68 ;
      RECT 52.15 1.92 52.35 2.12 ;
      RECT 50.71 3.04 50.91 3.24 ;
      RECT 44.575 2.935 44.775 3.135 ;
      RECT 43.795 0.9 43.995 1.1 ;
      RECT 43.565 3.04 43.765 3.24 ;
      RECT 43.085 2.315 43.285 2.515 ;
      RECT 42.085 7.125 42.285 7.325 ;
      RECT 41.485 3.04 41.685 3.24 ;
      RECT 39.925 2.48 40.125 2.68 ;
      RECT 39.545 3.6 39.745 3.8 ;
      RECT 39.045 2.48 39.245 2.68 ;
      RECT 38.085 2.48 38.285 2.68 ;
      RECT 37.365 2.48 37.565 2.68 ;
      RECT 36.365 1.92 36.565 2.12 ;
      RECT 34.925 3.04 35.125 3.24 ;
      RECT 28.8 2.935 29 3.135 ;
      RECT 28.02 0.9 28.22 1.1 ;
      RECT 27.79 3.04 27.99 3.24 ;
      RECT 27.31 2.315 27.51 2.515 ;
      RECT 26.31 7.125 26.51 7.325 ;
      RECT 25.71 3.04 25.91 3.24 ;
      RECT 24.15 2.48 24.35 2.68 ;
      RECT 23.77 3.6 23.97 3.8 ;
      RECT 23.27 2.48 23.47 2.68 ;
      RECT 22.31 2.48 22.51 2.68 ;
      RECT 21.59 2.48 21.79 2.68 ;
      RECT 20.59 1.92 20.79 2.12 ;
      RECT 19.15 3.04 19.35 3.24 ;
      RECT 13.02 2.935 13.22 3.135 ;
      RECT 12.24 0.9 12.44 1.1 ;
      RECT 12.01 3.04 12.21 3.24 ;
      RECT 11.53 2.315 11.73 2.515 ;
      RECT 10.53 7.125 10.73 7.325 ;
      RECT 9.93 3.04 10.13 3.24 ;
      RECT 8.37 2.48 8.57 2.68 ;
      RECT 7.99 3.6 8.19 3.8 ;
      RECT 7.49 2.48 7.69 2.68 ;
      RECT 6.53 2.48 6.73 2.68 ;
      RECT 5.81 2.48 6.01 2.68 ;
      RECT 4.81 1.92 5.01 2.12 ;
      RECT 3.37 3.04 3.57 3.24 ;
    LAYER met2 ;
      RECT 1.24 8.4 81.405 8.57 ;
      RECT 81.235 7.275 81.405 8.57 ;
      RECT 1.24 6.255 1.41 8.57 ;
      RECT 81.205 7.275 81.555 7.625 ;
      RECT 1.175 6.255 1.465 6.605 ;
      RECT 78.045 6.22 78.365 6.545 ;
      RECT 78.075 5.695 78.245 6.545 ;
      RECT 78.075 5.695 78.25 6.045 ;
      RECT 78.075 5.695 79.05 5.87 ;
      RECT 78.875 1.965 79.05 5.87 ;
      RECT 78.82 1.965 79.17 2.315 ;
      RECT 78.845 6.655 79.17 6.98 ;
      RECT 77.73 6.745 79.17 6.915 ;
      RECT 77.73 2.395 77.89 6.915 ;
      RECT 78.045 2.365 78.365 2.685 ;
      RECT 77.73 2.395 78.365 2.565 ;
      RECT 67.815 1.92 68.075 2.18 ;
      RECT 67.87 1.88 68.175 2.16 ;
      RECT 67.87 1.42 68.045 2.18 ;
      RECT 76.385 1.34 76.735 1.69 ;
      RECT 67.87 1.42 76.735 1.595 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 76.145 2.235 76.315 3.22 ;
      RECT 72.165 2.455 72.4 2.715 ;
      RECT 75.31 2.235 75.475 2.495 ;
      RECT 75.215 2.225 75.23 2.495 ;
      RECT 75.31 2.235 76.315 2.415 ;
      RECT 73.815 1.795 73.855 1.935 ;
      RECT 75.23 2.23 75.31 2.495 ;
      RECT 75.175 2.225 75.215 2.461 ;
      RECT 75.161 2.225 75.175 2.461 ;
      RECT 75.075 2.23 75.161 2.463 ;
      RECT 75.03 2.237 75.075 2.465 ;
      RECT 75 2.237 75.03 2.467 ;
      RECT 74.975 2.232 75 2.469 ;
      RECT 74.945 2.228 74.975 2.478 ;
      RECT 74.935 2.225 74.945 2.49 ;
      RECT 74.93 2.225 74.935 2.498 ;
      RECT 74.925 2.225 74.93 2.503 ;
      RECT 74.915 2.224 74.925 2.513 ;
      RECT 74.91 2.223 74.915 2.523 ;
      RECT 74.895 2.222 74.91 2.528 ;
      RECT 74.867 2.219 74.895 2.555 ;
      RECT 74.781 2.211 74.867 2.555 ;
      RECT 74.695 2.2 74.781 2.555 ;
      RECT 74.655 2.185 74.695 2.555 ;
      RECT 74.615 2.159 74.655 2.555 ;
      RECT 74.61 2.141 74.615 2.367 ;
      RECT 74.6 2.137 74.61 2.357 ;
      RECT 74.585 2.127 74.6 2.344 ;
      RECT 74.565 2.111 74.585 2.329 ;
      RECT 74.55 2.096 74.565 2.314 ;
      RECT 74.54 2.085 74.55 2.304 ;
      RECT 74.515 2.069 74.54 2.293 ;
      RECT 74.51 2.056 74.515 2.283 ;
      RECT 74.505 2.052 74.51 2.278 ;
      RECT 74.45 2.038 74.505 2.256 ;
      RECT 74.411 2.019 74.45 2.22 ;
      RECT 74.325 1.993 74.411 2.173 ;
      RECT 74.321 1.975 74.325 2.139 ;
      RECT 74.235 1.956 74.321 2.117 ;
      RECT 74.23 1.938 74.235 2.095 ;
      RECT 74.225 1.936 74.23 2.093 ;
      RECT 74.215 1.935 74.225 2.088 ;
      RECT 74.155 1.922 74.215 2.074 ;
      RECT 74.11 1.9 74.155 2.053 ;
      RECT 74.05 1.877 74.11 2.032 ;
      RECT 73.986 1.852 74.05 2.007 ;
      RECT 73.9 1.822 73.986 1.976 ;
      RECT 73.885 1.802 73.9 1.955 ;
      RECT 73.855 1.797 73.885 1.946 ;
      RECT 73.802 1.795 73.815 1.935 ;
      RECT 73.716 1.795 73.802 1.937 ;
      RECT 73.63 1.795 73.716 1.939 ;
      RECT 73.61 1.795 73.63 1.943 ;
      RECT 73.565 1.797 73.61 1.954 ;
      RECT 73.525 1.807 73.565 1.97 ;
      RECT 73.521 1.816 73.525 1.978 ;
      RECT 73.435 1.836 73.521 1.994 ;
      RECT 73.425 1.855 73.435 2.012 ;
      RECT 73.42 1.857 73.425 2.015 ;
      RECT 73.41 1.861 73.42 2.018 ;
      RECT 73.39 1.866 73.41 2.028 ;
      RECT 73.36 1.876 73.39 2.048 ;
      RECT 73.355 1.883 73.36 2.062 ;
      RECT 73.345 1.887 73.355 2.069 ;
      RECT 73.33 1.895 73.345 2.08 ;
      RECT 73.32 1.905 73.33 2.091 ;
      RECT 73.31 1.912 73.32 2.099 ;
      RECT 73.285 1.925 73.31 2.114 ;
      RECT 73.221 1.961 73.285 2.153 ;
      RECT 73.135 2.024 73.221 2.217 ;
      RECT 73.1 2.075 73.135 2.27 ;
      RECT 73.095 2.092 73.1 2.287 ;
      RECT 73.08 2.101 73.095 2.294 ;
      RECT 73.06 2.116 73.08 2.308 ;
      RECT 73.055 2.127 73.06 2.318 ;
      RECT 73.035 2.14 73.055 2.328 ;
      RECT 73.03 2.15 73.035 2.338 ;
      RECT 73.015 2.155 73.03 2.347 ;
      RECT 73.005 2.165 73.015 2.358 ;
      RECT 72.975 2.182 73.005 2.375 ;
      RECT 72.965 2.2 72.975 2.393 ;
      RECT 72.95 2.211 72.965 2.404 ;
      RECT 72.91 2.235 72.95 2.42 ;
      RECT 72.875 2.269 72.91 2.437 ;
      RECT 72.845 2.292 72.875 2.449 ;
      RECT 72.83 2.302 72.845 2.458 ;
      RECT 72.79 2.312 72.83 2.469 ;
      RECT 72.77 2.323 72.79 2.481 ;
      RECT 72.765 2.327 72.77 2.488 ;
      RECT 72.75 2.331 72.765 2.493 ;
      RECT 72.74 2.336 72.75 2.498 ;
      RECT 72.735 2.339 72.74 2.501 ;
      RECT 72.705 2.345 72.735 2.508 ;
      RECT 72.67 2.355 72.705 2.522 ;
      RECT 72.61 2.37 72.67 2.542 ;
      RECT 72.555 2.39 72.61 2.566 ;
      RECT 72.526 2.405 72.555 2.584 ;
      RECT 72.44 2.425 72.526 2.609 ;
      RECT 72.435 2.44 72.44 2.629 ;
      RECT 72.425 2.443 72.435 2.63 ;
      RECT 72.4 2.45 72.425 2.715 ;
      RECT 75.095 2.943 75.375 3.28 ;
      RECT 75.095 2.953 75.38 3.238 ;
      RECT 75.095 2.962 75.385 3.135 ;
      RECT 75.095 2.977 75.39 3.003 ;
      RECT 75.095 2.805 75.355 3.28 ;
      RECT 65.395 6.655 65.745 7.005 ;
      RECT 74.22 6.61 74.57 6.96 ;
      RECT 65.395 6.685 74.57 6.885 ;
      RECT 72.815 3.685 72.825 3.875 ;
      RECT 71.075 3.56 71.355 3.84 ;
      RECT 74.12 2.5 74.125 2.985 ;
      RECT 74.015 2.5 74.075 2.76 ;
      RECT 74.34 3.47 74.345 3.545 ;
      RECT 74.33 3.337 74.34 3.58 ;
      RECT 74.32 3.172 74.33 3.601 ;
      RECT 74.315 3.042 74.32 3.617 ;
      RECT 74.305 2.932 74.315 3.633 ;
      RECT 74.3 2.831 74.305 3.65 ;
      RECT 74.295 2.813 74.3 3.66 ;
      RECT 74.29 2.795 74.295 3.67 ;
      RECT 74.28 2.77 74.29 3.685 ;
      RECT 74.275 2.75 74.28 3.7 ;
      RECT 74.255 2.5 74.275 3.725 ;
      RECT 74.24 2.5 74.255 3.758 ;
      RECT 74.21 2.5 74.24 3.78 ;
      RECT 74.19 2.5 74.21 3.794 ;
      RECT 74.17 2.5 74.19 3.31 ;
      RECT 74.185 3.377 74.19 3.799 ;
      RECT 74.18 3.407 74.185 3.801 ;
      RECT 74.175 3.42 74.18 3.804 ;
      RECT 74.17 3.43 74.175 3.808 ;
      RECT 74.165 2.5 74.17 3.228 ;
      RECT 74.165 3.44 74.17 3.81 ;
      RECT 74.16 2.5 74.165 3.205 ;
      RECT 74.15 3.462 74.165 3.81 ;
      RECT 74.145 2.5 74.16 3.15 ;
      RECT 74.14 3.487 74.15 3.81 ;
      RECT 74.14 2.5 74.145 3.095 ;
      RECT 74.13 2.5 74.14 3.043 ;
      RECT 74.135 3.5 74.14 3.811 ;
      RECT 74.13 3.512 74.135 3.812 ;
      RECT 74.125 2.5 74.13 3.003 ;
      RECT 74.125 3.525 74.13 3.813 ;
      RECT 74.11 3.54 74.125 3.814 ;
      RECT 74.115 2.5 74.12 2.965 ;
      RECT 74.11 2.5 74.115 2.93 ;
      RECT 74.105 2.5 74.11 2.905 ;
      RECT 74.1 3.567 74.11 3.816 ;
      RECT 74.095 2.5 74.105 2.863 ;
      RECT 74.095 3.585 74.1 3.817 ;
      RECT 74.09 2.5 74.095 2.823 ;
      RECT 74.09 3.592 74.095 3.818 ;
      RECT 74.085 2.5 74.09 2.795 ;
      RECT 74.08 3.61 74.09 3.819 ;
      RECT 74.075 2.5 74.085 2.775 ;
      RECT 74.07 3.63 74.08 3.821 ;
      RECT 74.06 3.647 74.07 3.822 ;
      RECT 74.025 3.67 74.06 3.825 ;
      RECT 73.97 3.688 74.025 3.831 ;
      RECT 73.884 3.696 73.97 3.84 ;
      RECT 73.798 3.707 73.884 3.851 ;
      RECT 73.712 3.717 73.798 3.862 ;
      RECT 73.626 3.727 73.712 3.874 ;
      RECT 73.54 3.737 73.626 3.885 ;
      RECT 73.52 3.743 73.54 3.891 ;
      RECT 73.44 3.745 73.52 3.895 ;
      RECT 73.435 3.744 73.44 3.9 ;
      RECT 73.427 3.743 73.435 3.9 ;
      RECT 73.341 3.739 73.427 3.898 ;
      RECT 73.255 3.731 73.341 3.895 ;
      RECT 73.169 3.722 73.255 3.891 ;
      RECT 73.083 3.714 73.169 3.888 ;
      RECT 72.997 3.706 73.083 3.884 ;
      RECT 72.911 3.697 72.997 3.881 ;
      RECT 72.825 3.689 72.911 3.877 ;
      RECT 72.77 3.682 72.815 3.875 ;
      RECT 72.685 3.675 72.77 3.873 ;
      RECT 72.611 3.667 72.685 3.869 ;
      RECT 72.525 3.659 72.611 3.866 ;
      RECT 72.522 3.655 72.525 3.864 ;
      RECT 72.436 3.651 72.522 3.863 ;
      RECT 72.35 3.643 72.436 3.86 ;
      RECT 72.265 3.638 72.35 3.857 ;
      RECT 72.179 3.635 72.265 3.854 ;
      RECT 72.093 3.633 72.179 3.851 ;
      RECT 72.007 3.63 72.093 3.848 ;
      RECT 71.921 3.627 72.007 3.845 ;
      RECT 71.835 3.624 71.921 3.842 ;
      RECT 71.759 3.622 71.835 3.839 ;
      RECT 71.673 3.619 71.759 3.836 ;
      RECT 71.587 3.616 71.673 3.834 ;
      RECT 71.501 3.614 71.587 3.831 ;
      RECT 71.415 3.611 71.501 3.828 ;
      RECT 71.355 3.602 71.415 3.826 ;
      RECT 73.865 3.22 73.94 3.48 ;
      RECT 73.845 3.2 73.85 3.48 ;
      RECT 73.165 2.985 73.27 3.28 ;
      RECT 67.61 2.96 67.68 3.22 ;
      RECT 73.505 2.835 73.51 3.206 ;
      RECT 73.495 2.89 73.5 3.206 ;
      RECT 73.8 2.06 73.86 2.32 ;
      RECT 73.855 3.215 73.865 3.48 ;
      RECT 73.85 3.205 73.855 3.48 ;
      RECT 73.77 3.152 73.845 3.48 ;
      RECT 73.795 2.06 73.8 2.34 ;
      RECT 73.785 2.06 73.795 2.36 ;
      RECT 73.77 2.06 73.785 2.39 ;
      RECT 73.755 2.06 73.77 2.433 ;
      RECT 73.75 3.095 73.77 3.48 ;
      RECT 73.74 2.06 73.755 2.47 ;
      RECT 73.735 3.075 73.75 3.48 ;
      RECT 73.735 2.06 73.74 2.493 ;
      RECT 73.725 2.06 73.735 2.518 ;
      RECT 73.695 3.042 73.735 3.48 ;
      RECT 73.7 2.06 73.725 2.568 ;
      RECT 73.695 2.06 73.7 2.623 ;
      RECT 73.69 2.06 73.695 2.665 ;
      RECT 73.68 3.005 73.695 3.48 ;
      RECT 73.685 2.06 73.69 2.708 ;
      RECT 73.68 2.06 73.685 2.773 ;
      RECT 73.675 2.06 73.68 2.795 ;
      RECT 73.675 2.993 73.68 3.345 ;
      RECT 73.67 2.06 73.675 2.863 ;
      RECT 73.67 2.985 73.675 3.328 ;
      RECT 73.665 2.06 73.67 2.908 ;
      RECT 73.66 2.967 73.67 3.305 ;
      RECT 73.66 2.06 73.665 2.945 ;
      RECT 73.65 2.06 73.66 3.285 ;
      RECT 73.645 2.06 73.65 3.268 ;
      RECT 73.64 2.06 73.645 3.253 ;
      RECT 73.635 2.06 73.64 3.238 ;
      RECT 73.615 2.06 73.635 3.228 ;
      RECT 73.61 2.06 73.615 3.218 ;
      RECT 73.6 2.06 73.61 3.214 ;
      RECT 73.595 2.337 73.6 3.213 ;
      RECT 73.59 2.36 73.595 3.212 ;
      RECT 73.585 2.39 73.59 3.211 ;
      RECT 73.58 2.417 73.585 3.21 ;
      RECT 73.575 2.445 73.58 3.21 ;
      RECT 73.57 2.472 73.575 3.21 ;
      RECT 73.565 2.492 73.57 3.21 ;
      RECT 73.56 2.52 73.565 3.21 ;
      RECT 73.55 2.562 73.56 3.21 ;
      RECT 73.54 2.607 73.55 3.209 ;
      RECT 73.535 2.66 73.54 3.208 ;
      RECT 73.53 2.692 73.535 3.207 ;
      RECT 73.525 2.712 73.53 3.206 ;
      RECT 73.52 2.75 73.525 3.206 ;
      RECT 73.515 2.772 73.52 3.206 ;
      RECT 73.51 2.797 73.515 3.206 ;
      RECT 73.5 2.862 73.505 3.206 ;
      RECT 73.485 2.922 73.495 3.206 ;
      RECT 73.47 2.932 73.485 3.206 ;
      RECT 73.45 2.942 73.47 3.206 ;
      RECT 73.42 2.947 73.45 3.203 ;
      RECT 73.36 2.957 73.42 3.2 ;
      RECT 73.34 2.966 73.36 3.205 ;
      RECT 73.315 2.972 73.34 3.218 ;
      RECT 73.295 2.977 73.315 3.233 ;
      RECT 73.27 2.982 73.295 3.28 ;
      RECT 73.141 2.984 73.165 3.28 ;
      RECT 73.055 2.979 73.141 3.28 ;
      RECT 73.015 2.976 73.055 3.28 ;
      RECT 72.965 2.978 73.015 3.26 ;
      RECT 72.935 2.982 72.965 3.26 ;
      RECT 72.856 2.992 72.935 3.26 ;
      RECT 72.77 3.007 72.856 3.261 ;
      RECT 72.72 3.017 72.77 3.262 ;
      RECT 72.712 3.02 72.72 3.262 ;
      RECT 72.626 3.022 72.712 3.263 ;
      RECT 72.54 3.026 72.626 3.263 ;
      RECT 72.454 3.03 72.54 3.264 ;
      RECT 72.368 3.033 72.454 3.265 ;
      RECT 72.282 3.037 72.368 3.265 ;
      RECT 72.196 3.041 72.282 3.266 ;
      RECT 72.11 3.044 72.196 3.267 ;
      RECT 72.024 3.048 72.11 3.267 ;
      RECT 71.938 3.052 72.024 3.268 ;
      RECT 71.852 3.056 71.938 3.269 ;
      RECT 71.766 3.059 71.852 3.269 ;
      RECT 71.68 3.063 71.766 3.27 ;
      RECT 71.65 3.065 71.68 3.27 ;
      RECT 71.564 3.068 71.65 3.271 ;
      RECT 71.478 3.072 71.564 3.272 ;
      RECT 71.392 3.076 71.478 3.273 ;
      RECT 71.306 3.079 71.392 3.273 ;
      RECT 71.22 3.083 71.306 3.274 ;
      RECT 71.185 3.088 71.22 3.275 ;
      RECT 71.13 3.098 71.185 3.282 ;
      RECT 71.105 3.11 71.13 3.292 ;
      RECT 71.07 3.123 71.105 3.3 ;
      RECT 71.03 3.14 71.07 3.323 ;
      RECT 71.01 3.153 71.03 3.35 ;
      RECT 70.98 3.165 71.01 3.378 ;
      RECT 70.975 3.173 70.98 3.398 ;
      RECT 70.97 3.176 70.975 3.408 ;
      RECT 70.92 3.188 70.97 3.442 ;
      RECT 70.91 3.203 70.92 3.475 ;
      RECT 70.9 3.209 70.91 3.488 ;
      RECT 70.89 3.216 70.9 3.5 ;
      RECT 70.865 3.229 70.89 3.518 ;
      RECT 70.85 3.244 70.865 3.54 ;
      RECT 70.84 3.252 70.85 3.556 ;
      RECT 70.825 3.261 70.84 3.571 ;
      RECT 70.815 3.271 70.825 3.585 ;
      RECT 70.796 3.284 70.815 3.602 ;
      RECT 70.71 3.329 70.796 3.667 ;
      RECT 70.695 3.374 70.71 3.725 ;
      RECT 70.69 3.383 70.695 3.738 ;
      RECT 70.68 3.39 70.69 3.743 ;
      RECT 70.675 3.395 70.68 3.747 ;
      RECT 70.655 3.405 70.675 3.754 ;
      RECT 70.63 3.425 70.655 3.768 ;
      RECT 70.595 3.45 70.63 3.788 ;
      RECT 70.58 3.473 70.595 3.803 ;
      RECT 70.57 3.483 70.58 3.808 ;
      RECT 70.56 3.491 70.57 3.815 ;
      RECT 70.55 3.5 70.56 3.821 ;
      RECT 70.53 3.512 70.55 3.823 ;
      RECT 70.52 3.525 70.53 3.825 ;
      RECT 70.495 3.54 70.52 3.828 ;
      RECT 70.475 3.557 70.495 3.832 ;
      RECT 70.435 3.585 70.475 3.838 ;
      RECT 70.37 3.632 70.435 3.847 ;
      RECT 70.355 3.665 70.37 3.855 ;
      RECT 70.35 3.672 70.355 3.857 ;
      RECT 70.3 3.697 70.35 3.862 ;
      RECT 70.285 3.721 70.3 3.869 ;
      RECT 70.235 3.726 70.285 3.87 ;
      RECT 70.149 3.73 70.235 3.87 ;
      RECT 70.063 3.73 70.149 3.87 ;
      RECT 69.977 3.73 70.063 3.871 ;
      RECT 69.891 3.73 69.977 3.871 ;
      RECT 69.805 3.73 69.891 3.871 ;
      RECT 69.739 3.73 69.805 3.871 ;
      RECT 69.653 3.73 69.739 3.872 ;
      RECT 69.567 3.73 69.653 3.872 ;
      RECT 69.481 3.731 69.567 3.873 ;
      RECT 69.395 3.731 69.481 3.873 ;
      RECT 69.309 3.731 69.395 3.873 ;
      RECT 69.223 3.731 69.309 3.874 ;
      RECT 69.137 3.731 69.223 3.874 ;
      RECT 69.051 3.732 69.137 3.875 ;
      RECT 68.965 3.732 69.051 3.875 ;
      RECT 68.945 3.732 68.965 3.875 ;
      RECT 68.859 3.732 68.945 3.875 ;
      RECT 68.773 3.732 68.859 3.875 ;
      RECT 68.687 3.733 68.773 3.875 ;
      RECT 68.601 3.733 68.687 3.875 ;
      RECT 68.515 3.733 68.601 3.875 ;
      RECT 68.429 3.734 68.515 3.875 ;
      RECT 68.343 3.734 68.429 3.875 ;
      RECT 68.257 3.734 68.343 3.875 ;
      RECT 68.171 3.734 68.257 3.875 ;
      RECT 68.085 3.735 68.171 3.875 ;
      RECT 68.035 3.732 68.085 3.875 ;
      RECT 68.025 3.73 68.035 3.874 ;
      RECT 68.021 3.73 68.025 3.873 ;
      RECT 67.935 3.725 68.021 3.868 ;
      RECT 67.913 3.718 67.935 3.862 ;
      RECT 67.827 3.709 67.913 3.856 ;
      RECT 67.741 3.696 67.827 3.847 ;
      RECT 67.655 3.682 67.741 3.837 ;
      RECT 67.61 3.672 67.655 3.83 ;
      RECT 67.59 2.96 67.61 3.238 ;
      RECT 67.59 3.665 67.61 3.826 ;
      RECT 67.56 2.96 67.59 3.26 ;
      RECT 67.55 3.632 67.59 3.823 ;
      RECT 67.545 2.96 67.56 3.28 ;
      RECT 67.545 3.597 67.55 3.821 ;
      RECT 67.54 2.96 67.545 3.405 ;
      RECT 67.54 3.557 67.545 3.821 ;
      RECT 67.53 2.96 67.54 3.821 ;
      RECT 67.455 2.96 67.53 3.815 ;
      RECT 67.425 2.96 67.455 3.805 ;
      RECT 67.42 2.96 67.425 3.797 ;
      RECT 67.415 3.002 67.42 3.79 ;
      RECT 67.405 3.071 67.415 3.781 ;
      RECT 67.4 3.141 67.405 3.733 ;
      RECT 67.395 3.205 67.4 3.63 ;
      RECT 67.39 3.24 67.395 3.585 ;
      RECT 67.388 3.277 67.39 3.477 ;
      RECT 67.385 3.285 67.388 3.47 ;
      RECT 67.38 3.35 67.385 3.413 ;
      RECT 71.455 2.44 71.735 2.72 ;
      RECT 71.445 2.44 71.735 2.583 ;
      RECT 71.4 2.305 71.66 2.565 ;
      RECT 71.4 2.42 71.715 2.565 ;
      RECT 71.4 2.39 71.71 2.565 ;
      RECT 71.4 2.377 71.7 2.565 ;
      RECT 71.4 2.367 71.695 2.565 ;
      RECT 67.375 2.35 67.635 2.61 ;
      RECT 71.145 1.9 71.405 2.16 ;
      RECT 71.135 1.925 71.405 2.12 ;
      RECT 71.13 1.925 71.135 2.119 ;
      RECT 71.06 1.92 71.13 2.111 ;
      RECT 70.975 1.907 71.06 2.094 ;
      RECT 70.971 1.899 70.975 2.084 ;
      RECT 70.885 1.892 70.971 2.074 ;
      RECT 70.876 1.884 70.885 2.064 ;
      RECT 70.79 1.877 70.876 2.052 ;
      RECT 70.77 1.868 70.79 2.038 ;
      RECT 70.715 1.863 70.77 2.03 ;
      RECT 70.705 1.857 70.715 2.024 ;
      RECT 70.685 1.855 70.705 2.02 ;
      RECT 70.677 1.854 70.685 2.016 ;
      RECT 70.591 1.846 70.677 2.005 ;
      RECT 70.505 1.832 70.591 1.985 ;
      RECT 70.445 1.82 70.505 1.97 ;
      RECT 70.435 1.815 70.445 1.965 ;
      RECT 70.385 1.815 70.435 1.967 ;
      RECT 70.338 1.817 70.385 1.971 ;
      RECT 70.252 1.824 70.338 1.976 ;
      RECT 70.166 1.832 70.252 1.982 ;
      RECT 70.08 1.841 70.166 1.988 ;
      RECT 70.021 1.847 70.08 1.993 ;
      RECT 69.935 1.852 70.021 1.999 ;
      RECT 69.86 1.857 69.935 2.005 ;
      RECT 69.821 1.859 69.86 2.01 ;
      RECT 69.735 1.856 69.821 2.015 ;
      RECT 69.65 1.854 69.735 2.022 ;
      RECT 69.618 1.853 69.65 2.025 ;
      RECT 69.532 1.852 69.618 2.026 ;
      RECT 69.446 1.851 69.532 2.027 ;
      RECT 69.36 1.85 69.446 2.027 ;
      RECT 69.274 1.849 69.36 2.028 ;
      RECT 69.188 1.848 69.274 2.029 ;
      RECT 69.102 1.847 69.188 2.03 ;
      RECT 69.016 1.846 69.102 2.03 ;
      RECT 68.93 1.845 69.016 2.031 ;
      RECT 68.88 1.845 68.93 2.032 ;
      RECT 68.866 1.846 68.88 2.032 ;
      RECT 68.78 1.853 68.866 2.033 ;
      RECT 68.706 1.864 68.78 2.034 ;
      RECT 68.62 1.873 68.706 2.035 ;
      RECT 68.585 1.88 68.62 2.05 ;
      RECT 68.56 1.883 68.585 2.08 ;
      RECT 68.535 1.892 68.56 2.109 ;
      RECT 68.525 1.903 68.535 2.129 ;
      RECT 68.515 1.911 68.525 2.143 ;
      RECT 68.51 1.917 68.515 2.153 ;
      RECT 68.485 1.934 68.51 2.17 ;
      RECT 68.47 1.956 68.485 2.198 ;
      RECT 68.44 1.982 68.47 2.228 ;
      RECT 68.42 2.011 68.44 2.258 ;
      RECT 68.415 2.026 68.42 2.275 ;
      RECT 68.395 2.041 68.415 2.29 ;
      RECT 68.385 2.059 68.395 2.308 ;
      RECT 68.375 2.07 68.385 2.323 ;
      RECT 68.325 2.102 68.375 2.349 ;
      RECT 68.32 2.132 68.325 2.369 ;
      RECT 68.31 2.145 68.32 2.375 ;
      RECT 68.301 2.155 68.31 2.383 ;
      RECT 68.29 2.166 68.301 2.391 ;
      RECT 68.285 2.176 68.29 2.397 ;
      RECT 68.27 2.197 68.285 2.404 ;
      RECT 68.255 2.227 68.27 2.412 ;
      RECT 68.22 2.257 68.255 2.418 ;
      RECT 68.195 2.275 68.22 2.425 ;
      RECT 68.145 2.283 68.195 2.434 ;
      RECT 68.12 2.288 68.145 2.443 ;
      RECT 68.065 2.294 68.12 2.453 ;
      RECT 68.06 2.299 68.065 2.461 ;
      RECT 68.046 2.302 68.06 2.463 ;
      RECT 67.96 2.314 68.046 2.475 ;
      RECT 67.95 2.326 67.96 2.488 ;
      RECT 67.865 2.339 67.95 2.5 ;
      RECT 67.821 2.356 67.865 2.514 ;
      RECT 67.735 2.373 67.821 2.53 ;
      RECT 67.705 2.387 67.735 2.544 ;
      RECT 67.695 2.392 67.705 2.549 ;
      RECT 67.635 2.395 67.695 2.558 ;
      RECT 70.525 2.665 70.785 2.925 ;
      RECT 70.525 2.665 70.805 2.778 ;
      RECT 70.525 2.665 70.83 2.745 ;
      RECT 70.525 2.665 70.835 2.725 ;
      RECT 70.575 2.44 70.855 2.72 ;
      RECT 70.13 3.175 70.39 3.435 ;
      RECT 70.12 3.032 70.315 3.373 ;
      RECT 70.115 3.14 70.33 3.365 ;
      RECT 70.11 3.19 70.39 3.355 ;
      RECT 70.1 3.267 70.39 3.34 ;
      RECT 70.12 3.115 70.33 3.373 ;
      RECT 70.13 2.99 70.315 3.435 ;
      RECT 70.13 2.885 70.295 3.435 ;
      RECT 70.14 2.872 70.295 3.435 ;
      RECT 70.14 2.83 70.285 3.435 ;
      RECT 70.145 2.755 70.285 3.435 ;
      RECT 70.175 2.405 70.285 3.435 ;
      RECT 70.18 2.135 70.305 2.758 ;
      RECT 70.15 2.71 70.305 2.758 ;
      RECT 70.165 2.512 70.285 3.435 ;
      RECT 70.155 2.622 70.305 2.758 ;
      RECT 70.18 2.135 70.32 2.615 ;
      RECT 70.18 2.135 70.34 2.49 ;
      RECT 70.145 2.135 70.405 2.395 ;
      RECT 69.615 2.44 69.895 2.72 ;
      RECT 69.6 2.44 69.895 2.7 ;
      RECT 67.655 3.305 67.915 3.565 ;
      RECT 69.44 3.16 69.7 3.42 ;
      RECT 69.42 3.18 69.7 3.395 ;
      RECT 69.377 3.18 69.42 3.394 ;
      RECT 69.291 3.181 69.377 3.391 ;
      RECT 69.205 3.182 69.291 3.387 ;
      RECT 69.13 3.184 69.205 3.384 ;
      RECT 69.107 3.185 69.13 3.382 ;
      RECT 69.021 3.186 69.107 3.38 ;
      RECT 68.935 3.187 69.021 3.377 ;
      RECT 68.911 3.188 68.935 3.375 ;
      RECT 68.825 3.19 68.911 3.372 ;
      RECT 68.74 3.192 68.825 3.373 ;
      RECT 68.683 3.193 68.74 3.379 ;
      RECT 68.597 3.195 68.683 3.389 ;
      RECT 68.511 3.198 68.597 3.402 ;
      RECT 68.425 3.2 68.511 3.414 ;
      RECT 68.411 3.201 68.425 3.421 ;
      RECT 68.325 3.202 68.411 3.429 ;
      RECT 68.285 3.204 68.325 3.438 ;
      RECT 68.276 3.205 68.285 3.441 ;
      RECT 68.19 3.213 68.276 3.447 ;
      RECT 68.17 3.222 68.19 3.455 ;
      RECT 68.085 3.237 68.17 3.463 ;
      RECT 68.025 3.26 68.085 3.474 ;
      RECT 68.015 3.272 68.025 3.479 ;
      RECT 67.975 3.282 68.015 3.483 ;
      RECT 67.92 3.299 67.975 3.491 ;
      RECT 67.915 3.309 67.92 3.495 ;
      RECT 68.981 2.44 69.04 2.837 ;
      RECT 68.895 2.44 69.1 2.828 ;
      RECT 68.89 2.47 69.1 2.823 ;
      RECT 68.856 2.47 69.1 2.821 ;
      RECT 68.77 2.47 69.1 2.815 ;
      RECT 68.725 2.47 69.12 2.793 ;
      RECT 68.725 2.47 69.14 2.748 ;
      RECT 68.685 2.47 69.14 2.738 ;
      RECT 68.895 2.44 69.175 2.72 ;
      RECT 68.63 2.44 68.89 2.7 ;
      RECT 66.455 3 66.735 3.28 ;
      RECT 66.425 2.962 66.68 3.265 ;
      RECT 66.42 2.963 66.68 3.263 ;
      RECT 66.415 2.964 66.68 3.257 ;
      RECT 66.41 2.967 66.68 3.25 ;
      RECT 66.405 3 66.735 3.243 ;
      RECT 66.375 2.97 66.68 3.23 ;
      RECT 66.375 2.997 66.7 3.23 ;
      RECT 66.375 2.987 66.695 3.23 ;
      RECT 66.375 2.972 66.69 3.23 ;
      RECT 66.455 2.959 66.67 3.28 ;
      RECT 66.541 2.957 66.67 3.28 ;
      RECT 66.627 2.955 66.655 3.28 ;
      RECT 62.26 6.22 62.58 6.545 ;
      RECT 62.29 5.695 62.46 6.545 ;
      RECT 62.29 5.695 62.465 6.045 ;
      RECT 62.29 5.695 63.265 5.87 ;
      RECT 63.09 1.965 63.265 5.87 ;
      RECT 63.035 1.965 63.385 2.315 ;
      RECT 63.06 6.655 63.385 6.98 ;
      RECT 61.945 6.745 63.385 6.915 ;
      RECT 61.945 2.395 62.105 6.915 ;
      RECT 62.26 2.365 62.58 2.685 ;
      RECT 61.945 2.395 62.58 2.565 ;
      RECT 52.03 1.92 52.29 2.18 ;
      RECT 52.085 1.88 52.39 2.16 ;
      RECT 52.085 1.42 52.26 2.18 ;
      RECT 60.6 1.34 60.95 1.69 ;
      RECT 52.085 1.42 60.95 1.595 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 60.36 2.235 60.53 3.22 ;
      RECT 56.38 2.455 56.615 2.715 ;
      RECT 59.525 2.235 59.69 2.495 ;
      RECT 59.43 2.225 59.445 2.495 ;
      RECT 59.525 2.235 60.53 2.415 ;
      RECT 58.03 1.795 58.07 1.935 ;
      RECT 59.445 2.23 59.525 2.495 ;
      RECT 59.39 2.225 59.43 2.461 ;
      RECT 59.376 2.225 59.39 2.461 ;
      RECT 59.29 2.23 59.376 2.463 ;
      RECT 59.245 2.237 59.29 2.465 ;
      RECT 59.215 2.237 59.245 2.467 ;
      RECT 59.19 2.232 59.215 2.469 ;
      RECT 59.16 2.228 59.19 2.478 ;
      RECT 59.15 2.225 59.16 2.49 ;
      RECT 59.145 2.225 59.15 2.498 ;
      RECT 59.14 2.225 59.145 2.503 ;
      RECT 59.13 2.224 59.14 2.513 ;
      RECT 59.125 2.223 59.13 2.523 ;
      RECT 59.11 2.222 59.125 2.528 ;
      RECT 59.082 2.219 59.11 2.555 ;
      RECT 58.996 2.211 59.082 2.555 ;
      RECT 58.91 2.2 58.996 2.555 ;
      RECT 58.87 2.185 58.91 2.555 ;
      RECT 58.83 2.159 58.87 2.555 ;
      RECT 58.825 2.141 58.83 2.367 ;
      RECT 58.815 2.137 58.825 2.357 ;
      RECT 58.8 2.127 58.815 2.344 ;
      RECT 58.78 2.111 58.8 2.329 ;
      RECT 58.765 2.096 58.78 2.314 ;
      RECT 58.755 2.085 58.765 2.304 ;
      RECT 58.73 2.069 58.755 2.293 ;
      RECT 58.725 2.056 58.73 2.283 ;
      RECT 58.72 2.052 58.725 2.278 ;
      RECT 58.665 2.038 58.72 2.256 ;
      RECT 58.626 2.019 58.665 2.22 ;
      RECT 58.54 1.993 58.626 2.173 ;
      RECT 58.536 1.975 58.54 2.139 ;
      RECT 58.45 1.956 58.536 2.117 ;
      RECT 58.445 1.938 58.45 2.095 ;
      RECT 58.44 1.936 58.445 2.093 ;
      RECT 58.43 1.935 58.44 2.088 ;
      RECT 58.37 1.922 58.43 2.074 ;
      RECT 58.325 1.9 58.37 2.053 ;
      RECT 58.265 1.877 58.325 2.032 ;
      RECT 58.201 1.852 58.265 2.007 ;
      RECT 58.115 1.822 58.201 1.976 ;
      RECT 58.1 1.802 58.115 1.955 ;
      RECT 58.07 1.797 58.1 1.946 ;
      RECT 58.017 1.795 58.03 1.935 ;
      RECT 57.931 1.795 58.017 1.937 ;
      RECT 57.845 1.795 57.931 1.939 ;
      RECT 57.825 1.795 57.845 1.943 ;
      RECT 57.78 1.797 57.825 1.954 ;
      RECT 57.74 1.807 57.78 1.97 ;
      RECT 57.736 1.816 57.74 1.978 ;
      RECT 57.65 1.836 57.736 1.994 ;
      RECT 57.64 1.855 57.65 2.012 ;
      RECT 57.635 1.857 57.64 2.015 ;
      RECT 57.625 1.861 57.635 2.018 ;
      RECT 57.605 1.866 57.625 2.028 ;
      RECT 57.575 1.876 57.605 2.048 ;
      RECT 57.57 1.883 57.575 2.062 ;
      RECT 57.56 1.887 57.57 2.069 ;
      RECT 57.545 1.895 57.56 2.08 ;
      RECT 57.535 1.905 57.545 2.091 ;
      RECT 57.525 1.912 57.535 2.099 ;
      RECT 57.5 1.925 57.525 2.114 ;
      RECT 57.436 1.961 57.5 2.153 ;
      RECT 57.35 2.024 57.436 2.217 ;
      RECT 57.315 2.075 57.35 2.27 ;
      RECT 57.31 2.092 57.315 2.287 ;
      RECT 57.295 2.101 57.31 2.294 ;
      RECT 57.275 2.116 57.295 2.308 ;
      RECT 57.27 2.127 57.275 2.318 ;
      RECT 57.25 2.14 57.27 2.328 ;
      RECT 57.245 2.15 57.25 2.338 ;
      RECT 57.23 2.155 57.245 2.347 ;
      RECT 57.22 2.165 57.23 2.358 ;
      RECT 57.19 2.182 57.22 2.375 ;
      RECT 57.18 2.2 57.19 2.393 ;
      RECT 57.165 2.211 57.18 2.404 ;
      RECT 57.125 2.235 57.165 2.42 ;
      RECT 57.09 2.269 57.125 2.437 ;
      RECT 57.06 2.292 57.09 2.449 ;
      RECT 57.045 2.302 57.06 2.458 ;
      RECT 57.005 2.312 57.045 2.469 ;
      RECT 56.985 2.323 57.005 2.481 ;
      RECT 56.98 2.327 56.985 2.488 ;
      RECT 56.965 2.331 56.98 2.493 ;
      RECT 56.955 2.336 56.965 2.498 ;
      RECT 56.95 2.339 56.955 2.501 ;
      RECT 56.92 2.345 56.95 2.508 ;
      RECT 56.885 2.355 56.92 2.522 ;
      RECT 56.825 2.37 56.885 2.542 ;
      RECT 56.77 2.39 56.825 2.566 ;
      RECT 56.741 2.405 56.77 2.584 ;
      RECT 56.655 2.425 56.741 2.609 ;
      RECT 56.65 2.44 56.655 2.629 ;
      RECT 56.64 2.443 56.65 2.63 ;
      RECT 56.615 2.45 56.64 2.715 ;
      RECT 59.31 2.943 59.59 3.28 ;
      RECT 59.31 2.953 59.595 3.238 ;
      RECT 59.31 2.962 59.6 3.135 ;
      RECT 59.31 2.977 59.605 3.003 ;
      RECT 59.31 2.805 59.57 3.28 ;
      RECT 49.61 6.655 49.96 7.005 ;
      RECT 58.435 6.61 58.785 6.96 ;
      RECT 49.61 6.685 58.785 6.885 ;
      RECT 57.03 3.685 57.04 3.875 ;
      RECT 55.29 3.56 55.57 3.84 ;
      RECT 58.335 2.5 58.34 2.985 ;
      RECT 58.23 2.5 58.29 2.76 ;
      RECT 58.555 3.47 58.56 3.545 ;
      RECT 58.545 3.337 58.555 3.58 ;
      RECT 58.535 3.172 58.545 3.601 ;
      RECT 58.53 3.042 58.535 3.617 ;
      RECT 58.52 2.932 58.53 3.633 ;
      RECT 58.515 2.831 58.52 3.65 ;
      RECT 58.51 2.813 58.515 3.66 ;
      RECT 58.505 2.795 58.51 3.67 ;
      RECT 58.495 2.77 58.505 3.685 ;
      RECT 58.49 2.75 58.495 3.7 ;
      RECT 58.47 2.5 58.49 3.725 ;
      RECT 58.455 2.5 58.47 3.758 ;
      RECT 58.425 2.5 58.455 3.78 ;
      RECT 58.405 2.5 58.425 3.794 ;
      RECT 58.385 2.5 58.405 3.31 ;
      RECT 58.4 3.377 58.405 3.799 ;
      RECT 58.395 3.407 58.4 3.801 ;
      RECT 58.39 3.42 58.395 3.804 ;
      RECT 58.385 3.43 58.39 3.808 ;
      RECT 58.38 2.5 58.385 3.228 ;
      RECT 58.38 3.44 58.385 3.81 ;
      RECT 58.375 2.5 58.38 3.205 ;
      RECT 58.365 3.462 58.38 3.81 ;
      RECT 58.36 2.5 58.375 3.15 ;
      RECT 58.355 3.487 58.365 3.81 ;
      RECT 58.355 2.5 58.36 3.095 ;
      RECT 58.345 2.5 58.355 3.043 ;
      RECT 58.35 3.5 58.355 3.811 ;
      RECT 58.345 3.512 58.35 3.812 ;
      RECT 58.34 2.5 58.345 3.003 ;
      RECT 58.34 3.525 58.345 3.813 ;
      RECT 58.325 3.54 58.34 3.814 ;
      RECT 58.33 2.5 58.335 2.965 ;
      RECT 58.325 2.5 58.33 2.93 ;
      RECT 58.32 2.5 58.325 2.905 ;
      RECT 58.315 3.567 58.325 3.816 ;
      RECT 58.31 2.5 58.32 2.863 ;
      RECT 58.31 3.585 58.315 3.817 ;
      RECT 58.305 2.5 58.31 2.823 ;
      RECT 58.305 3.592 58.31 3.818 ;
      RECT 58.3 2.5 58.305 2.795 ;
      RECT 58.295 3.61 58.305 3.819 ;
      RECT 58.29 2.5 58.3 2.775 ;
      RECT 58.285 3.63 58.295 3.821 ;
      RECT 58.275 3.647 58.285 3.822 ;
      RECT 58.24 3.67 58.275 3.825 ;
      RECT 58.185 3.688 58.24 3.831 ;
      RECT 58.099 3.696 58.185 3.84 ;
      RECT 58.013 3.707 58.099 3.851 ;
      RECT 57.927 3.717 58.013 3.862 ;
      RECT 57.841 3.727 57.927 3.874 ;
      RECT 57.755 3.737 57.841 3.885 ;
      RECT 57.735 3.743 57.755 3.891 ;
      RECT 57.655 3.745 57.735 3.895 ;
      RECT 57.65 3.744 57.655 3.9 ;
      RECT 57.642 3.743 57.65 3.9 ;
      RECT 57.556 3.739 57.642 3.898 ;
      RECT 57.47 3.731 57.556 3.895 ;
      RECT 57.384 3.722 57.47 3.891 ;
      RECT 57.298 3.714 57.384 3.888 ;
      RECT 57.212 3.706 57.298 3.884 ;
      RECT 57.126 3.697 57.212 3.881 ;
      RECT 57.04 3.689 57.126 3.877 ;
      RECT 56.985 3.682 57.03 3.875 ;
      RECT 56.9 3.675 56.985 3.873 ;
      RECT 56.826 3.667 56.9 3.869 ;
      RECT 56.74 3.659 56.826 3.866 ;
      RECT 56.737 3.655 56.74 3.864 ;
      RECT 56.651 3.651 56.737 3.863 ;
      RECT 56.565 3.643 56.651 3.86 ;
      RECT 56.48 3.638 56.565 3.857 ;
      RECT 56.394 3.635 56.48 3.854 ;
      RECT 56.308 3.633 56.394 3.851 ;
      RECT 56.222 3.63 56.308 3.848 ;
      RECT 56.136 3.627 56.222 3.845 ;
      RECT 56.05 3.624 56.136 3.842 ;
      RECT 55.974 3.622 56.05 3.839 ;
      RECT 55.888 3.619 55.974 3.836 ;
      RECT 55.802 3.616 55.888 3.834 ;
      RECT 55.716 3.614 55.802 3.831 ;
      RECT 55.63 3.611 55.716 3.828 ;
      RECT 55.57 3.602 55.63 3.826 ;
      RECT 58.08 3.22 58.155 3.48 ;
      RECT 58.06 3.2 58.065 3.48 ;
      RECT 57.38 2.985 57.485 3.28 ;
      RECT 51.825 2.96 51.895 3.22 ;
      RECT 57.72 2.835 57.725 3.206 ;
      RECT 57.71 2.89 57.715 3.206 ;
      RECT 58.015 2.06 58.075 2.32 ;
      RECT 58.07 3.215 58.08 3.48 ;
      RECT 58.065 3.205 58.07 3.48 ;
      RECT 57.985 3.152 58.06 3.48 ;
      RECT 58.01 2.06 58.015 2.34 ;
      RECT 58 2.06 58.01 2.36 ;
      RECT 57.985 2.06 58 2.39 ;
      RECT 57.97 2.06 57.985 2.433 ;
      RECT 57.965 3.095 57.985 3.48 ;
      RECT 57.955 2.06 57.97 2.47 ;
      RECT 57.95 3.075 57.965 3.48 ;
      RECT 57.95 2.06 57.955 2.493 ;
      RECT 57.94 2.06 57.95 2.518 ;
      RECT 57.91 3.042 57.95 3.48 ;
      RECT 57.915 2.06 57.94 2.568 ;
      RECT 57.91 2.06 57.915 2.623 ;
      RECT 57.905 2.06 57.91 2.665 ;
      RECT 57.895 3.005 57.91 3.48 ;
      RECT 57.9 2.06 57.905 2.708 ;
      RECT 57.895 2.06 57.9 2.773 ;
      RECT 57.89 2.06 57.895 2.795 ;
      RECT 57.89 2.993 57.895 3.345 ;
      RECT 57.885 2.06 57.89 2.863 ;
      RECT 57.885 2.985 57.89 3.328 ;
      RECT 57.88 2.06 57.885 2.908 ;
      RECT 57.875 2.967 57.885 3.305 ;
      RECT 57.875 2.06 57.88 2.945 ;
      RECT 57.865 2.06 57.875 3.285 ;
      RECT 57.86 2.06 57.865 3.268 ;
      RECT 57.855 2.06 57.86 3.253 ;
      RECT 57.85 2.06 57.855 3.238 ;
      RECT 57.83 2.06 57.85 3.228 ;
      RECT 57.825 2.06 57.83 3.218 ;
      RECT 57.815 2.06 57.825 3.214 ;
      RECT 57.81 2.337 57.815 3.213 ;
      RECT 57.805 2.36 57.81 3.212 ;
      RECT 57.8 2.39 57.805 3.211 ;
      RECT 57.795 2.417 57.8 3.21 ;
      RECT 57.79 2.445 57.795 3.21 ;
      RECT 57.785 2.472 57.79 3.21 ;
      RECT 57.78 2.492 57.785 3.21 ;
      RECT 57.775 2.52 57.78 3.21 ;
      RECT 57.765 2.562 57.775 3.21 ;
      RECT 57.755 2.607 57.765 3.209 ;
      RECT 57.75 2.66 57.755 3.208 ;
      RECT 57.745 2.692 57.75 3.207 ;
      RECT 57.74 2.712 57.745 3.206 ;
      RECT 57.735 2.75 57.74 3.206 ;
      RECT 57.73 2.772 57.735 3.206 ;
      RECT 57.725 2.797 57.73 3.206 ;
      RECT 57.715 2.862 57.72 3.206 ;
      RECT 57.7 2.922 57.71 3.206 ;
      RECT 57.685 2.932 57.7 3.206 ;
      RECT 57.665 2.942 57.685 3.206 ;
      RECT 57.635 2.947 57.665 3.203 ;
      RECT 57.575 2.957 57.635 3.2 ;
      RECT 57.555 2.966 57.575 3.205 ;
      RECT 57.53 2.972 57.555 3.218 ;
      RECT 57.51 2.977 57.53 3.233 ;
      RECT 57.485 2.982 57.51 3.28 ;
      RECT 57.356 2.984 57.38 3.28 ;
      RECT 57.27 2.979 57.356 3.28 ;
      RECT 57.23 2.976 57.27 3.28 ;
      RECT 57.18 2.978 57.23 3.26 ;
      RECT 57.15 2.982 57.18 3.26 ;
      RECT 57.071 2.992 57.15 3.26 ;
      RECT 56.985 3.007 57.071 3.261 ;
      RECT 56.935 3.017 56.985 3.262 ;
      RECT 56.927 3.02 56.935 3.262 ;
      RECT 56.841 3.022 56.927 3.263 ;
      RECT 56.755 3.026 56.841 3.263 ;
      RECT 56.669 3.03 56.755 3.264 ;
      RECT 56.583 3.033 56.669 3.265 ;
      RECT 56.497 3.037 56.583 3.265 ;
      RECT 56.411 3.041 56.497 3.266 ;
      RECT 56.325 3.044 56.411 3.267 ;
      RECT 56.239 3.048 56.325 3.267 ;
      RECT 56.153 3.052 56.239 3.268 ;
      RECT 56.067 3.056 56.153 3.269 ;
      RECT 55.981 3.059 56.067 3.269 ;
      RECT 55.895 3.063 55.981 3.27 ;
      RECT 55.865 3.065 55.895 3.27 ;
      RECT 55.779 3.068 55.865 3.271 ;
      RECT 55.693 3.072 55.779 3.272 ;
      RECT 55.607 3.076 55.693 3.273 ;
      RECT 55.521 3.079 55.607 3.273 ;
      RECT 55.435 3.083 55.521 3.274 ;
      RECT 55.4 3.088 55.435 3.275 ;
      RECT 55.345 3.098 55.4 3.282 ;
      RECT 55.32 3.11 55.345 3.292 ;
      RECT 55.285 3.123 55.32 3.3 ;
      RECT 55.245 3.14 55.285 3.323 ;
      RECT 55.225 3.153 55.245 3.35 ;
      RECT 55.195 3.165 55.225 3.378 ;
      RECT 55.19 3.173 55.195 3.398 ;
      RECT 55.185 3.176 55.19 3.408 ;
      RECT 55.135 3.188 55.185 3.442 ;
      RECT 55.125 3.203 55.135 3.475 ;
      RECT 55.115 3.209 55.125 3.488 ;
      RECT 55.105 3.216 55.115 3.5 ;
      RECT 55.08 3.229 55.105 3.518 ;
      RECT 55.065 3.244 55.08 3.54 ;
      RECT 55.055 3.252 55.065 3.556 ;
      RECT 55.04 3.261 55.055 3.571 ;
      RECT 55.03 3.271 55.04 3.585 ;
      RECT 55.011 3.284 55.03 3.602 ;
      RECT 54.925 3.329 55.011 3.667 ;
      RECT 54.91 3.374 54.925 3.725 ;
      RECT 54.905 3.383 54.91 3.738 ;
      RECT 54.895 3.39 54.905 3.743 ;
      RECT 54.89 3.395 54.895 3.747 ;
      RECT 54.87 3.405 54.89 3.754 ;
      RECT 54.845 3.425 54.87 3.768 ;
      RECT 54.81 3.45 54.845 3.788 ;
      RECT 54.795 3.473 54.81 3.803 ;
      RECT 54.785 3.483 54.795 3.808 ;
      RECT 54.775 3.491 54.785 3.815 ;
      RECT 54.765 3.5 54.775 3.821 ;
      RECT 54.745 3.512 54.765 3.823 ;
      RECT 54.735 3.525 54.745 3.825 ;
      RECT 54.71 3.54 54.735 3.828 ;
      RECT 54.69 3.557 54.71 3.832 ;
      RECT 54.65 3.585 54.69 3.838 ;
      RECT 54.585 3.632 54.65 3.847 ;
      RECT 54.57 3.665 54.585 3.855 ;
      RECT 54.565 3.672 54.57 3.857 ;
      RECT 54.515 3.697 54.565 3.862 ;
      RECT 54.5 3.721 54.515 3.869 ;
      RECT 54.45 3.726 54.5 3.87 ;
      RECT 54.364 3.73 54.45 3.87 ;
      RECT 54.278 3.73 54.364 3.87 ;
      RECT 54.192 3.73 54.278 3.871 ;
      RECT 54.106 3.73 54.192 3.871 ;
      RECT 54.02 3.73 54.106 3.871 ;
      RECT 53.954 3.73 54.02 3.871 ;
      RECT 53.868 3.73 53.954 3.872 ;
      RECT 53.782 3.73 53.868 3.872 ;
      RECT 53.696 3.731 53.782 3.873 ;
      RECT 53.61 3.731 53.696 3.873 ;
      RECT 53.524 3.731 53.61 3.873 ;
      RECT 53.438 3.731 53.524 3.874 ;
      RECT 53.352 3.731 53.438 3.874 ;
      RECT 53.266 3.732 53.352 3.875 ;
      RECT 53.18 3.732 53.266 3.875 ;
      RECT 53.16 3.732 53.18 3.875 ;
      RECT 53.074 3.732 53.16 3.875 ;
      RECT 52.988 3.732 53.074 3.875 ;
      RECT 52.902 3.733 52.988 3.875 ;
      RECT 52.816 3.733 52.902 3.875 ;
      RECT 52.73 3.733 52.816 3.875 ;
      RECT 52.644 3.734 52.73 3.875 ;
      RECT 52.558 3.734 52.644 3.875 ;
      RECT 52.472 3.734 52.558 3.875 ;
      RECT 52.386 3.734 52.472 3.875 ;
      RECT 52.3 3.735 52.386 3.875 ;
      RECT 52.25 3.732 52.3 3.875 ;
      RECT 52.24 3.73 52.25 3.874 ;
      RECT 52.236 3.73 52.24 3.873 ;
      RECT 52.15 3.725 52.236 3.868 ;
      RECT 52.128 3.718 52.15 3.862 ;
      RECT 52.042 3.709 52.128 3.856 ;
      RECT 51.956 3.696 52.042 3.847 ;
      RECT 51.87 3.682 51.956 3.837 ;
      RECT 51.825 3.672 51.87 3.83 ;
      RECT 51.805 2.96 51.825 3.238 ;
      RECT 51.805 3.665 51.825 3.826 ;
      RECT 51.775 2.96 51.805 3.26 ;
      RECT 51.765 3.632 51.805 3.823 ;
      RECT 51.76 2.96 51.775 3.28 ;
      RECT 51.76 3.597 51.765 3.821 ;
      RECT 51.755 2.96 51.76 3.405 ;
      RECT 51.755 3.557 51.76 3.821 ;
      RECT 51.745 2.96 51.755 3.821 ;
      RECT 51.67 2.96 51.745 3.815 ;
      RECT 51.64 2.96 51.67 3.805 ;
      RECT 51.635 2.96 51.64 3.797 ;
      RECT 51.63 3.002 51.635 3.79 ;
      RECT 51.62 3.071 51.63 3.781 ;
      RECT 51.615 3.141 51.62 3.733 ;
      RECT 51.61 3.205 51.615 3.63 ;
      RECT 51.605 3.24 51.61 3.585 ;
      RECT 51.603 3.277 51.605 3.477 ;
      RECT 51.6 3.285 51.603 3.47 ;
      RECT 51.595 3.35 51.6 3.413 ;
      RECT 55.67 2.44 55.95 2.72 ;
      RECT 55.66 2.44 55.95 2.583 ;
      RECT 55.615 2.305 55.875 2.565 ;
      RECT 55.615 2.42 55.93 2.565 ;
      RECT 55.615 2.39 55.925 2.565 ;
      RECT 55.615 2.377 55.915 2.565 ;
      RECT 55.615 2.367 55.91 2.565 ;
      RECT 51.59 2.35 51.85 2.61 ;
      RECT 55.36 1.9 55.62 2.16 ;
      RECT 55.35 1.925 55.62 2.12 ;
      RECT 55.345 1.925 55.35 2.119 ;
      RECT 55.275 1.92 55.345 2.111 ;
      RECT 55.19 1.907 55.275 2.094 ;
      RECT 55.186 1.899 55.19 2.084 ;
      RECT 55.1 1.892 55.186 2.074 ;
      RECT 55.091 1.884 55.1 2.064 ;
      RECT 55.005 1.877 55.091 2.052 ;
      RECT 54.985 1.868 55.005 2.038 ;
      RECT 54.93 1.863 54.985 2.03 ;
      RECT 54.92 1.857 54.93 2.024 ;
      RECT 54.9 1.855 54.92 2.02 ;
      RECT 54.892 1.854 54.9 2.016 ;
      RECT 54.806 1.846 54.892 2.005 ;
      RECT 54.72 1.832 54.806 1.985 ;
      RECT 54.66 1.82 54.72 1.97 ;
      RECT 54.65 1.815 54.66 1.965 ;
      RECT 54.6 1.815 54.65 1.967 ;
      RECT 54.553 1.817 54.6 1.971 ;
      RECT 54.467 1.824 54.553 1.976 ;
      RECT 54.381 1.832 54.467 1.982 ;
      RECT 54.295 1.841 54.381 1.988 ;
      RECT 54.236 1.847 54.295 1.993 ;
      RECT 54.15 1.852 54.236 1.999 ;
      RECT 54.075 1.857 54.15 2.005 ;
      RECT 54.036 1.859 54.075 2.01 ;
      RECT 53.95 1.856 54.036 2.015 ;
      RECT 53.865 1.854 53.95 2.022 ;
      RECT 53.833 1.853 53.865 2.025 ;
      RECT 53.747 1.852 53.833 2.026 ;
      RECT 53.661 1.851 53.747 2.027 ;
      RECT 53.575 1.85 53.661 2.027 ;
      RECT 53.489 1.849 53.575 2.028 ;
      RECT 53.403 1.848 53.489 2.029 ;
      RECT 53.317 1.847 53.403 2.03 ;
      RECT 53.231 1.846 53.317 2.03 ;
      RECT 53.145 1.845 53.231 2.031 ;
      RECT 53.095 1.845 53.145 2.032 ;
      RECT 53.081 1.846 53.095 2.032 ;
      RECT 52.995 1.853 53.081 2.033 ;
      RECT 52.921 1.864 52.995 2.034 ;
      RECT 52.835 1.873 52.921 2.035 ;
      RECT 52.8 1.88 52.835 2.05 ;
      RECT 52.775 1.883 52.8 2.08 ;
      RECT 52.75 1.892 52.775 2.109 ;
      RECT 52.74 1.903 52.75 2.129 ;
      RECT 52.73 1.911 52.74 2.143 ;
      RECT 52.725 1.917 52.73 2.153 ;
      RECT 52.7 1.934 52.725 2.17 ;
      RECT 52.685 1.956 52.7 2.198 ;
      RECT 52.655 1.982 52.685 2.228 ;
      RECT 52.635 2.011 52.655 2.258 ;
      RECT 52.63 2.026 52.635 2.275 ;
      RECT 52.61 2.041 52.63 2.29 ;
      RECT 52.6 2.059 52.61 2.308 ;
      RECT 52.59 2.07 52.6 2.323 ;
      RECT 52.54 2.102 52.59 2.349 ;
      RECT 52.535 2.132 52.54 2.369 ;
      RECT 52.525 2.145 52.535 2.375 ;
      RECT 52.516 2.155 52.525 2.383 ;
      RECT 52.505 2.166 52.516 2.391 ;
      RECT 52.5 2.176 52.505 2.397 ;
      RECT 52.485 2.197 52.5 2.404 ;
      RECT 52.47 2.227 52.485 2.412 ;
      RECT 52.435 2.257 52.47 2.418 ;
      RECT 52.41 2.275 52.435 2.425 ;
      RECT 52.36 2.283 52.41 2.434 ;
      RECT 52.335 2.288 52.36 2.443 ;
      RECT 52.28 2.294 52.335 2.453 ;
      RECT 52.275 2.299 52.28 2.461 ;
      RECT 52.261 2.302 52.275 2.463 ;
      RECT 52.175 2.314 52.261 2.475 ;
      RECT 52.165 2.326 52.175 2.488 ;
      RECT 52.08 2.339 52.165 2.5 ;
      RECT 52.036 2.356 52.08 2.514 ;
      RECT 51.95 2.373 52.036 2.53 ;
      RECT 51.92 2.387 51.95 2.544 ;
      RECT 51.91 2.392 51.92 2.549 ;
      RECT 51.85 2.395 51.91 2.558 ;
      RECT 54.74 2.665 55 2.925 ;
      RECT 54.74 2.665 55.02 2.778 ;
      RECT 54.74 2.665 55.045 2.745 ;
      RECT 54.74 2.665 55.05 2.725 ;
      RECT 54.79 2.44 55.07 2.72 ;
      RECT 54.345 3.175 54.605 3.435 ;
      RECT 54.335 3.032 54.53 3.373 ;
      RECT 54.33 3.14 54.545 3.365 ;
      RECT 54.325 3.19 54.605 3.355 ;
      RECT 54.315 3.267 54.605 3.34 ;
      RECT 54.335 3.115 54.545 3.373 ;
      RECT 54.345 2.99 54.53 3.435 ;
      RECT 54.345 2.885 54.51 3.435 ;
      RECT 54.355 2.872 54.51 3.435 ;
      RECT 54.355 2.83 54.5 3.435 ;
      RECT 54.36 2.755 54.5 3.435 ;
      RECT 54.39 2.405 54.5 3.435 ;
      RECT 54.395 2.135 54.52 2.758 ;
      RECT 54.365 2.71 54.52 2.758 ;
      RECT 54.38 2.512 54.5 3.435 ;
      RECT 54.37 2.622 54.52 2.758 ;
      RECT 54.395 2.135 54.535 2.615 ;
      RECT 54.395 2.135 54.555 2.49 ;
      RECT 54.36 2.135 54.62 2.395 ;
      RECT 53.83 2.44 54.11 2.72 ;
      RECT 53.815 2.44 54.11 2.7 ;
      RECT 51.87 3.305 52.13 3.565 ;
      RECT 53.655 3.16 53.915 3.42 ;
      RECT 53.635 3.18 53.915 3.395 ;
      RECT 53.592 3.18 53.635 3.394 ;
      RECT 53.506 3.181 53.592 3.391 ;
      RECT 53.42 3.182 53.506 3.387 ;
      RECT 53.345 3.184 53.42 3.384 ;
      RECT 53.322 3.185 53.345 3.382 ;
      RECT 53.236 3.186 53.322 3.38 ;
      RECT 53.15 3.187 53.236 3.377 ;
      RECT 53.126 3.188 53.15 3.375 ;
      RECT 53.04 3.19 53.126 3.372 ;
      RECT 52.955 3.192 53.04 3.373 ;
      RECT 52.898 3.193 52.955 3.379 ;
      RECT 52.812 3.195 52.898 3.389 ;
      RECT 52.726 3.198 52.812 3.402 ;
      RECT 52.64 3.2 52.726 3.414 ;
      RECT 52.626 3.201 52.64 3.421 ;
      RECT 52.54 3.202 52.626 3.429 ;
      RECT 52.5 3.204 52.54 3.438 ;
      RECT 52.491 3.205 52.5 3.441 ;
      RECT 52.405 3.213 52.491 3.447 ;
      RECT 52.385 3.222 52.405 3.455 ;
      RECT 52.3 3.237 52.385 3.463 ;
      RECT 52.24 3.26 52.3 3.474 ;
      RECT 52.23 3.272 52.24 3.479 ;
      RECT 52.19 3.282 52.23 3.483 ;
      RECT 52.135 3.299 52.19 3.491 ;
      RECT 52.13 3.309 52.135 3.495 ;
      RECT 53.196 2.44 53.255 2.837 ;
      RECT 53.11 2.44 53.315 2.828 ;
      RECT 53.105 2.47 53.315 2.823 ;
      RECT 53.071 2.47 53.315 2.821 ;
      RECT 52.985 2.47 53.315 2.815 ;
      RECT 52.94 2.47 53.335 2.793 ;
      RECT 52.94 2.47 53.355 2.748 ;
      RECT 52.9 2.47 53.355 2.738 ;
      RECT 53.11 2.44 53.39 2.72 ;
      RECT 52.845 2.44 53.105 2.7 ;
      RECT 50.67 3 50.95 3.28 ;
      RECT 50.64 2.962 50.895 3.265 ;
      RECT 50.635 2.963 50.895 3.263 ;
      RECT 50.63 2.964 50.895 3.257 ;
      RECT 50.625 2.967 50.895 3.25 ;
      RECT 50.62 3 50.95 3.243 ;
      RECT 50.59 2.97 50.895 3.23 ;
      RECT 50.59 2.997 50.915 3.23 ;
      RECT 50.59 2.987 50.91 3.23 ;
      RECT 50.59 2.972 50.905 3.23 ;
      RECT 50.67 2.959 50.885 3.28 ;
      RECT 50.756 2.957 50.885 3.28 ;
      RECT 50.842 2.955 50.87 3.28 ;
      RECT 46.475 6.22 46.795 6.545 ;
      RECT 46.505 5.695 46.675 6.545 ;
      RECT 46.505 5.695 46.68 6.045 ;
      RECT 46.505 5.695 47.48 5.87 ;
      RECT 47.305 1.965 47.48 5.87 ;
      RECT 47.25 1.965 47.6 2.315 ;
      RECT 47.275 6.655 47.6 6.98 ;
      RECT 46.16 6.745 47.6 6.915 ;
      RECT 46.16 2.395 46.32 6.915 ;
      RECT 46.475 2.365 46.795 2.685 ;
      RECT 46.16 2.395 46.795 2.565 ;
      RECT 36.245 1.92 36.505 2.18 ;
      RECT 36.3 1.88 36.605 2.16 ;
      RECT 36.3 1.42 36.475 2.18 ;
      RECT 44.815 1.34 45.165 1.69 ;
      RECT 36.3 1.42 45.165 1.595 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 44.575 2.235 44.745 3.22 ;
      RECT 40.595 2.455 40.83 2.715 ;
      RECT 43.74 2.235 43.905 2.495 ;
      RECT 43.645 2.225 43.66 2.495 ;
      RECT 43.74 2.235 44.745 2.415 ;
      RECT 42.245 1.795 42.285 1.935 ;
      RECT 43.66 2.23 43.74 2.495 ;
      RECT 43.605 2.225 43.645 2.461 ;
      RECT 43.591 2.225 43.605 2.461 ;
      RECT 43.505 2.23 43.591 2.463 ;
      RECT 43.46 2.237 43.505 2.465 ;
      RECT 43.43 2.237 43.46 2.467 ;
      RECT 43.405 2.232 43.43 2.469 ;
      RECT 43.375 2.228 43.405 2.478 ;
      RECT 43.365 2.225 43.375 2.49 ;
      RECT 43.36 2.225 43.365 2.498 ;
      RECT 43.355 2.225 43.36 2.503 ;
      RECT 43.345 2.224 43.355 2.513 ;
      RECT 43.34 2.223 43.345 2.523 ;
      RECT 43.325 2.222 43.34 2.528 ;
      RECT 43.297 2.219 43.325 2.555 ;
      RECT 43.211 2.211 43.297 2.555 ;
      RECT 43.125 2.2 43.211 2.555 ;
      RECT 43.085 2.185 43.125 2.555 ;
      RECT 43.045 2.159 43.085 2.555 ;
      RECT 43.04 2.141 43.045 2.367 ;
      RECT 43.03 2.137 43.04 2.357 ;
      RECT 43.015 2.127 43.03 2.344 ;
      RECT 42.995 2.111 43.015 2.329 ;
      RECT 42.98 2.096 42.995 2.314 ;
      RECT 42.97 2.085 42.98 2.304 ;
      RECT 42.945 2.069 42.97 2.293 ;
      RECT 42.94 2.056 42.945 2.283 ;
      RECT 42.935 2.052 42.94 2.278 ;
      RECT 42.88 2.038 42.935 2.256 ;
      RECT 42.841 2.019 42.88 2.22 ;
      RECT 42.755 1.993 42.841 2.173 ;
      RECT 42.751 1.975 42.755 2.139 ;
      RECT 42.665 1.956 42.751 2.117 ;
      RECT 42.66 1.938 42.665 2.095 ;
      RECT 42.655 1.936 42.66 2.093 ;
      RECT 42.645 1.935 42.655 2.088 ;
      RECT 42.585 1.922 42.645 2.074 ;
      RECT 42.54 1.9 42.585 2.053 ;
      RECT 42.48 1.877 42.54 2.032 ;
      RECT 42.416 1.852 42.48 2.007 ;
      RECT 42.33 1.822 42.416 1.976 ;
      RECT 42.315 1.802 42.33 1.955 ;
      RECT 42.285 1.797 42.315 1.946 ;
      RECT 42.232 1.795 42.245 1.935 ;
      RECT 42.146 1.795 42.232 1.937 ;
      RECT 42.06 1.795 42.146 1.939 ;
      RECT 42.04 1.795 42.06 1.943 ;
      RECT 41.995 1.797 42.04 1.954 ;
      RECT 41.955 1.807 41.995 1.97 ;
      RECT 41.951 1.816 41.955 1.978 ;
      RECT 41.865 1.836 41.951 1.994 ;
      RECT 41.855 1.855 41.865 2.012 ;
      RECT 41.85 1.857 41.855 2.015 ;
      RECT 41.84 1.861 41.85 2.018 ;
      RECT 41.82 1.866 41.84 2.028 ;
      RECT 41.79 1.876 41.82 2.048 ;
      RECT 41.785 1.883 41.79 2.062 ;
      RECT 41.775 1.887 41.785 2.069 ;
      RECT 41.76 1.895 41.775 2.08 ;
      RECT 41.75 1.905 41.76 2.091 ;
      RECT 41.74 1.912 41.75 2.099 ;
      RECT 41.715 1.925 41.74 2.114 ;
      RECT 41.651 1.961 41.715 2.153 ;
      RECT 41.565 2.024 41.651 2.217 ;
      RECT 41.53 2.075 41.565 2.27 ;
      RECT 41.525 2.092 41.53 2.287 ;
      RECT 41.51 2.101 41.525 2.294 ;
      RECT 41.49 2.116 41.51 2.308 ;
      RECT 41.485 2.127 41.49 2.318 ;
      RECT 41.465 2.14 41.485 2.328 ;
      RECT 41.46 2.15 41.465 2.338 ;
      RECT 41.445 2.155 41.46 2.347 ;
      RECT 41.435 2.165 41.445 2.358 ;
      RECT 41.405 2.182 41.435 2.375 ;
      RECT 41.395 2.2 41.405 2.393 ;
      RECT 41.38 2.211 41.395 2.404 ;
      RECT 41.34 2.235 41.38 2.42 ;
      RECT 41.305 2.269 41.34 2.437 ;
      RECT 41.275 2.292 41.305 2.449 ;
      RECT 41.26 2.302 41.275 2.458 ;
      RECT 41.22 2.312 41.26 2.469 ;
      RECT 41.2 2.323 41.22 2.481 ;
      RECT 41.195 2.327 41.2 2.488 ;
      RECT 41.18 2.331 41.195 2.493 ;
      RECT 41.17 2.336 41.18 2.498 ;
      RECT 41.165 2.339 41.17 2.501 ;
      RECT 41.135 2.345 41.165 2.508 ;
      RECT 41.1 2.355 41.135 2.522 ;
      RECT 41.04 2.37 41.1 2.542 ;
      RECT 40.985 2.39 41.04 2.566 ;
      RECT 40.956 2.405 40.985 2.584 ;
      RECT 40.87 2.425 40.956 2.609 ;
      RECT 40.865 2.44 40.87 2.629 ;
      RECT 40.855 2.443 40.865 2.63 ;
      RECT 40.83 2.45 40.855 2.715 ;
      RECT 43.525 2.943 43.805 3.28 ;
      RECT 43.525 2.953 43.81 3.238 ;
      RECT 43.525 2.962 43.815 3.135 ;
      RECT 43.525 2.977 43.82 3.003 ;
      RECT 43.525 2.805 43.785 3.28 ;
      RECT 33.88 6.66 34.23 7.01 ;
      RECT 42.705 6.615 43.055 6.965 ;
      RECT 33.88 6.69 43.055 6.89 ;
      RECT 41.245 3.685 41.255 3.875 ;
      RECT 39.505 3.56 39.785 3.84 ;
      RECT 42.55 2.5 42.555 2.985 ;
      RECT 42.445 2.5 42.505 2.76 ;
      RECT 42.77 3.47 42.775 3.545 ;
      RECT 42.76 3.337 42.77 3.58 ;
      RECT 42.75 3.172 42.76 3.601 ;
      RECT 42.745 3.042 42.75 3.617 ;
      RECT 42.735 2.932 42.745 3.633 ;
      RECT 42.73 2.831 42.735 3.65 ;
      RECT 42.725 2.813 42.73 3.66 ;
      RECT 42.72 2.795 42.725 3.67 ;
      RECT 42.71 2.77 42.72 3.685 ;
      RECT 42.705 2.75 42.71 3.7 ;
      RECT 42.685 2.5 42.705 3.725 ;
      RECT 42.67 2.5 42.685 3.758 ;
      RECT 42.64 2.5 42.67 3.78 ;
      RECT 42.62 2.5 42.64 3.794 ;
      RECT 42.6 2.5 42.62 3.31 ;
      RECT 42.615 3.377 42.62 3.799 ;
      RECT 42.61 3.407 42.615 3.801 ;
      RECT 42.605 3.42 42.61 3.804 ;
      RECT 42.6 3.43 42.605 3.808 ;
      RECT 42.595 2.5 42.6 3.228 ;
      RECT 42.595 3.44 42.6 3.81 ;
      RECT 42.59 2.5 42.595 3.205 ;
      RECT 42.58 3.462 42.595 3.81 ;
      RECT 42.575 2.5 42.59 3.15 ;
      RECT 42.57 3.487 42.58 3.81 ;
      RECT 42.57 2.5 42.575 3.095 ;
      RECT 42.56 2.5 42.57 3.043 ;
      RECT 42.565 3.5 42.57 3.811 ;
      RECT 42.56 3.512 42.565 3.812 ;
      RECT 42.555 2.5 42.56 3.003 ;
      RECT 42.555 3.525 42.56 3.813 ;
      RECT 42.54 3.54 42.555 3.814 ;
      RECT 42.545 2.5 42.55 2.965 ;
      RECT 42.54 2.5 42.545 2.93 ;
      RECT 42.535 2.5 42.54 2.905 ;
      RECT 42.53 3.567 42.54 3.816 ;
      RECT 42.525 2.5 42.535 2.863 ;
      RECT 42.525 3.585 42.53 3.817 ;
      RECT 42.52 2.5 42.525 2.823 ;
      RECT 42.52 3.592 42.525 3.818 ;
      RECT 42.515 2.5 42.52 2.795 ;
      RECT 42.51 3.61 42.52 3.819 ;
      RECT 42.505 2.5 42.515 2.775 ;
      RECT 42.5 3.63 42.51 3.821 ;
      RECT 42.49 3.647 42.5 3.822 ;
      RECT 42.455 3.67 42.49 3.825 ;
      RECT 42.4 3.688 42.455 3.831 ;
      RECT 42.314 3.696 42.4 3.84 ;
      RECT 42.228 3.707 42.314 3.851 ;
      RECT 42.142 3.717 42.228 3.862 ;
      RECT 42.056 3.727 42.142 3.874 ;
      RECT 41.97 3.737 42.056 3.885 ;
      RECT 41.95 3.743 41.97 3.891 ;
      RECT 41.87 3.745 41.95 3.895 ;
      RECT 41.865 3.744 41.87 3.9 ;
      RECT 41.857 3.743 41.865 3.9 ;
      RECT 41.771 3.739 41.857 3.898 ;
      RECT 41.685 3.731 41.771 3.895 ;
      RECT 41.599 3.722 41.685 3.891 ;
      RECT 41.513 3.714 41.599 3.888 ;
      RECT 41.427 3.706 41.513 3.884 ;
      RECT 41.341 3.697 41.427 3.881 ;
      RECT 41.255 3.689 41.341 3.877 ;
      RECT 41.2 3.682 41.245 3.875 ;
      RECT 41.115 3.675 41.2 3.873 ;
      RECT 41.041 3.667 41.115 3.869 ;
      RECT 40.955 3.659 41.041 3.866 ;
      RECT 40.952 3.655 40.955 3.864 ;
      RECT 40.866 3.651 40.952 3.863 ;
      RECT 40.78 3.643 40.866 3.86 ;
      RECT 40.695 3.638 40.78 3.857 ;
      RECT 40.609 3.635 40.695 3.854 ;
      RECT 40.523 3.633 40.609 3.851 ;
      RECT 40.437 3.63 40.523 3.848 ;
      RECT 40.351 3.627 40.437 3.845 ;
      RECT 40.265 3.624 40.351 3.842 ;
      RECT 40.189 3.622 40.265 3.839 ;
      RECT 40.103 3.619 40.189 3.836 ;
      RECT 40.017 3.616 40.103 3.834 ;
      RECT 39.931 3.614 40.017 3.831 ;
      RECT 39.845 3.611 39.931 3.828 ;
      RECT 39.785 3.602 39.845 3.826 ;
      RECT 42.295 3.22 42.37 3.48 ;
      RECT 42.275 3.2 42.28 3.48 ;
      RECT 41.595 2.985 41.7 3.28 ;
      RECT 36.04 2.96 36.11 3.22 ;
      RECT 41.935 2.835 41.94 3.206 ;
      RECT 41.925 2.89 41.93 3.206 ;
      RECT 42.23 2.06 42.29 2.32 ;
      RECT 42.285 3.215 42.295 3.48 ;
      RECT 42.28 3.205 42.285 3.48 ;
      RECT 42.2 3.152 42.275 3.48 ;
      RECT 42.225 2.06 42.23 2.34 ;
      RECT 42.215 2.06 42.225 2.36 ;
      RECT 42.2 2.06 42.215 2.39 ;
      RECT 42.185 2.06 42.2 2.433 ;
      RECT 42.18 3.095 42.2 3.48 ;
      RECT 42.17 2.06 42.185 2.47 ;
      RECT 42.165 3.075 42.18 3.48 ;
      RECT 42.165 2.06 42.17 2.493 ;
      RECT 42.155 2.06 42.165 2.518 ;
      RECT 42.125 3.042 42.165 3.48 ;
      RECT 42.13 2.06 42.155 2.568 ;
      RECT 42.125 2.06 42.13 2.623 ;
      RECT 42.12 2.06 42.125 2.665 ;
      RECT 42.11 3.005 42.125 3.48 ;
      RECT 42.115 2.06 42.12 2.708 ;
      RECT 42.11 2.06 42.115 2.773 ;
      RECT 42.105 2.06 42.11 2.795 ;
      RECT 42.105 2.993 42.11 3.345 ;
      RECT 42.1 2.06 42.105 2.863 ;
      RECT 42.1 2.985 42.105 3.328 ;
      RECT 42.095 2.06 42.1 2.908 ;
      RECT 42.09 2.967 42.1 3.305 ;
      RECT 42.09 2.06 42.095 2.945 ;
      RECT 42.08 2.06 42.09 3.285 ;
      RECT 42.075 2.06 42.08 3.268 ;
      RECT 42.07 2.06 42.075 3.253 ;
      RECT 42.065 2.06 42.07 3.238 ;
      RECT 42.045 2.06 42.065 3.228 ;
      RECT 42.04 2.06 42.045 3.218 ;
      RECT 42.03 2.06 42.04 3.214 ;
      RECT 42.025 2.337 42.03 3.213 ;
      RECT 42.02 2.36 42.025 3.212 ;
      RECT 42.015 2.39 42.02 3.211 ;
      RECT 42.01 2.417 42.015 3.21 ;
      RECT 42.005 2.445 42.01 3.21 ;
      RECT 42 2.472 42.005 3.21 ;
      RECT 41.995 2.492 42 3.21 ;
      RECT 41.99 2.52 41.995 3.21 ;
      RECT 41.98 2.562 41.99 3.21 ;
      RECT 41.97 2.607 41.98 3.209 ;
      RECT 41.965 2.66 41.97 3.208 ;
      RECT 41.96 2.692 41.965 3.207 ;
      RECT 41.955 2.712 41.96 3.206 ;
      RECT 41.95 2.75 41.955 3.206 ;
      RECT 41.945 2.772 41.95 3.206 ;
      RECT 41.94 2.797 41.945 3.206 ;
      RECT 41.93 2.862 41.935 3.206 ;
      RECT 41.915 2.922 41.925 3.206 ;
      RECT 41.9 2.932 41.915 3.206 ;
      RECT 41.88 2.942 41.9 3.206 ;
      RECT 41.85 2.947 41.88 3.203 ;
      RECT 41.79 2.957 41.85 3.2 ;
      RECT 41.77 2.966 41.79 3.205 ;
      RECT 41.745 2.972 41.77 3.218 ;
      RECT 41.725 2.977 41.745 3.233 ;
      RECT 41.7 2.982 41.725 3.28 ;
      RECT 41.571 2.984 41.595 3.28 ;
      RECT 41.485 2.979 41.571 3.28 ;
      RECT 41.445 2.976 41.485 3.28 ;
      RECT 41.395 2.978 41.445 3.26 ;
      RECT 41.365 2.982 41.395 3.26 ;
      RECT 41.286 2.992 41.365 3.26 ;
      RECT 41.2 3.007 41.286 3.261 ;
      RECT 41.15 3.017 41.2 3.262 ;
      RECT 41.142 3.02 41.15 3.262 ;
      RECT 41.056 3.022 41.142 3.263 ;
      RECT 40.97 3.026 41.056 3.263 ;
      RECT 40.884 3.03 40.97 3.264 ;
      RECT 40.798 3.033 40.884 3.265 ;
      RECT 40.712 3.037 40.798 3.265 ;
      RECT 40.626 3.041 40.712 3.266 ;
      RECT 40.54 3.044 40.626 3.267 ;
      RECT 40.454 3.048 40.54 3.267 ;
      RECT 40.368 3.052 40.454 3.268 ;
      RECT 40.282 3.056 40.368 3.269 ;
      RECT 40.196 3.059 40.282 3.269 ;
      RECT 40.11 3.063 40.196 3.27 ;
      RECT 40.08 3.065 40.11 3.27 ;
      RECT 39.994 3.068 40.08 3.271 ;
      RECT 39.908 3.072 39.994 3.272 ;
      RECT 39.822 3.076 39.908 3.273 ;
      RECT 39.736 3.079 39.822 3.273 ;
      RECT 39.65 3.083 39.736 3.274 ;
      RECT 39.615 3.088 39.65 3.275 ;
      RECT 39.56 3.098 39.615 3.282 ;
      RECT 39.535 3.11 39.56 3.292 ;
      RECT 39.5 3.123 39.535 3.3 ;
      RECT 39.46 3.14 39.5 3.323 ;
      RECT 39.44 3.153 39.46 3.35 ;
      RECT 39.41 3.165 39.44 3.378 ;
      RECT 39.405 3.173 39.41 3.398 ;
      RECT 39.4 3.176 39.405 3.408 ;
      RECT 39.35 3.188 39.4 3.442 ;
      RECT 39.34 3.203 39.35 3.475 ;
      RECT 39.33 3.209 39.34 3.488 ;
      RECT 39.32 3.216 39.33 3.5 ;
      RECT 39.295 3.229 39.32 3.518 ;
      RECT 39.28 3.244 39.295 3.54 ;
      RECT 39.27 3.252 39.28 3.556 ;
      RECT 39.255 3.261 39.27 3.571 ;
      RECT 39.245 3.271 39.255 3.585 ;
      RECT 39.226 3.284 39.245 3.602 ;
      RECT 39.14 3.329 39.226 3.667 ;
      RECT 39.125 3.374 39.14 3.725 ;
      RECT 39.12 3.383 39.125 3.738 ;
      RECT 39.11 3.39 39.12 3.743 ;
      RECT 39.105 3.395 39.11 3.747 ;
      RECT 39.085 3.405 39.105 3.754 ;
      RECT 39.06 3.425 39.085 3.768 ;
      RECT 39.025 3.45 39.06 3.788 ;
      RECT 39.01 3.473 39.025 3.803 ;
      RECT 39 3.483 39.01 3.808 ;
      RECT 38.99 3.491 39 3.815 ;
      RECT 38.98 3.5 38.99 3.821 ;
      RECT 38.96 3.512 38.98 3.823 ;
      RECT 38.95 3.525 38.96 3.825 ;
      RECT 38.925 3.54 38.95 3.828 ;
      RECT 38.905 3.557 38.925 3.832 ;
      RECT 38.865 3.585 38.905 3.838 ;
      RECT 38.8 3.632 38.865 3.847 ;
      RECT 38.785 3.665 38.8 3.855 ;
      RECT 38.78 3.672 38.785 3.857 ;
      RECT 38.73 3.697 38.78 3.862 ;
      RECT 38.715 3.721 38.73 3.869 ;
      RECT 38.665 3.726 38.715 3.87 ;
      RECT 38.579 3.73 38.665 3.87 ;
      RECT 38.493 3.73 38.579 3.87 ;
      RECT 38.407 3.73 38.493 3.871 ;
      RECT 38.321 3.73 38.407 3.871 ;
      RECT 38.235 3.73 38.321 3.871 ;
      RECT 38.169 3.73 38.235 3.871 ;
      RECT 38.083 3.73 38.169 3.872 ;
      RECT 37.997 3.73 38.083 3.872 ;
      RECT 37.911 3.731 37.997 3.873 ;
      RECT 37.825 3.731 37.911 3.873 ;
      RECT 37.739 3.731 37.825 3.873 ;
      RECT 37.653 3.731 37.739 3.874 ;
      RECT 37.567 3.731 37.653 3.874 ;
      RECT 37.481 3.732 37.567 3.875 ;
      RECT 37.395 3.732 37.481 3.875 ;
      RECT 37.375 3.732 37.395 3.875 ;
      RECT 37.289 3.732 37.375 3.875 ;
      RECT 37.203 3.732 37.289 3.875 ;
      RECT 37.117 3.733 37.203 3.875 ;
      RECT 37.031 3.733 37.117 3.875 ;
      RECT 36.945 3.733 37.031 3.875 ;
      RECT 36.859 3.734 36.945 3.875 ;
      RECT 36.773 3.734 36.859 3.875 ;
      RECT 36.687 3.734 36.773 3.875 ;
      RECT 36.601 3.734 36.687 3.875 ;
      RECT 36.515 3.735 36.601 3.875 ;
      RECT 36.465 3.732 36.515 3.875 ;
      RECT 36.455 3.73 36.465 3.874 ;
      RECT 36.451 3.73 36.455 3.873 ;
      RECT 36.365 3.725 36.451 3.868 ;
      RECT 36.343 3.718 36.365 3.862 ;
      RECT 36.257 3.709 36.343 3.856 ;
      RECT 36.171 3.696 36.257 3.847 ;
      RECT 36.085 3.682 36.171 3.837 ;
      RECT 36.04 3.672 36.085 3.83 ;
      RECT 36.02 2.96 36.04 3.238 ;
      RECT 36.02 3.665 36.04 3.826 ;
      RECT 35.99 2.96 36.02 3.26 ;
      RECT 35.98 3.632 36.02 3.823 ;
      RECT 35.975 2.96 35.99 3.28 ;
      RECT 35.975 3.597 35.98 3.821 ;
      RECT 35.97 2.96 35.975 3.405 ;
      RECT 35.97 3.557 35.975 3.821 ;
      RECT 35.96 2.96 35.97 3.821 ;
      RECT 35.885 2.96 35.96 3.815 ;
      RECT 35.855 2.96 35.885 3.805 ;
      RECT 35.85 2.96 35.855 3.797 ;
      RECT 35.845 3.002 35.85 3.79 ;
      RECT 35.835 3.071 35.845 3.781 ;
      RECT 35.83 3.141 35.835 3.733 ;
      RECT 35.825 3.205 35.83 3.63 ;
      RECT 35.82 3.24 35.825 3.585 ;
      RECT 35.818 3.277 35.82 3.477 ;
      RECT 35.815 3.285 35.818 3.47 ;
      RECT 35.81 3.35 35.815 3.413 ;
      RECT 39.885 2.44 40.165 2.72 ;
      RECT 39.875 2.44 40.165 2.583 ;
      RECT 39.83 2.305 40.09 2.565 ;
      RECT 39.83 2.42 40.145 2.565 ;
      RECT 39.83 2.39 40.14 2.565 ;
      RECT 39.83 2.377 40.13 2.565 ;
      RECT 39.83 2.367 40.125 2.565 ;
      RECT 35.805 2.35 36.065 2.61 ;
      RECT 39.575 1.9 39.835 2.16 ;
      RECT 39.565 1.925 39.835 2.12 ;
      RECT 39.56 1.925 39.565 2.119 ;
      RECT 39.49 1.92 39.56 2.111 ;
      RECT 39.405 1.907 39.49 2.094 ;
      RECT 39.401 1.899 39.405 2.084 ;
      RECT 39.315 1.892 39.401 2.074 ;
      RECT 39.306 1.884 39.315 2.064 ;
      RECT 39.22 1.877 39.306 2.052 ;
      RECT 39.2 1.868 39.22 2.038 ;
      RECT 39.145 1.863 39.2 2.03 ;
      RECT 39.135 1.857 39.145 2.024 ;
      RECT 39.115 1.855 39.135 2.02 ;
      RECT 39.107 1.854 39.115 2.016 ;
      RECT 39.021 1.846 39.107 2.005 ;
      RECT 38.935 1.832 39.021 1.985 ;
      RECT 38.875 1.82 38.935 1.97 ;
      RECT 38.865 1.815 38.875 1.965 ;
      RECT 38.815 1.815 38.865 1.967 ;
      RECT 38.768 1.817 38.815 1.971 ;
      RECT 38.682 1.824 38.768 1.976 ;
      RECT 38.596 1.832 38.682 1.982 ;
      RECT 38.51 1.841 38.596 1.988 ;
      RECT 38.451 1.847 38.51 1.993 ;
      RECT 38.365 1.852 38.451 1.999 ;
      RECT 38.29 1.857 38.365 2.005 ;
      RECT 38.251 1.859 38.29 2.01 ;
      RECT 38.165 1.856 38.251 2.015 ;
      RECT 38.08 1.854 38.165 2.022 ;
      RECT 38.048 1.853 38.08 2.025 ;
      RECT 37.962 1.852 38.048 2.026 ;
      RECT 37.876 1.851 37.962 2.027 ;
      RECT 37.79 1.85 37.876 2.027 ;
      RECT 37.704 1.849 37.79 2.028 ;
      RECT 37.618 1.848 37.704 2.029 ;
      RECT 37.532 1.847 37.618 2.03 ;
      RECT 37.446 1.846 37.532 2.03 ;
      RECT 37.36 1.845 37.446 2.031 ;
      RECT 37.31 1.845 37.36 2.032 ;
      RECT 37.296 1.846 37.31 2.032 ;
      RECT 37.21 1.853 37.296 2.033 ;
      RECT 37.136 1.864 37.21 2.034 ;
      RECT 37.05 1.873 37.136 2.035 ;
      RECT 37.015 1.88 37.05 2.05 ;
      RECT 36.99 1.883 37.015 2.08 ;
      RECT 36.965 1.892 36.99 2.109 ;
      RECT 36.955 1.903 36.965 2.129 ;
      RECT 36.945 1.911 36.955 2.143 ;
      RECT 36.94 1.917 36.945 2.153 ;
      RECT 36.915 1.934 36.94 2.17 ;
      RECT 36.9 1.956 36.915 2.198 ;
      RECT 36.87 1.982 36.9 2.228 ;
      RECT 36.85 2.011 36.87 2.258 ;
      RECT 36.845 2.026 36.85 2.275 ;
      RECT 36.825 2.041 36.845 2.29 ;
      RECT 36.815 2.059 36.825 2.308 ;
      RECT 36.805 2.07 36.815 2.323 ;
      RECT 36.755 2.102 36.805 2.349 ;
      RECT 36.75 2.132 36.755 2.369 ;
      RECT 36.74 2.145 36.75 2.375 ;
      RECT 36.731 2.155 36.74 2.383 ;
      RECT 36.72 2.166 36.731 2.391 ;
      RECT 36.715 2.176 36.72 2.397 ;
      RECT 36.7 2.197 36.715 2.404 ;
      RECT 36.685 2.227 36.7 2.412 ;
      RECT 36.65 2.257 36.685 2.418 ;
      RECT 36.625 2.275 36.65 2.425 ;
      RECT 36.575 2.283 36.625 2.434 ;
      RECT 36.55 2.288 36.575 2.443 ;
      RECT 36.495 2.294 36.55 2.453 ;
      RECT 36.49 2.299 36.495 2.461 ;
      RECT 36.476 2.302 36.49 2.463 ;
      RECT 36.39 2.314 36.476 2.475 ;
      RECT 36.38 2.326 36.39 2.488 ;
      RECT 36.295 2.339 36.38 2.5 ;
      RECT 36.251 2.356 36.295 2.514 ;
      RECT 36.165 2.373 36.251 2.53 ;
      RECT 36.135 2.387 36.165 2.544 ;
      RECT 36.125 2.392 36.135 2.549 ;
      RECT 36.065 2.395 36.125 2.558 ;
      RECT 38.955 2.665 39.215 2.925 ;
      RECT 38.955 2.665 39.235 2.778 ;
      RECT 38.955 2.665 39.26 2.745 ;
      RECT 38.955 2.665 39.265 2.725 ;
      RECT 39.005 2.44 39.285 2.72 ;
      RECT 38.56 3.175 38.82 3.435 ;
      RECT 38.55 3.032 38.745 3.373 ;
      RECT 38.545 3.14 38.76 3.365 ;
      RECT 38.54 3.19 38.82 3.355 ;
      RECT 38.53 3.267 38.82 3.34 ;
      RECT 38.55 3.115 38.76 3.373 ;
      RECT 38.56 2.99 38.745 3.435 ;
      RECT 38.56 2.885 38.725 3.435 ;
      RECT 38.57 2.872 38.725 3.435 ;
      RECT 38.57 2.83 38.715 3.435 ;
      RECT 38.575 2.755 38.715 3.435 ;
      RECT 38.605 2.405 38.715 3.435 ;
      RECT 38.61 2.135 38.735 2.758 ;
      RECT 38.58 2.71 38.735 2.758 ;
      RECT 38.595 2.512 38.715 3.435 ;
      RECT 38.585 2.622 38.735 2.758 ;
      RECT 38.61 2.135 38.75 2.615 ;
      RECT 38.61 2.135 38.77 2.49 ;
      RECT 38.575 2.135 38.835 2.395 ;
      RECT 38.045 2.44 38.325 2.72 ;
      RECT 38.03 2.44 38.325 2.7 ;
      RECT 36.085 3.305 36.345 3.565 ;
      RECT 37.87 3.16 38.13 3.42 ;
      RECT 37.85 3.18 38.13 3.395 ;
      RECT 37.807 3.18 37.85 3.394 ;
      RECT 37.721 3.181 37.807 3.391 ;
      RECT 37.635 3.182 37.721 3.387 ;
      RECT 37.56 3.184 37.635 3.384 ;
      RECT 37.537 3.185 37.56 3.382 ;
      RECT 37.451 3.186 37.537 3.38 ;
      RECT 37.365 3.187 37.451 3.377 ;
      RECT 37.341 3.188 37.365 3.375 ;
      RECT 37.255 3.19 37.341 3.372 ;
      RECT 37.17 3.192 37.255 3.373 ;
      RECT 37.113 3.193 37.17 3.379 ;
      RECT 37.027 3.195 37.113 3.389 ;
      RECT 36.941 3.198 37.027 3.402 ;
      RECT 36.855 3.2 36.941 3.414 ;
      RECT 36.841 3.201 36.855 3.421 ;
      RECT 36.755 3.202 36.841 3.429 ;
      RECT 36.715 3.204 36.755 3.438 ;
      RECT 36.706 3.205 36.715 3.441 ;
      RECT 36.62 3.213 36.706 3.447 ;
      RECT 36.6 3.222 36.62 3.455 ;
      RECT 36.515 3.237 36.6 3.463 ;
      RECT 36.455 3.26 36.515 3.474 ;
      RECT 36.445 3.272 36.455 3.479 ;
      RECT 36.405 3.282 36.445 3.483 ;
      RECT 36.35 3.299 36.405 3.491 ;
      RECT 36.345 3.309 36.35 3.495 ;
      RECT 37.411 2.44 37.47 2.837 ;
      RECT 37.325 2.44 37.53 2.828 ;
      RECT 37.32 2.47 37.53 2.823 ;
      RECT 37.286 2.47 37.53 2.821 ;
      RECT 37.2 2.47 37.53 2.815 ;
      RECT 37.155 2.47 37.55 2.793 ;
      RECT 37.155 2.47 37.57 2.748 ;
      RECT 37.115 2.47 37.57 2.738 ;
      RECT 37.325 2.44 37.605 2.72 ;
      RECT 37.06 2.44 37.32 2.7 ;
      RECT 34.885 3 35.165 3.28 ;
      RECT 34.855 2.962 35.11 3.265 ;
      RECT 34.85 2.963 35.11 3.263 ;
      RECT 34.845 2.964 35.11 3.257 ;
      RECT 34.84 2.967 35.11 3.25 ;
      RECT 34.835 3 35.165 3.243 ;
      RECT 34.805 2.97 35.11 3.23 ;
      RECT 34.805 2.997 35.13 3.23 ;
      RECT 34.805 2.987 35.125 3.23 ;
      RECT 34.805 2.972 35.12 3.23 ;
      RECT 34.885 2.959 35.1 3.28 ;
      RECT 34.971 2.957 35.1 3.28 ;
      RECT 35.057 2.955 35.085 3.28 ;
      RECT 30.7 6.22 31.02 6.545 ;
      RECT 30.73 5.695 30.9 6.545 ;
      RECT 30.73 5.695 30.905 6.045 ;
      RECT 30.73 5.695 31.705 5.87 ;
      RECT 31.53 1.965 31.705 5.87 ;
      RECT 31.475 1.965 31.825 2.315 ;
      RECT 31.5 6.655 31.825 6.98 ;
      RECT 30.385 6.745 31.825 6.915 ;
      RECT 30.385 2.395 30.545 6.915 ;
      RECT 30.7 2.365 31.02 2.685 ;
      RECT 30.385 2.395 31.02 2.565 ;
      RECT 20.47 1.92 20.73 2.18 ;
      RECT 20.525 1.88 20.83 2.16 ;
      RECT 20.525 1.42 20.7 2.18 ;
      RECT 29.04 1.34 29.39 1.69 ;
      RECT 20.525 1.42 29.39 1.595 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 28.8 2.235 28.97 3.22 ;
      RECT 24.82 2.455 25.055 2.715 ;
      RECT 27.965 2.235 28.13 2.495 ;
      RECT 27.87 2.225 27.885 2.495 ;
      RECT 27.965 2.235 28.97 2.415 ;
      RECT 26.47 1.795 26.51 1.935 ;
      RECT 27.885 2.23 27.965 2.495 ;
      RECT 27.83 2.225 27.87 2.461 ;
      RECT 27.816 2.225 27.83 2.461 ;
      RECT 27.73 2.23 27.816 2.463 ;
      RECT 27.685 2.237 27.73 2.465 ;
      RECT 27.655 2.237 27.685 2.467 ;
      RECT 27.63 2.232 27.655 2.469 ;
      RECT 27.6 2.228 27.63 2.478 ;
      RECT 27.59 2.225 27.6 2.49 ;
      RECT 27.585 2.225 27.59 2.498 ;
      RECT 27.58 2.225 27.585 2.503 ;
      RECT 27.57 2.224 27.58 2.513 ;
      RECT 27.565 2.223 27.57 2.523 ;
      RECT 27.55 2.222 27.565 2.528 ;
      RECT 27.522 2.219 27.55 2.555 ;
      RECT 27.436 2.211 27.522 2.555 ;
      RECT 27.35 2.2 27.436 2.555 ;
      RECT 27.31 2.185 27.35 2.555 ;
      RECT 27.27 2.159 27.31 2.555 ;
      RECT 27.265 2.141 27.27 2.367 ;
      RECT 27.255 2.137 27.265 2.357 ;
      RECT 27.24 2.127 27.255 2.344 ;
      RECT 27.22 2.111 27.24 2.329 ;
      RECT 27.205 2.096 27.22 2.314 ;
      RECT 27.195 2.085 27.205 2.304 ;
      RECT 27.17 2.069 27.195 2.293 ;
      RECT 27.165 2.056 27.17 2.283 ;
      RECT 27.16 2.052 27.165 2.278 ;
      RECT 27.105 2.038 27.16 2.256 ;
      RECT 27.066 2.019 27.105 2.22 ;
      RECT 26.98 1.993 27.066 2.173 ;
      RECT 26.976 1.975 26.98 2.139 ;
      RECT 26.89 1.956 26.976 2.117 ;
      RECT 26.885 1.938 26.89 2.095 ;
      RECT 26.88 1.936 26.885 2.093 ;
      RECT 26.87 1.935 26.88 2.088 ;
      RECT 26.81 1.922 26.87 2.074 ;
      RECT 26.765 1.9 26.81 2.053 ;
      RECT 26.705 1.877 26.765 2.032 ;
      RECT 26.641 1.852 26.705 2.007 ;
      RECT 26.555 1.822 26.641 1.976 ;
      RECT 26.54 1.802 26.555 1.955 ;
      RECT 26.51 1.797 26.54 1.946 ;
      RECT 26.457 1.795 26.47 1.935 ;
      RECT 26.371 1.795 26.457 1.937 ;
      RECT 26.285 1.795 26.371 1.939 ;
      RECT 26.265 1.795 26.285 1.943 ;
      RECT 26.22 1.797 26.265 1.954 ;
      RECT 26.18 1.807 26.22 1.97 ;
      RECT 26.176 1.816 26.18 1.978 ;
      RECT 26.09 1.836 26.176 1.994 ;
      RECT 26.08 1.855 26.09 2.012 ;
      RECT 26.075 1.857 26.08 2.015 ;
      RECT 26.065 1.861 26.075 2.018 ;
      RECT 26.045 1.866 26.065 2.028 ;
      RECT 26.015 1.876 26.045 2.048 ;
      RECT 26.01 1.883 26.015 2.062 ;
      RECT 26 1.887 26.01 2.069 ;
      RECT 25.985 1.895 26 2.08 ;
      RECT 25.975 1.905 25.985 2.091 ;
      RECT 25.965 1.912 25.975 2.099 ;
      RECT 25.94 1.925 25.965 2.114 ;
      RECT 25.876 1.961 25.94 2.153 ;
      RECT 25.79 2.024 25.876 2.217 ;
      RECT 25.755 2.075 25.79 2.27 ;
      RECT 25.75 2.092 25.755 2.287 ;
      RECT 25.735 2.101 25.75 2.294 ;
      RECT 25.715 2.116 25.735 2.308 ;
      RECT 25.71 2.127 25.715 2.318 ;
      RECT 25.69 2.14 25.71 2.328 ;
      RECT 25.685 2.15 25.69 2.338 ;
      RECT 25.67 2.155 25.685 2.347 ;
      RECT 25.66 2.165 25.67 2.358 ;
      RECT 25.63 2.182 25.66 2.375 ;
      RECT 25.62 2.2 25.63 2.393 ;
      RECT 25.605 2.211 25.62 2.404 ;
      RECT 25.565 2.235 25.605 2.42 ;
      RECT 25.53 2.269 25.565 2.437 ;
      RECT 25.5 2.292 25.53 2.449 ;
      RECT 25.485 2.302 25.5 2.458 ;
      RECT 25.445 2.312 25.485 2.469 ;
      RECT 25.425 2.323 25.445 2.481 ;
      RECT 25.42 2.327 25.425 2.488 ;
      RECT 25.405 2.331 25.42 2.493 ;
      RECT 25.395 2.336 25.405 2.498 ;
      RECT 25.39 2.339 25.395 2.501 ;
      RECT 25.36 2.345 25.39 2.508 ;
      RECT 25.325 2.355 25.36 2.522 ;
      RECT 25.265 2.37 25.325 2.542 ;
      RECT 25.21 2.39 25.265 2.566 ;
      RECT 25.181 2.405 25.21 2.584 ;
      RECT 25.095 2.425 25.181 2.609 ;
      RECT 25.09 2.44 25.095 2.629 ;
      RECT 25.08 2.443 25.09 2.63 ;
      RECT 25.055 2.45 25.08 2.715 ;
      RECT 27.75 2.943 28.03 3.28 ;
      RECT 27.75 2.953 28.035 3.238 ;
      RECT 27.75 2.962 28.04 3.135 ;
      RECT 27.75 2.977 28.045 3.003 ;
      RECT 27.75 2.805 28.01 3.28 ;
      RECT 18.1 6.655 18.45 7.005 ;
      RECT 26.925 6.61 27.275 6.96 ;
      RECT 18.1 6.685 27.275 6.885 ;
      RECT 25.47 3.685 25.48 3.875 ;
      RECT 23.73 3.56 24.01 3.84 ;
      RECT 26.775 2.5 26.78 2.985 ;
      RECT 26.67 2.5 26.73 2.76 ;
      RECT 26.995 3.47 27 3.545 ;
      RECT 26.985 3.337 26.995 3.58 ;
      RECT 26.975 3.172 26.985 3.601 ;
      RECT 26.97 3.042 26.975 3.617 ;
      RECT 26.96 2.932 26.97 3.633 ;
      RECT 26.955 2.831 26.96 3.65 ;
      RECT 26.95 2.813 26.955 3.66 ;
      RECT 26.945 2.795 26.95 3.67 ;
      RECT 26.935 2.77 26.945 3.685 ;
      RECT 26.93 2.75 26.935 3.7 ;
      RECT 26.91 2.5 26.93 3.725 ;
      RECT 26.895 2.5 26.91 3.758 ;
      RECT 26.865 2.5 26.895 3.78 ;
      RECT 26.845 2.5 26.865 3.794 ;
      RECT 26.825 2.5 26.845 3.31 ;
      RECT 26.84 3.377 26.845 3.799 ;
      RECT 26.835 3.407 26.84 3.801 ;
      RECT 26.83 3.42 26.835 3.804 ;
      RECT 26.825 3.43 26.83 3.808 ;
      RECT 26.82 2.5 26.825 3.228 ;
      RECT 26.82 3.44 26.825 3.81 ;
      RECT 26.815 2.5 26.82 3.205 ;
      RECT 26.805 3.462 26.82 3.81 ;
      RECT 26.8 2.5 26.815 3.15 ;
      RECT 26.795 3.487 26.805 3.81 ;
      RECT 26.795 2.5 26.8 3.095 ;
      RECT 26.785 2.5 26.795 3.043 ;
      RECT 26.79 3.5 26.795 3.811 ;
      RECT 26.785 3.512 26.79 3.812 ;
      RECT 26.78 2.5 26.785 3.003 ;
      RECT 26.78 3.525 26.785 3.813 ;
      RECT 26.765 3.54 26.78 3.814 ;
      RECT 26.77 2.5 26.775 2.965 ;
      RECT 26.765 2.5 26.77 2.93 ;
      RECT 26.76 2.5 26.765 2.905 ;
      RECT 26.755 3.567 26.765 3.816 ;
      RECT 26.75 2.5 26.76 2.863 ;
      RECT 26.75 3.585 26.755 3.817 ;
      RECT 26.745 2.5 26.75 2.823 ;
      RECT 26.745 3.592 26.75 3.818 ;
      RECT 26.74 2.5 26.745 2.795 ;
      RECT 26.735 3.61 26.745 3.819 ;
      RECT 26.73 2.5 26.74 2.775 ;
      RECT 26.725 3.63 26.735 3.821 ;
      RECT 26.715 3.647 26.725 3.822 ;
      RECT 26.68 3.67 26.715 3.825 ;
      RECT 26.625 3.688 26.68 3.831 ;
      RECT 26.539 3.696 26.625 3.84 ;
      RECT 26.453 3.707 26.539 3.851 ;
      RECT 26.367 3.717 26.453 3.862 ;
      RECT 26.281 3.727 26.367 3.874 ;
      RECT 26.195 3.737 26.281 3.885 ;
      RECT 26.175 3.743 26.195 3.891 ;
      RECT 26.095 3.745 26.175 3.895 ;
      RECT 26.09 3.744 26.095 3.9 ;
      RECT 26.082 3.743 26.09 3.9 ;
      RECT 25.996 3.739 26.082 3.898 ;
      RECT 25.91 3.731 25.996 3.895 ;
      RECT 25.824 3.722 25.91 3.891 ;
      RECT 25.738 3.714 25.824 3.888 ;
      RECT 25.652 3.706 25.738 3.884 ;
      RECT 25.566 3.697 25.652 3.881 ;
      RECT 25.48 3.689 25.566 3.877 ;
      RECT 25.425 3.682 25.47 3.875 ;
      RECT 25.34 3.675 25.425 3.873 ;
      RECT 25.266 3.667 25.34 3.869 ;
      RECT 25.18 3.659 25.266 3.866 ;
      RECT 25.177 3.655 25.18 3.864 ;
      RECT 25.091 3.651 25.177 3.863 ;
      RECT 25.005 3.643 25.091 3.86 ;
      RECT 24.92 3.638 25.005 3.857 ;
      RECT 24.834 3.635 24.92 3.854 ;
      RECT 24.748 3.633 24.834 3.851 ;
      RECT 24.662 3.63 24.748 3.848 ;
      RECT 24.576 3.627 24.662 3.845 ;
      RECT 24.49 3.624 24.576 3.842 ;
      RECT 24.414 3.622 24.49 3.839 ;
      RECT 24.328 3.619 24.414 3.836 ;
      RECT 24.242 3.616 24.328 3.834 ;
      RECT 24.156 3.614 24.242 3.831 ;
      RECT 24.07 3.611 24.156 3.828 ;
      RECT 24.01 3.602 24.07 3.826 ;
      RECT 26.52 3.22 26.595 3.48 ;
      RECT 26.5 3.2 26.505 3.48 ;
      RECT 25.82 2.985 25.925 3.28 ;
      RECT 20.265 2.96 20.335 3.22 ;
      RECT 26.16 2.835 26.165 3.206 ;
      RECT 26.15 2.89 26.155 3.206 ;
      RECT 26.455 2.06 26.515 2.32 ;
      RECT 26.51 3.215 26.52 3.48 ;
      RECT 26.505 3.205 26.51 3.48 ;
      RECT 26.425 3.152 26.5 3.48 ;
      RECT 26.45 2.06 26.455 2.34 ;
      RECT 26.44 2.06 26.45 2.36 ;
      RECT 26.425 2.06 26.44 2.39 ;
      RECT 26.41 2.06 26.425 2.433 ;
      RECT 26.405 3.095 26.425 3.48 ;
      RECT 26.395 2.06 26.41 2.47 ;
      RECT 26.39 3.075 26.405 3.48 ;
      RECT 26.39 2.06 26.395 2.493 ;
      RECT 26.38 2.06 26.39 2.518 ;
      RECT 26.35 3.042 26.39 3.48 ;
      RECT 26.355 2.06 26.38 2.568 ;
      RECT 26.35 2.06 26.355 2.623 ;
      RECT 26.345 2.06 26.35 2.665 ;
      RECT 26.335 3.005 26.35 3.48 ;
      RECT 26.34 2.06 26.345 2.708 ;
      RECT 26.335 2.06 26.34 2.773 ;
      RECT 26.33 2.06 26.335 2.795 ;
      RECT 26.33 2.993 26.335 3.345 ;
      RECT 26.325 2.06 26.33 2.863 ;
      RECT 26.325 2.985 26.33 3.328 ;
      RECT 26.32 2.06 26.325 2.908 ;
      RECT 26.315 2.967 26.325 3.305 ;
      RECT 26.315 2.06 26.32 2.945 ;
      RECT 26.305 2.06 26.315 3.285 ;
      RECT 26.3 2.06 26.305 3.268 ;
      RECT 26.295 2.06 26.3 3.253 ;
      RECT 26.29 2.06 26.295 3.238 ;
      RECT 26.27 2.06 26.29 3.228 ;
      RECT 26.265 2.06 26.27 3.218 ;
      RECT 26.255 2.06 26.265 3.214 ;
      RECT 26.25 2.337 26.255 3.213 ;
      RECT 26.245 2.36 26.25 3.212 ;
      RECT 26.24 2.39 26.245 3.211 ;
      RECT 26.235 2.417 26.24 3.21 ;
      RECT 26.23 2.445 26.235 3.21 ;
      RECT 26.225 2.472 26.23 3.21 ;
      RECT 26.22 2.492 26.225 3.21 ;
      RECT 26.215 2.52 26.22 3.21 ;
      RECT 26.205 2.562 26.215 3.21 ;
      RECT 26.195 2.607 26.205 3.209 ;
      RECT 26.19 2.66 26.195 3.208 ;
      RECT 26.185 2.692 26.19 3.207 ;
      RECT 26.18 2.712 26.185 3.206 ;
      RECT 26.175 2.75 26.18 3.206 ;
      RECT 26.17 2.772 26.175 3.206 ;
      RECT 26.165 2.797 26.17 3.206 ;
      RECT 26.155 2.862 26.16 3.206 ;
      RECT 26.14 2.922 26.15 3.206 ;
      RECT 26.125 2.932 26.14 3.206 ;
      RECT 26.105 2.942 26.125 3.206 ;
      RECT 26.075 2.947 26.105 3.203 ;
      RECT 26.015 2.957 26.075 3.2 ;
      RECT 25.995 2.966 26.015 3.205 ;
      RECT 25.97 2.972 25.995 3.218 ;
      RECT 25.95 2.977 25.97 3.233 ;
      RECT 25.925 2.982 25.95 3.28 ;
      RECT 25.796 2.984 25.82 3.28 ;
      RECT 25.71 2.979 25.796 3.28 ;
      RECT 25.67 2.976 25.71 3.28 ;
      RECT 25.62 2.978 25.67 3.26 ;
      RECT 25.59 2.982 25.62 3.26 ;
      RECT 25.511 2.992 25.59 3.26 ;
      RECT 25.425 3.007 25.511 3.261 ;
      RECT 25.375 3.017 25.425 3.262 ;
      RECT 25.367 3.02 25.375 3.262 ;
      RECT 25.281 3.022 25.367 3.263 ;
      RECT 25.195 3.026 25.281 3.263 ;
      RECT 25.109 3.03 25.195 3.264 ;
      RECT 25.023 3.033 25.109 3.265 ;
      RECT 24.937 3.037 25.023 3.265 ;
      RECT 24.851 3.041 24.937 3.266 ;
      RECT 24.765 3.044 24.851 3.267 ;
      RECT 24.679 3.048 24.765 3.267 ;
      RECT 24.593 3.052 24.679 3.268 ;
      RECT 24.507 3.056 24.593 3.269 ;
      RECT 24.421 3.059 24.507 3.269 ;
      RECT 24.335 3.063 24.421 3.27 ;
      RECT 24.305 3.065 24.335 3.27 ;
      RECT 24.219 3.068 24.305 3.271 ;
      RECT 24.133 3.072 24.219 3.272 ;
      RECT 24.047 3.076 24.133 3.273 ;
      RECT 23.961 3.079 24.047 3.273 ;
      RECT 23.875 3.083 23.961 3.274 ;
      RECT 23.84 3.088 23.875 3.275 ;
      RECT 23.785 3.098 23.84 3.282 ;
      RECT 23.76 3.11 23.785 3.292 ;
      RECT 23.725 3.123 23.76 3.3 ;
      RECT 23.685 3.14 23.725 3.323 ;
      RECT 23.665 3.153 23.685 3.35 ;
      RECT 23.635 3.165 23.665 3.378 ;
      RECT 23.63 3.173 23.635 3.398 ;
      RECT 23.625 3.176 23.63 3.408 ;
      RECT 23.575 3.188 23.625 3.442 ;
      RECT 23.565 3.203 23.575 3.475 ;
      RECT 23.555 3.209 23.565 3.488 ;
      RECT 23.545 3.216 23.555 3.5 ;
      RECT 23.52 3.229 23.545 3.518 ;
      RECT 23.505 3.244 23.52 3.54 ;
      RECT 23.495 3.252 23.505 3.556 ;
      RECT 23.48 3.261 23.495 3.571 ;
      RECT 23.47 3.271 23.48 3.585 ;
      RECT 23.451 3.284 23.47 3.602 ;
      RECT 23.365 3.329 23.451 3.667 ;
      RECT 23.35 3.374 23.365 3.725 ;
      RECT 23.345 3.383 23.35 3.738 ;
      RECT 23.335 3.39 23.345 3.743 ;
      RECT 23.33 3.395 23.335 3.747 ;
      RECT 23.31 3.405 23.33 3.754 ;
      RECT 23.285 3.425 23.31 3.768 ;
      RECT 23.25 3.45 23.285 3.788 ;
      RECT 23.235 3.473 23.25 3.803 ;
      RECT 23.225 3.483 23.235 3.808 ;
      RECT 23.215 3.491 23.225 3.815 ;
      RECT 23.205 3.5 23.215 3.821 ;
      RECT 23.185 3.512 23.205 3.823 ;
      RECT 23.175 3.525 23.185 3.825 ;
      RECT 23.15 3.54 23.175 3.828 ;
      RECT 23.13 3.557 23.15 3.832 ;
      RECT 23.09 3.585 23.13 3.838 ;
      RECT 23.025 3.632 23.09 3.847 ;
      RECT 23.01 3.665 23.025 3.855 ;
      RECT 23.005 3.672 23.01 3.857 ;
      RECT 22.955 3.697 23.005 3.862 ;
      RECT 22.94 3.721 22.955 3.869 ;
      RECT 22.89 3.726 22.94 3.87 ;
      RECT 22.804 3.73 22.89 3.87 ;
      RECT 22.718 3.73 22.804 3.87 ;
      RECT 22.632 3.73 22.718 3.871 ;
      RECT 22.546 3.73 22.632 3.871 ;
      RECT 22.46 3.73 22.546 3.871 ;
      RECT 22.394 3.73 22.46 3.871 ;
      RECT 22.308 3.73 22.394 3.872 ;
      RECT 22.222 3.73 22.308 3.872 ;
      RECT 22.136 3.731 22.222 3.873 ;
      RECT 22.05 3.731 22.136 3.873 ;
      RECT 21.964 3.731 22.05 3.873 ;
      RECT 21.878 3.731 21.964 3.874 ;
      RECT 21.792 3.731 21.878 3.874 ;
      RECT 21.706 3.732 21.792 3.875 ;
      RECT 21.62 3.732 21.706 3.875 ;
      RECT 21.6 3.732 21.62 3.875 ;
      RECT 21.514 3.732 21.6 3.875 ;
      RECT 21.428 3.732 21.514 3.875 ;
      RECT 21.342 3.733 21.428 3.875 ;
      RECT 21.256 3.733 21.342 3.875 ;
      RECT 21.17 3.733 21.256 3.875 ;
      RECT 21.084 3.734 21.17 3.875 ;
      RECT 20.998 3.734 21.084 3.875 ;
      RECT 20.912 3.734 20.998 3.875 ;
      RECT 20.826 3.734 20.912 3.875 ;
      RECT 20.74 3.735 20.826 3.875 ;
      RECT 20.69 3.732 20.74 3.875 ;
      RECT 20.68 3.73 20.69 3.874 ;
      RECT 20.676 3.73 20.68 3.873 ;
      RECT 20.59 3.725 20.676 3.868 ;
      RECT 20.568 3.718 20.59 3.862 ;
      RECT 20.482 3.709 20.568 3.856 ;
      RECT 20.396 3.696 20.482 3.847 ;
      RECT 20.31 3.682 20.396 3.837 ;
      RECT 20.265 3.672 20.31 3.83 ;
      RECT 20.245 2.96 20.265 3.238 ;
      RECT 20.245 3.665 20.265 3.826 ;
      RECT 20.215 2.96 20.245 3.26 ;
      RECT 20.205 3.632 20.245 3.823 ;
      RECT 20.2 2.96 20.215 3.28 ;
      RECT 20.2 3.597 20.205 3.821 ;
      RECT 20.195 2.96 20.2 3.405 ;
      RECT 20.195 3.557 20.2 3.821 ;
      RECT 20.185 2.96 20.195 3.821 ;
      RECT 20.11 2.96 20.185 3.815 ;
      RECT 20.08 2.96 20.11 3.805 ;
      RECT 20.075 2.96 20.08 3.797 ;
      RECT 20.07 3.002 20.075 3.79 ;
      RECT 20.06 3.071 20.07 3.781 ;
      RECT 20.055 3.141 20.06 3.733 ;
      RECT 20.05 3.205 20.055 3.63 ;
      RECT 20.045 3.24 20.05 3.585 ;
      RECT 20.043 3.277 20.045 3.477 ;
      RECT 20.04 3.285 20.043 3.47 ;
      RECT 20.035 3.35 20.04 3.413 ;
      RECT 24.11 2.44 24.39 2.72 ;
      RECT 24.1 2.44 24.39 2.583 ;
      RECT 24.055 2.305 24.315 2.565 ;
      RECT 24.055 2.42 24.37 2.565 ;
      RECT 24.055 2.39 24.365 2.565 ;
      RECT 24.055 2.377 24.355 2.565 ;
      RECT 24.055 2.367 24.35 2.565 ;
      RECT 20.03 2.35 20.29 2.61 ;
      RECT 23.8 1.9 24.06 2.16 ;
      RECT 23.79 1.925 24.06 2.12 ;
      RECT 23.785 1.925 23.79 2.119 ;
      RECT 23.715 1.92 23.785 2.111 ;
      RECT 23.63 1.907 23.715 2.094 ;
      RECT 23.626 1.899 23.63 2.084 ;
      RECT 23.54 1.892 23.626 2.074 ;
      RECT 23.531 1.884 23.54 2.064 ;
      RECT 23.445 1.877 23.531 2.052 ;
      RECT 23.425 1.868 23.445 2.038 ;
      RECT 23.37 1.863 23.425 2.03 ;
      RECT 23.36 1.857 23.37 2.024 ;
      RECT 23.34 1.855 23.36 2.02 ;
      RECT 23.332 1.854 23.34 2.016 ;
      RECT 23.246 1.846 23.332 2.005 ;
      RECT 23.16 1.832 23.246 1.985 ;
      RECT 23.1 1.82 23.16 1.97 ;
      RECT 23.09 1.815 23.1 1.965 ;
      RECT 23.04 1.815 23.09 1.967 ;
      RECT 22.993 1.817 23.04 1.971 ;
      RECT 22.907 1.824 22.993 1.976 ;
      RECT 22.821 1.832 22.907 1.982 ;
      RECT 22.735 1.841 22.821 1.988 ;
      RECT 22.676 1.847 22.735 1.993 ;
      RECT 22.59 1.852 22.676 1.999 ;
      RECT 22.515 1.857 22.59 2.005 ;
      RECT 22.476 1.859 22.515 2.01 ;
      RECT 22.39 1.856 22.476 2.015 ;
      RECT 22.305 1.854 22.39 2.022 ;
      RECT 22.273 1.853 22.305 2.025 ;
      RECT 22.187 1.852 22.273 2.026 ;
      RECT 22.101 1.851 22.187 2.027 ;
      RECT 22.015 1.85 22.101 2.027 ;
      RECT 21.929 1.849 22.015 2.028 ;
      RECT 21.843 1.848 21.929 2.029 ;
      RECT 21.757 1.847 21.843 2.03 ;
      RECT 21.671 1.846 21.757 2.03 ;
      RECT 21.585 1.845 21.671 2.031 ;
      RECT 21.535 1.845 21.585 2.032 ;
      RECT 21.521 1.846 21.535 2.032 ;
      RECT 21.435 1.853 21.521 2.033 ;
      RECT 21.361 1.864 21.435 2.034 ;
      RECT 21.275 1.873 21.361 2.035 ;
      RECT 21.24 1.88 21.275 2.05 ;
      RECT 21.215 1.883 21.24 2.08 ;
      RECT 21.19 1.892 21.215 2.109 ;
      RECT 21.18 1.903 21.19 2.129 ;
      RECT 21.17 1.911 21.18 2.143 ;
      RECT 21.165 1.917 21.17 2.153 ;
      RECT 21.14 1.934 21.165 2.17 ;
      RECT 21.125 1.956 21.14 2.198 ;
      RECT 21.095 1.982 21.125 2.228 ;
      RECT 21.075 2.011 21.095 2.258 ;
      RECT 21.07 2.026 21.075 2.275 ;
      RECT 21.05 2.041 21.07 2.29 ;
      RECT 21.04 2.059 21.05 2.308 ;
      RECT 21.03 2.07 21.04 2.323 ;
      RECT 20.98 2.102 21.03 2.349 ;
      RECT 20.975 2.132 20.98 2.369 ;
      RECT 20.965 2.145 20.975 2.375 ;
      RECT 20.956 2.155 20.965 2.383 ;
      RECT 20.945 2.166 20.956 2.391 ;
      RECT 20.94 2.176 20.945 2.397 ;
      RECT 20.925 2.197 20.94 2.404 ;
      RECT 20.91 2.227 20.925 2.412 ;
      RECT 20.875 2.257 20.91 2.418 ;
      RECT 20.85 2.275 20.875 2.425 ;
      RECT 20.8 2.283 20.85 2.434 ;
      RECT 20.775 2.288 20.8 2.443 ;
      RECT 20.72 2.294 20.775 2.453 ;
      RECT 20.715 2.299 20.72 2.461 ;
      RECT 20.701 2.302 20.715 2.463 ;
      RECT 20.615 2.314 20.701 2.475 ;
      RECT 20.605 2.326 20.615 2.488 ;
      RECT 20.52 2.339 20.605 2.5 ;
      RECT 20.476 2.356 20.52 2.514 ;
      RECT 20.39 2.373 20.476 2.53 ;
      RECT 20.36 2.387 20.39 2.544 ;
      RECT 20.35 2.392 20.36 2.549 ;
      RECT 20.29 2.395 20.35 2.558 ;
      RECT 23.18 2.665 23.44 2.925 ;
      RECT 23.18 2.665 23.46 2.778 ;
      RECT 23.18 2.665 23.485 2.745 ;
      RECT 23.18 2.665 23.49 2.725 ;
      RECT 23.23 2.44 23.51 2.72 ;
      RECT 22.785 3.175 23.045 3.435 ;
      RECT 22.775 3.032 22.97 3.373 ;
      RECT 22.77 3.14 22.985 3.365 ;
      RECT 22.765 3.19 23.045 3.355 ;
      RECT 22.755 3.267 23.045 3.34 ;
      RECT 22.775 3.115 22.985 3.373 ;
      RECT 22.785 2.99 22.97 3.435 ;
      RECT 22.785 2.885 22.95 3.435 ;
      RECT 22.795 2.872 22.95 3.435 ;
      RECT 22.795 2.83 22.94 3.435 ;
      RECT 22.8 2.755 22.94 3.435 ;
      RECT 22.83 2.405 22.94 3.435 ;
      RECT 22.835 2.135 22.96 2.758 ;
      RECT 22.805 2.71 22.96 2.758 ;
      RECT 22.82 2.512 22.94 3.435 ;
      RECT 22.81 2.622 22.96 2.758 ;
      RECT 22.835 2.135 22.975 2.615 ;
      RECT 22.835 2.135 22.995 2.49 ;
      RECT 22.8 2.135 23.06 2.395 ;
      RECT 22.27 2.44 22.55 2.72 ;
      RECT 22.255 2.44 22.55 2.7 ;
      RECT 20.31 3.305 20.57 3.565 ;
      RECT 22.095 3.16 22.355 3.42 ;
      RECT 22.075 3.18 22.355 3.395 ;
      RECT 22.032 3.18 22.075 3.394 ;
      RECT 21.946 3.181 22.032 3.391 ;
      RECT 21.86 3.182 21.946 3.387 ;
      RECT 21.785 3.184 21.86 3.384 ;
      RECT 21.762 3.185 21.785 3.382 ;
      RECT 21.676 3.186 21.762 3.38 ;
      RECT 21.59 3.187 21.676 3.377 ;
      RECT 21.566 3.188 21.59 3.375 ;
      RECT 21.48 3.19 21.566 3.372 ;
      RECT 21.395 3.192 21.48 3.373 ;
      RECT 21.338 3.193 21.395 3.379 ;
      RECT 21.252 3.195 21.338 3.389 ;
      RECT 21.166 3.198 21.252 3.402 ;
      RECT 21.08 3.2 21.166 3.414 ;
      RECT 21.066 3.201 21.08 3.421 ;
      RECT 20.98 3.202 21.066 3.429 ;
      RECT 20.94 3.204 20.98 3.438 ;
      RECT 20.931 3.205 20.94 3.441 ;
      RECT 20.845 3.213 20.931 3.447 ;
      RECT 20.825 3.222 20.845 3.455 ;
      RECT 20.74 3.237 20.825 3.463 ;
      RECT 20.68 3.26 20.74 3.474 ;
      RECT 20.67 3.272 20.68 3.479 ;
      RECT 20.63 3.282 20.67 3.483 ;
      RECT 20.575 3.299 20.63 3.491 ;
      RECT 20.57 3.309 20.575 3.495 ;
      RECT 21.636 2.44 21.695 2.837 ;
      RECT 21.55 2.44 21.755 2.828 ;
      RECT 21.545 2.47 21.755 2.823 ;
      RECT 21.511 2.47 21.755 2.821 ;
      RECT 21.425 2.47 21.755 2.815 ;
      RECT 21.38 2.47 21.775 2.793 ;
      RECT 21.38 2.47 21.795 2.748 ;
      RECT 21.34 2.47 21.795 2.738 ;
      RECT 21.55 2.44 21.83 2.72 ;
      RECT 21.285 2.44 21.545 2.7 ;
      RECT 19.11 3 19.39 3.28 ;
      RECT 19.08 2.962 19.335 3.265 ;
      RECT 19.075 2.963 19.335 3.263 ;
      RECT 19.07 2.964 19.335 3.257 ;
      RECT 19.065 2.967 19.335 3.25 ;
      RECT 19.06 3 19.39 3.243 ;
      RECT 19.03 2.97 19.335 3.23 ;
      RECT 19.03 2.997 19.355 3.23 ;
      RECT 19.03 2.987 19.35 3.23 ;
      RECT 19.03 2.972 19.345 3.23 ;
      RECT 19.11 2.959 19.325 3.28 ;
      RECT 19.196 2.957 19.325 3.28 ;
      RECT 19.282 2.955 19.31 3.28 ;
      RECT 14.92 6.22 15.24 6.545 ;
      RECT 14.95 5.695 15.12 6.545 ;
      RECT 14.95 5.695 15.125 6.045 ;
      RECT 14.95 5.695 15.925 5.87 ;
      RECT 15.75 1.965 15.925 5.87 ;
      RECT 15.695 1.965 16.045 2.315 ;
      RECT 15.72 6.655 16.045 6.98 ;
      RECT 14.605 6.745 16.045 6.915 ;
      RECT 14.605 2.395 14.765 6.915 ;
      RECT 14.92 2.365 15.24 2.685 ;
      RECT 14.605 2.395 15.24 2.565 ;
      RECT 4.69 1.92 4.95 2.18 ;
      RECT 4.745 1.88 5.05 2.16 ;
      RECT 4.745 1.42 4.92 2.18 ;
      RECT 13.26 1.34 13.61 1.69 ;
      RECT 4.745 1.42 13.61 1.595 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 13.02 2.235 13.19 3.22 ;
      RECT 9.04 2.455 9.275 2.715 ;
      RECT 12.185 2.235 12.35 2.495 ;
      RECT 12.09 2.225 12.105 2.495 ;
      RECT 12.185 2.235 13.19 2.415 ;
      RECT 10.69 1.795 10.73 1.935 ;
      RECT 12.105 2.23 12.185 2.495 ;
      RECT 12.05 2.225 12.09 2.461 ;
      RECT 12.036 2.225 12.05 2.461 ;
      RECT 11.95 2.23 12.036 2.463 ;
      RECT 11.905 2.237 11.95 2.465 ;
      RECT 11.875 2.237 11.905 2.467 ;
      RECT 11.85 2.232 11.875 2.469 ;
      RECT 11.82 2.228 11.85 2.478 ;
      RECT 11.81 2.225 11.82 2.49 ;
      RECT 11.805 2.225 11.81 2.498 ;
      RECT 11.8 2.225 11.805 2.503 ;
      RECT 11.79 2.224 11.8 2.513 ;
      RECT 11.785 2.223 11.79 2.523 ;
      RECT 11.77 2.222 11.785 2.528 ;
      RECT 11.742 2.219 11.77 2.555 ;
      RECT 11.656 2.211 11.742 2.555 ;
      RECT 11.57 2.2 11.656 2.555 ;
      RECT 11.53 2.185 11.57 2.555 ;
      RECT 11.49 2.159 11.53 2.555 ;
      RECT 11.485 2.141 11.49 2.367 ;
      RECT 11.475 2.137 11.485 2.357 ;
      RECT 11.46 2.127 11.475 2.344 ;
      RECT 11.44 2.111 11.46 2.329 ;
      RECT 11.425 2.096 11.44 2.314 ;
      RECT 11.415 2.085 11.425 2.304 ;
      RECT 11.39 2.069 11.415 2.293 ;
      RECT 11.385 2.056 11.39 2.283 ;
      RECT 11.38 2.052 11.385 2.278 ;
      RECT 11.325 2.038 11.38 2.256 ;
      RECT 11.286 2.019 11.325 2.22 ;
      RECT 11.2 1.993 11.286 2.173 ;
      RECT 11.196 1.975 11.2 2.139 ;
      RECT 11.11 1.956 11.196 2.117 ;
      RECT 11.105 1.938 11.11 2.095 ;
      RECT 11.1 1.936 11.105 2.093 ;
      RECT 11.09 1.935 11.1 2.088 ;
      RECT 11.03 1.922 11.09 2.074 ;
      RECT 10.985 1.9 11.03 2.053 ;
      RECT 10.925 1.877 10.985 2.032 ;
      RECT 10.861 1.852 10.925 2.007 ;
      RECT 10.775 1.822 10.861 1.976 ;
      RECT 10.76 1.802 10.775 1.955 ;
      RECT 10.73 1.797 10.76 1.946 ;
      RECT 10.677 1.795 10.69 1.935 ;
      RECT 10.591 1.795 10.677 1.937 ;
      RECT 10.505 1.795 10.591 1.939 ;
      RECT 10.485 1.795 10.505 1.943 ;
      RECT 10.44 1.797 10.485 1.954 ;
      RECT 10.4 1.807 10.44 1.97 ;
      RECT 10.396 1.816 10.4 1.978 ;
      RECT 10.31 1.836 10.396 1.994 ;
      RECT 10.3 1.855 10.31 2.012 ;
      RECT 10.295 1.857 10.3 2.015 ;
      RECT 10.285 1.861 10.295 2.018 ;
      RECT 10.265 1.866 10.285 2.028 ;
      RECT 10.235 1.876 10.265 2.048 ;
      RECT 10.23 1.883 10.235 2.062 ;
      RECT 10.22 1.887 10.23 2.069 ;
      RECT 10.205 1.895 10.22 2.08 ;
      RECT 10.195 1.905 10.205 2.091 ;
      RECT 10.185 1.912 10.195 2.099 ;
      RECT 10.16 1.925 10.185 2.114 ;
      RECT 10.096 1.961 10.16 2.153 ;
      RECT 10.01 2.024 10.096 2.217 ;
      RECT 9.975 2.075 10.01 2.27 ;
      RECT 9.97 2.092 9.975 2.287 ;
      RECT 9.955 2.101 9.97 2.294 ;
      RECT 9.935 2.116 9.955 2.308 ;
      RECT 9.93 2.127 9.935 2.318 ;
      RECT 9.91 2.14 9.93 2.328 ;
      RECT 9.905 2.15 9.91 2.338 ;
      RECT 9.89 2.155 9.905 2.347 ;
      RECT 9.88 2.165 9.89 2.358 ;
      RECT 9.85 2.182 9.88 2.375 ;
      RECT 9.84 2.2 9.85 2.393 ;
      RECT 9.825 2.211 9.84 2.404 ;
      RECT 9.785 2.235 9.825 2.42 ;
      RECT 9.75 2.269 9.785 2.437 ;
      RECT 9.72 2.292 9.75 2.449 ;
      RECT 9.705 2.302 9.72 2.458 ;
      RECT 9.665 2.312 9.705 2.469 ;
      RECT 9.645 2.323 9.665 2.481 ;
      RECT 9.64 2.327 9.645 2.488 ;
      RECT 9.625 2.331 9.64 2.493 ;
      RECT 9.615 2.336 9.625 2.498 ;
      RECT 9.61 2.339 9.615 2.501 ;
      RECT 9.58 2.345 9.61 2.508 ;
      RECT 9.545 2.355 9.58 2.522 ;
      RECT 9.485 2.37 9.545 2.542 ;
      RECT 9.43 2.39 9.485 2.566 ;
      RECT 9.401 2.405 9.43 2.584 ;
      RECT 9.315 2.425 9.401 2.609 ;
      RECT 9.31 2.44 9.315 2.629 ;
      RECT 9.3 2.443 9.31 2.63 ;
      RECT 9.275 2.45 9.3 2.715 ;
      RECT 11.97 2.943 12.25 3.28 ;
      RECT 11.97 2.953 12.255 3.238 ;
      RECT 11.97 2.962 12.26 3.135 ;
      RECT 11.97 2.977 12.265 3.003 ;
      RECT 11.97 2.805 12.23 3.28 ;
      RECT 1.55 6.995 1.84 7.345 ;
      RECT 1.55 7.085 2.955 7.255 ;
      RECT 2.785 6.685 2.955 7.255 ;
      RECT 11.115 6.605 11.465 6.955 ;
      RECT 2.785 6.685 11.465 6.855 ;
      RECT 9.69 3.685 9.7 3.875 ;
      RECT 7.95 3.56 8.23 3.84 ;
      RECT 10.995 2.5 11 2.985 ;
      RECT 10.89 2.5 10.95 2.76 ;
      RECT 11.215 3.47 11.22 3.545 ;
      RECT 11.205 3.337 11.215 3.58 ;
      RECT 11.195 3.172 11.205 3.601 ;
      RECT 11.19 3.042 11.195 3.617 ;
      RECT 11.18 2.932 11.19 3.633 ;
      RECT 11.175 2.831 11.18 3.65 ;
      RECT 11.17 2.813 11.175 3.66 ;
      RECT 11.165 2.795 11.17 3.67 ;
      RECT 11.155 2.77 11.165 3.685 ;
      RECT 11.15 2.75 11.155 3.7 ;
      RECT 11.13 2.5 11.15 3.725 ;
      RECT 11.115 2.5 11.13 3.758 ;
      RECT 11.085 2.5 11.115 3.78 ;
      RECT 11.065 2.5 11.085 3.794 ;
      RECT 11.045 2.5 11.065 3.31 ;
      RECT 11.06 3.377 11.065 3.799 ;
      RECT 11.055 3.407 11.06 3.801 ;
      RECT 11.05 3.42 11.055 3.804 ;
      RECT 11.045 3.43 11.05 3.808 ;
      RECT 11.04 2.5 11.045 3.228 ;
      RECT 11.04 3.44 11.045 3.81 ;
      RECT 11.035 2.5 11.04 3.205 ;
      RECT 11.025 3.462 11.04 3.81 ;
      RECT 11.02 2.5 11.035 3.15 ;
      RECT 11.015 3.487 11.025 3.81 ;
      RECT 11.015 2.5 11.02 3.095 ;
      RECT 11.005 2.5 11.015 3.043 ;
      RECT 11.01 3.5 11.015 3.811 ;
      RECT 11.005 3.512 11.01 3.812 ;
      RECT 11 2.5 11.005 3.003 ;
      RECT 11 3.525 11.005 3.813 ;
      RECT 10.985 3.54 11 3.814 ;
      RECT 10.99 2.5 10.995 2.965 ;
      RECT 10.985 2.5 10.99 2.93 ;
      RECT 10.98 2.5 10.985 2.905 ;
      RECT 10.975 3.567 10.985 3.816 ;
      RECT 10.97 2.5 10.98 2.863 ;
      RECT 10.97 3.585 10.975 3.817 ;
      RECT 10.965 2.5 10.97 2.823 ;
      RECT 10.965 3.592 10.97 3.818 ;
      RECT 10.96 2.5 10.965 2.795 ;
      RECT 10.955 3.61 10.965 3.819 ;
      RECT 10.95 2.5 10.96 2.775 ;
      RECT 10.945 3.63 10.955 3.821 ;
      RECT 10.935 3.647 10.945 3.822 ;
      RECT 10.9 3.67 10.935 3.825 ;
      RECT 10.845 3.688 10.9 3.831 ;
      RECT 10.759 3.696 10.845 3.84 ;
      RECT 10.673 3.707 10.759 3.851 ;
      RECT 10.587 3.717 10.673 3.862 ;
      RECT 10.501 3.727 10.587 3.874 ;
      RECT 10.415 3.737 10.501 3.885 ;
      RECT 10.395 3.743 10.415 3.891 ;
      RECT 10.315 3.745 10.395 3.895 ;
      RECT 10.31 3.744 10.315 3.9 ;
      RECT 10.302 3.743 10.31 3.9 ;
      RECT 10.216 3.739 10.302 3.898 ;
      RECT 10.13 3.731 10.216 3.895 ;
      RECT 10.044 3.722 10.13 3.891 ;
      RECT 9.958 3.714 10.044 3.888 ;
      RECT 9.872 3.706 9.958 3.884 ;
      RECT 9.786 3.697 9.872 3.881 ;
      RECT 9.7 3.689 9.786 3.877 ;
      RECT 9.645 3.682 9.69 3.875 ;
      RECT 9.56 3.675 9.645 3.873 ;
      RECT 9.486 3.667 9.56 3.869 ;
      RECT 9.4 3.659 9.486 3.866 ;
      RECT 9.397 3.655 9.4 3.864 ;
      RECT 9.311 3.651 9.397 3.863 ;
      RECT 9.225 3.643 9.311 3.86 ;
      RECT 9.14 3.638 9.225 3.857 ;
      RECT 9.054 3.635 9.14 3.854 ;
      RECT 8.968 3.633 9.054 3.851 ;
      RECT 8.882 3.63 8.968 3.848 ;
      RECT 8.796 3.627 8.882 3.845 ;
      RECT 8.71 3.624 8.796 3.842 ;
      RECT 8.634 3.622 8.71 3.839 ;
      RECT 8.548 3.619 8.634 3.836 ;
      RECT 8.462 3.616 8.548 3.834 ;
      RECT 8.376 3.614 8.462 3.831 ;
      RECT 8.29 3.611 8.376 3.828 ;
      RECT 8.23 3.602 8.29 3.826 ;
      RECT 10.74 3.22 10.815 3.48 ;
      RECT 10.72 3.2 10.725 3.48 ;
      RECT 10.04 2.985 10.145 3.28 ;
      RECT 4.485 2.96 4.555 3.22 ;
      RECT 10.38 2.835 10.385 3.206 ;
      RECT 10.37 2.89 10.375 3.206 ;
      RECT 10.675 2.06 10.735 2.32 ;
      RECT 10.73 3.215 10.74 3.48 ;
      RECT 10.725 3.205 10.73 3.48 ;
      RECT 10.645 3.152 10.72 3.48 ;
      RECT 10.67 2.06 10.675 2.34 ;
      RECT 10.66 2.06 10.67 2.36 ;
      RECT 10.645 2.06 10.66 2.39 ;
      RECT 10.63 2.06 10.645 2.433 ;
      RECT 10.625 3.095 10.645 3.48 ;
      RECT 10.615 2.06 10.63 2.47 ;
      RECT 10.61 3.075 10.625 3.48 ;
      RECT 10.61 2.06 10.615 2.493 ;
      RECT 10.6 2.06 10.61 2.518 ;
      RECT 10.57 3.042 10.61 3.48 ;
      RECT 10.575 2.06 10.6 2.568 ;
      RECT 10.57 2.06 10.575 2.623 ;
      RECT 10.565 2.06 10.57 2.665 ;
      RECT 10.555 3.005 10.57 3.48 ;
      RECT 10.56 2.06 10.565 2.708 ;
      RECT 10.555 2.06 10.56 2.773 ;
      RECT 10.55 2.06 10.555 2.795 ;
      RECT 10.55 2.993 10.555 3.345 ;
      RECT 10.545 2.06 10.55 2.863 ;
      RECT 10.545 2.985 10.55 3.328 ;
      RECT 10.54 2.06 10.545 2.908 ;
      RECT 10.535 2.967 10.545 3.305 ;
      RECT 10.535 2.06 10.54 2.945 ;
      RECT 10.525 2.06 10.535 3.285 ;
      RECT 10.52 2.06 10.525 3.268 ;
      RECT 10.515 2.06 10.52 3.253 ;
      RECT 10.51 2.06 10.515 3.238 ;
      RECT 10.49 2.06 10.51 3.228 ;
      RECT 10.485 2.06 10.49 3.218 ;
      RECT 10.475 2.06 10.485 3.214 ;
      RECT 10.47 2.337 10.475 3.213 ;
      RECT 10.465 2.36 10.47 3.212 ;
      RECT 10.46 2.39 10.465 3.211 ;
      RECT 10.455 2.417 10.46 3.21 ;
      RECT 10.45 2.445 10.455 3.21 ;
      RECT 10.445 2.472 10.45 3.21 ;
      RECT 10.44 2.492 10.445 3.21 ;
      RECT 10.435 2.52 10.44 3.21 ;
      RECT 10.425 2.562 10.435 3.21 ;
      RECT 10.415 2.607 10.425 3.209 ;
      RECT 10.41 2.66 10.415 3.208 ;
      RECT 10.405 2.692 10.41 3.207 ;
      RECT 10.4 2.712 10.405 3.206 ;
      RECT 10.395 2.75 10.4 3.206 ;
      RECT 10.39 2.772 10.395 3.206 ;
      RECT 10.385 2.797 10.39 3.206 ;
      RECT 10.375 2.862 10.38 3.206 ;
      RECT 10.36 2.922 10.37 3.206 ;
      RECT 10.345 2.932 10.36 3.206 ;
      RECT 10.325 2.942 10.345 3.206 ;
      RECT 10.295 2.947 10.325 3.203 ;
      RECT 10.235 2.957 10.295 3.2 ;
      RECT 10.215 2.966 10.235 3.205 ;
      RECT 10.19 2.972 10.215 3.218 ;
      RECT 10.17 2.977 10.19 3.233 ;
      RECT 10.145 2.982 10.17 3.28 ;
      RECT 10.016 2.984 10.04 3.28 ;
      RECT 9.93 2.979 10.016 3.28 ;
      RECT 9.89 2.976 9.93 3.28 ;
      RECT 9.84 2.978 9.89 3.26 ;
      RECT 9.81 2.982 9.84 3.26 ;
      RECT 9.731 2.992 9.81 3.26 ;
      RECT 9.645 3.007 9.731 3.261 ;
      RECT 9.595 3.017 9.645 3.262 ;
      RECT 9.587 3.02 9.595 3.262 ;
      RECT 9.501 3.022 9.587 3.263 ;
      RECT 9.415 3.026 9.501 3.263 ;
      RECT 9.329 3.03 9.415 3.264 ;
      RECT 9.243 3.033 9.329 3.265 ;
      RECT 9.157 3.037 9.243 3.265 ;
      RECT 9.071 3.041 9.157 3.266 ;
      RECT 8.985 3.044 9.071 3.267 ;
      RECT 8.899 3.048 8.985 3.267 ;
      RECT 8.813 3.052 8.899 3.268 ;
      RECT 8.727 3.056 8.813 3.269 ;
      RECT 8.641 3.059 8.727 3.269 ;
      RECT 8.555 3.063 8.641 3.27 ;
      RECT 8.525 3.065 8.555 3.27 ;
      RECT 8.439 3.068 8.525 3.271 ;
      RECT 8.353 3.072 8.439 3.272 ;
      RECT 8.267 3.076 8.353 3.273 ;
      RECT 8.181 3.079 8.267 3.273 ;
      RECT 8.095 3.083 8.181 3.274 ;
      RECT 8.06 3.088 8.095 3.275 ;
      RECT 8.005 3.098 8.06 3.282 ;
      RECT 7.98 3.11 8.005 3.292 ;
      RECT 7.945 3.123 7.98 3.3 ;
      RECT 7.905 3.14 7.945 3.323 ;
      RECT 7.885 3.153 7.905 3.35 ;
      RECT 7.855 3.165 7.885 3.378 ;
      RECT 7.85 3.173 7.855 3.398 ;
      RECT 7.845 3.176 7.85 3.408 ;
      RECT 7.795 3.188 7.845 3.442 ;
      RECT 7.785 3.203 7.795 3.475 ;
      RECT 7.775 3.209 7.785 3.488 ;
      RECT 7.765 3.216 7.775 3.5 ;
      RECT 7.74 3.229 7.765 3.518 ;
      RECT 7.725 3.244 7.74 3.54 ;
      RECT 7.715 3.252 7.725 3.556 ;
      RECT 7.7 3.261 7.715 3.571 ;
      RECT 7.69 3.271 7.7 3.585 ;
      RECT 7.671 3.284 7.69 3.602 ;
      RECT 7.585 3.329 7.671 3.667 ;
      RECT 7.57 3.374 7.585 3.725 ;
      RECT 7.565 3.383 7.57 3.738 ;
      RECT 7.555 3.39 7.565 3.743 ;
      RECT 7.55 3.395 7.555 3.747 ;
      RECT 7.53 3.405 7.55 3.754 ;
      RECT 7.505 3.425 7.53 3.768 ;
      RECT 7.47 3.45 7.505 3.788 ;
      RECT 7.455 3.473 7.47 3.803 ;
      RECT 7.445 3.483 7.455 3.808 ;
      RECT 7.435 3.491 7.445 3.815 ;
      RECT 7.425 3.5 7.435 3.821 ;
      RECT 7.405 3.512 7.425 3.823 ;
      RECT 7.395 3.525 7.405 3.825 ;
      RECT 7.37 3.54 7.395 3.828 ;
      RECT 7.35 3.557 7.37 3.832 ;
      RECT 7.31 3.585 7.35 3.838 ;
      RECT 7.245 3.632 7.31 3.847 ;
      RECT 7.23 3.665 7.245 3.855 ;
      RECT 7.225 3.672 7.23 3.857 ;
      RECT 7.175 3.697 7.225 3.862 ;
      RECT 7.16 3.721 7.175 3.869 ;
      RECT 7.11 3.726 7.16 3.87 ;
      RECT 7.024 3.73 7.11 3.87 ;
      RECT 6.938 3.73 7.024 3.87 ;
      RECT 6.852 3.73 6.938 3.871 ;
      RECT 6.766 3.73 6.852 3.871 ;
      RECT 6.68 3.73 6.766 3.871 ;
      RECT 6.614 3.73 6.68 3.871 ;
      RECT 6.528 3.73 6.614 3.872 ;
      RECT 6.442 3.73 6.528 3.872 ;
      RECT 6.356 3.731 6.442 3.873 ;
      RECT 6.27 3.731 6.356 3.873 ;
      RECT 6.184 3.731 6.27 3.873 ;
      RECT 6.098 3.731 6.184 3.874 ;
      RECT 6.012 3.731 6.098 3.874 ;
      RECT 5.926 3.732 6.012 3.875 ;
      RECT 5.84 3.732 5.926 3.875 ;
      RECT 5.82 3.732 5.84 3.875 ;
      RECT 5.734 3.732 5.82 3.875 ;
      RECT 5.648 3.732 5.734 3.875 ;
      RECT 5.562 3.733 5.648 3.875 ;
      RECT 5.476 3.733 5.562 3.875 ;
      RECT 5.39 3.733 5.476 3.875 ;
      RECT 5.304 3.734 5.39 3.875 ;
      RECT 5.218 3.734 5.304 3.875 ;
      RECT 5.132 3.734 5.218 3.875 ;
      RECT 5.046 3.734 5.132 3.875 ;
      RECT 4.96 3.735 5.046 3.875 ;
      RECT 4.91 3.732 4.96 3.875 ;
      RECT 4.9 3.73 4.91 3.874 ;
      RECT 4.896 3.73 4.9 3.873 ;
      RECT 4.81 3.725 4.896 3.868 ;
      RECT 4.788 3.718 4.81 3.862 ;
      RECT 4.702 3.709 4.788 3.856 ;
      RECT 4.616 3.696 4.702 3.847 ;
      RECT 4.53 3.682 4.616 3.837 ;
      RECT 4.485 3.672 4.53 3.83 ;
      RECT 4.465 2.96 4.485 3.238 ;
      RECT 4.465 3.665 4.485 3.826 ;
      RECT 4.435 2.96 4.465 3.26 ;
      RECT 4.425 3.632 4.465 3.823 ;
      RECT 4.42 2.96 4.435 3.28 ;
      RECT 4.42 3.597 4.425 3.821 ;
      RECT 4.415 2.96 4.42 3.405 ;
      RECT 4.415 3.557 4.42 3.821 ;
      RECT 4.405 2.96 4.415 3.821 ;
      RECT 4.33 2.96 4.405 3.815 ;
      RECT 4.3 2.96 4.33 3.805 ;
      RECT 4.295 2.96 4.3 3.797 ;
      RECT 4.29 3.002 4.295 3.79 ;
      RECT 4.28 3.071 4.29 3.781 ;
      RECT 4.275 3.141 4.28 3.733 ;
      RECT 4.27 3.205 4.275 3.63 ;
      RECT 4.265 3.24 4.27 3.585 ;
      RECT 4.263 3.277 4.265 3.477 ;
      RECT 4.26 3.285 4.263 3.47 ;
      RECT 4.255 3.35 4.26 3.413 ;
      RECT 8.33 2.44 8.61 2.72 ;
      RECT 8.32 2.44 8.61 2.583 ;
      RECT 8.275 2.305 8.535 2.565 ;
      RECT 8.275 2.42 8.59 2.565 ;
      RECT 8.275 2.39 8.585 2.565 ;
      RECT 8.275 2.377 8.575 2.565 ;
      RECT 8.275 2.367 8.57 2.565 ;
      RECT 4.25 2.35 4.51 2.61 ;
      RECT 8.02 1.9 8.28 2.16 ;
      RECT 8.01 1.925 8.28 2.12 ;
      RECT 8.005 1.925 8.01 2.119 ;
      RECT 7.935 1.92 8.005 2.111 ;
      RECT 7.85 1.907 7.935 2.094 ;
      RECT 7.846 1.899 7.85 2.084 ;
      RECT 7.76 1.892 7.846 2.074 ;
      RECT 7.751 1.884 7.76 2.064 ;
      RECT 7.665 1.877 7.751 2.052 ;
      RECT 7.645 1.868 7.665 2.038 ;
      RECT 7.59 1.863 7.645 2.03 ;
      RECT 7.58 1.857 7.59 2.024 ;
      RECT 7.56 1.855 7.58 2.02 ;
      RECT 7.552 1.854 7.56 2.016 ;
      RECT 7.466 1.846 7.552 2.005 ;
      RECT 7.38 1.832 7.466 1.985 ;
      RECT 7.32 1.82 7.38 1.97 ;
      RECT 7.31 1.815 7.32 1.965 ;
      RECT 7.26 1.815 7.31 1.967 ;
      RECT 7.213 1.817 7.26 1.971 ;
      RECT 7.127 1.824 7.213 1.976 ;
      RECT 7.041 1.832 7.127 1.982 ;
      RECT 6.955 1.841 7.041 1.988 ;
      RECT 6.896 1.847 6.955 1.993 ;
      RECT 6.81 1.852 6.896 1.999 ;
      RECT 6.735 1.857 6.81 2.005 ;
      RECT 6.696 1.859 6.735 2.01 ;
      RECT 6.61 1.856 6.696 2.015 ;
      RECT 6.525 1.854 6.61 2.022 ;
      RECT 6.493 1.853 6.525 2.025 ;
      RECT 6.407 1.852 6.493 2.026 ;
      RECT 6.321 1.851 6.407 2.027 ;
      RECT 6.235 1.85 6.321 2.027 ;
      RECT 6.149 1.849 6.235 2.028 ;
      RECT 6.063 1.848 6.149 2.029 ;
      RECT 5.977 1.847 6.063 2.03 ;
      RECT 5.891 1.846 5.977 2.03 ;
      RECT 5.805 1.845 5.891 2.031 ;
      RECT 5.755 1.845 5.805 2.032 ;
      RECT 5.741 1.846 5.755 2.032 ;
      RECT 5.655 1.853 5.741 2.033 ;
      RECT 5.581 1.864 5.655 2.034 ;
      RECT 5.495 1.873 5.581 2.035 ;
      RECT 5.46 1.88 5.495 2.05 ;
      RECT 5.435 1.883 5.46 2.08 ;
      RECT 5.41 1.892 5.435 2.109 ;
      RECT 5.4 1.903 5.41 2.129 ;
      RECT 5.39 1.911 5.4 2.143 ;
      RECT 5.385 1.917 5.39 2.153 ;
      RECT 5.36 1.934 5.385 2.17 ;
      RECT 5.345 1.956 5.36 2.198 ;
      RECT 5.315 1.982 5.345 2.228 ;
      RECT 5.295 2.011 5.315 2.258 ;
      RECT 5.29 2.026 5.295 2.275 ;
      RECT 5.27 2.041 5.29 2.29 ;
      RECT 5.26 2.059 5.27 2.308 ;
      RECT 5.25 2.07 5.26 2.323 ;
      RECT 5.2 2.102 5.25 2.349 ;
      RECT 5.195 2.132 5.2 2.369 ;
      RECT 5.185 2.145 5.195 2.375 ;
      RECT 5.176 2.155 5.185 2.383 ;
      RECT 5.165 2.166 5.176 2.391 ;
      RECT 5.16 2.176 5.165 2.397 ;
      RECT 5.145 2.197 5.16 2.404 ;
      RECT 5.13 2.227 5.145 2.412 ;
      RECT 5.095 2.257 5.13 2.418 ;
      RECT 5.07 2.275 5.095 2.425 ;
      RECT 5.02 2.283 5.07 2.434 ;
      RECT 4.995 2.288 5.02 2.443 ;
      RECT 4.94 2.294 4.995 2.453 ;
      RECT 4.935 2.299 4.94 2.461 ;
      RECT 4.921 2.302 4.935 2.463 ;
      RECT 4.835 2.314 4.921 2.475 ;
      RECT 4.825 2.326 4.835 2.488 ;
      RECT 4.74 2.339 4.825 2.5 ;
      RECT 4.696 2.356 4.74 2.514 ;
      RECT 4.61 2.373 4.696 2.53 ;
      RECT 4.58 2.387 4.61 2.544 ;
      RECT 4.57 2.392 4.58 2.549 ;
      RECT 4.51 2.395 4.57 2.558 ;
      RECT 7.4 2.665 7.66 2.925 ;
      RECT 7.4 2.665 7.68 2.778 ;
      RECT 7.4 2.665 7.705 2.745 ;
      RECT 7.4 2.665 7.71 2.725 ;
      RECT 7.45 2.44 7.73 2.72 ;
      RECT 7.005 3.175 7.265 3.435 ;
      RECT 6.995 3.032 7.19 3.373 ;
      RECT 6.99 3.14 7.205 3.365 ;
      RECT 6.985 3.19 7.265 3.355 ;
      RECT 6.975 3.267 7.265 3.34 ;
      RECT 6.995 3.115 7.205 3.373 ;
      RECT 7.005 2.99 7.19 3.435 ;
      RECT 7.005 2.885 7.17 3.435 ;
      RECT 7.015 2.872 7.17 3.435 ;
      RECT 7.015 2.83 7.16 3.435 ;
      RECT 7.02 2.755 7.16 3.435 ;
      RECT 7.05 2.405 7.16 3.435 ;
      RECT 7.055 2.135 7.18 2.758 ;
      RECT 7.025 2.71 7.18 2.758 ;
      RECT 7.04 2.512 7.16 3.435 ;
      RECT 7.03 2.622 7.18 2.758 ;
      RECT 7.055 2.135 7.195 2.615 ;
      RECT 7.055 2.135 7.215 2.49 ;
      RECT 7.02 2.135 7.28 2.395 ;
      RECT 6.49 2.44 6.77 2.72 ;
      RECT 6.475 2.44 6.77 2.7 ;
      RECT 4.53 3.305 4.79 3.565 ;
      RECT 6.315 3.16 6.575 3.42 ;
      RECT 6.295 3.18 6.575 3.395 ;
      RECT 6.252 3.18 6.295 3.394 ;
      RECT 6.166 3.181 6.252 3.391 ;
      RECT 6.08 3.182 6.166 3.387 ;
      RECT 6.005 3.184 6.08 3.384 ;
      RECT 5.982 3.185 6.005 3.382 ;
      RECT 5.896 3.186 5.982 3.38 ;
      RECT 5.81 3.187 5.896 3.377 ;
      RECT 5.786 3.188 5.81 3.375 ;
      RECT 5.7 3.19 5.786 3.372 ;
      RECT 5.615 3.192 5.7 3.373 ;
      RECT 5.558 3.193 5.615 3.379 ;
      RECT 5.472 3.195 5.558 3.389 ;
      RECT 5.386 3.198 5.472 3.402 ;
      RECT 5.3 3.2 5.386 3.414 ;
      RECT 5.286 3.201 5.3 3.421 ;
      RECT 5.2 3.202 5.286 3.429 ;
      RECT 5.16 3.204 5.2 3.438 ;
      RECT 5.151 3.205 5.16 3.441 ;
      RECT 5.065 3.213 5.151 3.447 ;
      RECT 5.045 3.222 5.065 3.455 ;
      RECT 4.96 3.237 5.045 3.463 ;
      RECT 4.9 3.26 4.96 3.474 ;
      RECT 4.89 3.272 4.9 3.479 ;
      RECT 4.85 3.282 4.89 3.483 ;
      RECT 4.795 3.299 4.85 3.491 ;
      RECT 4.79 3.309 4.795 3.495 ;
      RECT 5.856 2.44 5.915 2.837 ;
      RECT 5.77 2.44 5.975 2.828 ;
      RECT 5.765 2.47 5.975 2.823 ;
      RECT 5.731 2.47 5.975 2.821 ;
      RECT 5.645 2.47 5.975 2.815 ;
      RECT 5.6 2.47 5.995 2.793 ;
      RECT 5.6 2.47 6.015 2.748 ;
      RECT 5.56 2.47 6.015 2.738 ;
      RECT 5.77 2.44 6.05 2.72 ;
      RECT 5.505 2.44 5.765 2.7 ;
      RECT 3.33 3 3.61 3.28 ;
      RECT 3.3 2.962 3.555 3.265 ;
      RECT 3.295 2.963 3.555 3.263 ;
      RECT 3.29 2.964 3.555 3.257 ;
      RECT 3.285 2.967 3.555 3.25 ;
      RECT 3.28 3 3.61 3.243 ;
      RECT 3.25 2.97 3.555 3.23 ;
      RECT 3.25 2.997 3.575 3.23 ;
      RECT 3.25 2.987 3.57 3.23 ;
      RECT 3.25 2.972 3.565 3.23 ;
      RECT 3.33 2.959 3.545 3.28 ;
      RECT 3.416 2.957 3.545 3.28 ;
      RECT 3.502 2.955 3.53 3.28 ;
      RECT 75.28 0.815 75.65 1.185 ;
      RECT 73.57 7.04 73.94 7.41 ;
      RECT 59.495 0.815 59.865 1.185 ;
      RECT 57.785 7.04 58.155 7.41 ;
      RECT 43.71 0.815 44.08 1.185 ;
      RECT 42 7.04 42.37 7.41 ;
      RECT 27.935 0.815 28.305 1.185 ;
      RECT 26.225 7.04 26.595 7.41 ;
      RECT 12.155 0.815 12.525 1.185 ;
      RECT 10.445 7.04 10.815 7.41 ;
    LAYER via1 ;
      RECT 81.305 7.375 81.455 7.525 ;
      RECT 78.935 6.74 79.085 6.89 ;
      RECT 78.92 2.065 79.07 2.215 ;
      RECT 78.13 2.45 78.28 2.6 ;
      RECT 78.13 6.325 78.28 6.475 ;
      RECT 76.485 1.44 76.635 1.59 ;
      RECT 76.17 2.96 76.32 3.11 ;
      RECT 75.39 0.925 75.54 1.075 ;
      RECT 75.27 2.29 75.42 2.44 ;
      RECT 75.15 2.86 75.3 3.01 ;
      RECT 74.32 6.71 74.47 6.86 ;
      RECT 74.07 2.555 74.22 2.705 ;
      RECT 73.735 3.275 73.885 3.425 ;
      RECT 73.68 7.15 73.83 7.3 ;
      RECT 73.655 2.115 73.805 2.265 ;
      RECT 72.22 2.51 72.37 2.66 ;
      RECT 71.455 2.36 71.605 2.51 ;
      RECT 71.2 1.955 71.35 2.105 ;
      RECT 70.58 2.72 70.73 2.87 ;
      RECT 70.2 2.19 70.35 2.34 ;
      RECT 70.185 3.23 70.335 3.38 ;
      RECT 69.655 2.495 69.805 2.645 ;
      RECT 69.495 3.215 69.645 3.365 ;
      RECT 68.685 2.495 68.835 2.645 ;
      RECT 67.87 1.975 68.02 2.125 ;
      RECT 67.71 3.36 67.86 3.51 ;
      RECT 67.475 3.015 67.625 3.165 ;
      RECT 67.43 2.405 67.58 2.555 ;
      RECT 66.43 3.025 66.58 3.175 ;
      RECT 65.495 6.755 65.645 6.905 ;
      RECT 63.15 6.74 63.3 6.89 ;
      RECT 63.135 2.065 63.285 2.215 ;
      RECT 62.345 2.45 62.495 2.6 ;
      RECT 62.345 6.325 62.495 6.475 ;
      RECT 60.7 1.44 60.85 1.59 ;
      RECT 60.385 2.96 60.535 3.11 ;
      RECT 59.605 0.925 59.755 1.075 ;
      RECT 59.485 2.29 59.635 2.44 ;
      RECT 59.365 2.86 59.515 3.01 ;
      RECT 58.535 6.71 58.685 6.86 ;
      RECT 58.285 2.555 58.435 2.705 ;
      RECT 57.95 3.275 58.1 3.425 ;
      RECT 57.895 7.15 58.045 7.3 ;
      RECT 57.87 2.115 58.02 2.265 ;
      RECT 56.435 2.51 56.585 2.66 ;
      RECT 55.67 2.36 55.82 2.51 ;
      RECT 55.415 1.955 55.565 2.105 ;
      RECT 54.795 2.72 54.945 2.87 ;
      RECT 54.415 2.19 54.565 2.34 ;
      RECT 54.4 3.23 54.55 3.38 ;
      RECT 53.87 2.495 54.02 2.645 ;
      RECT 53.71 3.215 53.86 3.365 ;
      RECT 52.9 2.495 53.05 2.645 ;
      RECT 52.085 1.975 52.235 2.125 ;
      RECT 51.925 3.36 52.075 3.51 ;
      RECT 51.69 3.015 51.84 3.165 ;
      RECT 51.645 2.405 51.795 2.555 ;
      RECT 50.645 3.025 50.795 3.175 ;
      RECT 49.71 6.755 49.86 6.905 ;
      RECT 47.365 6.74 47.515 6.89 ;
      RECT 47.35 2.065 47.5 2.215 ;
      RECT 46.56 2.45 46.71 2.6 ;
      RECT 46.56 6.325 46.71 6.475 ;
      RECT 44.915 1.44 45.065 1.59 ;
      RECT 44.6 2.96 44.75 3.11 ;
      RECT 43.82 0.925 43.97 1.075 ;
      RECT 43.7 2.29 43.85 2.44 ;
      RECT 43.58 2.86 43.73 3.01 ;
      RECT 42.805 6.715 42.955 6.865 ;
      RECT 42.5 2.555 42.65 2.705 ;
      RECT 42.165 3.275 42.315 3.425 ;
      RECT 42.11 7.15 42.26 7.3 ;
      RECT 42.085 2.115 42.235 2.265 ;
      RECT 40.65 2.51 40.8 2.66 ;
      RECT 39.885 2.36 40.035 2.51 ;
      RECT 39.63 1.955 39.78 2.105 ;
      RECT 39.01 2.72 39.16 2.87 ;
      RECT 38.63 2.19 38.78 2.34 ;
      RECT 38.615 3.23 38.765 3.38 ;
      RECT 38.085 2.495 38.235 2.645 ;
      RECT 37.925 3.215 38.075 3.365 ;
      RECT 37.115 2.495 37.265 2.645 ;
      RECT 36.3 1.975 36.45 2.125 ;
      RECT 36.14 3.36 36.29 3.51 ;
      RECT 35.905 3.015 36.055 3.165 ;
      RECT 35.86 2.405 36.01 2.555 ;
      RECT 34.86 3.025 35.01 3.175 ;
      RECT 33.98 6.76 34.13 6.91 ;
      RECT 31.59 6.74 31.74 6.89 ;
      RECT 31.575 2.065 31.725 2.215 ;
      RECT 30.785 2.45 30.935 2.6 ;
      RECT 30.785 6.325 30.935 6.475 ;
      RECT 29.14 1.44 29.29 1.59 ;
      RECT 28.825 2.96 28.975 3.11 ;
      RECT 28.045 0.925 28.195 1.075 ;
      RECT 27.925 2.29 28.075 2.44 ;
      RECT 27.805 2.86 27.955 3.01 ;
      RECT 27.025 6.71 27.175 6.86 ;
      RECT 26.725 2.555 26.875 2.705 ;
      RECT 26.39 3.275 26.54 3.425 ;
      RECT 26.335 7.15 26.485 7.3 ;
      RECT 26.31 2.115 26.46 2.265 ;
      RECT 24.875 2.51 25.025 2.66 ;
      RECT 24.11 2.36 24.26 2.51 ;
      RECT 23.855 1.955 24.005 2.105 ;
      RECT 23.235 2.72 23.385 2.87 ;
      RECT 22.855 2.19 23.005 2.34 ;
      RECT 22.84 3.23 22.99 3.38 ;
      RECT 22.31 2.495 22.46 2.645 ;
      RECT 22.15 3.215 22.3 3.365 ;
      RECT 21.34 2.495 21.49 2.645 ;
      RECT 20.525 1.975 20.675 2.125 ;
      RECT 20.365 3.36 20.515 3.51 ;
      RECT 20.13 3.015 20.28 3.165 ;
      RECT 20.085 2.405 20.235 2.555 ;
      RECT 19.085 3.025 19.235 3.175 ;
      RECT 18.2 6.755 18.35 6.905 ;
      RECT 15.81 6.74 15.96 6.89 ;
      RECT 15.795 2.065 15.945 2.215 ;
      RECT 15.005 2.45 15.155 2.6 ;
      RECT 15.005 6.325 15.155 6.475 ;
      RECT 13.36 1.44 13.51 1.59 ;
      RECT 13.045 2.96 13.195 3.11 ;
      RECT 12.265 0.925 12.415 1.075 ;
      RECT 12.145 2.29 12.295 2.44 ;
      RECT 12.025 2.86 12.175 3.01 ;
      RECT 11.215 6.705 11.365 6.855 ;
      RECT 10.945 2.555 11.095 2.705 ;
      RECT 10.61 3.275 10.76 3.425 ;
      RECT 10.555 7.15 10.705 7.3 ;
      RECT 10.53 2.115 10.68 2.265 ;
      RECT 9.095 2.51 9.245 2.66 ;
      RECT 8.33 2.36 8.48 2.51 ;
      RECT 8.075 1.955 8.225 2.105 ;
      RECT 7.455 2.72 7.605 2.87 ;
      RECT 7.075 2.19 7.225 2.34 ;
      RECT 7.06 3.23 7.21 3.38 ;
      RECT 6.53 2.495 6.68 2.645 ;
      RECT 6.37 3.215 6.52 3.365 ;
      RECT 5.56 2.495 5.71 2.645 ;
      RECT 4.745 1.975 4.895 2.125 ;
      RECT 4.585 3.36 4.735 3.51 ;
      RECT 4.35 3.015 4.5 3.165 ;
      RECT 4.305 2.405 4.455 2.555 ;
      RECT 3.305 3.025 3.455 3.175 ;
      RECT 1.62 7.095 1.77 7.245 ;
      RECT 1.245 6.355 1.395 6.505 ;
    LAYER met1 ;
      RECT 66.18 1.26 75.84 1.74 ;
      RECT 50.395 1.26 60.055 1.74 ;
      RECT 34.61 1.26 44.27 1.74 ;
      RECT 18.835 1.26 28.495 1.74 ;
      RECT 3.055 1.26 12.715 1.74 ;
      RECT 66.18 1.26 75.895 1.59 ;
      RECT 50.395 1.26 60.11 1.59 ;
      RECT 34.61 1.26 44.325 1.59 ;
      RECT 18.835 1.26 28.55 1.59 ;
      RECT 3.055 1.26 12.77 1.59 ;
      RECT 66.295 0 76.01 1.585 ;
      RECT 50.51 0 60.225 1.585 ;
      RECT 34.725 0 44.44 1.585 ;
      RECT 18.95 0 28.665 1.585 ;
      RECT 3.17 0 12.885 1.585 ;
      RECT 0 0 81.775 0.305 ;
      RECT 81.17 7.77 81.46 8 ;
      RECT 81.23 6.29 81.4 8 ;
      RECT 81.205 7.275 81.555 7.625 ;
      RECT 81.17 6.29 81.46 6.52 ;
      RECT 80.765 2.395 80.87 2.965 ;
      RECT 80.765 2.73 81.09 2.96 ;
      RECT 80.765 2.76 81.26 2.93 ;
      RECT 80.765 2.395 80.955 2.96 ;
      RECT 80.18 2.36 80.47 2.59 ;
      RECT 80.18 2.395 80.955 2.565 ;
      RECT 80.24 0.88 80.41 2.59 ;
      RECT 80.18 0.88 80.47 1.11 ;
      RECT 80.18 7.77 80.47 8 ;
      RECT 80.24 6.29 80.41 8 ;
      RECT 80.18 6.29 80.47 6.52 ;
      RECT 80.18 6.325 81.035 6.485 ;
      RECT 80.865 5.92 81.035 6.485 ;
      RECT 80.18 6.32 80.575 6.485 ;
      RECT 80.8 5.92 81.09 6.15 ;
      RECT 80.8 5.95 81.26 6.12 ;
      RECT 79.81 2.73 80.1 2.96 ;
      RECT 79.81 2.76 80.27 2.93 ;
      RECT 79.875 1.655 80.04 2.96 ;
      RECT 78.39 1.625 78.68 1.855 ;
      RECT 78.39 1.655 80.04 1.825 ;
      RECT 78.45 0.885 78.62 1.855 ;
      RECT 78.39 0.885 78.68 1.115 ;
      RECT 78.39 7.765 78.68 7.995 ;
      RECT 78.45 7.025 78.62 7.995 ;
      RECT 78.45 7.12 80.04 7.29 ;
      RECT 79.87 5.92 80.04 7.29 ;
      RECT 78.39 7.025 78.68 7.255 ;
      RECT 79.81 5.92 80.1 6.15 ;
      RECT 79.81 5.95 80.27 6.12 ;
      RECT 78.82 1.965 79.17 2.315 ;
      RECT 76.485 2.025 79.17 2.195 ;
      RECT 76.485 1.34 76.655 2.195 ;
      RECT 76.385 1.34 76.735 1.69 ;
      RECT 78.845 6.655 79.17 6.98 ;
      RECT 74.22 6.61 74.57 6.96 ;
      RECT 78.82 6.655 79.17 6.885 ;
      RECT 74.04 6.655 74.57 6.885 ;
      RECT 73.87 6.685 79.17 6.855 ;
      RECT 78.045 2.365 78.365 2.685 ;
      RECT 78.015 2.365 78.365 2.595 ;
      RECT 77.845 2.395 78.365 2.565 ;
      RECT 78.045 6.255 78.365 6.545 ;
      RECT 78.015 6.285 78.365 6.515 ;
      RECT 77.845 6.315 78.365 6.485 ;
      RECT 74.68 2.465 74.865 2.675 ;
      RECT 74.67 2.47 74.88 2.668 ;
      RECT 74.67 2.47 74.966 2.645 ;
      RECT 74.67 2.47 75.025 2.62 ;
      RECT 74.67 2.47 75.08 2.6 ;
      RECT 74.67 2.47 75.09 2.588 ;
      RECT 74.67 2.47 75.285 2.527 ;
      RECT 74.67 2.47 75.315 2.51 ;
      RECT 74.67 2.47 75.335 2.5 ;
      RECT 75.215 2.235 75.475 2.495 ;
      RECT 75.2 2.325 75.215 2.542 ;
      RECT 74.735 2.457 75.475 2.495 ;
      RECT 75.186 2.336 75.2 2.548 ;
      RECT 74.775 2.45 75.475 2.495 ;
      RECT 75.1 2.376 75.186 2.567 ;
      RECT 75.025 2.437 75.475 2.495 ;
      RECT 75.095 2.412 75.1 2.584 ;
      RECT 75.08 2.422 75.475 2.495 ;
      RECT 75.09 2.417 75.095 2.586 ;
      RECT 75.385 2.922 75.39 3.014 ;
      RECT 75.38 2.9 75.385 3.031 ;
      RECT 75.375 2.89 75.38 3.043 ;
      RECT 75.365 2.881 75.375 3.053 ;
      RECT 75.36 2.876 75.365 3.061 ;
      RECT 75.355 2.735 75.36 3.064 ;
      RECT 75.321 2.735 75.355 3.075 ;
      RECT 75.235 2.735 75.321 3.11 ;
      RECT 75.155 2.735 75.235 3.158 ;
      RECT 75.126 2.735 75.155 3.182 ;
      RECT 75.04 2.735 75.126 3.188 ;
      RECT 75.035 2.919 75.04 3.193 ;
      RECT 75 2.93 75.035 3.196 ;
      RECT 74.975 2.945 75 3.2 ;
      RECT 74.961 2.954 74.975 3.202 ;
      RECT 74.875 2.981 74.961 3.208 ;
      RECT 74.81 3.022 74.875 3.217 ;
      RECT 74.795 3.042 74.81 3.222 ;
      RECT 74.765 3.052 74.795 3.225 ;
      RECT 74.76 3.062 74.765 3.228 ;
      RECT 74.73 3.067 74.76 3.23 ;
      RECT 74.71 3.072 74.73 3.234 ;
      RECT 74.625 3.075 74.71 3.241 ;
      RECT 74.61 3.072 74.625 3.247 ;
      RECT 74.6 3.069 74.61 3.249 ;
      RECT 74.58 3.066 74.6 3.251 ;
      RECT 74.56 3.062 74.58 3.252 ;
      RECT 74.545 3.058 74.56 3.254 ;
      RECT 74.535 3.055 74.545 3.255 ;
      RECT 74.495 3.049 74.535 3.253 ;
      RECT 74.485 3.044 74.495 3.251 ;
      RECT 74.47 3.041 74.485 3.247 ;
      RECT 74.445 3.036 74.47 3.24 ;
      RECT 74.395 3.027 74.445 3.228 ;
      RECT 74.325 3.013 74.395 3.21 ;
      RECT 74.267 2.998 74.325 3.192 ;
      RECT 74.181 2.981 74.267 3.172 ;
      RECT 74.095 2.96 74.181 3.147 ;
      RECT 74.045 2.945 74.095 3.128 ;
      RECT 74.041 2.939 74.045 3.12 ;
      RECT 73.955 2.929 74.041 3.107 ;
      RECT 73.92 2.914 73.955 3.09 ;
      RECT 73.905 2.907 73.92 3.083 ;
      RECT 73.845 2.895 73.905 3.071 ;
      RECT 73.825 2.882 73.845 3.059 ;
      RECT 73.785 2.873 73.825 3.051 ;
      RECT 73.78 2.865 73.785 3.044 ;
      RECT 73.7 2.855 73.78 3.03 ;
      RECT 73.685 2.842 73.7 3.015 ;
      RECT 73.68 2.84 73.685 3.013 ;
      RECT 73.601 2.828 73.68 3 ;
      RECT 73.515 2.803 73.601 2.975 ;
      RECT 73.5 2.772 73.515 2.96 ;
      RECT 73.485 2.747 73.5 2.956 ;
      RECT 73.47 2.74 73.485 2.952 ;
      RECT 73.295 2.745 73.3 2.948 ;
      RECT 73.29 2.75 73.295 2.943 ;
      RECT 73.3 2.74 73.47 2.95 ;
      RECT 74.015 2.5 74.12 2.76 ;
      RECT 74.83 2.025 74.835 2.25 ;
      RECT 74.96 2.025 75.015 2.235 ;
      RECT 75.015 2.03 75.025 2.228 ;
      RECT 74.921 2.025 74.96 2.238 ;
      RECT 74.835 2.025 74.921 2.245 ;
      RECT 74.815 2.03 74.83 2.251 ;
      RECT 74.805 2.07 74.815 2.253 ;
      RECT 74.775 2.08 74.805 2.255 ;
      RECT 74.77 2.085 74.775 2.257 ;
      RECT 74.745 2.09 74.77 2.259 ;
      RECT 74.73 2.095 74.745 2.261 ;
      RECT 74.715 2.097 74.73 2.263 ;
      RECT 74.71 2.102 74.715 2.265 ;
      RECT 74.66 2.11 74.71 2.268 ;
      RECT 74.635 2.119 74.66 2.273 ;
      RECT 74.625 2.126 74.635 2.278 ;
      RECT 74.62 2.129 74.625 2.282 ;
      RECT 74.6 2.132 74.62 2.291 ;
      RECT 74.57 2.14 74.6 2.311 ;
      RECT 74.541 2.153 74.57 2.333 ;
      RECT 74.455 2.187 74.541 2.377 ;
      RECT 74.45 2.213 74.455 2.415 ;
      RECT 74.445 2.217 74.45 2.424 ;
      RECT 74.41 2.23 74.445 2.457 ;
      RECT 74.4 2.244 74.41 2.495 ;
      RECT 74.395 2.248 74.4 2.508 ;
      RECT 74.39 2.252 74.395 2.513 ;
      RECT 74.38 2.26 74.39 2.525 ;
      RECT 74.375 2.267 74.38 2.54 ;
      RECT 74.35 2.28 74.375 2.565 ;
      RECT 74.31 2.309 74.35 2.62 ;
      RECT 74.295 2.334 74.31 2.675 ;
      RECT 74.285 2.345 74.295 2.698 ;
      RECT 74.28 2.352 74.285 2.71 ;
      RECT 74.275 2.356 74.28 2.718 ;
      RECT 74.22 2.384 74.275 2.76 ;
      RECT 74.2 2.42 74.22 2.76 ;
      RECT 74.185 2.435 74.2 2.76 ;
      RECT 74.13 2.467 74.185 2.76 ;
      RECT 74.12 2.497 74.13 2.76 ;
      RECT 73.73 2.112 73.915 2.35 ;
      RECT 73.715 2.114 73.925 2.345 ;
      RECT 73.6 2.06 73.86 2.32 ;
      RECT 73.595 2.097 73.86 2.274 ;
      RECT 73.59 2.107 73.86 2.271 ;
      RECT 73.585 2.147 73.925 2.265 ;
      RECT 73.58 2.18 73.925 2.255 ;
      RECT 73.59 2.122 73.94 2.193 ;
      RECT 73.887 3.22 73.9 3.75 ;
      RECT 73.801 3.22 73.9 3.749 ;
      RECT 73.801 3.22 73.905 3.748 ;
      RECT 73.715 3.22 73.905 3.746 ;
      RECT 73.71 3.22 73.905 3.743 ;
      RECT 73.71 3.22 73.915 3.741 ;
      RECT 73.705 3.512 73.915 3.738 ;
      RECT 73.705 3.522 73.92 3.735 ;
      RECT 73.705 3.59 73.925 3.731 ;
      RECT 73.695 3.595 73.925 3.73 ;
      RECT 73.695 3.687 73.93 3.727 ;
      RECT 73.68 3.22 73.94 3.48 ;
      RECT 73.61 7.765 73.9 7.995 ;
      RECT 73.67 7.025 73.84 7.995 ;
      RECT 73.585 7.055 73.925 7.4 ;
      RECT 73.61 7.025 73.9 7.4 ;
      RECT 72.91 2.21 72.955 3.745 ;
      RECT 73.11 2.21 73.14 2.425 ;
      RECT 71.485 1.95 71.605 2.16 ;
      RECT 71.145 1.9 71.405 2.16 ;
      RECT 71.145 1.945 71.44 2.15 ;
      RECT 73.15 2.226 73.155 2.28 ;
      RECT 73.145 2.219 73.15 2.413 ;
      RECT 73.14 2.213 73.145 2.42 ;
      RECT 73.095 2.21 73.11 2.433 ;
      RECT 73.09 2.21 73.095 2.455 ;
      RECT 73.085 2.21 73.09 2.503 ;
      RECT 73.08 2.21 73.085 2.523 ;
      RECT 73.07 2.21 73.08 2.63 ;
      RECT 73.065 2.21 73.07 2.693 ;
      RECT 73.06 2.21 73.065 2.75 ;
      RECT 73.055 2.21 73.06 2.758 ;
      RECT 73.04 2.21 73.055 2.865 ;
      RECT 73.03 2.21 73.04 3 ;
      RECT 73.02 2.21 73.03 3.11 ;
      RECT 73.01 2.21 73.02 3.167 ;
      RECT 73.005 2.21 73.01 3.207 ;
      RECT 73 2.21 73.005 3.243 ;
      RECT 72.99 2.21 73 3.283 ;
      RECT 72.985 2.21 72.99 3.325 ;
      RECT 72.965 2.21 72.985 3.39 ;
      RECT 72.97 3.535 72.975 3.715 ;
      RECT 72.965 3.517 72.97 3.723 ;
      RECT 72.96 2.21 72.965 3.453 ;
      RECT 72.96 3.497 72.965 3.73 ;
      RECT 72.955 2.21 72.96 3.74 ;
      RECT 72.9 2.21 72.91 2.51 ;
      RECT 72.905 2.757 72.91 3.745 ;
      RECT 72.9 2.822 72.905 3.745 ;
      RECT 72.895 2.211 72.9 2.5 ;
      RECT 72.89 2.887 72.9 3.745 ;
      RECT 72.885 2.212 72.895 2.49 ;
      RECT 72.875 3 72.89 3.745 ;
      RECT 72.88 2.213 72.885 2.48 ;
      RECT 72.86 2.214 72.88 2.458 ;
      RECT 72.865 3.097 72.875 3.745 ;
      RECT 72.86 3.172 72.865 3.745 ;
      RECT 72.85 2.213 72.86 2.435 ;
      RECT 72.855 3.215 72.86 3.745 ;
      RECT 72.85 3.242 72.855 3.745 ;
      RECT 72.84 2.211 72.85 2.423 ;
      RECT 72.845 3.285 72.85 3.745 ;
      RECT 72.84 3.312 72.845 3.745 ;
      RECT 72.83 2.21 72.84 2.41 ;
      RECT 72.835 3.327 72.84 3.745 ;
      RECT 72.795 3.385 72.835 3.745 ;
      RECT 72.825 2.209 72.83 2.395 ;
      RECT 72.82 2.207 72.825 2.388 ;
      RECT 72.81 2.204 72.82 2.378 ;
      RECT 72.805 2.201 72.81 2.363 ;
      RECT 72.79 2.197 72.805 2.356 ;
      RECT 72.785 3.44 72.795 3.745 ;
      RECT 72.785 2.194 72.79 2.351 ;
      RECT 72.77 2.19 72.785 2.345 ;
      RECT 72.78 3.457 72.785 3.745 ;
      RECT 72.77 3.52 72.78 3.745 ;
      RECT 72.69 2.175 72.77 2.325 ;
      RECT 72.765 3.527 72.77 3.74 ;
      RECT 72.76 3.535 72.765 3.73 ;
      RECT 72.68 2.161 72.69 2.309 ;
      RECT 72.665 2.157 72.68 2.307 ;
      RECT 72.655 2.152 72.665 2.303 ;
      RECT 72.63 2.145 72.655 2.295 ;
      RECT 72.625 2.14 72.63 2.29 ;
      RECT 72.615 2.14 72.625 2.288 ;
      RECT 72.605 2.138 72.615 2.286 ;
      RECT 72.575 2.13 72.605 2.28 ;
      RECT 72.56 2.122 72.575 2.273 ;
      RECT 72.54 2.117 72.56 2.266 ;
      RECT 72.535 2.113 72.54 2.261 ;
      RECT 72.505 2.106 72.535 2.255 ;
      RECT 72.48 2.097 72.505 2.245 ;
      RECT 72.45 2.09 72.48 2.237 ;
      RECT 72.425 2.08 72.45 2.228 ;
      RECT 72.41 2.072 72.425 2.222 ;
      RECT 72.385 2.067 72.41 2.217 ;
      RECT 72.375 2.063 72.385 2.212 ;
      RECT 72.355 2.058 72.375 2.207 ;
      RECT 72.32 2.053 72.355 2.2 ;
      RECT 72.26 2.048 72.32 2.193 ;
      RECT 72.247 2.044 72.26 2.191 ;
      RECT 72.161 2.039 72.247 2.188 ;
      RECT 72.075 2.029 72.161 2.184 ;
      RECT 72.034 2.022 72.075 2.181 ;
      RECT 71.948 2.015 72.034 2.178 ;
      RECT 71.862 2.005 71.948 2.174 ;
      RECT 71.776 1.995 71.862 2.169 ;
      RECT 71.69 1.985 71.776 2.165 ;
      RECT 71.68 1.97 71.69 2.163 ;
      RECT 71.67 1.955 71.68 2.163 ;
      RECT 71.605 1.95 71.67 2.162 ;
      RECT 71.44 1.947 71.485 2.155 ;
      RECT 72.685 2.852 72.69 3.043 ;
      RECT 72.68 2.847 72.685 3.05 ;
      RECT 72.666 2.845 72.68 3.056 ;
      RECT 72.58 2.845 72.666 3.058 ;
      RECT 72.576 2.845 72.58 3.061 ;
      RECT 72.49 2.845 72.576 3.079 ;
      RECT 72.48 2.85 72.49 3.098 ;
      RECT 72.47 2.905 72.48 3.102 ;
      RECT 72.445 2.92 72.47 3.109 ;
      RECT 72.405 2.94 72.445 3.122 ;
      RECT 72.4 2.952 72.405 3.132 ;
      RECT 72.385 2.958 72.4 3.137 ;
      RECT 72.38 2.963 72.385 3.141 ;
      RECT 72.36 2.97 72.38 3.146 ;
      RECT 72.29 2.995 72.36 3.163 ;
      RECT 72.25 3.023 72.29 3.183 ;
      RECT 72.245 3.033 72.25 3.191 ;
      RECT 72.225 3.04 72.245 3.193 ;
      RECT 72.22 3.047 72.225 3.196 ;
      RECT 72.19 3.055 72.22 3.199 ;
      RECT 72.185 3.06 72.19 3.203 ;
      RECT 72.111 3.064 72.185 3.211 ;
      RECT 72.025 3.073 72.111 3.227 ;
      RECT 72.021 3.078 72.025 3.236 ;
      RECT 71.935 3.083 72.021 3.246 ;
      RECT 71.895 3.091 71.935 3.258 ;
      RECT 71.845 3.097 71.895 3.265 ;
      RECT 71.76 3.106 71.845 3.28 ;
      RECT 71.685 3.117 71.76 3.298 ;
      RECT 71.65 3.124 71.685 3.308 ;
      RECT 71.575 3.132 71.65 3.313 ;
      RECT 71.52 3.141 71.575 3.313 ;
      RECT 71.495 3.146 71.52 3.311 ;
      RECT 71.485 3.149 71.495 3.309 ;
      RECT 71.45 3.151 71.485 3.307 ;
      RECT 71.42 3.153 71.45 3.303 ;
      RECT 71.375 3.152 71.42 3.299 ;
      RECT 71.355 3.147 71.375 3.296 ;
      RECT 71.305 3.132 71.355 3.293 ;
      RECT 71.295 3.117 71.305 3.288 ;
      RECT 71.245 3.102 71.295 3.278 ;
      RECT 71.195 3.077 71.245 3.258 ;
      RECT 71.185 3.062 71.195 3.24 ;
      RECT 71.18 3.06 71.185 3.234 ;
      RECT 71.16 3.055 71.18 3.229 ;
      RECT 71.155 3.047 71.16 3.223 ;
      RECT 71.14 3.041 71.155 3.216 ;
      RECT 71.135 3.036 71.14 3.208 ;
      RECT 71.115 3.031 71.135 3.2 ;
      RECT 71.1 3.024 71.115 3.193 ;
      RECT 71.085 3.018 71.1 3.184 ;
      RECT 71.08 3.012 71.085 3.177 ;
      RECT 71.035 2.987 71.08 3.163 ;
      RECT 71.02 2.957 71.035 3.145 ;
      RECT 71.005 2.94 71.02 3.136 ;
      RECT 70.98 2.92 71.005 3.124 ;
      RECT 70.94 2.89 70.98 3.104 ;
      RECT 70.93 2.86 70.94 3.089 ;
      RECT 70.915 2.85 70.93 3.082 ;
      RECT 70.86 2.815 70.915 3.061 ;
      RECT 70.845 2.778 70.86 3.04 ;
      RECT 70.835 2.765 70.845 3.032 ;
      RECT 70.785 2.735 70.835 3.014 ;
      RECT 70.77 2.665 70.785 2.995 ;
      RECT 70.725 2.665 70.77 2.978 ;
      RECT 70.7 2.665 70.725 2.96 ;
      RECT 70.69 2.665 70.7 2.953 ;
      RECT 70.611 2.665 70.69 2.946 ;
      RECT 70.525 2.665 70.611 2.938 ;
      RECT 70.51 2.697 70.525 2.933 ;
      RECT 70.435 2.707 70.51 2.929 ;
      RECT 70.415 2.717 70.435 2.924 ;
      RECT 70.39 2.717 70.415 2.921 ;
      RECT 70.38 2.707 70.39 2.92 ;
      RECT 70.37 2.68 70.38 2.919 ;
      RECT 70.33 2.675 70.37 2.917 ;
      RECT 70.285 2.675 70.33 2.913 ;
      RECT 70.26 2.675 70.285 2.908 ;
      RECT 70.21 2.675 70.26 2.895 ;
      RECT 70.17 2.68 70.18 2.88 ;
      RECT 70.18 2.675 70.21 2.885 ;
      RECT 72.165 2.455 72.425 2.715 ;
      RECT 72.16 2.477 72.425 2.673 ;
      RECT 71.4 2.305 71.62 2.67 ;
      RECT 71.382 2.392 71.62 2.669 ;
      RECT 71.365 2.397 71.62 2.666 ;
      RECT 71.365 2.397 71.64 2.665 ;
      RECT 71.335 2.407 71.64 2.663 ;
      RECT 71.33 2.422 71.64 2.659 ;
      RECT 71.33 2.422 71.645 2.658 ;
      RECT 71.325 2.48 71.645 2.656 ;
      RECT 71.325 2.48 71.655 2.653 ;
      RECT 71.32 2.545 71.655 2.648 ;
      RECT 71.4 2.305 71.66 2.565 ;
      RECT 70.145 2.135 70.405 2.395 ;
      RECT 70.145 2.178 70.491 2.369 ;
      RECT 70.145 2.178 70.535 2.368 ;
      RECT 70.145 2.178 70.555 2.366 ;
      RECT 70.145 2.178 70.655 2.365 ;
      RECT 70.145 2.178 70.675 2.363 ;
      RECT 70.145 2.178 70.685 2.358 ;
      RECT 70.555 2.145 70.745 2.355 ;
      RECT 70.555 2.147 70.75 2.353 ;
      RECT 70.545 2.152 70.755 2.345 ;
      RECT 70.491 2.176 70.755 2.345 ;
      RECT 70.535 2.17 70.545 2.367 ;
      RECT 70.545 2.15 70.75 2.353 ;
      RECT 69.5 3.21 69.705 3.44 ;
      RECT 69.44 3.16 69.495 3.42 ;
      RECT 69.5 3.16 69.7 3.44 ;
      RECT 70.47 3.475 70.475 3.502 ;
      RECT 70.46 3.385 70.47 3.507 ;
      RECT 70.455 3.307 70.46 3.513 ;
      RECT 70.445 3.297 70.455 3.52 ;
      RECT 70.44 3.287 70.445 3.526 ;
      RECT 70.43 3.282 70.44 3.528 ;
      RECT 70.415 3.274 70.43 3.536 ;
      RECT 70.4 3.265 70.415 3.548 ;
      RECT 70.39 3.257 70.4 3.558 ;
      RECT 70.355 3.175 70.39 3.576 ;
      RECT 70.32 3.175 70.355 3.595 ;
      RECT 70.305 3.175 70.32 3.603 ;
      RECT 70.25 3.175 70.305 3.603 ;
      RECT 70.216 3.175 70.25 3.594 ;
      RECT 70.13 3.175 70.216 3.57 ;
      RECT 70.12 3.235 70.13 3.552 ;
      RECT 70.08 3.237 70.12 3.543 ;
      RECT 70.075 3.239 70.08 3.533 ;
      RECT 70.055 3.241 70.075 3.528 ;
      RECT 70.045 3.244 70.055 3.523 ;
      RECT 70.035 3.245 70.045 3.518 ;
      RECT 70.011 3.246 70.035 3.51 ;
      RECT 69.925 3.251 70.011 3.488 ;
      RECT 69.87 3.25 69.925 3.461 ;
      RECT 69.855 3.243 69.87 3.448 ;
      RECT 69.82 3.238 69.855 3.444 ;
      RECT 69.765 3.23 69.82 3.443 ;
      RECT 69.705 3.217 69.765 3.441 ;
      RECT 69.495 3.16 69.5 3.428 ;
      RECT 69.57 2.53 69.755 2.74 ;
      RECT 69.56 2.535 69.77 2.733 ;
      RECT 69.6 2.44 69.86 2.7 ;
      RECT 69.555 2.597 69.86 2.623 ;
      RECT 68.9 2.39 68.905 3.19 ;
      RECT 68.845 2.44 68.875 3.19 ;
      RECT 68.835 2.44 68.84 2.75 ;
      RECT 68.82 2.44 68.825 2.745 ;
      RECT 68.365 2.485 68.38 2.7 ;
      RECT 68.295 2.485 68.38 2.695 ;
      RECT 69.56 2.065 69.63 2.275 ;
      RECT 69.63 2.072 69.64 2.27 ;
      RECT 69.526 2.065 69.56 2.282 ;
      RECT 69.44 2.065 69.526 2.306 ;
      RECT 69.43 2.07 69.44 2.325 ;
      RECT 69.425 2.082 69.43 2.328 ;
      RECT 69.41 2.097 69.425 2.332 ;
      RECT 69.405 2.115 69.41 2.336 ;
      RECT 69.365 2.125 69.405 2.345 ;
      RECT 69.35 2.132 69.365 2.357 ;
      RECT 69.335 2.137 69.35 2.362 ;
      RECT 69.32 2.14 69.335 2.367 ;
      RECT 69.31 2.142 69.32 2.371 ;
      RECT 69.275 2.149 69.31 2.379 ;
      RECT 69.24 2.157 69.275 2.393 ;
      RECT 69.23 2.163 69.24 2.402 ;
      RECT 69.225 2.165 69.23 2.404 ;
      RECT 69.205 2.168 69.225 2.41 ;
      RECT 69.175 2.175 69.205 2.421 ;
      RECT 69.165 2.181 69.175 2.428 ;
      RECT 69.14 2.184 69.165 2.435 ;
      RECT 69.13 2.188 69.14 2.443 ;
      RECT 69.125 2.189 69.13 2.465 ;
      RECT 69.12 2.19 69.125 2.48 ;
      RECT 69.115 2.191 69.12 2.495 ;
      RECT 69.11 2.192 69.115 2.51 ;
      RECT 69.105 2.193 69.11 2.54 ;
      RECT 69.095 2.195 69.105 2.573 ;
      RECT 69.08 2.199 69.095 2.62 ;
      RECT 69.07 2.202 69.08 2.665 ;
      RECT 69.065 2.205 69.07 2.693 ;
      RECT 69.055 2.207 69.065 2.72 ;
      RECT 69.05 2.21 69.055 2.755 ;
      RECT 69.02 2.215 69.05 2.813 ;
      RECT 69.015 2.22 69.02 2.898 ;
      RECT 69.01 2.222 69.015 2.933 ;
      RECT 69.005 2.224 69.01 3.015 ;
      RECT 69 2.226 69.005 3.103 ;
      RECT 68.99 2.228 69 3.185 ;
      RECT 68.975 2.242 68.99 3.19 ;
      RECT 68.94 2.287 68.975 3.19 ;
      RECT 68.93 2.327 68.94 3.19 ;
      RECT 68.915 2.355 68.93 3.19 ;
      RECT 68.91 2.372 68.915 3.19 ;
      RECT 68.905 2.38 68.91 3.19 ;
      RECT 68.895 2.395 68.9 3.19 ;
      RECT 68.89 2.402 68.895 3.19 ;
      RECT 68.88 2.422 68.89 3.19 ;
      RECT 68.875 2.435 68.88 3.19 ;
      RECT 68.84 2.44 68.845 2.775 ;
      RECT 68.825 2.83 68.845 3.19 ;
      RECT 68.825 2.44 68.835 2.748 ;
      RECT 68.82 2.87 68.825 3.19 ;
      RECT 68.77 2.44 68.82 2.743 ;
      RECT 68.815 2.907 68.82 3.19 ;
      RECT 68.805 2.93 68.815 3.19 ;
      RECT 68.8 2.975 68.805 3.19 ;
      RECT 68.79 2.985 68.8 3.183 ;
      RECT 68.716 2.44 68.77 2.737 ;
      RECT 68.63 2.44 68.716 2.73 ;
      RECT 68.581 2.487 68.63 2.723 ;
      RECT 68.495 2.495 68.581 2.716 ;
      RECT 68.48 2.492 68.495 2.711 ;
      RECT 68.466 2.485 68.48 2.71 ;
      RECT 68.38 2.485 68.466 2.705 ;
      RECT 68.285 2.49 68.295 2.69 ;
      RECT 67.875 1.92 67.89 2.32 ;
      RECT 68.07 1.92 68.075 2.18 ;
      RECT 67.815 1.92 67.86 2.18 ;
      RECT 68.27 3.225 68.275 3.43 ;
      RECT 68.265 3.215 68.27 3.435 ;
      RECT 68.26 3.202 68.265 3.44 ;
      RECT 68.255 3.182 68.26 3.44 ;
      RECT 68.23 3.135 68.255 3.44 ;
      RECT 68.195 3.05 68.23 3.44 ;
      RECT 68.19 2.987 68.195 3.44 ;
      RECT 68.185 2.972 68.19 3.44 ;
      RECT 68.17 2.932 68.185 3.44 ;
      RECT 68.165 2.907 68.17 3.44 ;
      RECT 68.155 2.89 68.165 3.44 ;
      RECT 68.12 2.812 68.155 3.44 ;
      RECT 68.115 2.755 68.12 3.44 ;
      RECT 68.11 2.742 68.115 3.44 ;
      RECT 68.1 2.72 68.11 3.44 ;
      RECT 68.09 2.685 68.1 3.44 ;
      RECT 68.08 2.655 68.09 3.44 ;
      RECT 68.07 2.57 68.08 3.083 ;
      RECT 68.077 3.215 68.08 3.44 ;
      RECT 68.075 3.225 68.077 3.44 ;
      RECT 68.065 3.235 68.075 3.435 ;
      RECT 68.06 1.92 68.07 2.315 ;
      RECT 68.065 2.447 68.07 3.058 ;
      RECT 68.06 2.345 68.065 3.041 ;
      RECT 68.05 1.92 68.06 3.017 ;
      RECT 68.045 1.92 68.05 2.988 ;
      RECT 68.04 1.92 68.045 2.978 ;
      RECT 68.02 1.92 68.04 2.94 ;
      RECT 68.015 1.92 68.02 2.898 ;
      RECT 68.01 1.92 68.015 2.878 ;
      RECT 67.98 1.92 68.01 2.828 ;
      RECT 67.97 1.92 67.98 2.775 ;
      RECT 67.965 1.92 67.97 2.748 ;
      RECT 67.96 1.92 67.965 2.733 ;
      RECT 67.95 1.92 67.96 2.71 ;
      RECT 67.94 1.92 67.95 2.685 ;
      RECT 67.935 1.92 67.94 2.625 ;
      RECT 67.925 1.92 67.935 2.563 ;
      RECT 67.92 1.92 67.925 2.483 ;
      RECT 67.915 1.92 67.92 2.448 ;
      RECT 67.91 1.92 67.915 2.423 ;
      RECT 67.905 1.92 67.91 2.408 ;
      RECT 67.9 1.92 67.905 2.378 ;
      RECT 67.895 1.92 67.9 2.355 ;
      RECT 67.89 1.92 67.895 2.328 ;
      RECT 67.86 1.92 67.875 2.315 ;
      RECT 67.015 3.455 67.2 3.665 ;
      RECT 67.005 3.46 67.215 3.658 ;
      RECT 67.005 3.46 67.235 3.63 ;
      RECT 67.005 3.46 67.25 3.609 ;
      RECT 67.005 3.46 67.265 3.607 ;
      RECT 67.005 3.46 67.275 3.606 ;
      RECT 67.005 3.46 67.305 3.603 ;
      RECT 67.655 3.305 67.915 3.565 ;
      RECT 67.615 3.352 67.915 3.548 ;
      RECT 67.606 3.36 67.615 3.551 ;
      RECT 67.2 3.453 67.915 3.548 ;
      RECT 67.52 3.378 67.606 3.558 ;
      RECT 67.215 3.45 67.915 3.548 ;
      RECT 67.461 3.4 67.52 3.57 ;
      RECT 67.235 3.446 67.915 3.548 ;
      RECT 67.375 3.412 67.461 3.581 ;
      RECT 67.25 3.442 67.915 3.548 ;
      RECT 67.32 3.425 67.375 3.593 ;
      RECT 67.265 3.44 67.915 3.548 ;
      RECT 67.305 3.431 67.32 3.599 ;
      RECT 67.275 3.436 67.915 3.548 ;
      RECT 67.42 2.96 67.68 3.22 ;
      RECT 67.42 2.98 67.79 3.19 ;
      RECT 67.42 2.985 67.8 3.185 ;
      RECT 67.611 2.399 67.69 2.63 ;
      RECT 67.525 2.402 67.74 2.625 ;
      RECT 67.52 2.402 67.74 2.62 ;
      RECT 67.52 2.407 67.75 2.618 ;
      RECT 67.495 2.407 67.75 2.615 ;
      RECT 67.495 2.415 67.76 2.613 ;
      RECT 67.375 2.35 67.635 2.61 ;
      RECT 67.375 2.397 67.685 2.61 ;
      RECT 66.63 2.97 66.635 3.23 ;
      RECT 66.46 2.74 66.465 3.23 ;
      RECT 66.345 2.98 66.35 3.205 ;
      RECT 67.055 2.075 67.06 2.285 ;
      RECT 67.06 2.08 67.075 2.28 ;
      RECT 66.995 2.075 67.055 2.293 ;
      RECT 66.98 2.075 66.995 2.303 ;
      RECT 66.93 2.075 66.98 2.32 ;
      RECT 66.91 2.075 66.93 2.343 ;
      RECT 66.895 2.075 66.91 2.355 ;
      RECT 66.875 2.075 66.895 2.365 ;
      RECT 66.865 2.08 66.875 2.374 ;
      RECT 66.86 2.09 66.865 2.379 ;
      RECT 66.855 2.102 66.86 2.383 ;
      RECT 66.845 2.125 66.855 2.388 ;
      RECT 66.84 2.14 66.845 2.392 ;
      RECT 66.835 2.157 66.84 2.395 ;
      RECT 66.83 2.165 66.835 2.398 ;
      RECT 66.82 2.17 66.83 2.402 ;
      RECT 66.815 2.177 66.82 2.407 ;
      RECT 66.805 2.182 66.815 2.411 ;
      RECT 66.78 2.194 66.805 2.422 ;
      RECT 66.76 2.211 66.78 2.438 ;
      RECT 66.735 2.228 66.76 2.46 ;
      RECT 66.7 2.251 66.735 2.518 ;
      RECT 66.68 2.273 66.7 2.58 ;
      RECT 66.675 2.283 66.68 2.615 ;
      RECT 66.665 2.29 66.675 2.653 ;
      RECT 66.66 2.297 66.665 2.673 ;
      RECT 66.655 2.308 66.66 2.71 ;
      RECT 66.65 2.316 66.655 2.775 ;
      RECT 66.64 2.327 66.65 2.828 ;
      RECT 66.635 2.345 66.64 2.898 ;
      RECT 66.63 2.355 66.635 2.935 ;
      RECT 66.625 2.365 66.63 3.23 ;
      RECT 66.62 2.377 66.625 3.23 ;
      RECT 66.615 2.387 66.62 3.23 ;
      RECT 66.605 2.397 66.615 3.23 ;
      RECT 66.595 2.42 66.605 3.23 ;
      RECT 66.58 2.455 66.595 3.23 ;
      RECT 66.54 2.517 66.58 3.23 ;
      RECT 66.535 2.57 66.54 3.23 ;
      RECT 66.51 2.605 66.535 3.23 ;
      RECT 66.495 2.65 66.51 3.23 ;
      RECT 66.49 2.672 66.495 3.23 ;
      RECT 66.48 2.685 66.49 3.23 ;
      RECT 66.47 2.71 66.48 3.23 ;
      RECT 66.465 2.732 66.47 3.23 ;
      RECT 66.44 2.77 66.46 3.23 ;
      RECT 66.4 2.827 66.44 3.23 ;
      RECT 66.395 2.877 66.4 3.23 ;
      RECT 66.39 2.895 66.395 3.23 ;
      RECT 66.385 2.907 66.39 3.23 ;
      RECT 66.375 2.925 66.385 3.23 ;
      RECT 66.365 2.945 66.375 3.205 ;
      RECT 66.36 2.962 66.365 3.205 ;
      RECT 66.35 2.975 66.36 3.205 ;
      RECT 66.32 2.985 66.345 3.205 ;
      RECT 66.31 2.992 66.32 3.205 ;
      RECT 66.295 3.002 66.31 3.2 ;
      RECT 65.385 7.77 65.675 8 ;
      RECT 65.445 6.29 65.615 8 ;
      RECT 65.395 6.655 65.745 7.005 ;
      RECT 65.385 6.29 65.675 6.52 ;
      RECT 64.98 2.395 65.085 2.965 ;
      RECT 64.98 2.73 65.305 2.96 ;
      RECT 64.98 2.76 65.475 2.93 ;
      RECT 64.98 2.395 65.17 2.96 ;
      RECT 64.395 2.36 64.685 2.59 ;
      RECT 64.395 2.395 65.17 2.565 ;
      RECT 64.455 0.88 64.625 2.59 ;
      RECT 64.395 0.88 64.685 1.11 ;
      RECT 64.395 7.77 64.685 8 ;
      RECT 64.455 6.29 64.625 8 ;
      RECT 64.395 6.29 64.685 6.52 ;
      RECT 64.395 6.325 65.25 6.485 ;
      RECT 65.08 5.92 65.25 6.485 ;
      RECT 64.395 6.32 64.79 6.485 ;
      RECT 65.015 5.92 65.305 6.15 ;
      RECT 65.015 5.95 65.475 6.12 ;
      RECT 64.025 2.73 64.315 2.96 ;
      RECT 64.025 2.76 64.485 2.93 ;
      RECT 64.09 1.655 64.255 2.96 ;
      RECT 62.605 1.625 62.895 1.855 ;
      RECT 62.605 1.655 64.255 1.825 ;
      RECT 62.665 0.885 62.835 1.855 ;
      RECT 62.605 0.885 62.895 1.115 ;
      RECT 62.605 7.765 62.895 7.995 ;
      RECT 62.665 7.025 62.835 7.995 ;
      RECT 62.665 7.12 64.255 7.29 ;
      RECT 64.085 5.92 64.255 7.29 ;
      RECT 62.605 7.025 62.895 7.255 ;
      RECT 64.025 5.92 64.315 6.15 ;
      RECT 64.025 5.95 64.485 6.12 ;
      RECT 63.035 1.965 63.385 2.315 ;
      RECT 60.7 2.025 63.385 2.195 ;
      RECT 60.7 1.34 60.87 2.195 ;
      RECT 60.6 1.34 60.95 1.69 ;
      RECT 63.06 6.655 63.385 6.98 ;
      RECT 58.435 6.61 58.785 6.96 ;
      RECT 63.035 6.655 63.385 6.885 ;
      RECT 58.255 6.655 58.785 6.885 ;
      RECT 58.085 6.685 63.385 6.855 ;
      RECT 62.26 2.365 62.58 2.685 ;
      RECT 62.23 2.365 62.58 2.595 ;
      RECT 62.06 2.395 62.58 2.565 ;
      RECT 62.26 6.255 62.58 6.545 ;
      RECT 62.23 6.285 62.58 6.515 ;
      RECT 62.06 6.315 62.58 6.485 ;
      RECT 58.895 2.465 59.08 2.675 ;
      RECT 58.885 2.47 59.095 2.668 ;
      RECT 58.885 2.47 59.181 2.645 ;
      RECT 58.885 2.47 59.24 2.62 ;
      RECT 58.885 2.47 59.295 2.6 ;
      RECT 58.885 2.47 59.305 2.588 ;
      RECT 58.885 2.47 59.5 2.527 ;
      RECT 58.885 2.47 59.53 2.51 ;
      RECT 58.885 2.47 59.55 2.5 ;
      RECT 59.43 2.235 59.69 2.495 ;
      RECT 59.415 2.325 59.43 2.542 ;
      RECT 58.95 2.457 59.69 2.495 ;
      RECT 59.401 2.336 59.415 2.548 ;
      RECT 58.99 2.45 59.69 2.495 ;
      RECT 59.315 2.376 59.401 2.567 ;
      RECT 59.24 2.437 59.69 2.495 ;
      RECT 59.31 2.412 59.315 2.584 ;
      RECT 59.295 2.422 59.69 2.495 ;
      RECT 59.305 2.417 59.31 2.586 ;
      RECT 59.6 2.922 59.605 3.014 ;
      RECT 59.595 2.9 59.6 3.031 ;
      RECT 59.59 2.89 59.595 3.043 ;
      RECT 59.58 2.881 59.59 3.053 ;
      RECT 59.575 2.876 59.58 3.061 ;
      RECT 59.57 2.735 59.575 3.064 ;
      RECT 59.536 2.735 59.57 3.075 ;
      RECT 59.45 2.735 59.536 3.11 ;
      RECT 59.37 2.735 59.45 3.158 ;
      RECT 59.341 2.735 59.37 3.182 ;
      RECT 59.255 2.735 59.341 3.188 ;
      RECT 59.25 2.919 59.255 3.193 ;
      RECT 59.215 2.93 59.25 3.196 ;
      RECT 59.19 2.945 59.215 3.2 ;
      RECT 59.176 2.954 59.19 3.202 ;
      RECT 59.09 2.981 59.176 3.208 ;
      RECT 59.025 3.022 59.09 3.217 ;
      RECT 59.01 3.042 59.025 3.222 ;
      RECT 58.98 3.052 59.01 3.225 ;
      RECT 58.975 3.062 58.98 3.228 ;
      RECT 58.945 3.067 58.975 3.23 ;
      RECT 58.925 3.072 58.945 3.234 ;
      RECT 58.84 3.075 58.925 3.241 ;
      RECT 58.825 3.072 58.84 3.247 ;
      RECT 58.815 3.069 58.825 3.249 ;
      RECT 58.795 3.066 58.815 3.251 ;
      RECT 58.775 3.062 58.795 3.252 ;
      RECT 58.76 3.058 58.775 3.254 ;
      RECT 58.75 3.055 58.76 3.255 ;
      RECT 58.71 3.049 58.75 3.253 ;
      RECT 58.7 3.044 58.71 3.251 ;
      RECT 58.685 3.041 58.7 3.247 ;
      RECT 58.66 3.036 58.685 3.24 ;
      RECT 58.61 3.027 58.66 3.228 ;
      RECT 58.54 3.013 58.61 3.21 ;
      RECT 58.482 2.998 58.54 3.192 ;
      RECT 58.396 2.981 58.482 3.172 ;
      RECT 58.31 2.96 58.396 3.147 ;
      RECT 58.26 2.945 58.31 3.128 ;
      RECT 58.256 2.939 58.26 3.12 ;
      RECT 58.17 2.929 58.256 3.107 ;
      RECT 58.135 2.914 58.17 3.09 ;
      RECT 58.12 2.907 58.135 3.083 ;
      RECT 58.06 2.895 58.12 3.071 ;
      RECT 58.04 2.882 58.06 3.059 ;
      RECT 58 2.873 58.04 3.051 ;
      RECT 57.995 2.865 58 3.044 ;
      RECT 57.915 2.855 57.995 3.03 ;
      RECT 57.9 2.842 57.915 3.015 ;
      RECT 57.895 2.84 57.9 3.013 ;
      RECT 57.816 2.828 57.895 3 ;
      RECT 57.73 2.803 57.816 2.975 ;
      RECT 57.715 2.772 57.73 2.96 ;
      RECT 57.7 2.747 57.715 2.956 ;
      RECT 57.685 2.74 57.7 2.952 ;
      RECT 57.51 2.745 57.515 2.948 ;
      RECT 57.505 2.75 57.51 2.943 ;
      RECT 57.515 2.74 57.685 2.95 ;
      RECT 58.23 2.5 58.335 2.76 ;
      RECT 59.045 2.025 59.05 2.25 ;
      RECT 59.175 2.025 59.23 2.235 ;
      RECT 59.23 2.03 59.24 2.228 ;
      RECT 59.136 2.025 59.175 2.238 ;
      RECT 59.05 2.025 59.136 2.245 ;
      RECT 59.03 2.03 59.045 2.251 ;
      RECT 59.02 2.07 59.03 2.253 ;
      RECT 58.99 2.08 59.02 2.255 ;
      RECT 58.985 2.085 58.99 2.257 ;
      RECT 58.96 2.09 58.985 2.259 ;
      RECT 58.945 2.095 58.96 2.261 ;
      RECT 58.93 2.097 58.945 2.263 ;
      RECT 58.925 2.102 58.93 2.265 ;
      RECT 58.875 2.11 58.925 2.268 ;
      RECT 58.85 2.119 58.875 2.273 ;
      RECT 58.84 2.126 58.85 2.278 ;
      RECT 58.835 2.129 58.84 2.282 ;
      RECT 58.815 2.132 58.835 2.291 ;
      RECT 58.785 2.14 58.815 2.311 ;
      RECT 58.756 2.153 58.785 2.333 ;
      RECT 58.67 2.187 58.756 2.377 ;
      RECT 58.665 2.213 58.67 2.415 ;
      RECT 58.66 2.217 58.665 2.424 ;
      RECT 58.625 2.23 58.66 2.457 ;
      RECT 58.615 2.244 58.625 2.495 ;
      RECT 58.61 2.248 58.615 2.508 ;
      RECT 58.605 2.252 58.61 2.513 ;
      RECT 58.595 2.26 58.605 2.525 ;
      RECT 58.59 2.267 58.595 2.54 ;
      RECT 58.565 2.28 58.59 2.565 ;
      RECT 58.525 2.309 58.565 2.62 ;
      RECT 58.51 2.334 58.525 2.675 ;
      RECT 58.5 2.345 58.51 2.698 ;
      RECT 58.495 2.352 58.5 2.71 ;
      RECT 58.49 2.356 58.495 2.718 ;
      RECT 58.435 2.384 58.49 2.76 ;
      RECT 58.415 2.42 58.435 2.76 ;
      RECT 58.4 2.435 58.415 2.76 ;
      RECT 58.345 2.467 58.4 2.76 ;
      RECT 58.335 2.497 58.345 2.76 ;
      RECT 57.945 2.112 58.13 2.35 ;
      RECT 57.93 2.114 58.14 2.345 ;
      RECT 57.815 2.06 58.075 2.32 ;
      RECT 57.81 2.097 58.075 2.274 ;
      RECT 57.805 2.107 58.075 2.271 ;
      RECT 57.8 2.147 58.14 2.265 ;
      RECT 57.795 2.18 58.14 2.255 ;
      RECT 57.805 2.122 58.155 2.193 ;
      RECT 58.102 3.22 58.115 3.75 ;
      RECT 58.016 3.22 58.115 3.749 ;
      RECT 58.016 3.22 58.12 3.748 ;
      RECT 57.93 3.22 58.12 3.746 ;
      RECT 57.925 3.22 58.12 3.743 ;
      RECT 57.925 3.22 58.13 3.741 ;
      RECT 57.92 3.512 58.13 3.738 ;
      RECT 57.92 3.522 58.135 3.735 ;
      RECT 57.92 3.59 58.14 3.731 ;
      RECT 57.91 3.595 58.14 3.73 ;
      RECT 57.91 3.687 58.145 3.727 ;
      RECT 57.895 3.22 58.155 3.48 ;
      RECT 57.825 7.765 58.115 7.995 ;
      RECT 57.885 7.025 58.055 7.995 ;
      RECT 57.8 7.055 58.14 7.4 ;
      RECT 57.825 7.025 58.115 7.4 ;
      RECT 57.125 2.21 57.17 3.745 ;
      RECT 57.325 2.21 57.355 2.425 ;
      RECT 55.7 1.95 55.82 2.16 ;
      RECT 55.36 1.9 55.62 2.16 ;
      RECT 55.36 1.945 55.655 2.15 ;
      RECT 57.365 2.226 57.37 2.28 ;
      RECT 57.36 2.219 57.365 2.413 ;
      RECT 57.355 2.213 57.36 2.42 ;
      RECT 57.31 2.21 57.325 2.433 ;
      RECT 57.305 2.21 57.31 2.455 ;
      RECT 57.3 2.21 57.305 2.503 ;
      RECT 57.295 2.21 57.3 2.523 ;
      RECT 57.285 2.21 57.295 2.63 ;
      RECT 57.28 2.21 57.285 2.693 ;
      RECT 57.275 2.21 57.28 2.75 ;
      RECT 57.27 2.21 57.275 2.758 ;
      RECT 57.255 2.21 57.27 2.865 ;
      RECT 57.245 2.21 57.255 3 ;
      RECT 57.235 2.21 57.245 3.11 ;
      RECT 57.225 2.21 57.235 3.167 ;
      RECT 57.22 2.21 57.225 3.207 ;
      RECT 57.215 2.21 57.22 3.243 ;
      RECT 57.205 2.21 57.215 3.283 ;
      RECT 57.2 2.21 57.205 3.325 ;
      RECT 57.18 2.21 57.2 3.39 ;
      RECT 57.185 3.535 57.19 3.715 ;
      RECT 57.18 3.517 57.185 3.723 ;
      RECT 57.175 2.21 57.18 3.453 ;
      RECT 57.175 3.497 57.18 3.73 ;
      RECT 57.17 2.21 57.175 3.74 ;
      RECT 57.115 2.21 57.125 2.51 ;
      RECT 57.12 2.757 57.125 3.745 ;
      RECT 57.115 2.822 57.12 3.745 ;
      RECT 57.11 2.211 57.115 2.5 ;
      RECT 57.105 2.887 57.115 3.745 ;
      RECT 57.1 2.212 57.11 2.49 ;
      RECT 57.09 3 57.105 3.745 ;
      RECT 57.095 2.213 57.1 2.48 ;
      RECT 57.075 2.214 57.095 2.458 ;
      RECT 57.08 3.097 57.09 3.745 ;
      RECT 57.075 3.172 57.08 3.745 ;
      RECT 57.065 2.213 57.075 2.435 ;
      RECT 57.07 3.215 57.075 3.745 ;
      RECT 57.065 3.242 57.07 3.745 ;
      RECT 57.055 2.211 57.065 2.423 ;
      RECT 57.06 3.285 57.065 3.745 ;
      RECT 57.055 3.312 57.06 3.745 ;
      RECT 57.045 2.21 57.055 2.41 ;
      RECT 57.05 3.327 57.055 3.745 ;
      RECT 57.01 3.385 57.05 3.745 ;
      RECT 57.04 2.209 57.045 2.395 ;
      RECT 57.035 2.207 57.04 2.388 ;
      RECT 57.025 2.204 57.035 2.378 ;
      RECT 57.02 2.201 57.025 2.363 ;
      RECT 57.005 2.197 57.02 2.356 ;
      RECT 57 3.44 57.01 3.745 ;
      RECT 57 2.194 57.005 2.351 ;
      RECT 56.985 2.19 57 2.345 ;
      RECT 56.995 3.457 57 3.745 ;
      RECT 56.985 3.52 56.995 3.745 ;
      RECT 56.905 2.175 56.985 2.325 ;
      RECT 56.98 3.527 56.985 3.74 ;
      RECT 56.975 3.535 56.98 3.73 ;
      RECT 56.895 2.161 56.905 2.309 ;
      RECT 56.88 2.157 56.895 2.307 ;
      RECT 56.87 2.152 56.88 2.303 ;
      RECT 56.845 2.145 56.87 2.295 ;
      RECT 56.84 2.14 56.845 2.29 ;
      RECT 56.83 2.14 56.84 2.288 ;
      RECT 56.82 2.138 56.83 2.286 ;
      RECT 56.79 2.13 56.82 2.28 ;
      RECT 56.775 2.122 56.79 2.273 ;
      RECT 56.755 2.117 56.775 2.266 ;
      RECT 56.75 2.113 56.755 2.261 ;
      RECT 56.72 2.106 56.75 2.255 ;
      RECT 56.695 2.097 56.72 2.245 ;
      RECT 56.665 2.09 56.695 2.237 ;
      RECT 56.64 2.08 56.665 2.228 ;
      RECT 56.625 2.072 56.64 2.222 ;
      RECT 56.6 2.067 56.625 2.217 ;
      RECT 56.59 2.063 56.6 2.212 ;
      RECT 56.57 2.058 56.59 2.207 ;
      RECT 56.535 2.053 56.57 2.2 ;
      RECT 56.475 2.048 56.535 2.193 ;
      RECT 56.462 2.044 56.475 2.191 ;
      RECT 56.376 2.039 56.462 2.188 ;
      RECT 56.29 2.029 56.376 2.184 ;
      RECT 56.249 2.022 56.29 2.181 ;
      RECT 56.163 2.015 56.249 2.178 ;
      RECT 56.077 2.005 56.163 2.174 ;
      RECT 55.991 1.995 56.077 2.169 ;
      RECT 55.905 1.985 55.991 2.165 ;
      RECT 55.895 1.97 55.905 2.163 ;
      RECT 55.885 1.955 55.895 2.163 ;
      RECT 55.82 1.95 55.885 2.162 ;
      RECT 55.655 1.947 55.7 2.155 ;
      RECT 56.9 2.852 56.905 3.043 ;
      RECT 56.895 2.847 56.9 3.05 ;
      RECT 56.881 2.845 56.895 3.056 ;
      RECT 56.795 2.845 56.881 3.058 ;
      RECT 56.791 2.845 56.795 3.061 ;
      RECT 56.705 2.845 56.791 3.079 ;
      RECT 56.695 2.85 56.705 3.098 ;
      RECT 56.685 2.905 56.695 3.102 ;
      RECT 56.66 2.92 56.685 3.109 ;
      RECT 56.62 2.94 56.66 3.122 ;
      RECT 56.615 2.952 56.62 3.132 ;
      RECT 56.6 2.958 56.615 3.137 ;
      RECT 56.595 2.963 56.6 3.141 ;
      RECT 56.575 2.97 56.595 3.146 ;
      RECT 56.505 2.995 56.575 3.163 ;
      RECT 56.465 3.023 56.505 3.183 ;
      RECT 56.46 3.033 56.465 3.191 ;
      RECT 56.44 3.04 56.46 3.193 ;
      RECT 56.435 3.047 56.44 3.196 ;
      RECT 56.405 3.055 56.435 3.199 ;
      RECT 56.4 3.06 56.405 3.203 ;
      RECT 56.326 3.064 56.4 3.211 ;
      RECT 56.24 3.073 56.326 3.227 ;
      RECT 56.236 3.078 56.24 3.236 ;
      RECT 56.15 3.083 56.236 3.246 ;
      RECT 56.11 3.091 56.15 3.258 ;
      RECT 56.06 3.097 56.11 3.265 ;
      RECT 55.975 3.106 56.06 3.28 ;
      RECT 55.9 3.117 55.975 3.298 ;
      RECT 55.865 3.124 55.9 3.308 ;
      RECT 55.79 3.132 55.865 3.313 ;
      RECT 55.735 3.141 55.79 3.313 ;
      RECT 55.71 3.146 55.735 3.311 ;
      RECT 55.7 3.149 55.71 3.309 ;
      RECT 55.665 3.151 55.7 3.307 ;
      RECT 55.635 3.153 55.665 3.303 ;
      RECT 55.59 3.152 55.635 3.299 ;
      RECT 55.57 3.147 55.59 3.296 ;
      RECT 55.52 3.132 55.57 3.293 ;
      RECT 55.51 3.117 55.52 3.288 ;
      RECT 55.46 3.102 55.51 3.278 ;
      RECT 55.41 3.077 55.46 3.258 ;
      RECT 55.4 3.062 55.41 3.24 ;
      RECT 55.395 3.06 55.4 3.234 ;
      RECT 55.375 3.055 55.395 3.229 ;
      RECT 55.37 3.047 55.375 3.223 ;
      RECT 55.355 3.041 55.37 3.216 ;
      RECT 55.35 3.036 55.355 3.208 ;
      RECT 55.33 3.031 55.35 3.2 ;
      RECT 55.315 3.024 55.33 3.193 ;
      RECT 55.3 3.018 55.315 3.184 ;
      RECT 55.295 3.012 55.3 3.177 ;
      RECT 55.25 2.987 55.295 3.163 ;
      RECT 55.235 2.957 55.25 3.145 ;
      RECT 55.22 2.94 55.235 3.136 ;
      RECT 55.195 2.92 55.22 3.124 ;
      RECT 55.155 2.89 55.195 3.104 ;
      RECT 55.145 2.86 55.155 3.089 ;
      RECT 55.13 2.85 55.145 3.082 ;
      RECT 55.075 2.815 55.13 3.061 ;
      RECT 55.06 2.778 55.075 3.04 ;
      RECT 55.05 2.765 55.06 3.032 ;
      RECT 55 2.735 55.05 3.014 ;
      RECT 54.985 2.665 55 2.995 ;
      RECT 54.94 2.665 54.985 2.978 ;
      RECT 54.915 2.665 54.94 2.96 ;
      RECT 54.905 2.665 54.915 2.953 ;
      RECT 54.826 2.665 54.905 2.946 ;
      RECT 54.74 2.665 54.826 2.938 ;
      RECT 54.725 2.697 54.74 2.933 ;
      RECT 54.65 2.707 54.725 2.929 ;
      RECT 54.63 2.717 54.65 2.924 ;
      RECT 54.605 2.717 54.63 2.921 ;
      RECT 54.595 2.707 54.605 2.92 ;
      RECT 54.585 2.68 54.595 2.919 ;
      RECT 54.545 2.675 54.585 2.917 ;
      RECT 54.5 2.675 54.545 2.913 ;
      RECT 54.475 2.675 54.5 2.908 ;
      RECT 54.425 2.675 54.475 2.895 ;
      RECT 54.385 2.68 54.395 2.88 ;
      RECT 54.395 2.675 54.425 2.885 ;
      RECT 56.38 2.455 56.64 2.715 ;
      RECT 56.375 2.477 56.64 2.673 ;
      RECT 55.615 2.305 55.835 2.67 ;
      RECT 55.597 2.392 55.835 2.669 ;
      RECT 55.58 2.397 55.835 2.666 ;
      RECT 55.58 2.397 55.855 2.665 ;
      RECT 55.55 2.407 55.855 2.663 ;
      RECT 55.545 2.422 55.855 2.659 ;
      RECT 55.545 2.422 55.86 2.658 ;
      RECT 55.54 2.48 55.86 2.656 ;
      RECT 55.54 2.48 55.87 2.653 ;
      RECT 55.535 2.545 55.87 2.648 ;
      RECT 55.615 2.305 55.875 2.565 ;
      RECT 54.36 2.135 54.62 2.395 ;
      RECT 54.36 2.178 54.706 2.369 ;
      RECT 54.36 2.178 54.75 2.368 ;
      RECT 54.36 2.178 54.77 2.366 ;
      RECT 54.36 2.178 54.87 2.365 ;
      RECT 54.36 2.178 54.89 2.363 ;
      RECT 54.36 2.178 54.9 2.358 ;
      RECT 54.77 2.145 54.96 2.355 ;
      RECT 54.77 2.147 54.965 2.353 ;
      RECT 54.76 2.152 54.97 2.345 ;
      RECT 54.706 2.176 54.97 2.345 ;
      RECT 54.75 2.17 54.76 2.367 ;
      RECT 54.76 2.15 54.965 2.353 ;
      RECT 53.715 3.21 53.92 3.44 ;
      RECT 53.655 3.16 53.71 3.42 ;
      RECT 53.715 3.16 53.915 3.44 ;
      RECT 54.685 3.475 54.69 3.502 ;
      RECT 54.675 3.385 54.685 3.507 ;
      RECT 54.67 3.307 54.675 3.513 ;
      RECT 54.66 3.297 54.67 3.52 ;
      RECT 54.655 3.287 54.66 3.526 ;
      RECT 54.645 3.282 54.655 3.528 ;
      RECT 54.63 3.274 54.645 3.536 ;
      RECT 54.615 3.265 54.63 3.548 ;
      RECT 54.605 3.257 54.615 3.558 ;
      RECT 54.57 3.175 54.605 3.576 ;
      RECT 54.535 3.175 54.57 3.595 ;
      RECT 54.52 3.175 54.535 3.603 ;
      RECT 54.465 3.175 54.52 3.603 ;
      RECT 54.431 3.175 54.465 3.594 ;
      RECT 54.345 3.175 54.431 3.57 ;
      RECT 54.335 3.235 54.345 3.552 ;
      RECT 54.295 3.237 54.335 3.543 ;
      RECT 54.29 3.239 54.295 3.533 ;
      RECT 54.27 3.241 54.29 3.528 ;
      RECT 54.26 3.244 54.27 3.523 ;
      RECT 54.25 3.245 54.26 3.518 ;
      RECT 54.226 3.246 54.25 3.51 ;
      RECT 54.14 3.251 54.226 3.488 ;
      RECT 54.085 3.25 54.14 3.461 ;
      RECT 54.07 3.243 54.085 3.448 ;
      RECT 54.035 3.238 54.07 3.444 ;
      RECT 53.98 3.23 54.035 3.443 ;
      RECT 53.92 3.217 53.98 3.441 ;
      RECT 53.71 3.16 53.715 3.428 ;
      RECT 53.785 2.53 53.97 2.74 ;
      RECT 53.775 2.535 53.985 2.733 ;
      RECT 53.815 2.44 54.075 2.7 ;
      RECT 53.77 2.597 54.075 2.623 ;
      RECT 53.115 2.39 53.12 3.19 ;
      RECT 53.06 2.44 53.09 3.19 ;
      RECT 53.05 2.44 53.055 2.75 ;
      RECT 53.035 2.44 53.04 2.745 ;
      RECT 52.58 2.485 52.595 2.7 ;
      RECT 52.51 2.485 52.595 2.695 ;
      RECT 53.775 2.065 53.845 2.275 ;
      RECT 53.845 2.072 53.855 2.27 ;
      RECT 53.741 2.065 53.775 2.282 ;
      RECT 53.655 2.065 53.741 2.306 ;
      RECT 53.645 2.07 53.655 2.325 ;
      RECT 53.64 2.082 53.645 2.328 ;
      RECT 53.625 2.097 53.64 2.332 ;
      RECT 53.62 2.115 53.625 2.336 ;
      RECT 53.58 2.125 53.62 2.345 ;
      RECT 53.565 2.132 53.58 2.357 ;
      RECT 53.55 2.137 53.565 2.362 ;
      RECT 53.535 2.14 53.55 2.367 ;
      RECT 53.525 2.142 53.535 2.371 ;
      RECT 53.49 2.149 53.525 2.379 ;
      RECT 53.455 2.157 53.49 2.393 ;
      RECT 53.445 2.163 53.455 2.402 ;
      RECT 53.44 2.165 53.445 2.404 ;
      RECT 53.42 2.168 53.44 2.41 ;
      RECT 53.39 2.175 53.42 2.421 ;
      RECT 53.38 2.181 53.39 2.428 ;
      RECT 53.355 2.184 53.38 2.435 ;
      RECT 53.345 2.188 53.355 2.443 ;
      RECT 53.34 2.189 53.345 2.465 ;
      RECT 53.335 2.19 53.34 2.48 ;
      RECT 53.33 2.191 53.335 2.495 ;
      RECT 53.325 2.192 53.33 2.51 ;
      RECT 53.32 2.193 53.325 2.54 ;
      RECT 53.31 2.195 53.32 2.573 ;
      RECT 53.295 2.199 53.31 2.62 ;
      RECT 53.285 2.202 53.295 2.665 ;
      RECT 53.28 2.205 53.285 2.693 ;
      RECT 53.27 2.207 53.28 2.72 ;
      RECT 53.265 2.21 53.27 2.755 ;
      RECT 53.235 2.215 53.265 2.813 ;
      RECT 53.23 2.22 53.235 2.898 ;
      RECT 53.225 2.222 53.23 2.933 ;
      RECT 53.22 2.224 53.225 3.015 ;
      RECT 53.215 2.226 53.22 3.103 ;
      RECT 53.205 2.228 53.215 3.185 ;
      RECT 53.19 2.242 53.205 3.19 ;
      RECT 53.155 2.287 53.19 3.19 ;
      RECT 53.145 2.327 53.155 3.19 ;
      RECT 53.13 2.355 53.145 3.19 ;
      RECT 53.125 2.372 53.13 3.19 ;
      RECT 53.12 2.38 53.125 3.19 ;
      RECT 53.11 2.395 53.115 3.19 ;
      RECT 53.105 2.402 53.11 3.19 ;
      RECT 53.095 2.422 53.105 3.19 ;
      RECT 53.09 2.435 53.095 3.19 ;
      RECT 53.055 2.44 53.06 2.775 ;
      RECT 53.04 2.83 53.06 3.19 ;
      RECT 53.04 2.44 53.05 2.748 ;
      RECT 53.035 2.87 53.04 3.19 ;
      RECT 52.985 2.44 53.035 2.743 ;
      RECT 53.03 2.907 53.035 3.19 ;
      RECT 53.02 2.93 53.03 3.19 ;
      RECT 53.015 2.975 53.02 3.19 ;
      RECT 53.005 2.985 53.015 3.183 ;
      RECT 52.931 2.44 52.985 2.737 ;
      RECT 52.845 2.44 52.931 2.73 ;
      RECT 52.796 2.487 52.845 2.723 ;
      RECT 52.71 2.495 52.796 2.716 ;
      RECT 52.695 2.492 52.71 2.711 ;
      RECT 52.681 2.485 52.695 2.71 ;
      RECT 52.595 2.485 52.681 2.705 ;
      RECT 52.5 2.49 52.51 2.69 ;
      RECT 52.09 1.92 52.105 2.32 ;
      RECT 52.285 1.92 52.29 2.18 ;
      RECT 52.03 1.92 52.075 2.18 ;
      RECT 52.485 3.225 52.49 3.43 ;
      RECT 52.48 3.215 52.485 3.435 ;
      RECT 52.475 3.202 52.48 3.44 ;
      RECT 52.47 3.182 52.475 3.44 ;
      RECT 52.445 3.135 52.47 3.44 ;
      RECT 52.41 3.05 52.445 3.44 ;
      RECT 52.405 2.987 52.41 3.44 ;
      RECT 52.4 2.972 52.405 3.44 ;
      RECT 52.385 2.932 52.4 3.44 ;
      RECT 52.38 2.907 52.385 3.44 ;
      RECT 52.37 2.89 52.38 3.44 ;
      RECT 52.335 2.812 52.37 3.44 ;
      RECT 52.33 2.755 52.335 3.44 ;
      RECT 52.325 2.742 52.33 3.44 ;
      RECT 52.315 2.72 52.325 3.44 ;
      RECT 52.305 2.685 52.315 3.44 ;
      RECT 52.295 2.655 52.305 3.44 ;
      RECT 52.285 2.57 52.295 3.083 ;
      RECT 52.292 3.215 52.295 3.44 ;
      RECT 52.29 3.225 52.292 3.44 ;
      RECT 52.28 3.235 52.29 3.435 ;
      RECT 52.275 1.92 52.285 2.315 ;
      RECT 52.28 2.447 52.285 3.058 ;
      RECT 52.275 2.345 52.28 3.041 ;
      RECT 52.265 1.92 52.275 3.017 ;
      RECT 52.26 1.92 52.265 2.988 ;
      RECT 52.255 1.92 52.26 2.978 ;
      RECT 52.235 1.92 52.255 2.94 ;
      RECT 52.23 1.92 52.235 2.898 ;
      RECT 52.225 1.92 52.23 2.878 ;
      RECT 52.195 1.92 52.225 2.828 ;
      RECT 52.185 1.92 52.195 2.775 ;
      RECT 52.18 1.92 52.185 2.748 ;
      RECT 52.175 1.92 52.18 2.733 ;
      RECT 52.165 1.92 52.175 2.71 ;
      RECT 52.155 1.92 52.165 2.685 ;
      RECT 52.15 1.92 52.155 2.625 ;
      RECT 52.14 1.92 52.15 2.563 ;
      RECT 52.135 1.92 52.14 2.483 ;
      RECT 52.13 1.92 52.135 2.448 ;
      RECT 52.125 1.92 52.13 2.423 ;
      RECT 52.12 1.92 52.125 2.408 ;
      RECT 52.115 1.92 52.12 2.378 ;
      RECT 52.11 1.92 52.115 2.355 ;
      RECT 52.105 1.92 52.11 2.328 ;
      RECT 52.075 1.92 52.09 2.315 ;
      RECT 51.23 3.455 51.415 3.665 ;
      RECT 51.22 3.46 51.43 3.658 ;
      RECT 51.22 3.46 51.45 3.63 ;
      RECT 51.22 3.46 51.465 3.609 ;
      RECT 51.22 3.46 51.48 3.607 ;
      RECT 51.22 3.46 51.49 3.606 ;
      RECT 51.22 3.46 51.52 3.603 ;
      RECT 51.87 3.305 52.13 3.565 ;
      RECT 51.83 3.352 52.13 3.548 ;
      RECT 51.821 3.36 51.83 3.551 ;
      RECT 51.415 3.453 52.13 3.548 ;
      RECT 51.735 3.378 51.821 3.558 ;
      RECT 51.43 3.45 52.13 3.548 ;
      RECT 51.676 3.4 51.735 3.57 ;
      RECT 51.45 3.446 52.13 3.548 ;
      RECT 51.59 3.412 51.676 3.581 ;
      RECT 51.465 3.442 52.13 3.548 ;
      RECT 51.535 3.425 51.59 3.593 ;
      RECT 51.48 3.44 52.13 3.548 ;
      RECT 51.52 3.431 51.535 3.599 ;
      RECT 51.49 3.436 52.13 3.548 ;
      RECT 51.635 2.96 51.895 3.22 ;
      RECT 51.635 2.98 52.005 3.19 ;
      RECT 51.635 2.985 52.015 3.185 ;
      RECT 51.826 2.399 51.905 2.63 ;
      RECT 51.74 2.402 51.955 2.625 ;
      RECT 51.735 2.402 51.955 2.62 ;
      RECT 51.735 2.407 51.965 2.618 ;
      RECT 51.71 2.407 51.965 2.615 ;
      RECT 51.71 2.415 51.975 2.613 ;
      RECT 51.59 2.35 51.85 2.61 ;
      RECT 51.59 2.397 51.9 2.61 ;
      RECT 50.845 2.97 50.85 3.23 ;
      RECT 50.675 2.74 50.68 3.23 ;
      RECT 50.56 2.98 50.565 3.205 ;
      RECT 51.27 2.075 51.275 2.285 ;
      RECT 51.275 2.08 51.29 2.28 ;
      RECT 51.21 2.075 51.27 2.293 ;
      RECT 51.195 2.075 51.21 2.303 ;
      RECT 51.145 2.075 51.195 2.32 ;
      RECT 51.125 2.075 51.145 2.343 ;
      RECT 51.11 2.075 51.125 2.355 ;
      RECT 51.09 2.075 51.11 2.365 ;
      RECT 51.08 2.08 51.09 2.374 ;
      RECT 51.075 2.09 51.08 2.379 ;
      RECT 51.07 2.102 51.075 2.383 ;
      RECT 51.06 2.125 51.07 2.388 ;
      RECT 51.055 2.14 51.06 2.392 ;
      RECT 51.05 2.157 51.055 2.395 ;
      RECT 51.045 2.165 51.05 2.398 ;
      RECT 51.035 2.17 51.045 2.402 ;
      RECT 51.03 2.177 51.035 2.407 ;
      RECT 51.02 2.182 51.03 2.411 ;
      RECT 50.995 2.194 51.02 2.422 ;
      RECT 50.975 2.211 50.995 2.438 ;
      RECT 50.95 2.228 50.975 2.46 ;
      RECT 50.915 2.251 50.95 2.518 ;
      RECT 50.895 2.273 50.915 2.58 ;
      RECT 50.89 2.283 50.895 2.615 ;
      RECT 50.88 2.29 50.89 2.653 ;
      RECT 50.875 2.297 50.88 2.673 ;
      RECT 50.87 2.308 50.875 2.71 ;
      RECT 50.865 2.316 50.87 2.775 ;
      RECT 50.855 2.327 50.865 2.828 ;
      RECT 50.85 2.345 50.855 2.898 ;
      RECT 50.845 2.355 50.85 2.935 ;
      RECT 50.84 2.365 50.845 3.23 ;
      RECT 50.835 2.377 50.84 3.23 ;
      RECT 50.83 2.387 50.835 3.23 ;
      RECT 50.82 2.397 50.83 3.23 ;
      RECT 50.81 2.42 50.82 3.23 ;
      RECT 50.795 2.455 50.81 3.23 ;
      RECT 50.755 2.517 50.795 3.23 ;
      RECT 50.75 2.57 50.755 3.23 ;
      RECT 50.725 2.605 50.75 3.23 ;
      RECT 50.71 2.65 50.725 3.23 ;
      RECT 50.705 2.672 50.71 3.23 ;
      RECT 50.695 2.685 50.705 3.23 ;
      RECT 50.685 2.71 50.695 3.23 ;
      RECT 50.68 2.732 50.685 3.23 ;
      RECT 50.655 2.77 50.675 3.23 ;
      RECT 50.615 2.827 50.655 3.23 ;
      RECT 50.61 2.877 50.615 3.23 ;
      RECT 50.605 2.895 50.61 3.23 ;
      RECT 50.6 2.907 50.605 3.23 ;
      RECT 50.59 2.925 50.6 3.23 ;
      RECT 50.58 2.945 50.59 3.205 ;
      RECT 50.575 2.962 50.58 3.205 ;
      RECT 50.565 2.975 50.575 3.205 ;
      RECT 50.535 2.985 50.56 3.205 ;
      RECT 50.525 2.992 50.535 3.205 ;
      RECT 50.51 3.002 50.525 3.2 ;
      RECT 49.6 7.77 49.89 8 ;
      RECT 49.66 6.29 49.83 8 ;
      RECT 49.61 6.655 49.96 7.005 ;
      RECT 49.6 6.29 49.89 6.52 ;
      RECT 49.195 2.395 49.3 2.965 ;
      RECT 49.195 2.73 49.52 2.96 ;
      RECT 49.195 2.76 49.69 2.93 ;
      RECT 49.195 2.395 49.385 2.96 ;
      RECT 48.61 2.36 48.9 2.59 ;
      RECT 48.61 2.395 49.385 2.565 ;
      RECT 48.67 0.88 48.84 2.59 ;
      RECT 48.61 0.88 48.9 1.11 ;
      RECT 48.61 7.77 48.9 8 ;
      RECT 48.67 6.29 48.84 8 ;
      RECT 48.61 6.29 48.9 6.52 ;
      RECT 48.61 6.325 49.465 6.485 ;
      RECT 49.295 5.92 49.465 6.485 ;
      RECT 48.61 6.32 49.005 6.485 ;
      RECT 49.23 5.92 49.52 6.15 ;
      RECT 49.23 5.95 49.69 6.12 ;
      RECT 48.24 2.73 48.53 2.96 ;
      RECT 48.24 2.76 48.7 2.93 ;
      RECT 48.305 1.655 48.47 2.96 ;
      RECT 46.82 1.625 47.11 1.855 ;
      RECT 46.82 1.655 48.47 1.825 ;
      RECT 46.88 0.885 47.05 1.855 ;
      RECT 46.82 0.885 47.11 1.115 ;
      RECT 46.82 7.765 47.11 7.995 ;
      RECT 46.88 7.025 47.05 7.995 ;
      RECT 46.88 7.12 48.47 7.29 ;
      RECT 48.3 5.92 48.47 7.29 ;
      RECT 46.82 7.025 47.11 7.255 ;
      RECT 48.24 5.92 48.53 6.15 ;
      RECT 48.24 5.95 48.7 6.12 ;
      RECT 47.25 1.965 47.6 2.315 ;
      RECT 44.915 2.025 47.6 2.195 ;
      RECT 44.915 1.34 45.085 2.195 ;
      RECT 44.815 1.34 45.165 1.69 ;
      RECT 47.275 6.655 47.6 6.98 ;
      RECT 42.705 6.615 43.055 6.965 ;
      RECT 47.25 6.655 47.6 6.885 ;
      RECT 42.47 6.655 43.055 6.885 ;
      RECT 42.3 6.685 47.6 6.855 ;
      RECT 46.475 2.365 46.795 2.685 ;
      RECT 46.445 2.365 46.795 2.595 ;
      RECT 46.275 2.395 46.795 2.565 ;
      RECT 46.475 6.255 46.795 6.545 ;
      RECT 46.445 6.285 46.795 6.515 ;
      RECT 46.275 6.315 46.795 6.485 ;
      RECT 43.11 2.465 43.295 2.675 ;
      RECT 43.1 2.47 43.31 2.668 ;
      RECT 43.1 2.47 43.396 2.645 ;
      RECT 43.1 2.47 43.455 2.62 ;
      RECT 43.1 2.47 43.51 2.6 ;
      RECT 43.1 2.47 43.52 2.588 ;
      RECT 43.1 2.47 43.715 2.527 ;
      RECT 43.1 2.47 43.745 2.51 ;
      RECT 43.1 2.47 43.765 2.5 ;
      RECT 43.645 2.235 43.905 2.495 ;
      RECT 43.63 2.325 43.645 2.542 ;
      RECT 43.165 2.457 43.905 2.495 ;
      RECT 43.616 2.336 43.63 2.548 ;
      RECT 43.205 2.45 43.905 2.495 ;
      RECT 43.53 2.376 43.616 2.567 ;
      RECT 43.455 2.437 43.905 2.495 ;
      RECT 43.525 2.412 43.53 2.584 ;
      RECT 43.51 2.422 43.905 2.495 ;
      RECT 43.52 2.417 43.525 2.586 ;
      RECT 43.815 2.922 43.82 3.014 ;
      RECT 43.81 2.9 43.815 3.031 ;
      RECT 43.805 2.89 43.81 3.043 ;
      RECT 43.795 2.881 43.805 3.053 ;
      RECT 43.79 2.876 43.795 3.061 ;
      RECT 43.785 2.735 43.79 3.064 ;
      RECT 43.751 2.735 43.785 3.075 ;
      RECT 43.665 2.735 43.751 3.11 ;
      RECT 43.585 2.735 43.665 3.158 ;
      RECT 43.556 2.735 43.585 3.182 ;
      RECT 43.47 2.735 43.556 3.188 ;
      RECT 43.465 2.919 43.47 3.193 ;
      RECT 43.43 2.93 43.465 3.196 ;
      RECT 43.405 2.945 43.43 3.2 ;
      RECT 43.391 2.954 43.405 3.202 ;
      RECT 43.305 2.981 43.391 3.208 ;
      RECT 43.24 3.022 43.305 3.217 ;
      RECT 43.225 3.042 43.24 3.222 ;
      RECT 43.195 3.052 43.225 3.225 ;
      RECT 43.19 3.062 43.195 3.228 ;
      RECT 43.16 3.067 43.19 3.23 ;
      RECT 43.14 3.072 43.16 3.234 ;
      RECT 43.055 3.075 43.14 3.241 ;
      RECT 43.04 3.072 43.055 3.247 ;
      RECT 43.03 3.069 43.04 3.249 ;
      RECT 43.01 3.066 43.03 3.251 ;
      RECT 42.99 3.062 43.01 3.252 ;
      RECT 42.975 3.058 42.99 3.254 ;
      RECT 42.965 3.055 42.975 3.255 ;
      RECT 42.925 3.049 42.965 3.253 ;
      RECT 42.915 3.044 42.925 3.251 ;
      RECT 42.9 3.041 42.915 3.247 ;
      RECT 42.875 3.036 42.9 3.24 ;
      RECT 42.825 3.027 42.875 3.228 ;
      RECT 42.755 3.013 42.825 3.21 ;
      RECT 42.697 2.998 42.755 3.192 ;
      RECT 42.611 2.981 42.697 3.172 ;
      RECT 42.525 2.96 42.611 3.147 ;
      RECT 42.475 2.945 42.525 3.128 ;
      RECT 42.471 2.939 42.475 3.12 ;
      RECT 42.385 2.929 42.471 3.107 ;
      RECT 42.35 2.914 42.385 3.09 ;
      RECT 42.335 2.907 42.35 3.083 ;
      RECT 42.275 2.895 42.335 3.071 ;
      RECT 42.255 2.882 42.275 3.059 ;
      RECT 42.215 2.873 42.255 3.051 ;
      RECT 42.21 2.865 42.215 3.044 ;
      RECT 42.13 2.855 42.21 3.03 ;
      RECT 42.115 2.842 42.13 3.015 ;
      RECT 42.11 2.84 42.115 3.013 ;
      RECT 42.031 2.828 42.11 3 ;
      RECT 41.945 2.803 42.031 2.975 ;
      RECT 41.93 2.772 41.945 2.96 ;
      RECT 41.915 2.747 41.93 2.956 ;
      RECT 41.9 2.74 41.915 2.952 ;
      RECT 41.725 2.745 41.73 2.948 ;
      RECT 41.72 2.75 41.725 2.943 ;
      RECT 41.73 2.74 41.9 2.95 ;
      RECT 42.445 2.5 42.55 2.76 ;
      RECT 43.26 2.025 43.265 2.25 ;
      RECT 43.39 2.025 43.445 2.235 ;
      RECT 43.445 2.03 43.455 2.228 ;
      RECT 43.351 2.025 43.39 2.238 ;
      RECT 43.265 2.025 43.351 2.245 ;
      RECT 43.245 2.03 43.26 2.251 ;
      RECT 43.235 2.07 43.245 2.253 ;
      RECT 43.205 2.08 43.235 2.255 ;
      RECT 43.2 2.085 43.205 2.257 ;
      RECT 43.175 2.09 43.2 2.259 ;
      RECT 43.16 2.095 43.175 2.261 ;
      RECT 43.145 2.097 43.16 2.263 ;
      RECT 43.14 2.102 43.145 2.265 ;
      RECT 43.09 2.11 43.14 2.268 ;
      RECT 43.065 2.119 43.09 2.273 ;
      RECT 43.055 2.126 43.065 2.278 ;
      RECT 43.05 2.129 43.055 2.282 ;
      RECT 43.03 2.132 43.05 2.291 ;
      RECT 43 2.14 43.03 2.311 ;
      RECT 42.971 2.153 43 2.333 ;
      RECT 42.885 2.187 42.971 2.377 ;
      RECT 42.88 2.213 42.885 2.415 ;
      RECT 42.875 2.217 42.88 2.424 ;
      RECT 42.84 2.23 42.875 2.457 ;
      RECT 42.83 2.244 42.84 2.495 ;
      RECT 42.825 2.248 42.83 2.508 ;
      RECT 42.82 2.252 42.825 2.513 ;
      RECT 42.81 2.26 42.82 2.525 ;
      RECT 42.805 2.267 42.81 2.54 ;
      RECT 42.78 2.28 42.805 2.565 ;
      RECT 42.74 2.309 42.78 2.62 ;
      RECT 42.725 2.334 42.74 2.675 ;
      RECT 42.715 2.345 42.725 2.698 ;
      RECT 42.71 2.352 42.715 2.71 ;
      RECT 42.705 2.356 42.71 2.718 ;
      RECT 42.65 2.384 42.705 2.76 ;
      RECT 42.63 2.42 42.65 2.76 ;
      RECT 42.615 2.435 42.63 2.76 ;
      RECT 42.56 2.467 42.615 2.76 ;
      RECT 42.55 2.497 42.56 2.76 ;
      RECT 42.16 2.112 42.345 2.35 ;
      RECT 42.145 2.114 42.355 2.345 ;
      RECT 42.03 2.06 42.29 2.32 ;
      RECT 42.025 2.097 42.29 2.274 ;
      RECT 42.02 2.107 42.29 2.271 ;
      RECT 42.015 2.147 42.355 2.265 ;
      RECT 42.01 2.18 42.355 2.255 ;
      RECT 42.02 2.122 42.37 2.193 ;
      RECT 42.317 3.22 42.33 3.75 ;
      RECT 42.231 3.22 42.33 3.749 ;
      RECT 42.231 3.22 42.335 3.748 ;
      RECT 42.145 3.22 42.335 3.746 ;
      RECT 42.14 3.22 42.335 3.743 ;
      RECT 42.14 3.22 42.345 3.741 ;
      RECT 42.135 3.512 42.345 3.738 ;
      RECT 42.135 3.522 42.35 3.735 ;
      RECT 42.135 3.59 42.355 3.731 ;
      RECT 42.125 3.595 42.355 3.73 ;
      RECT 42.125 3.687 42.36 3.727 ;
      RECT 42.11 3.22 42.37 3.48 ;
      RECT 42.04 7.765 42.33 7.995 ;
      RECT 42.1 7.025 42.27 7.995 ;
      RECT 42.015 7.055 42.355 7.4 ;
      RECT 42.04 7.025 42.33 7.4 ;
      RECT 41.34 2.21 41.385 3.745 ;
      RECT 41.54 2.21 41.57 2.425 ;
      RECT 39.915 1.95 40.035 2.16 ;
      RECT 39.575 1.9 39.835 2.16 ;
      RECT 39.575 1.945 39.87 2.15 ;
      RECT 41.58 2.226 41.585 2.28 ;
      RECT 41.575 2.219 41.58 2.413 ;
      RECT 41.57 2.213 41.575 2.42 ;
      RECT 41.525 2.21 41.54 2.433 ;
      RECT 41.52 2.21 41.525 2.455 ;
      RECT 41.515 2.21 41.52 2.503 ;
      RECT 41.51 2.21 41.515 2.523 ;
      RECT 41.5 2.21 41.51 2.63 ;
      RECT 41.495 2.21 41.5 2.693 ;
      RECT 41.49 2.21 41.495 2.75 ;
      RECT 41.485 2.21 41.49 2.758 ;
      RECT 41.47 2.21 41.485 2.865 ;
      RECT 41.46 2.21 41.47 3 ;
      RECT 41.45 2.21 41.46 3.11 ;
      RECT 41.44 2.21 41.45 3.167 ;
      RECT 41.435 2.21 41.44 3.207 ;
      RECT 41.43 2.21 41.435 3.243 ;
      RECT 41.42 2.21 41.43 3.283 ;
      RECT 41.415 2.21 41.42 3.325 ;
      RECT 41.395 2.21 41.415 3.39 ;
      RECT 41.4 3.535 41.405 3.715 ;
      RECT 41.395 3.517 41.4 3.723 ;
      RECT 41.39 2.21 41.395 3.453 ;
      RECT 41.39 3.497 41.395 3.73 ;
      RECT 41.385 2.21 41.39 3.74 ;
      RECT 41.33 2.21 41.34 2.51 ;
      RECT 41.335 2.757 41.34 3.745 ;
      RECT 41.33 2.822 41.335 3.745 ;
      RECT 41.325 2.211 41.33 2.5 ;
      RECT 41.32 2.887 41.33 3.745 ;
      RECT 41.315 2.212 41.325 2.49 ;
      RECT 41.305 3 41.32 3.745 ;
      RECT 41.31 2.213 41.315 2.48 ;
      RECT 41.29 2.214 41.31 2.458 ;
      RECT 41.295 3.097 41.305 3.745 ;
      RECT 41.29 3.172 41.295 3.745 ;
      RECT 41.28 2.213 41.29 2.435 ;
      RECT 41.285 3.215 41.29 3.745 ;
      RECT 41.28 3.242 41.285 3.745 ;
      RECT 41.27 2.211 41.28 2.423 ;
      RECT 41.275 3.285 41.28 3.745 ;
      RECT 41.27 3.312 41.275 3.745 ;
      RECT 41.26 2.21 41.27 2.41 ;
      RECT 41.265 3.327 41.27 3.745 ;
      RECT 41.225 3.385 41.265 3.745 ;
      RECT 41.255 2.209 41.26 2.395 ;
      RECT 41.25 2.207 41.255 2.388 ;
      RECT 41.24 2.204 41.25 2.378 ;
      RECT 41.235 2.201 41.24 2.363 ;
      RECT 41.22 2.197 41.235 2.356 ;
      RECT 41.215 3.44 41.225 3.745 ;
      RECT 41.215 2.194 41.22 2.351 ;
      RECT 41.2 2.19 41.215 2.345 ;
      RECT 41.21 3.457 41.215 3.745 ;
      RECT 41.2 3.52 41.21 3.745 ;
      RECT 41.12 2.175 41.2 2.325 ;
      RECT 41.195 3.527 41.2 3.74 ;
      RECT 41.19 3.535 41.195 3.73 ;
      RECT 41.11 2.161 41.12 2.309 ;
      RECT 41.095 2.157 41.11 2.307 ;
      RECT 41.085 2.152 41.095 2.303 ;
      RECT 41.06 2.145 41.085 2.295 ;
      RECT 41.055 2.14 41.06 2.29 ;
      RECT 41.045 2.14 41.055 2.288 ;
      RECT 41.035 2.138 41.045 2.286 ;
      RECT 41.005 2.13 41.035 2.28 ;
      RECT 40.99 2.122 41.005 2.273 ;
      RECT 40.97 2.117 40.99 2.266 ;
      RECT 40.965 2.113 40.97 2.261 ;
      RECT 40.935 2.106 40.965 2.255 ;
      RECT 40.91 2.097 40.935 2.245 ;
      RECT 40.88 2.09 40.91 2.237 ;
      RECT 40.855 2.08 40.88 2.228 ;
      RECT 40.84 2.072 40.855 2.222 ;
      RECT 40.815 2.067 40.84 2.217 ;
      RECT 40.805 2.063 40.815 2.212 ;
      RECT 40.785 2.058 40.805 2.207 ;
      RECT 40.75 2.053 40.785 2.2 ;
      RECT 40.69 2.048 40.75 2.193 ;
      RECT 40.677 2.044 40.69 2.191 ;
      RECT 40.591 2.039 40.677 2.188 ;
      RECT 40.505 2.029 40.591 2.184 ;
      RECT 40.464 2.022 40.505 2.181 ;
      RECT 40.378 2.015 40.464 2.178 ;
      RECT 40.292 2.005 40.378 2.174 ;
      RECT 40.206 1.995 40.292 2.169 ;
      RECT 40.12 1.985 40.206 2.165 ;
      RECT 40.11 1.97 40.12 2.163 ;
      RECT 40.1 1.955 40.11 2.163 ;
      RECT 40.035 1.95 40.1 2.162 ;
      RECT 39.87 1.947 39.915 2.155 ;
      RECT 41.115 2.852 41.12 3.043 ;
      RECT 41.11 2.847 41.115 3.05 ;
      RECT 41.096 2.845 41.11 3.056 ;
      RECT 41.01 2.845 41.096 3.058 ;
      RECT 41.006 2.845 41.01 3.061 ;
      RECT 40.92 2.845 41.006 3.079 ;
      RECT 40.91 2.85 40.92 3.098 ;
      RECT 40.9 2.905 40.91 3.102 ;
      RECT 40.875 2.92 40.9 3.109 ;
      RECT 40.835 2.94 40.875 3.122 ;
      RECT 40.83 2.952 40.835 3.132 ;
      RECT 40.815 2.958 40.83 3.137 ;
      RECT 40.81 2.963 40.815 3.141 ;
      RECT 40.79 2.97 40.81 3.146 ;
      RECT 40.72 2.995 40.79 3.163 ;
      RECT 40.68 3.023 40.72 3.183 ;
      RECT 40.675 3.033 40.68 3.191 ;
      RECT 40.655 3.04 40.675 3.193 ;
      RECT 40.65 3.047 40.655 3.196 ;
      RECT 40.62 3.055 40.65 3.199 ;
      RECT 40.615 3.06 40.62 3.203 ;
      RECT 40.541 3.064 40.615 3.211 ;
      RECT 40.455 3.073 40.541 3.227 ;
      RECT 40.451 3.078 40.455 3.236 ;
      RECT 40.365 3.083 40.451 3.246 ;
      RECT 40.325 3.091 40.365 3.258 ;
      RECT 40.275 3.097 40.325 3.265 ;
      RECT 40.19 3.106 40.275 3.28 ;
      RECT 40.115 3.117 40.19 3.298 ;
      RECT 40.08 3.124 40.115 3.308 ;
      RECT 40.005 3.132 40.08 3.313 ;
      RECT 39.95 3.141 40.005 3.313 ;
      RECT 39.925 3.146 39.95 3.311 ;
      RECT 39.915 3.149 39.925 3.309 ;
      RECT 39.88 3.151 39.915 3.307 ;
      RECT 39.85 3.153 39.88 3.303 ;
      RECT 39.805 3.152 39.85 3.299 ;
      RECT 39.785 3.147 39.805 3.296 ;
      RECT 39.735 3.132 39.785 3.293 ;
      RECT 39.725 3.117 39.735 3.288 ;
      RECT 39.675 3.102 39.725 3.278 ;
      RECT 39.625 3.077 39.675 3.258 ;
      RECT 39.615 3.062 39.625 3.24 ;
      RECT 39.61 3.06 39.615 3.234 ;
      RECT 39.59 3.055 39.61 3.229 ;
      RECT 39.585 3.047 39.59 3.223 ;
      RECT 39.57 3.041 39.585 3.216 ;
      RECT 39.565 3.036 39.57 3.208 ;
      RECT 39.545 3.031 39.565 3.2 ;
      RECT 39.53 3.024 39.545 3.193 ;
      RECT 39.515 3.018 39.53 3.184 ;
      RECT 39.51 3.012 39.515 3.177 ;
      RECT 39.465 2.987 39.51 3.163 ;
      RECT 39.45 2.957 39.465 3.145 ;
      RECT 39.435 2.94 39.45 3.136 ;
      RECT 39.41 2.92 39.435 3.124 ;
      RECT 39.37 2.89 39.41 3.104 ;
      RECT 39.36 2.86 39.37 3.089 ;
      RECT 39.345 2.85 39.36 3.082 ;
      RECT 39.29 2.815 39.345 3.061 ;
      RECT 39.275 2.778 39.29 3.04 ;
      RECT 39.265 2.765 39.275 3.032 ;
      RECT 39.215 2.735 39.265 3.014 ;
      RECT 39.2 2.665 39.215 2.995 ;
      RECT 39.155 2.665 39.2 2.978 ;
      RECT 39.13 2.665 39.155 2.96 ;
      RECT 39.12 2.665 39.13 2.953 ;
      RECT 39.041 2.665 39.12 2.946 ;
      RECT 38.955 2.665 39.041 2.938 ;
      RECT 38.94 2.697 38.955 2.933 ;
      RECT 38.865 2.707 38.94 2.929 ;
      RECT 38.845 2.717 38.865 2.924 ;
      RECT 38.82 2.717 38.845 2.921 ;
      RECT 38.81 2.707 38.82 2.92 ;
      RECT 38.8 2.68 38.81 2.919 ;
      RECT 38.76 2.675 38.8 2.917 ;
      RECT 38.715 2.675 38.76 2.913 ;
      RECT 38.69 2.675 38.715 2.908 ;
      RECT 38.64 2.675 38.69 2.895 ;
      RECT 38.6 2.68 38.61 2.88 ;
      RECT 38.61 2.675 38.64 2.885 ;
      RECT 40.595 2.455 40.855 2.715 ;
      RECT 40.59 2.477 40.855 2.673 ;
      RECT 39.83 2.305 40.05 2.67 ;
      RECT 39.812 2.392 40.05 2.669 ;
      RECT 39.795 2.397 40.05 2.666 ;
      RECT 39.795 2.397 40.07 2.665 ;
      RECT 39.765 2.407 40.07 2.663 ;
      RECT 39.76 2.422 40.07 2.659 ;
      RECT 39.76 2.422 40.075 2.658 ;
      RECT 39.755 2.48 40.075 2.656 ;
      RECT 39.755 2.48 40.085 2.653 ;
      RECT 39.75 2.545 40.085 2.648 ;
      RECT 39.83 2.305 40.09 2.565 ;
      RECT 38.575 2.135 38.835 2.395 ;
      RECT 38.575 2.178 38.921 2.369 ;
      RECT 38.575 2.178 38.965 2.368 ;
      RECT 38.575 2.178 38.985 2.366 ;
      RECT 38.575 2.178 39.085 2.365 ;
      RECT 38.575 2.178 39.105 2.363 ;
      RECT 38.575 2.178 39.115 2.358 ;
      RECT 38.985 2.145 39.175 2.355 ;
      RECT 38.985 2.147 39.18 2.353 ;
      RECT 38.975 2.152 39.185 2.345 ;
      RECT 38.921 2.176 39.185 2.345 ;
      RECT 38.965 2.17 38.975 2.367 ;
      RECT 38.975 2.15 39.18 2.353 ;
      RECT 37.93 3.21 38.135 3.44 ;
      RECT 37.87 3.16 37.925 3.42 ;
      RECT 37.93 3.16 38.13 3.44 ;
      RECT 38.9 3.475 38.905 3.502 ;
      RECT 38.89 3.385 38.9 3.507 ;
      RECT 38.885 3.307 38.89 3.513 ;
      RECT 38.875 3.297 38.885 3.52 ;
      RECT 38.87 3.287 38.875 3.526 ;
      RECT 38.86 3.282 38.87 3.528 ;
      RECT 38.845 3.274 38.86 3.536 ;
      RECT 38.83 3.265 38.845 3.548 ;
      RECT 38.82 3.257 38.83 3.558 ;
      RECT 38.785 3.175 38.82 3.576 ;
      RECT 38.75 3.175 38.785 3.595 ;
      RECT 38.735 3.175 38.75 3.603 ;
      RECT 38.68 3.175 38.735 3.603 ;
      RECT 38.646 3.175 38.68 3.594 ;
      RECT 38.56 3.175 38.646 3.57 ;
      RECT 38.55 3.235 38.56 3.552 ;
      RECT 38.51 3.237 38.55 3.543 ;
      RECT 38.505 3.239 38.51 3.533 ;
      RECT 38.485 3.241 38.505 3.528 ;
      RECT 38.475 3.244 38.485 3.523 ;
      RECT 38.465 3.245 38.475 3.518 ;
      RECT 38.441 3.246 38.465 3.51 ;
      RECT 38.355 3.251 38.441 3.488 ;
      RECT 38.3 3.25 38.355 3.461 ;
      RECT 38.285 3.243 38.3 3.448 ;
      RECT 38.25 3.238 38.285 3.444 ;
      RECT 38.195 3.23 38.25 3.443 ;
      RECT 38.135 3.217 38.195 3.441 ;
      RECT 37.925 3.16 37.93 3.428 ;
      RECT 38 2.53 38.185 2.74 ;
      RECT 37.99 2.535 38.2 2.733 ;
      RECT 38.03 2.44 38.29 2.7 ;
      RECT 37.985 2.597 38.29 2.623 ;
      RECT 37.33 2.39 37.335 3.19 ;
      RECT 37.275 2.44 37.305 3.19 ;
      RECT 37.265 2.44 37.27 2.75 ;
      RECT 37.25 2.44 37.255 2.745 ;
      RECT 36.795 2.485 36.81 2.7 ;
      RECT 36.725 2.485 36.81 2.695 ;
      RECT 37.99 2.065 38.06 2.275 ;
      RECT 38.06 2.072 38.07 2.27 ;
      RECT 37.956 2.065 37.99 2.282 ;
      RECT 37.87 2.065 37.956 2.306 ;
      RECT 37.86 2.07 37.87 2.325 ;
      RECT 37.855 2.082 37.86 2.328 ;
      RECT 37.84 2.097 37.855 2.332 ;
      RECT 37.835 2.115 37.84 2.336 ;
      RECT 37.795 2.125 37.835 2.345 ;
      RECT 37.78 2.132 37.795 2.357 ;
      RECT 37.765 2.137 37.78 2.362 ;
      RECT 37.75 2.14 37.765 2.367 ;
      RECT 37.74 2.142 37.75 2.371 ;
      RECT 37.705 2.149 37.74 2.379 ;
      RECT 37.67 2.157 37.705 2.393 ;
      RECT 37.66 2.163 37.67 2.402 ;
      RECT 37.655 2.165 37.66 2.404 ;
      RECT 37.635 2.168 37.655 2.41 ;
      RECT 37.605 2.175 37.635 2.421 ;
      RECT 37.595 2.181 37.605 2.428 ;
      RECT 37.57 2.184 37.595 2.435 ;
      RECT 37.56 2.188 37.57 2.443 ;
      RECT 37.555 2.189 37.56 2.465 ;
      RECT 37.55 2.19 37.555 2.48 ;
      RECT 37.545 2.191 37.55 2.495 ;
      RECT 37.54 2.192 37.545 2.51 ;
      RECT 37.535 2.193 37.54 2.54 ;
      RECT 37.525 2.195 37.535 2.573 ;
      RECT 37.51 2.199 37.525 2.62 ;
      RECT 37.5 2.202 37.51 2.665 ;
      RECT 37.495 2.205 37.5 2.693 ;
      RECT 37.485 2.207 37.495 2.72 ;
      RECT 37.48 2.21 37.485 2.755 ;
      RECT 37.45 2.215 37.48 2.813 ;
      RECT 37.445 2.22 37.45 2.898 ;
      RECT 37.44 2.222 37.445 2.933 ;
      RECT 37.435 2.224 37.44 3.015 ;
      RECT 37.43 2.226 37.435 3.103 ;
      RECT 37.42 2.228 37.43 3.185 ;
      RECT 37.405 2.242 37.42 3.19 ;
      RECT 37.37 2.287 37.405 3.19 ;
      RECT 37.36 2.327 37.37 3.19 ;
      RECT 37.345 2.355 37.36 3.19 ;
      RECT 37.34 2.372 37.345 3.19 ;
      RECT 37.335 2.38 37.34 3.19 ;
      RECT 37.325 2.395 37.33 3.19 ;
      RECT 37.32 2.402 37.325 3.19 ;
      RECT 37.31 2.422 37.32 3.19 ;
      RECT 37.305 2.435 37.31 3.19 ;
      RECT 37.27 2.44 37.275 2.775 ;
      RECT 37.255 2.83 37.275 3.19 ;
      RECT 37.255 2.44 37.265 2.748 ;
      RECT 37.25 2.87 37.255 3.19 ;
      RECT 37.2 2.44 37.25 2.743 ;
      RECT 37.245 2.907 37.25 3.19 ;
      RECT 37.235 2.93 37.245 3.19 ;
      RECT 37.23 2.975 37.235 3.19 ;
      RECT 37.22 2.985 37.23 3.183 ;
      RECT 37.146 2.44 37.2 2.737 ;
      RECT 37.06 2.44 37.146 2.73 ;
      RECT 37.011 2.487 37.06 2.723 ;
      RECT 36.925 2.495 37.011 2.716 ;
      RECT 36.91 2.492 36.925 2.711 ;
      RECT 36.896 2.485 36.91 2.71 ;
      RECT 36.81 2.485 36.896 2.705 ;
      RECT 36.715 2.49 36.725 2.69 ;
      RECT 36.305 1.92 36.32 2.32 ;
      RECT 36.5 1.92 36.505 2.18 ;
      RECT 36.245 1.92 36.29 2.18 ;
      RECT 36.7 3.225 36.705 3.43 ;
      RECT 36.695 3.215 36.7 3.435 ;
      RECT 36.69 3.202 36.695 3.44 ;
      RECT 36.685 3.182 36.69 3.44 ;
      RECT 36.66 3.135 36.685 3.44 ;
      RECT 36.625 3.05 36.66 3.44 ;
      RECT 36.62 2.987 36.625 3.44 ;
      RECT 36.615 2.972 36.62 3.44 ;
      RECT 36.6 2.932 36.615 3.44 ;
      RECT 36.595 2.907 36.6 3.44 ;
      RECT 36.585 2.89 36.595 3.44 ;
      RECT 36.55 2.812 36.585 3.44 ;
      RECT 36.545 2.755 36.55 3.44 ;
      RECT 36.54 2.742 36.545 3.44 ;
      RECT 36.53 2.72 36.54 3.44 ;
      RECT 36.52 2.685 36.53 3.44 ;
      RECT 36.51 2.655 36.52 3.44 ;
      RECT 36.5 2.57 36.51 3.083 ;
      RECT 36.507 3.215 36.51 3.44 ;
      RECT 36.505 3.225 36.507 3.44 ;
      RECT 36.495 3.235 36.505 3.435 ;
      RECT 36.49 1.92 36.5 2.315 ;
      RECT 36.495 2.447 36.5 3.058 ;
      RECT 36.49 2.345 36.495 3.041 ;
      RECT 36.48 1.92 36.49 3.017 ;
      RECT 36.475 1.92 36.48 2.988 ;
      RECT 36.47 1.92 36.475 2.978 ;
      RECT 36.45 1.92 36.47 2.94 ;
      RECT 36.445 1.92 36.45 2.898 ;
      RECT 36.44 1.92 36.445 2.878 ;
      RECT 36.41 1.92 36.44 2.828 ;
      RECT 36.4 1.92 36.41 2.775 ;
      RECT 36.395 1.92 36.4 2.748 ;
      RECT 36.39 1.92 36.395 2.733 ;
      RECT 36.38 1.92 36.39 2.71 ;
      RECT 36.37 1.92 36.38 2.685 ;
      RECT 36.365 1.92 36.37 2.625 ;
      RECT 36.355 1.92 36.365 2.563 ;
      RECT 36.35 1.92 36.355 2.483 ;
      RECT 36.345 1.92 36.35 2.448 ;
      RECT 36.34 1.92 36.345 2.423 ;
      RECT 36.335 1.92 36.34 2.408 ;
      RECT 36.33 1.92 36.335 2.378 ;
      RECT 36.325 1.92 36.33 2.355 ;
      RECT 36.32 1.92 36.325 2.328 ;
      RECT 36.29 1.92 36.305 2.315 ;
      RECT 35.445 3.455 35.63 3.665 ;
      RECT 35.435 3.46 35.645 3.658 ;
      RECT 35.435 3.46 35.665 3.63 ;
      RECT 35.435 3.46 35.68 3.609 ;
      RECT 35.435 3.46 35.695 3.607 ;
      RECT 35.435 3.46 35.705 3.606 ;
      RECT 35.435 3.46 35.735 3.603 ;
      RECT 36.085 3.305 36.345 3.565 ;
      RECT 36.045 3.352 36.345 3.548 ;
      RECT 36.036 3.36 36.045 3.551 ;
      RECT 35.63 3.453 36.345 3.548 ;
      RECT 35.95 3.378 36.036 3.558 ;
      RECT 35.645 3.45 36.345 3.548 ;
      RECT 35.891 3.4 35.95 3.57 ;
      RECT 35.665 3.446 36.345 3.548 ;
      RECT 35.805 3.412 35.891 3.581 ;
      RECT 35.68 3.442 36.345 3.548 ;
      RECT 35.75 3.425 35.805 3.593 ;
      RECT 35.695 3.44 36.345 3.548 ;
      RECT 35.735 3.431 35.75 3.599 ;
      RECT 35.705 3.436 36.345 3.548 ;
      RECT 35.85 2.96 36.11 3.22 ;
      RECT 35.85 2.98 36.22 3.19 ;
      RECT 35.85 2.985 36.23 3.185 ;
      RECT 36.041 2.399 36.12 2.63 ;
      RECT 35.955 2.402 36.17 2.625 ;
      RECT 35.95 2.402 36.17 2.62 ;
      RECT 35.95 2.407 36.18 2.618 ;
      RECT 35.925 2.407 36.18 2.615 ;
      RECT 35.925 2.415 36.19 2.613 ;
      RECT 35.805 2.35 36.065 2.61 ;
      RECT 35.805 2.397 36.115 2.61 ;
      RECT 35.06 2.97 35.065 3.23 ;
      RECT 34.89 2.74 34.895 3.23 ;
      RECT 34.775 2.98 34.78 3.205 ;
      RECT 35.485 2.075 35.49 2.285 ;
      RECT 35.49 2.08 35.505 2.28 ;
      RECT 35.425 2.075 35.485 2.293 ;
      RECT 35.41 2.075 35.425 2.303 ;
      RECT 35.36 2.075 35.41 2.32 ;
      RECT 35.34 2.075 35.36 2.343 ;
      RECT 35.325 2.075 35.34 2.355 ;
      RECT 35.305 2.075 35.325 2.365 ;
      RECT 35.295 2.08 35.305 2.374 ;
      RECT 35.29 2.09 35.295 2.379 ;
      RECT 35.285 2.102 35.29 2.383 ;
      RECT 35.275 2.125 35.285 2.388 ;
      RECT 35.27 2.14 35.275 2.392 ;
      RECT 35.265 2.157 35.27 2.395 ;
      RECT 35.26 2.165 35.265 2.398 ;
      RECT 35.25 2.17 35.26 2.402 ;
      RECT 35.245 2.177 35.25 2.407 ;
      RECT 35.235 2.182 35.245 2.411 ;
      RECT 35.21 2.194 35.235 2.422 ;
      RECT 35.19 2.211 35.21 2.438 ;
      RECT 35.165 2.228 35.19 2.46 ;
      RECT 35.13 2.251 35.165 2.518 ;
      RECT 35.11 2.273 35.13 2.58 ;
      RECT 35.105 2.283 35.11 2.615 ;
      RECT 35.095 2.29 35.105 2.653 ;
      RECT 35.09 2.297 35.095 2.673 ;
      RECT 35.085 2.308 35.09 2.71 ;
      RECT 35.08 2.316 35.085 2.775 ;
      RECT 35.07 2.327 35.08 2.828 ;
      RECT 35.065 2.345 35.07 2.898 ;
      RECT 35.06 2.355 35.065 2.935 ;
      RECT 35.055 2.365 35.06 3.23 ;
      RECT 35.05 2.377 35.055 3.23 ;
      RECT 35.045 2.387 35.05 3.23 ;
      RECT 35.035 2.397 35.045 3.23 ;
      RECT 35.025 2.42 35.035 3.23 ;
      RECT 35.01 2.455 35.025 3.23 ;
      RECT 34.97 2.517 35.01 3.23 ;
      RECT 34.965 2.57 34.97 3.23 ;
      RECT 34.94 2.605 34.965 3.23 ;
      RECT 34.925 2.65 34.94 3.23 ;
      RECT 34.92 2.672 34.925 3.23 ;
      RECT 34.91 2.685 34.92 3.23 ;
      RECT 34.9 2.71 34.91 3.23 ;
      RECT 34.895 2.732 34.9 3.23 ;
      RECT 34.87 2.77 34.89 3.23 ;
      RECT 34.83 2.827 34.87 3.23 ;
      RECT 34.825 2.877 34.83 3.23 ;
      RECT 34.82 2.895 34.825 3.23 ;
      RECT 34.815 2.907 34.82 3.23 ;
      RECT 34.805 2.925 34.815 3.23 ;
      RECT 34.795 2.945 34.805 3.205 ;
      RECT 34.79 2.962 34.795 3.205 ;
      RECT 34.78 2.975 34.79 3.205 ;
      RECT 34.75 2.985 34.775 3.205 ;
      RECT 34.74 2.992 34.75 3.205 ;
      RECT 34.725 3.002 34.74 3.2 ;
      RECT 33.825 7.77 34.115 8 ;
      RECT 33.885 6.29 34.055 8 ;
      RECT 33.875 6.66 34.23 7.015 ;
      RECT 33.825 6.29 34.115 6.52 ;
      RECT 33.42 2.395 33.525 2.965 ;
      RECT 33.42 2.73 33.745 2.96 ;
      RECT 33.42 2.76 33.915 2.93 ;
      RECT 33.42 2.395 33.61 2.96 ;
      RECT 32.835 2.36 33.125 2.59 ;
      RECT 32.835 2.395 33.61 2.565 ;
      RECT 32.895 0.88 33.065 2.59 ;
      RECT 32.835 0.88 33.125 1.11 ;
      RECT 32.835 7.77 33.125 8 ;
      RECT 32.895 6.29 33.065 8 ;
      RECT 32.835 6.29 33.125 6.52 ;
      RECT 32.835 6.325 33.69 6.485 ;
      RECT 33.52 5.92 33.69 6.485 ;
      RECT 32.835 6.32 33.23 6.485 ;
      RECT 33.455 5.92 33.745 6.15 ;
      RECT 33.455 5.95 33.915 6.12 ;
      RECT 32.465 2.73 32.755 2.96 ;
      RECT 32.465 2.76 32.925 2.93 ;
      RECT 32.53 1.655 32.695 2.96 ;
      RECT 31.045 1.625 31.335 1.855 ;
      RECT 31.045 1.655 32.695 1.825 ;
      RECT 31.105 0.885 31.275 1.855 ;
      RECT 31.045 0.885 31.335 1.115 ;
      RECT 31.045 7.765 31.335 7.995 ;
      RECT 31.105 7.025 31.275 7.995 ;
      RECT 31.105 7.12 32.695 7.29 ;
      RECT 32.525 5.92 32.695 7.29 ;
      RECT 31.045 7.025 31.335 7.255 ;
      RECT 32.465 5.92 32.755 6.15 ;
      RECT 32.465 5.95 32.925 6.12 ;
      RECT 31.475 1.965 31.825 2.315 ;
      RECT 29.14 2.025 31.825 2.195 ;
      RECT 29.14 1.34 29.31 2.195 ;
      RECT 29.04 1.34 29.39 1.69 ;
      RECT 31.5 6.655 31.825 6.98 ;
      RECT 26.925 6.61 27.275 6.96 ;
      RECT 31.475 6.655 31.825 6.885 ;
      RECT 26.695 6.655 27.275 6.885 ;
      RECT 26.525 6.685 31.825 6.855 ;
      RECT 30.7 2.365 31.02 2.685 ;
      RECT 30.67 2.365 31.02 2.595 ;
      RECT 30.5 2.395 31.02 2.565 ;
      RECT 30.7 6.255 31.02 6.545 ;
      RECT 30.67 6.285 31.02 6.515 ;
      RECT 30.5 6.315 31.02 6.485 ;
      RECT 27.335 2.465 27.52 2.675 ;
      RECT 27.325 2.47 27.535 2.668 ;
      RECT 27.325 2.47 27.621 2.645 ;
      RECT 27.325 2.47 27.68 2.62 ;
      RECT 27.325 2.47 27.735 2.6 ;
      RECT 27.325 2.47 27.745 2.588 ;
      RECT 27.325 2.47 27.94 2.527 ;
      RECT 27.325 2.47 27.97 2.51 ;
      RECT 27.325 2.47 27.99 2.5 ;
      RECT 27.87 2.235 28.13 2.495 ;
      RECT 27.855 2.325 27.87 2.542 ;
      RECT 27.39 2.457 28.13 2.495 ;
      RECT 27.841 2.336 27.855 2.548 ;
      RECT 27.43 2.45 28.13 2.495 ;
      RECT 27.755 2.376 27.841 2.567 ;
      RECT 27.68 2.437 28.13 2.495 ;
      RECT 27.75 2.412 27.755 2.584 ;
      RECT 27.735 2.422 28.13 2.495 ;
      RECT 27.745 2.417 27.75 2.586 ;
      RECT 28.04 2.922 28.045 3.014 ;
      RECT 28.035 2.9 28.04 3.031 ;
      RECT 28.03 2.89 28.035 3.043 ;
      RECT 28.02 2.881 28.03 3.053 ;
      RECT 28.015 2.876 28.02 3.061 ;
      RECT 28.01 2.735 28.015 3.064 ;
      RECT 27.976 2.735 28.01 3.075 ;
      RECT 27.89 2.735 27.976 3.11 ;
      RECT 27.81 2.735 27.89 3.158 ;
      RECT 27.781 2.735 27.81 3.182 ;
      RECT 27.695 2.735 27.781 3.188 ;
      RECT 27.69 2.919 27.695 3.193 ;
      RECT 27.655 2.93 27.69 3.196 ;
      RECT 27.63 2.945 27.655 3.2 ;
      RECT 27.616 2.954 27.63 3.202 ;
      RECT 27.53 2.981 27.616 3.208 ;
      RECT 27.465 3.022 27.53 3.217 ;
      RECT 27.45 3.042 27.465 3.222 ;
      RECT 27.42 3.052 27.45 3.225 ;
      RECT 27.415 3.062 27.42 3.228 ;
      RECT 27.385 3.067 27.415 3.23 ;
      RECT 27.365 3.072 27.385 3.234 ;
      RECT 27.28 3.075 27.365 3.241 ;
      RECT 27.265 3.072 27.28 3.247 ;
      RECT 27.255 3.069 27.265 3.249 ;
      RECT 27.235 3.066 27.255 3.251 ;
      RECT 27.215 3.062 27.235 3.252 ;
      RECT 27.2 3.058 27.215 3.254 ;
      RECT 27.19 3.055 27.2 3.255 ;
      RECT 27.15 3.049 27.19 3.253 ;
      RECT 27.14 3.044 27.15 3.251 ;
      RECT 27.125 3.041 27.14 3.247 ;
      RECT 27.1 3.036 27.125 3.24 ;
      RECT 27.05 3.027 27.1 3.228 ;
      RECT 26.98 3.013 27.05 3.21 ;
      RECT 26.922 2.998 26.98 3.192 ;
      RECT 26.836 2.981 26.922 3.172 ;
      RECT 26.75 2.96 26.836 3.147 ;
      RECT 26.7 2.945 26.75 3.128 ;
      RECT 26.696 2.939 26.7 3.12 ;
      RECT 26.61 2.929 26.696 3.107 ;
      RECT 26.575 2.914 26.61 3.09 ;
      RECT 26.56 2.907 26.575 3.083 ;
      RECT 26.5 2.895 26.56 3.071 ;
      RECT 26.48 2.882 26.5 3.059 ;
      RECT 26.44 2.873 26.48 3.051 ;
      RECT 26.435 2.865 26.44 3.044 ;
      RECT 26.355 2.855 26.435 3.03 ;
      RECT 26.34 2.842 26.355 3.015 ;
      RECT 26.335 2.84 26.34 3.013 ;
      RECT 26.256 2.828 26.335 3 ;
      RECT 26.17 2.803 26.256 2.975 ;
      RECT 26.155 2.772 26.17 2.96 ;
      RECT 26.14 2.747 26.155 2.956 ;
      RECT 26.125 2.74 26.14 2.952 ;
      RECT 25.95 2.745 25.955 2.948 ;
      RECT 25.945 2.75 25.95 2.943 ;
      RECT 25.955 2.74 26.125 2.95 ;
      RECT 26.67 2.5 26.775 2.76 ;
      RECT 27.485 2.025 27.49 2.25 ;
      RECT 27.615 2.025 27.67 2.235 ;
      RECT 27.67 2.03 27.68 2.228 ;
      RECT 27.576 2.025 27.615 2.238 ;
      RECT 27.49 2.025 27.576 2.245 ;
      RECT 27.47 2.03 27.485 2.251 ;
      RECT 27.46 2.07 27.47 2.253 ;
      RECT 27.43 2.08 27.46 2.255 ;
      RECT 27.425 2.085 27.43 2.257 ;
      RECT 27.4 2.09 27.425 2.259 ;
      RECT 27.385 2.095 27.4 2.261 ;
      RECT 27.37 2.097 27.385 2.263 ;
      RECT 27.365 2.102 27.37 2.265 ;
      RECT 27.315 2.11 27.365 2.268 ;
      RECT 27.29 2.119 27.315 2.273 ;
      RECT 27.28 2.126 27.29 2.278 ;
      RECT 27.275 2.129 27.28 2.282 ;
      RECT 27.255 2.132 27.275 2.291 ;
      RECT 27.225 2.14 27.255 2.311 ;
      RECT 27.196 2.153 27.225 2.333 ;
      RECT 27.11 2.187 27.196 2.377 ;
      RECT 27.105 2.213 27.11 2.415 ;
      RECT 27.1 2.217 27.105 2.424 ;
      RECT 27.065 2.23 27.1 2.457 ;
      RECT 27.055 2.244 27.065 2.495 ;
      RECT 27.05 2.248 27.055 2.508 ;
      RECT 27.045 2.252 27.05 2.513 ;
      RECT 27.035 2.26 27.045 2.525 ;
      RECT 27.03 2.267 27.035 2.54 ;
      RECT 27.005 2.28 27.03 2.565 ;
      RECT 26.965 2.309 27.005 2.62 ;
      RECT 26.95 2.334 26.965 2.675 ;
      RECT 26.94 2.345 26.95 2.698 ;
      RECT 26.935 2.352 26.94 2.71 ;
      RECT 26.93 2.356 26.935 2.718 ;
      RECT 26.875 2.384 26.93 2.76 ;
      RECT 26.855 2.42 26.875 2.76 ;
      RECT 26.84 2.435 26.855 2.76 ;
      RECT 26.785 2.467 26.84 2.76 ;
      RECT 26.775 2.497 26.785 2.76 ;
      RECT 26.385 2.112 26.57 2.35 ;
      RECT 26.37 2.114 26.58 2.345 ;
      RECT 26.255 2.06 26.515 2.32 ;
      RECT 26.25 2.097 26.515 2.274 ;
      RECT 26.245 2.107 26.515 2.271 ;
      RECT 26.24 2.147 26.58 2.265 ;
      RECT 26.235 2.18 26.58 2.255 ;
      RECT 26.245 2.122 26.595 2.193 ;
      RECT 26.542 3.22 26.555 3.75 ;
      RECT 26.456 3.22 26.555 3.749 ;
      RECT 26.456 3.22 26.56 3.748 ;
      RECT 26.37 3.22 26.56 3.746 ;
      RECT 26.365 3.22 26.56 3.743 ;
      RECT 26.365 3.22 26.57 3.741 ;
      RECT 26.36 3.512 26.57 3.738 ;
      RECT 26.36 3.522 26.575 3.735 ;
      RECT 26.36 3.59 26.58 3.731 ;
      RECT 26.35 3.595 26.58 3.73 ;
      RECT 26.35 3.687 26.585 3.727 ;
      RECT 26.335 3.22 26.595 3.48 ;
      RECT 26.265 7.765 26.555 7.995 ;
      RECT 26.325 7.025 26.495 7.995 ;
      RECT 26.24 7.055 26.58 7.4 ;
      RECT 26.265 7.025 26.555 7.4 ;
      RECT 25.565 2.21 25.61 3.745 ;
      RECT 25.765 2.21 25.795 2.425 ;
      RECT 24.14 1.95 24.26 2.16 ;
      RECT 23.8 1.9 24.06 2.16 ;
      RECT 23.8 1.945 24.095 2.15 ;
      RECT 25.805 2.226 25.81 2.28 ;
      RECT 25.8 2.219 25.805 2.413 ;
      RECT 25.795 2.213 25.8 2.42 ;
      RECT 25.75 2.21 25.765 2.433 ;
      RECT 25.745 2.21 25.75 2.455 ;
      RECT 25.74 2.21 25.745 2.503 ;
      RECT 25.735 2.21 25.74 2.523 ;
      RECT 25.725 2.21 25.735 2.63 ;
      RECT 25.72 2.21 25.725 2.693 ;
      RECT 25.715 2.21 25.72 2.75 ;
      RECT 25.71 2.21 25.715 2.758 ;
      RECT 25.695 2.21 25.71 2.865 ;
      RECT 25.685 2.21 25.695 3 ;
      RECT 25.675 2.21 25.685 3.11 ;
      RECT 25.665 2.21 25.675 3.167 ;
      RECT 25.66 2.21 25.665 3.207 ;
      RECT 25.655 2.21 25.66 3.243 ;
      RECT 25.645 2.21 25.655 3.283 ;
      RECT 25.64 2.21 25.645 3.325 ;
      RECT 25.62 2.21 25.64 3.39 ;
      RECT 25.625 3.535 25.63 3.715 ;
      RECT 25.62 3.517 25.625 3.723 ;
      RECT 25.615 2.21 25.62 3.453 ;
      RECT 25.615 3.497 25.62 3.73 ;
      RECT 25.61 2.21 25.615 3.74 ;
      RECT 25.555 2.21 25.565 2.51 ;
      RECT 25.56 2.757 25.565 3.745 ;
      RECT 25.555 2.822 25.56 3.745 ;
      RECT 25.55 2.211 25.555 2.5 ;
      RECT 25.545 2.887 25.555 3.745 ;
      RECT 25.54 2.212 25.55 2.49 ;
      RECT 25.53 3 25.545 3.745 ;
      RECT 25.535 2.213 25.54 2.48 ;
      RECT 25.515 2.214 25.535 2.458 ;
      RECT 25.52 3.097 25.53 3.745 ;
      RECT 25.515 3.172 25.52 3.745 ;
      RECT 25.505 2.213 25.515 2.435 ;
      RECT 25.51 3.215 25.515 3.745 ;
      RECT 25.505 3.242 25.51 3.745 ;
      RECT 25.495 2.211 25.505 2.423 ;
      RECT 25.5 3.285 25.505 3.745 ;
      RECT 25.495 3.312 25.5 3.745 ;
      RECT 25.485 2.21 25.495 2.41 ;
      RECT 25.49 3.327 25.495 3.745 ;
      RECT 25.45 3.385 25.49 3.745 ;
      RECT 25.48 2.209 25.485 2.395 ;
      RECT 25.475 2.207 25.48 2.388 ;
      RECT 25.465 2.204 25.475 2.378 ;
      RECT 25.46 2.201 25.465 2.363 ;
      RECT 25.445 2.197 25.46 2.356 ;
      RECT 25.44 3.44 25.45 3.745 ;
      RECT 25.44 2.194 25.445 2.351 ;
      RECT 25.425 2.19 25.44 2.345 ;
      RECT 25.435 3.457 25.44 3.745 ;
      RECT 25.425 3.52 25.435 3.745 ;
      RECT 25.345 2.175 25.425 2.325 ;
      RECT 25.42 3.527 25.425 3.74 ;
      RECT 25.415 3.535 25.42 3.73 ;
      RECT 25.335 2.161 25.345 2.309 ;
      RECT 25.32 2.157 25.335 2.307 ;
      RECT 25.31 2.152 25.32 2.303 ;
      RECT 25.285 2.145 25.31 2.295 ;
      RECT 25.28 2.14 25.285 2.29 ;
      RECT 25.27 2.14 25.28 2.288 ;
      RECT 25.26 2.138 25.27 2.286 ;
      RECT 25.23 2.13 25.26 2.28 ;
      RECT 25.215 2.122 25.23 2.273 ;
      RECT 25.195 2.117 25.215 2.266 ;
      RECT 25.19 2.113 25.195 2.261 ;
      RECT 25.16 2.106 25.19 2.255 ;
      RECT 25.135 2.097 25.16 2.245 ;
      RECT 25.105 2.09 25.135 2.237 ;
      RECT 25.08 2.08 25.105 2.228 ;
      RECT 25.065 2.072 25.08 2.222 ;
      RECT 25.04 2.067 25.065 2.217 ;
      RECT 25.03 2.063 25.04 2.212 ;
      RECT 25.01 2.058 25.03 2.207 ;
      RECT 24.975 2.053 25.01 2.2 ;
      RECT 24.915 2.048 24.975 2.193 ;
      RECT 24.902 2.044 24.915 2.191 ;
      RECT 24.816 2.039 24.902 2.188 ;
      RECT 24.73 2.029 24.816 2.184 ;
      RECT 24.689 2.022 24.73 2.181 ;
      RECT 24.603 2.015 24.689 2.178 ;
      RECT 24.517 2.005 24.603 2.174 ;
      RECT 24.431 1.995 24.517 2.169 ;
      RECT 24.345 1.985 24.431 2.165 ;
      RECT 24.335 1.97 24.345 2.163 ;
      RECT 24.325 1.955 24.335 2.163 ;
      RECT 24.26 1.95 24.325 2.162 ;
      RECT 24.095 1.947 24.14 2.155 ;
      RECT 25.34 2.852 25.345 3.043 ;
      RECT 25.335 2.847 25.34 3.05 ;
      RECT 25.321 2.845 25.335 3.056 ;
      RECT 25.235 2.845 25.321 3.058 ;
      RECT 25.231 2.845 25.235 3.061 ;
      RECT 25.145 2.845 25.231 3.079 ;
      RECT 25.135 2.85 25.145 3.098 ;
      RECT 25.125 2.905 25.135 3.102 ;
      RECT 25.1 2.92 25.125 3.109 ;
      RECT 25.06 2.94 25.1 3.122 ;
      RECT 25.055 2.952 25.06 3.132 ;
      RECT 25.04 2.958 25.055 3.137 ;
      RECT 25.035 2.963 25.04 3.141 ;
      RECT 25.015 2.97 25.035 3.146 ;
      RECT 24.945 2.995 25.015 3.163 ;
      RECT 24.905 3.023 24.945 3.183 ;
      RECT 24.9 3.033 24.905 3.191 ;
      RECT 24.88 3.04 24.9 3.193 ;
      RECT 24.875 3.047 24.88 3.196 ;
      RECT 24.845 3.055 24.875 3.199 ;
      RECT 24.84 3.06 24.845 3.203 ;
      RECT 24.766 3.064 24.84 3.211 ;
      RECT 24.68 3.073 24.766 3.227 ;
      RECT 24.676 3.078 24.68 3.236 ;
      RECT 24.59 3.083 24.676 3.246 ;
      RECT 24.55 3.091 24.59 3.258 ;
      RECT 24.5 3.097 24.55 3.265 ;
      RECT 24.415 3.106 24.5 3.28 ;
      RECT 24.34 3.117 24.415 3.298 ;
      RECT 24.305 3.124 24.34 3.308 ;
      RECT 24.23 3.132 24.305 3.313 ;
      RECT 24.175 3.141 24.23 3.313 ;
      RECT 24.15 3.146 24.175 3.311 ;
      RECT 24.14 3.149 24.15 3.309 ;
      RECT 24.105 3.151 24.14 3.307 ;
      RECT 24.075 3.153 24.105 3.303 ;
      RECT 24.03 3.152 24.075 3.299 ;
      RECT 24.01 3.147 24.03 3.296 ;
      RECT 23.96 3.132 24.01 3.293 ;
      RECT 23.95 3.117 23.96 3.288 ;
      RECT 23.9 3.102 23.95 3.278 ;
      RECT 23.85 3.077 23.9 3.258 ;
      RECT 23.84 3.062 23.85 3.24 ;
      RECT 23.835 3.06 23.84 3.234 ;
      RECT 23.815 3.055 23.835 3.229 ;
      RECT 23.81 3.047 23.815 3.223 ;
      RECT 23.795 3.041 23.81 3.216 ;
      RECT 23.79 3.036 23.795 3.208 ;
      RECT 23.77 3.031 23.79 3.2 ;
      RECT 23.755 3.024 23.77 3.193 ;
      RECT 23.74 3.018 23.755 3.184 ;
      RECT 23.735 3.012 23.74 3.177 ;
      RECT 23.69 2.987 23.735 3.163 ;
      RECT 23.675 2.957 23.69 3.145 ;
      RECT 23.66 2.94 23.675 3.136 ;
      RECT 23.635 2.92 23.66 3.124 ;
      RECT 23.595 2.89 23.635 3.104 ;
      RECT 23.585 2.86 23.595 3.089 ;
      RECT 23.57 2.85 23.585 3.082 ;
      RECT 23.515 2.815 23.57 3.061 ;
      RECT 23.5 2.778 23.515 3.04 ;
      RECT 23.49 2.765 23.5 3.032 ;
      RECT 23.44 2.735 23.49 3.014 ;
      RECT 23.425 2.665 23.44 2.995 ;
      RECT 23.38 2.665 23.425 2.978 ;
      RECT 23.355 2.665 23.38 2.96 ;
      RECT 23.345 2.665 23.355 2.953 ;
      RECT 23.266 2.665 23.345 2.946 ;
      RECT 23.18 2.665 23.266 2.938 ;
      RECT 23.165 2.697 23.18 2.933 ;
      RECT 23.09 2.707 23.165 2.929 ;
      RECT 23.07 2.717 23.09 2.924 ;
      RECT 23.045 2.717 23.07 2.921 ;
      RECT 23.035 2.707 23.045 2.92 ;
      RECT 23.025 2.68 23.035 2.919 ;
      RECT 22.985 2.675 23.025 2.917 ;
      RECT 22.94 2.675 22.985 2.913 ;
      RECT 22.915 2.675 22.94 2.908 ;
      RECT 22.865 2.675 22.915 2.895 ;
      RECT 22.825 2.68 22.835 2.88 ;
      RECT 22.835 2.675 22.865 2.885 ;
      RECT 24.82 2.455 25.08 2.715 ;
      RECT 24.815 2.477 25.08 2.673 ;
      RECT 24.055 2.305 24.275 2.67 ;
      RECT 24.037 2.392 24.275 2.669 ;
      RECT 24.02 2.397 24.275 2.666 ;
      RECT 24.02 2.397 24.295 2.665 ;
      RECT 23.99 2.407 24.295 2.663 ;
      RECT 23.985 2.422 24.295 2.659 ;
      RECT 23.985 2.422 24.3 2.658 ;
      RECT 23.98 2.48 24.3 2.656 ;
      RECT 23.98 2.48 24.31 2.653 ;
      RECT 23.975 2.545 24.31 2.648 ;
      RECT 24.055 2.305 24.315 2.565 ;
      RECT 22.8 2.135 23.06 2.395 ;
      RECT 22.8 2.178 23.146 2.369 ;
      RECT 22.8 2.178 23.19 2.368 ;
      RECT 22.8 2.178 23.21 2.366 ;
      RECT 22.8 2.178 23.31 2.365 ;
      RECT 22.8 2.178 23.33 2.363 ;
      RECT 22.8 2.178 23.34 2.358 ;
      RECT 23.21 2.145 23.4 2.355 ;
      RECT 23.21 2.147 23.405 2.353 ;
      RECT 23.2 2.152 23.41 2.345 ;
      RECT 23.146 2.176 23.41 2.345 ;
      RECT 23.19 2.17 23.2 2.367 ;
      RECT 23.2 2.15 23.405 2.353 ;
      RECT 22.155 3.21 22.36 3.44 ;
      RECT 22.095 3.16 22.15 3.42 ;
      RECT 22.155 3.16 22.355 3.44 ;
      RECT 23.125 3.475 23.13 3.502 ;
      RECT 23.115 3.385 23.125 3.507 ;
      RECT 23.11 3.307 23.115 3.513 ;
      RECT 23.1 3.297 23.11 3.52 ;
      RECT 23.095 3.287 23.1 3.526 ;
      RECT 23.085 3.282 23.095 3.528 ;
      RECT 23.07 3.274 23.085 3.536 ;
      RECT 23.055 3.265 23.07 3.548 ;
      RECT 23.045 3.257 23.055 3.558 ;
      RECT 23.01 3.175 23.045 3.576 ;
      RECT 22.975 3.175 23.01 3.595 ;
      RECT 22.96 3.175 22.975 3.603 ;
      RECT 22.905 3.175 22.96 3.603 ;
      RECT 22.871 3.175 22.905 3.594 ;
      RECT 22.785 3.175 22.871 3.57 ;
      RECT 22.775 3.235 22.785 3.552 ;
      RECT 22.735 3.237 22.775 3.543 ;
      RECT 22.73 3.239 22.735 3.533 ;
      RECT 22.71 3.241 22.73 3.528 ;
      RECT 22.7 3.244 22.71 3.523 ;
      RECT 22.69 3.245 22.7 3.518 ;
      RECT 22.666 3.246 22.69 3.51 ;
      RECT 22.58 3.251 22.666 3.488 ;
      RECT 22.525 3.25 22.58 3.461 ;
      RECT 22.51 3.243 22.525 3.448 ;
      RECT 22.475 3.238 22.51 3.444 ;
      RECT 22.42 3.23 22.475 3.443 ;
      RECT 22.36 3.217 22.42 3.441 ;
      RECT 22.15 3.16 22.155 3.428 ;
      RECT 22.225 2.53 22.41 2.74 ;
      RECT 22.215 2.535 22.425 2.733 ;
      RECT 22.255 2.44 22.515 2.7 ;
      RECT 22.21 2.597 22.515 2.623 ;
      RECT 21.555 2.39 21.56 3.19 ;
      RECT 21.5 2.44 21.53 3.19 ;
      RECT 21.49 2.44 21.495 2.75 ;
      RECT 21.475 2.44 21.48 2.745 ;
      RECT 21.02 2.485 21.035 2.7 ;
      RECT 20.95 2.485 21.035 2.695 ;
      RECT 22.215 2.065 22.285 2.275 ;
      RECT 22.285 2.072 22.295 2.27 ;
      RECT 22.181 2.065 22.215 2.282 ;
      RECT 22.095 2.065 22.181 2.306 ;
      RECT 22.085 2.07 22.095 2.325 ;
      RECT 22.08 2.082 22.085 2.328 ;
      RECT 22.065 2.097 22.08 2.332 ;
      RECT 22.06 2.115 22.065 2.336 ;
      RECT 22.02 2.125 22.06 2.345 ;
      RECT 22.005 2.132 22.02 2.357 ;
      RECT 21.99 2.137 22.005 2.362 ;
      RECT 21.975 2.14 21.99 2.367 ;
      RECT 21.965 2.142 21.975 2.371 ;
      RECT 21.93 2.149 21.965 2.379 ;
      RECT 21.895 2.157 21.93 2.393 ;
      RECT 21.885 2.163 21.895 2.402 ;
      RECT 21.88 2.165 21.885 2.404 ;
      RECT 21.86 2.168 21.88 2.41 ;
      RECT 21.83 2.175 21.86 2.421 ;
      RECT 21.82 2.181 21.83 2.428 ;
      RECT 21.795 2.184 21.82 2.435 ;
      RECT 21.785 2.188 21.795 2.443 ;
      RECT 21.78 2.189 21.785 2.465 ;
      RECT 21.775 2.19 21.78 2.48 ;
      RECT 21.77 2.191 21.775 2.495 ;
      RECT 21.765 2.192 21.77 2.51 ;
      RECT 21.76 2.193 21.765 2.54 ;
      RECT 21.75 2.195 21.76 2.573 ;
      RECT 21.735 2.199 21.75 2.62 ;
      RECT 21.725 2.202 21.735 2.665 ;
      RECT 21.72 2.205 21.725 2.693 ;
      RECT 21.71 2.207 21.72 2.72 ;
      RECT 21.705 2.21 21.71 2.755 ;
      RECT 21.675 2.215 21.705 2.813 ;
      RECT 21.67 2.22 21.675 2.898 ;
      RECT 21.665 2.222 21.67 2.933 ;
      RECT 21.66 2.224 21.665 3.015 ;
      RECT 21.655 2.226 21.66 3.103 ;
      RECT 21.645 2.228 21.655 3.185 ;
      RECT 21.63 2.242 21.645 3.19 ;
      RECT 21.595 2.287 21.63 3.19 ;
      RECT 21.585 2.327 21.595 3.19 ;
      RECT 21.57 2.355 21.585 3.19 ;
      RECT 21.565 2.372 21.57 3.19 ;
      RECT 21.56 2.38 21.565 3.19 ;
      RECT 21.55 2.395 21.555 3.19 ;
      RECT 21.545 2.402 21.55 3.19 ;
      RECT 21.535 2.422 21.545 3.19 ;
      RECT 21.53 2.435 21.535 3.19 ;
      RECT 21.495 2.44 21.5 2.775 ;
      RECT 21.48 2.83 21.5 3.19 ;
      RECT 21.48 2.44 21.49 2.748 ;
      RECT 21.475 2.87 21.48 3.19 ;
      RECT 21.425 2.44 21.475 2.743 ;
      RECT 21.47 2.907 21.475 3.19 ;
      RECT 21.46 2.93 21.47 3.19 ;
      RECT 21.455 2.975 21.46 3.19 ;
      RECT 21.445 2.985 21.455 3.183 ;
      RECT 21.371 2.44 21.425 2.737 ;
      RECT 21.285 2.44 21.371 2.73 ;
      RECT 21.236 2.487 21.285 2.723 ;
      RECT 21.15 2.495 21.236 2.716 ;
      RECT 21.135 2.492 21.15 2.711 ;
      RECT 21.121 2.485 21.135 2.71 ;
      RECT 21.035 2.485 21.121 2.705 ;
      RECT 20.94 2.49 20.95 2.69 ;
      RECT 20.53 1.92 20.545 2.32 ;
      RECT 20.725 1.92 20.73 2.18 ;
      RECT 20.47 1.92 20.515 2.18 ;
      RECT 20.925 3.225 20.93 3.43 ;
      RECT 20.92 3.215 20.925 3.435 ;
      RECT 20.915 3.202 20.92 3.44 ;
      RECT 20.91 3.182 20.915 3.44 ;
      RECT 20.885 3.135 20.91 3.44 ;
      RECT 20.85 3.05 20.885 3.44 ;
      RECT 20.845 2.987 20.85 3.44 ;
      RECT 20.84 2.972 20.845 3.44 ;
      RECT 20.825 2.932 20.84 3.44 ;
      RECT 20.82 2.907 20.825 3.44 ;
      RECT 20.81 2.89 20.82 3.44 ;
      RECT 20.775 2.812 20.81 3.44 ;
      RECT 20.77 2.755 20.775 3.44 ;
      RECT 20.765 2.742 20.77 3.44 ;
      RECT 20.755 2.72 20.765 3.44 ;
      RECT 20.745 2.685 20.755 3.44 ;
      RECT 20.735 2.655 20.745 3.44 ;
      RECT 20.725 2.57 20.735 3.083 ;
      RECT 20.732 3.215 20.735 3.44 ;
      RECT 20.73 3.225 20.732 3.44 ;
      RECT 20.72 3.235 20.73 3.435 ;
      RECT 20.715 1.92 20.725 2.315 ;
      RECT 20.72 2.447 20.725 3.058 ;
      RECT 20.715 2.345 20.72 3.041 ;
      RECT 20.705 1.92 20.715 3.017 ;
      RECT 20.7 1.92 20.705 2.988 ;
      RECT 20.695 1.92 20.7 2.978 ;
      RECT 20.675 1.92 20.695 2.94 ;
      RECT 20.67 1.92 20.675 2.898 ;
      RECT 20.665 1.92 20.67 2.878 ;
      RECT 20.635 1.92 20.665 2.828 ;
      RECT 20.625 1.92 20.635 2.775 ;
      RECT 20.62 1.92 20.625 2.748 ;
      RECT 20.615 1.92 20.62 2.733 ;
      RECT 20.605 1.92 20.615 2.71 ;
      RECT 20.595 1.92 20.605 2.685 ;
      RECT 20.59 1.92 20.595 2.625 ;
      RECT 20.58 1.92 20.59 2.563 ;
      RECT 20.575 1.92 20.58 2.483 ;
      RECT 20.57 1.92 20.575 2.448 ;
      RECT 20.565 1.92 20.57 2.423 ;
      RECT 20.56 1.92 20.565 2.408 ;
      RECT 20.555 1.92 20.56 2.378 ;
      RECT 20.55 1.92 20.555 2.355 ;
      RECT 20.545 1.92 20.55 2.328 ;
      RECT 20.515 1.92 20.53 2.315 ;
      RECT 19.67 3.455 19.855 3.665 ;
      RECT 19.66 3.46 19.87 3.658 ;
      RECT 19.66 3.46 19.89 3.63 ;
      RECT 19.66 3.46 19.905 3.609 ;
      RECT 19.66 3.46 19.92 3.607 ;
      RECT 19.66 3.46 19.93 3.606 ;
      RECT 19.66 3.46 19.96 3.603 ;
      RECT 20.31 3.305 20.57 3.565 ;
      RECT 20.27 3.352 20.57 3.548 ;
      RECT 20.261 3.36 20.27 3.551 ;
      RECT 19.855 3.453 20.57 3.548 ;
      RECT 20.175 3.378 20.261 3.558 ;
      RECT 19.87 3.45 20.57 3.548 ;
      RECT 20.116 3.4 20.175 3.57 ;
      RECT 19.89 3.446 20.57 3.548 ;
      RECT 20.03 3.412 20.116 3.581 ;
      RECT 19.905 3.442 20.57 3.548 ;
      RECT 19.975 3.425 20.03 3.593 ;
      RECT 19.92 3.44 20.57 3.548 ;
      RECT 19.96 3.431 19.975 3.599 ;
      RECT 19.93 3.436 20.57 3.548 ;
      RECT 20.075 2.96 20.335 3.22 ;
      RECT 20.075 2.98 20.445 3.19 ;
      RECT 20.075 2.985 20.455 3.185 ;
      RECT 20.266 2.399 20.345 2.63 ;
      RECT 20.18 2.402 20.395 2.625 ;
      RECT 20.175 2.402 20.395 2.62 ;
      RECT 20.175 2.407 20.405 2.618 ;
      RECT 20.15 2.407 20.405 2.615 ;
      RECT 20.15 2.415 20.415 2.613 ;
      RECT 20.03 2.35 20.29 2.61 ;
      RECT 20.03 2.397 20.34 2.61 ;
      RECT 19.285 2.97 19.29 3.23 ;
      RECT 19.115 2.74 19.12 3.23 ;
      RECT 19 2.98 19.005 3.205 ;
      RECT 19.71 2.075 19.715 2.285 ;
      RECT 19.715 2.08 19.73 2.28 ;
      RECT 19.65 2.075 19.71 2.293 ;
      RECT 19.635 2.075 19.65 2.303 ;
      RECT 19.585 2.075 19.635 2.32 ;
      RECT 19.565 2.075 19.585 2.343 ;
      RECT 19.55 2.075 19.565 2.355 ;
      RECT 19.53 2.075 19.55 2.365 ;
      RECT 19.52 2.08 19.53 2.374 ;
      RECT 19.515 2.09 19.52 2.379 ;
      RECT 19.51 2.102 19.515 2.383 ;
      RECT 19.5 2.125 19.51 2.388 ;
      RECT 19.495 2.14 19.5 2.392 ;
      RECT 19.49 2.157 19.495 2.395 ;
      RECT 19.485 2.165 19.49 2.398 ;
      RECT 19.475 2.17 19.485 2.402 ;
      RECT 19.47 2.177 19.475 2.407 ;
      RECT 19.46 2.182 19.47 2.411 ;
      RECT 19.435 2.194 19.46 2.422 ;
      RECT 19.415 2.211 19.435 2.438 ;
      RECT 19.39 2.228 19.415 2.46 ;
      RECT 19.355 2.251 19.39 2.518 ;
      RECT 19.335 2.273 19.355 2.58 ;
      RECT 19.33 2.283 19.335 2.615 ;
      RECT 19.32 2.29 19.33 2.653 ;
      RECT 19.315 2.297 19.32 2.673 ;
      RECT 19.31 2.308 19.315 2.71 ;
      RECT 19.305 2.316 19.31 2.775 ;
      RECT 19.295 2.327 19.305 2.828 ;
      RECT 19.29 2.345 19.295 2.898 ;
      RECT 19.285 2.355 19.29 2.935 ;
      RECT 19.28 2.365 19.285 3.23 ;
      RECT 19.275 2.377 19.28 3.23 ;
      RECT 19.27 2.387 19.275 3.23 ;
      RECT 19.26 2.397 19.27 3.23 ;
      RECT 19.25 2.42 19.26 3.23 ;
      RECT 19.235 2.455 19.25 3.23 ;
      RECT 19.195 2.517 19.235 3.23 ;
      RECT 19.19 2.57 19.195 3.23 ;
      RECT 19.165 2.605 19.19 3.23 ;
      RECT 19.15 2.65 19.165 3.23 ;
      RECT 19.145 2.672 19.15 3.23 ;
      RECT 19.135 2.685 19.145 3.23 ;
      RECT 19.125 2.71 19.135 3.23 ;
      RECT 19.12 2.732 19.125 3.23 ;
      RECT 19.095 2.77 19.115 3.23 ;
      RECT 19.055 2.827 19.095 3.23 ;
      RECT 19.05 2.877 19.055 3.23 ;
      RECT 19.045 2.895 19.05 3.23 ;
      RECT 19.04 2.907 19.045 3.23 ;
      RECT 19.03 2.925 19.04 3.23 ;
      RECT 19.02 2.945 19.03 3.205 ;
      RECT 19.015 2.962 19.02 3.205 ;
      RECT 19.005 2.975 19.015 3.205 ;
      RECT 18.975 2.985 19 3.205 ;
      RECT 18.965 2.992 18.975 3.205 ;
      RECT 18.95 3.002 18.965 3.2 ;
      RECT 18.045 7.77 18.335 8 ;
      RECT 18.105 6.29 18.275 8 ;
      RECT 18.1 6.655 18.45 7.005 ;
      RECT 18.045 6.29 18.335 6.52 ;
      RECT 17.64 2.395 17.745 2.965 ;
      RECT 17.64 2.73 17.965 2.96 ;
      RECT 17.64 2.76 18.135 2.93 ;
      RECT 17.64 2.395 17.83 2.96 ;
      RECT 17.055 2.36 17.345 2.59 ;
      RECT 17.055 2.395 17.83 2.565 ;
      RECT 17.115 0.88 17.285 2.59 ;
      RECT 17.055 0.88 17.345 1.11 ;
      RECT 17.055 7.77 17.345 8 ;
      RECT 17.115 6.29 17.285 8 ;
      RECT 17.055 6.29 17.345 6.52 ;
      RECT 17.055 6.325 17.91 6.485 ;
      RECT 17.74 5.92 17.91 6.485 ;
      RECT 17.055 6.32 17.45 6.485 ;
      RECT 17.675 5.92 17.965 6.15 ;
      RECT 17.675 5.95 18.135 6.12 ;
      RECT 16.685 2.73 16.975 2.96 ;
      RECT 16.685 2.76 17.145 2.93 ;
      RECT 16.75 1.655 16.915 2.96 ;
      RECT 15.265 1.625 15.555 1.855 ;
      RECT 15.265 1.655 16.915 1.825 ;
      RECT 15.325 0.885 15.495 1.855 ;
      RECT 15.265 0.885 15.555 1.115 ;
      RECT 15.265 7.765 15.555 7.995 ;
      RECT 15.325 7.025 15.495 7.995 ;
      RECT 15.325 7.12 16.915 7.29 ;
      RECT 16.745 5.92 16.915 7.29 ;
      RECT 15.265 7.025 15.555 7.255 ;
      RECT 16.685 5.92 16.975 6.15 ;
      RECT 16.685 5.95 17.145 6.12 ;
      RECT 15.695 1.965 16.045 2.315 ;
      RECT 13.36 2.025 16.045 2.195 ;
      RECT 13.36 1.34 13.53 2.195 ;
      RECT 13.26 1.34 13.61 1.69 ;
      RECT 15.72 6.655 16.045 6.98 ;
      RECT 11.115 6.605 11.465 6.955 ;
      RECT 15.695 6.655 16.045 6.885 ;
      RECT 10.915 6.655 11.465 6.885 ;
      RECT 10.745 6.685 16.045 6.855 ;
      RECT 14.92 2.365 15.24 2.685 ;
      RECT 14.89 2.365 15.24 2.595 ;
      RECT 14.72 2.395 15.24 2.565 ;
      RECT 14.92 6.255 15.24 6.545 ;
      RECT 14.89 6.285 15.24 6.515 ;
      RECT 14.72 6.315 15.24 6.485 ;
      RECT 11.555 2.465 11.74 2.675 ;
      RECT 11.545 2.47 11.755 2.668 ;
      RECT 11.545 2.47 11.841 2.645 ;
      RECT 11.545 2.47 11.9 2.62 ;
      RECT 11.545 2.47 11.955 2.6 ;
      RECT 11.545 2.47 11.965 2.588 ;
      RECT 11.545 2.47 12.16 2.527 ;
      RECT 11.545 2.47 12.19 2.51 ;
      RECT 11.545 2.47 12.21 2.5 ;
      RECT 12.09 2.235 12.35 2.495 ;
      RECT 12.075 2.325 12.09 2.542 ;
      RECT 11.61 2.457 12.35 2.495 ;
      RECT 12.061 2.336 12.075 2.548 ;
      RECT 11.65 2.45 12.35 2.495 ;
      RECT 11.975 2.376 12.061 2.567 ;
      RECT 11.9 2.437 12.35 2.495 ;
      RECT 11.97 2.412 11.975 2.584 ;
      RECT 11.955 2.422 12.35 2.495 ;
      RECT 11.965 2.417 11.97 2.586 ;
      RECT 12.26 2.922 12.265 3.014 ;
      RECT 12.255 2.9 12.26 3.031 ;
      RECT 12.25 2.89 12.255 3.043 ;
      RECT 12.24 2.881 12.25 3.053 ;
      RECT 12.235 2.876 12.24 3.061 ;
      RECT 12.23 2.735 12.235 3.064 ;
      RECT 12.196 2.735 12.23 3.075 ;
      RECT 12.11 2.735 12.196 3.11 ;
      RECT 12.03 2.735 12.11 3.158 ;
      RECT 12.001 2.735 12.03 3.182 ;
      RECT 11.915 2.735 12.001 3.188 ;
      RECT 11.91 2.919 11.915 3.193 ;
      RECT 11.875 2.93 11.91 3.196 ;
      RECT 11.85 2.945 11.875 3.2 ;
      RECT 11.836 2.954 11.85 3.202 ;
      RECT 11.75 2.981 11.836 3.208 ;
      RECT 11.685 3.022 11.75 3.217 ;
      RECT 11.67 3.042 11.685 3.222 ;
      RECT 11.64 3.052 11.67 3.225 ;
      RECT 11.635 3.062 11.64 3.228 ;
      RECT 11.605 3.067 11.635 3.23 ;
      RECT 11.585 3.072 11.605 3.234 ;
      RECT 11.5 3.075 11.585 3.241 ;
      RECT 11.485 3.072 11.5 3.247 ;
      RECT 11.475 3.069 11.485 3.249 ;
      RECT 11.455 3.066 11.475 3.251 ;
      RECT 11.435 3.062 11.455 3.252 ;
      RECT 11.42 3.058 11.435 3.254 ;
      RECT 11.41 3.055 11.42 3.255 ;
      RECT 11.37 3.049 11.41 3.253 ;
      RECT 11.36 3.044 11.37 3.251 ;
      RECT 11.345 3.041 11.36 3.247 ;
      RECT 11.32 3.036 11.345 3.24 ;
      RECT 11.27 3.027 11.32 3.228 ;
      RECT 11.2 3.013 11.27 3.21 ;
      RECT 11.142 2.998 11.2 3.192 ;
      RECT 11.056 2.981 11.142 3.172 ;
      RECT 10.97 2.96 11.056 3.147 ;
      RECT 10.92 2.945 10.97 3.128 ;
      RECT 10.916 2.939 10.92 3.12 ;
      RECT 10.83 2.929 10.916 3.107 ;
      RECT 10.795 2.914 10.83 3.09 ;
      RECT 10.78 2.907 10.795 3.083 ;
      RECT 10.72 2.895 10.78 3.071 ;
      RECT 10.7 2.882 10.72 3.059 ;
      RECT 10.66 2.873 10.7 3.051 ;
      RECT 10.655 2.865 10.66 3.044 ;
      RECT 10.575 2.855 10.655 3.03 ;
      RECT 10.56 2.842 10.575 3.015 ;
      RECT 10.555 2.84 10.56 3.013 ;
      RECT 10.476 2.828 10.555 3 ;
      RECT 10.39 2.803 10.476 2.975 ;
      RECT 10.375 2.772 10.39 2.96 ;
      RECT 10.36 2.747 10.375 2.956 ;
      RECT 10.345 2.74 10.36 2.952 ;
      RECT 10.17 2.745 10.175 2.948 ;
      RECT 10.165 2.75 10.17 2.943 ;
      RECT 10.175 2.74 10.345 2.95 ;
      RECT 10.89 2.5 10.995 2.76 ;
      RECT 11.705 2.025 11.71 2.25 ;
      RECT 11.835 2.025 11.89 2.235 ;
      RECT 11.89 2.03 11.9 2.228 ;
      RECT 11.796 2.025 11.835 2.238 ;
      RECT 11.71 2.025 11.796 2.245 ;
      RECT 11.69 2.03 11.705 2.251 ;
      RECT 11.68 2.07 11.69 2.253 ;
      RECT 11.65 2.08 11.68 2.255 ;
      RECT 11.645 2.085 11.65 2.257 ;
      RECT 11.62 2.09 11.645 2.259 ;
      RECT 11.605 2.095 11.62 2.261 ;
      RECT 11.59 2.097 11.605 2.263 ;
      RECT 11.585 2.102 11.59 2.265 ;
      RECT 11.535 2.11 11.585 2.268 ;
      RECT 11.51 2.119 11.535 2.273 ;
      RECT 11.5 2.126 11.51 2.278 ;
      RECT 11.495 2.129 11.5 2.282 ;
      RECT 11.475 2.132 11.495 2.291 ;
      RECT 11.445 2.14 11.475 2.311 ;
      RECT 11.416 2.153 11.445 2.333 ;
      RECT 11.33 2.187 11.416 2.377 ;
      RECT 11.325 2.213 11.33 2.415 ;
      RECT 11.32 2.217 11.325 2.424 ;
      RECT 11.285 2.23 11.32 2.457 ;
      RECT 11.275 2.244 11.285 2.495 ;
      RECT 11.27 2.248 11.275 2.508 ;
      RECT 11.265 2.252 11.27 2.513 ;
      RECT 11.255 2.26 11.265 2.525 ;
      RECT 11.25 2.267 11.255 2.54 ;
      RECT 11.225 2.28 11.25 2.565 ;
      RECT 11.185 2.309 11.225 2.62 ;
      RECT 11.17 2.334 11.185 2.675 ;
      RECT 11.16 2.345 11.17 2.698 ;
      RECT 11.155 2.352 11.16 2.71 ;
      RECT 11.15 2.356 11.155 2.718 ;
      RECT 11.095 2.384 11.15 2.76 ;
      RECT 11.075 2.42 11.095 2.76 ;
      RECT 11.06 2.435 11.075 2.76 ;
      RECT 11.005 2.467 11.06 2.76 ;
      RECT 10.995 2.497 11.005 2.76 ;
      RECT 10.605 2.112 10.79 2.35 ;
      RECT 10.59 2.114 10.8 2.345 ;
      RECT 10.475 2.06 10.735 2.32 ;
      RECT 10.47 2.097 10.735 2.274 ;
      RECT 10.465 2.107 10.735 2.271 ;
      RECT 10.46 2.147 10.8 2.265 ;
      RECT 10.455 2.18 10.8 2.255 ;
      RECT 10.465 2.122 10.815 2.193 ;
      RECT 10.762 3.22 10.775 3.75 ;
      RECT 10.676 3.22 10.775 3.749 ;
      RECT 10.676 3.22 10.78 3.748 ;
      RECT 10.59 3.22 10.78 3.746 ;
      RECT 10.585 3.22 10.78 3.743 ;
      RECT 10.585 3.22 10.79 3.741 ;
      RECT 10.58 3.512 10.79 3.738 ;
      RECT 10.58 3.522 10.795 3.735 ;
      RECT 10.58 3.59 10.8 3.731 ;
      RECT 10.57 3.595 10.8 3.73 ;
      RECT 10.57 3.687 10.805 3.727 ;
      RECT 10.555 3.22 10.815 3.48 ;
      RECT 10.485 7.765 10.775 7.995 ;
      RECT 10.545 7.025 10.715 7.995 ;
      RECT 10.46 7.055 10.8 7.4 ;
      RECT 10.485 7.025 10.775 7.4 ;
      RECT 9.785 2.21 9.83 3.745 ;
      RECT 9.985 2.21 10.015 2.425 ;
      RECT 8.36 1.95 8.48 2.16 ;
      RECT 8.02 1.9 8.28 2.16 ;
      RECT 8.02 1.945 8.315 2.15 ;
      RECT 10.025 2.226 10.03 2.28 ;
      RECT 10.02 2.219 10.025 2.413 ;
      RECT 10.015 2.213 10.02 2.42 ;
      RECT 9.97 2.21 9.985 2.433 ;
      RECT 9.965 2.21 9.97 2.455 ;
      RECT 9.96 2.21 9.965 2.503 ;
      RECT 9.955 2.21 9.96 2.523 ;
      RECT 9.945 2.21 9.955 2.63 ;
      RECT 9.94 2.21 9.945 2.693 ;
      RECT 9.935 2.21 9.94 2.75 ;
      RECT 9.93 2.21 9.935 2.758 ;
      RECT 9.915 2.21 9.93 2.865 ;
      RECT 9.905 2.21 9.915 3 ;
      RECT 9.895 2.21 9.905 3.11 ;
      RECT 9.885 2.21 9.895 3.167 ;
      RECT 9.88 2.21 9.885 3.207 ;
      RECT 9.875 2.21 9.88 3.243 ;
      RECT 9.865 2.21 9.875 3.283 ;
      RECT 9.86 2.21 9.865 3.325 ;
      RECT 9.84 2.21 9.86 3.39 ;
      RECT 9.845 3.535 9.85 3.715 ;
      RECT 9.84 3.517 9.845 3.723 ;
      RECT 9.835 2.21 9.84 3.453 ;
      RECT 9.835 3.497 9.84 3.73 ;
      RECT 9.83 2.21 9.835 3.74 ;
      RECT 9.775 2.21 9.785 2.51 ;
      RECT 9.78 2.757 9.785 3.745 ;
      RECT 9.775 2.822 9.78 3.745 ;
      RECT 9.77 2.211 9.775 2.5 ;
      RECT 9.765 2.887 9.775 3.745 ;
      RECT 9.76 2.212 9.77 2.49 ;
      RECT 9.75 3 9.765 3.745 ;
      RECT 9.755 2.213 9.76 2.48 ;
      RECT 9.735 2.214 9.755 2.458 ;
      RECT 9.74 3.097 9.75 3.745 ;
      RECT 9.735 3.172 9.74 3.745 ;
      RECT 9.725 2.213 9.735 2.435 ;
      RECT 9.73 3.215 9.735 3.745 ;
      RECT 9.725 3.242 9.73 3.745 ;
      RECT 9.715 2.211 9.725 2.423 ;
      RECT 9.72 3.285 9.725 3.745 ;
      RECT 9.715 3.312 9.72 3.745 ;
      RECT 9.705 2.21 9.715 2.41 ;
      RECT 9.71 3.327 9.715 3.745 ;
      RECT 9.67 3.385 9.71 3.745 ;
      RECT 9.7 2.209 9.705 2.395 ;
      RECT 9.695 2.207 9.7 2.388 ;
      RECT 9.685 2.204 9.695 2.378 ;
      RECT 9.68 2.201 9.685 2.363 ;
      RECT 9.665 2.197 9.68 2.356 ;
      RECT 9.66 3.44 9.67 3.745 ;
      RECT 9.66 2.194 9.665 2.351 ;
      RECT 9.645 2.19 9.66 2.345 ;
      RECT 9.655 3.457 9.66 3.745 ;
      RECT 9.645 3.52 9.655 3.745 ;
      RECT 9.565 2.175 9.645 2.325 ;
      RECT 9.64 3.527 9.645 3.74 ;
      RECT 9.635 3.535 9.64 3.73 ;
      RECT 9.555 2.161 9.565 2.309 ;
      RECT 9.54 2.157 9.555 2.307 ;
      RECT 9.53 2.152 9.54 2.303 ;
      RECT 9.505 2.145 9.53 2.295 ;
      RECT 9.5 2.14 9.505 2.29 ;
      RECT 9.49 2.14 9.5 2.288 ;
      RECT 9.48 2.138 9.49 2.286 ;
      RECT 9.45 2.13 9.48 2.28 ;
      RECT 9.435 2.122 9.45 2.273 ;
      RECT 9.415 2.117 9.435 2.266 ;
      RECT 9.41 2.113 9.415 2.261 ;
      RECT 9.38 2.106 9.41 2.255 ;
      RECT 9.355 2.097 9.38 2.245 ;
      RECT 9.325 2.09 9.355 2.237 ;
      RECT 9.3 2.08 9.325 2.228 ;
      RECT 9.285 2.072 9.3 2.222 ;
      RECT 9.26 2.067 9.285 2.217 ;
      RECT 9.25 2.063 9.26 2.212 ;
      RECT 9.23 2.058 9.25 2.207 ;
      RECT 9.195 2.053 9.23 2.2 ;
      RECT 9.135 2.048 9.195 2.193 ;
      RECT 9.122 2.044 9.135 2.191 ;
      RECT 9.036 2.039 9.122 2.188 ;
      RECT 8.95 2.029 9.036 2.184 ;
      RECT 8.909 2.022 8.95 2.181 ;
      RECT 8.823 2.015 8.909 2.178 ;
      RECT 8.737 2.005 8.823 2.174 ;
      RECT 8.651 1.995 8.737 2.169 ;
      RECT 8.565 1.985 8.651 2.165 ;
      RECT 8.555 1.97 8.565 2.163 ;
      RECT 8.545 1.955 8.555 2.163 ;
      RECT 8.48 1.95 8.545 2.162 ;
      RECT 8.315 1.947 8.36 2.155 ;
      RECT 9.56 2.852 9.565 3.043 ;
      RECT 9.555 2.847 9.56 3.05 ;
      RECT 9.541 2.845 9.555 3.056 ;
      RECT 9.455 2.845 9.541 3.058 ;
      RECT 9.451 2.845 9.455 3.061 ;
      RECT 9.365 2.845 9.451 3.079 ;
      RECT 9.355 2.85 9.365 3.098 ;
      RECT 9.345 2.905 9.355 3.102 ;
      RECT 9.32 2.92 9.345 3.109 ;
      RECT 9.28 2.94 9.32 3.122 ;
      RECT 9.275 2.952 9.28 3.132 ;
      RECT 9.26 2.958 9.275 3.137 ;
      RECT 9.255 2.963 9.26 3.141 ;
      RECT 9.235 2.97 9.255 3.146 ;
      RECT 9.165 2.995 9.235 3.163 ;
      RECT 9.125 3.023 9.165 3.183 ;
      RECT 9.12 3.033 9.125 3.191 ;
      RECT 9.1 3.04 9.12 3.193 ;
      RECT 9.095 3.047 9.1 3.196 ;
      RECT 9.065 3.055 9.095 3.199 ;
      RECT 9.06 3.06 9.065 3.203 ;
      RECT 8.986 3.064 9.06 3.211 ;
      RECT 8.9 3.073 8.986 3.227 ;
      RECT 8.896 3.078 8.9 3.236 ;
      RECT 8.81 3.083 8.896 3.246 ;
      RECT 8.77 3.091 8.81 3.258 ;
      RECT 8.72 3.097 8.77 3.265 ;
      RECT 8.635 3.106 8.72 3.28 ;
      RECT 8.56 3.117 8.635 3.298 ;
      RECT 8.525 3.124 8.56 3.308 ;
      RECT 8.45 3.132 8.525 3.313 ;
      RECT 8.395 3.141 8.45 3.313 ;
      RECT 8.37 3.146 8.395 3.311 ;
      RECT 8.36 3.149 8.37 3.309 ;
      RECT 8.325 3.151 8.36 3.307 ;
      RECT 8.295 3.153 8.325 3.303 ;
      RECT 8.25 3.152 8.295 3.299 ;
      RECT 8.23 3.147 8.25 3.296 ;
      RECT 8.18 3.132 8.23 3.293 ;
      RECT 8.17 3.117 8.18 3.288 ;
      RECT 8.12 3.102 8.17 3.278 ;
      RECT 8.07 3.077 8.12 3.258 ;
      RECT 8.06 3.062 8.07 3.24 ;
      RECT 8.055 3.06 8.06 3.234 ;
      RECT 8.035 3.055 8.055 3.229 ;
      RECT 8.03 3.047 8.035 3.223 ;
      RECT 8.015 3.041 8.03 3.216 ;
      RECT 8.01 3.036 8.015 3.208 ;
      RECT 7.99 3.031 8.01 3.2 ;
      RECT 7.975 3.024 7.99 3.193 ;
      RECT 7.96 3.018 7.975 3.184 ;
      RECT 7.955 3.012 7.96 3.177 ;
      RECT 7.91 2.987 7.955 3.163 ;
      RECT 7.895 2.957 7.91 3.145 ;
      RECT 7.88 2.94 7.895 3.136 ;
      RECT 7.855 2.92 7.88 3.124 ;
      RECT 7.815 2.89 7.855 3.104 ;
      RECT 7.805 2.86 7.815 3.089 ;
      RECT 7.79 2.85 7.805 3.082 ;
      RECT 7.735 2.815 7.79 3.061 ;
      RECT 7.72 2.778 7.735 3.04 ;
      RECT 7.71 2.765 7.72 3.032 ;
      RECT 7.66 2.735 7.71 3.014 ;
      RECT 7.645 2.665 7.66 2.995 ;
      RECT 7.6 2.665 7.645 2.978 ;
      RECT 7.575 2.665 7.6 2.96 ;
      RECT 7.565 2.665 7.575 2.953 ;
      RECT 7.486 2.665 7.565 2.946 ;
      RECT 7.4 2.665 7.486 2.938 ;
      RECT 7.385 2.697 7.4 2.933 ;
      RECT 7.31 2.707 7.385 2.929 ;
      RECT 7.29 2.717 7.31 2.924 ;
      RECT 7.265 2.717 7.29 2.921 ;
      RECT 7.255 2.707 7.265 2.92 ;
      RECT 7.245 2.68 7.255 2.919 ;
      RECT 7.205 2.675 7.245 2.917 ;
      RECT 7.16 2.675 7.205 2.913 ;
      RECT 7.135 2.675 7.16 2.908 ;
      RECT 7.085 2.675 7.135 2.895 ;
      RECT 7.045 2.68 7.055 2.88 ;
      RECT 7.055 2.675 7.085 2.885 ;
      RECT 9.04 2.455 9.3 2.715 ;
      RECT 9.035 2.477 9.3 2.673 ;
      RECT 8.275 2.305 8.495 2.67 ;
      RECT 8.257 2.392 8.495 2.669 ;
      RECT 8.24 2.397 8.495 2.666 ;
      RECT 8.24 2.397 8.515 2.665 ;
      RECT 8.21 2.407 8.515 2.663 ;
      RECT 8.205 2.422 8.515 2.659 ;
      RECT 8.205 2.422 8.52 2.658 ;
      RECT 8.2 2.48 8.52 2.656 ;
      RECT 8.2 2.48 8.53 2.653 ;
      RECT 8.195 2.545 8.53 2.648 ;
      RECT 8.275 2.305 8.535 2.565 ;
      RECT 7.02 2.135 7.28 2.395 ;
      RECT 7.02 2.178 7.366 2.369 ;
      RECT 7.02 2.178 7.41 2.368 ;
      RECT 7.02 2.178 7.43 2.366 ;
      RECT 7.02 2.178 7.53 2.365 ;
      RECT 7.02 2.178 7.55 2.363 ;
      RECT 7.02 2.178 7.56 2.358 ;
      RECT 7.43 2.145 7.62 2.355 ;
      RECT 7.43 2.147 7.625 2.353 ;
      RECT 7.42 2.152 7.63 2.345 ;
      RECT 7.366 2.176 7.63 2.345 ;
      RECT 7.41 2.17 7.42 2.367 ;
      RECT 7.42 2.15 7.625 2.353 ;
      RECT 6.375 3.21 6.58 3.44 ;
      RECT 6.315 3.16 6.37 3.42 ;
      RECT 6.375 3.16 6.575 3.44 ;
      RECT 7.345 3.475 7.35 3.502 ;
      RECT 7.335 3.385 7.345 3.507 ;
      RECT 7.33 3.307 7.335 3.513 ;
      RECT 7.32 3.297 7.33 3.52 ;
      RECT 7.315 3.287 7.32 3.526 ;
      RECT 7.305 3.282 7.315 3.528 ;
      RECT 7.29 3.274 7.305 3.536 ;
      RECT 7.275 3.265 7.29 3.548 ;
      RECT 7.265 3.257 7.275 3.558 ;
      RECT 7.23 3.175 7.265 3.576 ;
      RECT 7.195 3.175 7.23 3.595 ;
      RECT 7.18 3.175 7.195 3.603 ;
      RECT 7.125 3.175 7.18 3.603 ;
      RECT 7.091 3.175 7.125 3.594 ;
      RECT 7.005 3.175 7.091 3.57 ;
      RECT 6.995 3.235 7.005 3.552 ;
      RECT 6.955 3.237 6.995 3.543 ;
      RECT 6.95 3.239 6.955 3.533 ;
      RECT 6.93 3.241 6.95 3.528 ;
      RECT 6.92 3.244 6.93 3.523 ;
      RECT 6.91 3.245 6.92 3.518 ;
      RECT 6.886 3.246 6.91 3.51 ;
      RECT 6.8 3.251 6.886 3.488 ;
      RECT 6.745 3.25 6.8 3.461 ;
      RECT 6.73 3.243 6.745 3.448 ;
      RECT 6.695 3.238 6.73 3.444 ;
      RECT 6.64 3.23 6.695 3.443 ;
      RECT 6.58 3.217 6.64 3.441 ;
      RECT 6.37 3.16 6.375 3.428 ;
      RECT 6.445 2.53 6.63 2.74 ;
      RECT 6.435 2.535 6.645 2.733 ;
      RECT 6.475 2.44 6.735 2.7 ;
      RECT 6.43 2.597 6.735 2.623 ;
      RECT 5.775 2.39 5.78 3.19 ;
      RECT 5.72 2.44 5.75 3.19 ;
      RECT 5.71 2.44 5.715 2.75 ;
      RECT 5.695 2.44 5.7 2.745 ;
      RECT 5.24 2.485 5.255 2.7 ;
      RECT 5.17 2.485 5.255 2.695 ;
      RECT 6.435 2.065 6.505 2.275 ;
      RECT 6.505 2.072 6.515 2.27 ;
      RECT 6.401 2.065 6.435 2.282 ;
      RECT 6.315 2.065 6.401 2.306 ;
      RECT 6.305 2.07 6.315 2.325 ;
      RECT 6.3 2.082 6.305 2.328 ;
      RECT 6.285 2.097 6.3 2.332 ;
      RECT 6.28 2.115 6.285 2.336 ;
      RECT 6.24 2.125 6.28 2.345 ;
      RECT 6.225 2.132 6.24 2.357 ;
      RECT 6.21 2.137 6.225 2.362 ;
      RECT 6.195 2.14 6.21 2.367 ;
      RECT 6.185 2.142 6.195 2.371 ;
      RECT 6.15 2.149 6.185 2.379 ;
      RECT 6.115 2.157 6.15 2.393 ;
      RECT 6.105 2.163 6.115 2.402 ;
      RECT 6.1 2.165 6.105 2.404 ;
      RECT 6.08 2.168 6.1 2.41 ;
      RECT 6.05 2.175 6.08 2.421 ;
      RECT 6.04 2.181 6.05 2.428 ;
      RECT 6.015 2.184 6.04 2.435 ;
      RECT 6.005 2.188 6.015 2.443 ;
      RECT 6 2.189 6.005 2.465 ;
      RECT 5.995 2.19 6 2.48 ;
      RECT 5.99 2.191 5.995 2.495 ;
      RECT 5.985 2.192 5.99 2.51 ;
      RECT 5.98 2.193 5.985 2.54 ;
      RECT 5.97 2.195 5.98 2.573 ;
      RECT 5.955 2.199 5.97 2.62 ;
      RECT 5.945 2.202 5.955 2.665 ;
      RECT 5.94 2.205 5.945 2.693 ;
      RECT 5.93 2.207 5.94 2.72 ;
      RECT 5.925 2.21 5.93 2.755 ;
      RECT 5.895 2.215 5.925 2.813 ;
      RECT 5.89 2.22 5.895 2.898 ;
      RECT 5.885 2.222 5.89 2.933 ;
      RECT 5.88 2.224 5.885 3.015 ;
      RECT 5.875 2.226 5.88 3.103 ;
      RECT 5.865 2.228 5.875 3.185 ;
      RECT 5.85 2.242 5.865 3.19 ;
      RECT 5.815 2.287 5.85 3.19 ;
      RECT 5.805 2.327 5.815 3.19 ;
      RECT 5.79 2.355 5.805 3.19 ;
      RECT 5.785 2.372 5.79 3.19 ;
      RECT 5.78 2.38 5.785 3.19 ;
      RECT 5.77 2.395 5.775 3.19 ;
      RECT 5.765 2.402 5.77 3.19 ;
      RECT 5.755 2.422 5.765 3.19 ;
      RECT 5.75 2.435 5.755 3.19 ;
      RECT 5.715 2.44 5.72 2.775 ;
      RECT 5.7 2.83 5.72 3.19 ;
      RECT 5.7 2.44 5.71 2.748 ;
      RECT 5.695 2.87 5.7 3.19 ;
      RECT 5.645 2.44 5.695 2.743 ;
      RECT 5.69 2.907 5.695 3.19 ;
      RECT 5.68 2.93 5.69 3.19 ;
      RECT 5.675 2.975 5.68 3.19 ;
      RECT 5.665 2.985 5.675 3.183 ;
      RECT 5.591 2.44 5.645 2.737 ;
      RECT 5.505 2.44 5.591 2.73 ;
      RECT 5.456 2.487 5.505 2.723 ;
      RECT 5.37 2.495 5.456 2.716 ;
      RECT 5.355 2.492 5.37 2.711 ;
      RECT 5.341 2.485 5.355 2.71 ;
      RECT 5.255 2.485 5.341 2.705 ;
      RECT 5.16 2.49 5.17 2.69 ;
      RECT 4.75 1.92 4.765 2.32 ;
      RECT 4.945 1.92 4.95 2.18 ;
      RECT 4.69 1.92 4.735 2.18 ;
      RECT 5.145 3.225 5.15 3.43 ;
      RECT 5.14 3.215 5.145 3.435 ;
      RECT 5.135 3.202 5.14 3.44 ;
      RECT 5.13 3.182 5.135 3.44 ;
      RECT 5.105 3.135 5.13 3.44 ;
      RECT 5.07 3.05 5.105 3.44 ;
      RECT 5.065 2.987 5.07 3.44 ;
      RECT 5.06 2.972 5.065 3.44 ;
      RECT 5.045 2.932 5.06 3.44 ;
      RECT 5.04 2.907 5.045 3.44 ;
      RECT 5.03 2.89 5.04 3.44 ;
      RECT 4.995 2.812 5.03 3.44 ;
      RECT 4.99 2.755 4.995 3.44 ;
      RECT 4.985 2.742 4.99 3.44 ;
      RECT 4.975 2.72 4.985 3.44 ;
      RECT 4.965 2.685 4.975 3.44 ;
      RECT 4.955 2.655 4.965 3.44 ;
      RECT 4.945 2.57 4.955 3.083 ;
      RECT 4.952 3.215 4.955 3.44 ;
      RECT 4.95 3.225 4.952 3.44 ;
      RECT 4.94 3.235 4.95 3.435 ;
      RECT 4.935 1.92 4.945 2.315 ;
      RECT 4.94 2.447 4.945 3.058 ;
      RECT 4.935 2.345 4.94 3.041 ;
      RECT 4.925 1.92 4.935 3.017 ;
      RECT 4.92 1.92 4.925 2.988 ;
      RECT 4.915 1.92 4.92 2.978 ;
      RECT 4.895 1.92 4.915 2.94 ;
      RECT 4.89 1.92 4.895 2.898 ;
      RECT 4.885 1.92 4.89 2.878 ;
      RECT 4.855 1.92 4.885 2.828 ;
      RECT 4.845 1.92 4.855 2.775 ;
      RECT 4.84 1.92 4.845 2.748 ;
      RECT 4.835 1.92 4.84 2.733 ;
      RECT 4.825 1.92 4.835 2.71 ;
      RECT 4.815 1.92 4.825 2.685 ;
      RECT 4.81 1.92 4.815 2.625 ;
      RECT 4.8 1.92 4.81 2.563 ;
      RECT 4.795 1.92 4.8 2.483 ;
      RECT 4.79 1.92 4.795 2.448 ;
      RECT 4.785 1.92 4.79 2.423 ;
      RECT 4.78 1.92 4.785 2.408 ;
      RECT 4.775 1.92 4.78 2.378 ;
      RECT 4.77 1.92 4.775 2.355 ;
      RECT 4.765 1.92 4.77 2.328 ;
      RECT 4.735 1.92 4.75 2.315 ;
      RECT 3.89 3.455 4.075 3.665 ;
      RECT 3.88 3.46 4.09 3.658 ;
      RECT 3.88 3.46 4.11 3.63 ;
      RECT 3.88 3.46 4.125 3.609 ;
      RECT 3.88 3.46 4.14 3.607 ;
      RECT 3.88 3.46 4.15 3.606 ;
      RECT 3.88 3.46 4.18 3.603 ;
      RECT 4.53 3.305 4.79 3.565 ;
      RECT 4.49 3.352 4.79 3.548 ;
      RECT 4.481 3.36 4.49 3.551 ;
      RECT 4.075 3.453 4.79 3.548 ;
      RECT 4.395 3.378 4.481 3.558 ;
      RECT 4.09 3.45 4.79 3.548 ;
      RECT 4.336 3.4 4.395 3.57 ;
      RECT 4.11 3.446 4.79 3.548 ;
      RECT 4.25 3.412 4.336 3.581 ;
      RECT 4.125 3.442 4.79 3.548 ;
      RECT 4.195 3.425 4.25 3.593 ;
      RECT 4.14 3.44 4.79 3.548 ;
      RECT 4.18 3.431 4.195 3.599 ;
      RECT 4.15 3.436 4.79 3.548 ;
      RECT 4.295 2.96 4.555 3.22 ;
      RECT 4.295 2.98 4.665 3.19 ;
      RECT 4.295 2.985 4.675 3.185 ;
      RECT 4.486 2.399 4.565 2.63 ;
      RECT 4.4 2.402 4.615 2.625 ;
      RECT 4.395 2.402 4.615 2.62 ;
      RECT 4.395 2.407 4.625 2.618 ;
      RECT 4.37 2.407 4.625 2.615 ;
      RECT 4.37 2.415 4.635 2.613 ;
      RECT 4.25 2.35 4.51 2.61 ;
      RECT 4.25 2.397 4.56 2.61 ;
      RECT 3.505 2.97 3.51 3.23 ;
      RECT 3.335 2.74 3.34 3.23 ;
      RECT 3.22 2.98 3.225 3.205 ;
      RECT 3.93 2.075 3.935 2.285 ;
      RECT 3.935 2.08 3.95 2.28 ;
      RECT 3.87 2.075 3.93 2.293 ;
      RECT 3.855 2.075 3.87 2.303 ;
      RECT 3.805 2.075 3.855 2.32 ;
      RECT 3.785 2.075 3.805 2.343 ;
      RECT 3.77 2.075 3.785 2.355 ;
      RECT 3.75 2.075 3.77 2.365 ;
      RECT 3.74 2.08 3.75 2.374 ;
      RECT 3.735 2.09 3.74 2.379 ;
      RECT 3.73 2.102 3.735 2.383 ;
      RECT 3.72 2.125 3.73 2.388 ;
      RECT 3.715 2.14 3.72 2.392 ;
      RECT 3.71 2.157 3.715 2.395 ;
      RECT 3.705 2.165 3.71 2.398 ;
      RECT 3.695 2.17 3.705 2.402 ;
      RECT 3.69 2.177 3.695 2.407 ;
      RECT 3.68 2.182 3.69 2.411 ;
      RECT 3.655 2.194 3.68 2.422 ;
      RECT 3.635 2.211 3.655 2.438 ;
      RECT 3.61 2.228 3.635 2.46 ;
      RECT 3.575 2.251 3.61 2.518 ;
      RECT 3.555 2.273 3.575 2.58 ;
      RECT 3.55 2.283 3.555 2.615 ;
      RECT 3.54 2.29 3.55 2.653 ;
      RECT 3.535 2.297 3.54 2.673 ;
      RECT 3.53 2.308 3.535 2.71 ;
      RECT 3.525 2.316 3.53 2.775 ;
      RECT 3.515 2.327 3.525 2.828 ;
      RECT 3.51 2.345 3.515 2.898 ;
      RECT 3.505 2.355 3.51 2.935 ;
      RECT 3.5 2.365 3.505 3.23 ;
      RECT 3.495 2.377 3.5 3.23 ;
      RECT 3.49 2.387 3.495 3.23 ;
      RECT 3.48 2.397 3.49 3.23 ;
      RECT 3.47 2.42 3.48 3.23 ;
      RECT 3.455 2.455 3.47 3.23 ;
      RECT 3.415 2.517 3.455 3.23 ;
      RECT 3.41 2.57 3.415 3.23 ;
      RECT 3.385 2.605 3.41 3.23 ;
      RECT 3.37 2.65 3.385 3.23 ;
      RECT 3.365 2.672 3.37 3.23 ;
      RECT 3.355 2.685 3.365 3.23 ;
      RECT 3.345 2.71 3.355 3.23 ;
      RECT 3.34 2.732 3.345 3.23 ;
      RECT 3.315 2.77 3.335 3.23 ;
      RECT 3.275 2.827 3.315 3.23 ;
      RECT 3.27 2.877 3.275 3.23 ;
      RECT 3.265 2.895 3.27 3.23 ;
      RECT 3.26 2.907 3.265 3.23 ;
      RECT 3.25 2.925 3.26 3.23 ;
      RECT 3.24 2.945 3.25 3.205 ;
      RECT 3.235 2.962 3.24 3.205 ;
      RECT 3.225 2.975 3.235 3.205 ;
      RECT 3.195 2.985 3.22 3.205 ;
      RECT 3.185 2.992 3.195 3.205 ;
      RECT 3.17 3.002 3.185 3.2 ;
      RECT 1.55 7.765 1.84 7.995 ;
      RECT 1.61 7.025 1.78 7.995 ;
      RECT 1.52 7.025 1.87 7.315 ;
      RECT 1.145 6.285 1.495 6.575 ;
      RECT 1.005 6.315 1.495 6.485 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 12.935 2.85 13.305 3.22 ;
    LAYER mcon ;
      RECT 81.23 6.32 81.4 6.49 ;
      RECT 81.235 6.315 81.405 6.485 ;
      RECT 65.445 6.32 65.615 6.49 ;
      RECT 65.45 6.315 65.62 6.485 ;
      RECT 49.66 6.32 49.83 6.49 ;
      RECT 49.665 6.315 49.835 6.485 ;
      RECT 33.885 6.32 34.055 6.49 ;
      RECT 33.89 6.315 34.06 6.485 ;
      RECT 18.105 6.32 18.275 6.49 ;
      RECT 18.11 6.315 18.28 6.485 ;
      RECT 81.23 7.8 81.4 7.97 ;
      RECT 80.88 0.1 81.05 0.27 ;
      RECT 80.86 2.76 81.03 2.93 ;
      RECT 80.86 5.95 81.03 6.12 ;
      RECT 80.24 0.91 80.41 1.08 ;
      RECT 80.24 2.39 80.41 2.56 ;
      RECT 80.24 6.32 80.41 6.49 ;
      RECT 80.24 7.8 80.41 7.97 ;
      RECT 79.89 0.1 80.06 0.27 ;
      RECT 79.87 2.76 80.04 2.93 ;
      RECT 79.87 5.95 80.04 6.12 ;
      RECT 79.19 0.105 79.36 0.275 ;
      RECT 78.88 2.025 79.05 2.195 ;
      RECT 78.88 6.685 79.05 6.855 ;
      RECT 78.51 0.105 78.68 0.275 ;
      RECT 78.45 0.915 78.62 1.085 ;
      RECT 78.45 1.655 78.62 1.825 ;
      RECT 78.45 7.055 78.62 7.225 ;
      RECT 78.45 7.795 78.62 7.965 ;
      RECT 78.075 2.395 78.245 2.565 ;
      RECT 78.075 6.315 78.245 6.485 ;
      RECT 77.83 0.105 78 0.275 ;
      RECT 77.15 0.105 77.32 0.275 ;
      RECT 75.525 1.415 75.695 1.585 ;
      RECT 75.155 2.875 75.325 3.045 ;
      RECT 75.065 1.415 75.235 1.585 ;
      RECT 74.835 2.045 75.005 2.215 ;
      RECT 74.69 2.485 74.86 2.655 ;
      RECT 74.605 1.415 74.775 1.585 ;
      RECT 74.145 1.415 74.315 1.585 ;
      RECT 74.1 6.685 74.27 6.855 ;
      RECT 74.08 2.525 74.25 2.695 ;
      RECT 73.735 2.16 73.905 2.33 ;
      RECT 73.725 3.52 73.895 3.69 ;
      RECT 73.685 1.415 73.855 1.585 ;
      RECT 73.67 7.055 73.84 7.225 ;
      RECT 73.67 7.795 73.84 7.965 ;
      RECT 73.31 2.76 73.48 2.93 ;
      RECT 73.225 1.415 73.395 1.585 ;
      RECT 72.96 2.235 73.13 2.405 ;
      RECT 72.78 3.55 72.95 3.72 ;
      RECT 72.765 1.415 72.935 1.585 ;
      RECT 72.5 2.865 72.67 3.035 ;
      RECT 72.305 1.415 72.475 1.585 ;
      RECT 72.18 2.49 72.35 2.66 ;
      RECT 71.845 1.415 72.015 1.585 ;
      RECT 71.49 1.97 71.66 2.14 ;
      RECT 71.415 2.44 71.585 2.61 ;
      RECT 71.385 1.415 71.555 1.585 ;
      RECT 70.925 1.415 71.095 1.585 ;
      RECT 70.565 2.165 70.735 2.335 ;
      RECT 70.465 1.415 70.635 1.585 ;
      RECT 70.225 3.36 70.395 3.53 ;
      RECT 70.19 2.695 70.36 2.865 ;
      RECT 70.005 1.415 70.175 1.585 ;
      RECT 69.58 2.55 69.75 2.72 ;
      RECT 69.545 1.415 69.715 1.585 ;
      RECT 69.51 3.25 69.68 3.42 ;
      RECT 69.45 2.085 69.62 2.255 ;
      RECT 69.085 1.415 69.255 1.585 ;
      RECT 68.81 3 68.98 3.17 ;
      RECT 68.625 1.415 68.795 1.585 ;
      RECT 68.305 2.505 68.475 2.675 ;
      RECT 68.165 1.415 68.335 1.585 ;
      RECT 68.085 3.25 68.255 3.42 ;
      RECT 67.88 2.13 68.05 2.3 ;
      RECT 67.705 1.415 67.875 1.585 ;
      RECT 67.61 3 67.78 3.17 ;
      RECT 67.57 2.43 67.74 2.6 ;
      RECT 67.245 1.415 67.415 1.585 ;
      RECT 67.025 3.475 67.195 3.645 ;
      RECT 66.885 2.095 67.055 2.265 ;
      RECT 66.785 1.415 66.955 1.585 ;
      RECT 66.325 1.415 66.495 1.585 ;
      RECT 66.315 3.015 66.485 3.185 ;
      RECT 65.445 7.8 65.615 7.97 ;
      RECT 65.095 0.1 65.265 0.27 ;
      RECT 65.075 2.76 65.245 2.93 ;
      RECT 65.075 5.95 65.245 6.12 ;
      RECT 64.455 0.91 64.625 1.08 ;
      RECT 64.455 2.39 64.625 2.56 ;
      RECT 64.455 6.32 64.625 6.49 ;
      RECT 64.455 7.8 64.625 7.97 ;
      RECT 64.105 0.1 64.275 0.27 ;
      RECT 64.085 2.76 64.255 2.93 ;
      RECT 64.085 5.95 64.255 6.12 ;
      RECT 63.405 0.105 63.575 0.275 ;
      RECT 63.095 2.025 63.265 2.195 ;
      RECT 63.095 6.685 63.265 6.855 ;
      RECT 62.725 0.105 62.895 0.275 ;
      RECT 62.665 0.915 62.835 1.085 ;
      RECT 62.665 1.655 62.835 1.825 ;
      RECT 62.665 7.055 62.835 7.225 ;
      RECT 62.665 7.795 62.835 7.965 ;
      RECT 62.29 2.395 62.46 2.565 ;
      RECT 62.29 6.315 62.46 6.485 ;
      RECT 62.045 0.105 62.215 0.275 ;
      RECT 61.365 0.105 61.535 0.275 ;
      RECT 59.74 1.415 59.91 1.585 ;
      RECT 59.37 2.875 59.54 3.045 ;
      RECT 59.28 1.415 59.45 1.585 ;
      RECT 59.05 2.045 59.22 2.215 ;
      RECT 58.905 2.485 59.075 2.655 ;
      RECT 58.82 1.415 58.99 1.585 ;
      RECT 58.36 1.415 58.53 1.585 ;
      RECT 58.315 6.685 58.485 6.855 ;
      RECT 58.295 2.525 58.465 2.695 ;
      RECT 57.95 2.16 58.12 2.33 ;
      RECT 57.94 3.52 58.11 3.69 ;
      RECT 57.9 1.415 58.07 1.585 ;
      RECT 57.885 7.055 58.055 7.225 ;
      RECT 57.885 7.795 58.055 7.965 ;
      RECT 57.525 2.76 57.695 2.93 ;
      RECT 57.44 1.415 57.61 1.585 ;
      RECT 57.175 2.235 57.345 2.405 ;
      RECT 56.995 3.55 57.165 3.72 ;
      RECT 56.98 1.415 57.15 1.585 ;
      RECT 56.715 2.865 56.885 3.035 ;
      RECT 56.52 1.415 56.69 1.585 ;
      RECT 56.395 2.49 56.565 2.66 ;
      RECT 56.06 1.415 56.23 1.585 ;
      RECT 55.705 1.97 55.875 2.14 ;
      RECT 55.63 2.44 55.8 2.61 ;
      RECT 55.6 1.415 55.77 1.585 ;
      RECT 55.14 1.415 55.31 1.585 ;
      RECT 54.78 2.165 54.95 2.335 ;
      RECT 54.68 1.415 54.85 1.585 ;
      RECT 54.44 3.36 54.61 3.53 ;
      RECT 54.405 2.695 54.575 2.865 ;
      RECT 54.22 1.415 54.39 1.585 ;
      RECT 53.795 2.55 53.965 2.72 ;
      RECT 53.76 1.415 53.93 1.585 ;
      RECT 53.725 3.25 53.895 3.42 ;
      RECT 53.665 2.085 53.835 2.255 ;
      RECT 53.3 1.415 53.47 1.585 ;
      RECT 53.025 3 53.195 3.17 ;
      RECT 52.84 1.415 53.01 1.585 ;
      RECT 52.52 2.505 52.69 2.675 ;
      RECT 52.38 1.415 52.55 1.585 ;
      RECT 52.3 3.25 52.47 3.42 ;
      RECT 52.095 2.13 52.265 2.3 ;
      RECT 51.92 1.415 52.09 1.585 ;
      RECT 51.825 3 51.995 3.17 ;
      RECT 51.785 2.43 51.955 2.6 ;
      RECT 51.46 1.415 51.63 1.585 ;
      RECT 51.24 3.475 51.41 3.645 ;
      RECT 51.1 2.095 51.27 2.265 ;
      RECT 51 1.415 51.17 1.585 ;
      RECT 50.54 1.415 50.71 1.585 ;
      RECT 50.53 3.015 50.7 3.185 ;
      RECT 49.66 7.8 49.83 7.97 ;
      RECT 49.31 0.1 49.48 0.27 ;
      RECT 49.29 2.76 49.46 2.93 ;
      RECT 49.29 5.95 49.46 6.12 ;
      RECT 48.67 0.91 48.84 1.08 ;
      RECT 48.67 2.39 48.84 2.56 ;
      RECT 48.67 6.32 48.84 6.49 ;
      RECT 48.67 7.8 48.84 7.97 ;
      RECT 48.32 0.1 48.49 0.27 ;
      RECT 48.3 2.76 48.47 2.93 ;
      RECT 48.3 5.95 48.47 6.12 ;
      RECT 47.62 0.105 47.79 0.275 ;
      RECT 47.31 2.025 47.48 2.195 ;
      RECT 47.31 6.685 47.48 6.855 ;
      RECT 46.94 0.105 47.11 0.275 ;
      RECT 46.88 0.915 47.05 1.085 ;
      RECT 46.88 1.655 47.05 1.825 ;
      RECT 46.88 7.055 47.05 7.225 ;
      RECT 46.88 7.795 47.05 7.965 ;
      RECT 46.505 2.395 46.675 2.565 ;
      RECT 46.505 6.315 46.675 6.485 ;
      RECT 46.26 0.105 46.43 0.275 ;
      RECT 45.58 0.105 45.75 0.275 ;
      RECT 43.955 1.415 44.125 1.585 ;
      RECT 43.585 2.875 43.755 3.045 ;
      RECT 43.495 1.415 43.665 1.585 ;
      RECT 43.265 2.045 43.435 2.215 ;
      RECT 43.12 2.485 43.29 2.655 ;
      RECT 43.035 1.415 43.205 1.585 ;
      RECT 42.575 1.415 42.745 1.585 ;
      RECT 42.53 6.685 42.7 6.855 ;
      RECT 42.51 2.525 42.68 2.695 ;
      RECT 42.165 2.16 42.335 2.33 ;
      RECT 42.155 3.52 42.325 3.69 ;
      RECT 42.115 1.415 42.285 1.585 ;
      RECT 42.1 7.055 42.27 7.225 ;
      RECT 42.1 7.795 42.27 7.965 ;
      RECT 41.74 2.76 41.91 2.93 ;
      RECT 41.655 1.415 41.825 1.585 ;
      RECT 41.39 2.235 41.56 2.405 ;
      RECT 41.21 3.55 41.38 3.72 ;
      RECT 41.195 1.415 41.365 1.585 ;
      RECT 40.93 2.865 41.1 3.035 ;
      RECT 40.735 1.415 40.905 1.585 ;
      RECT 40.61 2.49 40.78 2.66 ;
      RECT 40.275 1.415 40.445 1.585 ;
      RECT 39.92 1.97 40.09 2.14 ;
      RECT 39.845 2.44 40.015 2.61 ;
      RECT 39.815 1.415 39.985 1.585 ;
      RECT 39.355 1.415 39.525 1.585 ;
      RECT 38.995 2.165 39.165 2.335 ;
      RECT 38.895 1.415 39.065 1.585 ;
      RECT 38.655 3.36 38.825 3.53 ;
      RECT 38.62 2.695 38.79 2.865 ;
      RECT 38.435 1.415 38.605 1.585 ;
      RECT 38.01 2.55 38.18 2.72 ;
      RECT 37.975 1.415 38.145 1.585 ;
      RECT 37.94 3.25 38.11 3.42 ;
      RECT 37.88 2.085 38.05 2.255 ;
      RECT 37.515 1.415 37.685 1.585 ;
      RECT 37.24 3 37.41 3.17 ;
      RECT 37.055 1.415 37.225 1.585 ;
      RECT 36.735 2.505 36.905 2.675 ;
      RECT 36.595 1.415 36.765 1.585 ;
      RECT 36.515 3.25 36.685 3.42 ;
      RECT 36.31 2.13 36.48 2.3 ;
      RECT 36.135 1.415 36.305 1.585 ;
      RECT 36.04 3 36.21 3.17 ;
      RECT 36 2.43 36.17 2.6 ;
      RECT 35.675 1.415 35.845 1.585 ;
      RECT 35.455 3.475 35.625 3.645 ;
      RECT 35.315 2.095 35.485 2.265 ;
      RECT 35.215 1.415 35.385 1.585 ;
      RECT 34.755 1.415 34.925 1.585 ;
      RECT 34.745 3.015 34.915 3.185 ;
      RECT 33.885 7.8 34.055 7.97 ;
      RECT 33.535 0.1 33.705 0.27 ;
      RECT 33.515 2.76 33.685 2.93 ;
      RECT 33.515 5.95 33.685 6.12 ;
      RECT 32.895 0.91 33.065 1.08 ;
      RECT 32.895 2.39 33.065 2.56 ;
      RECT 32.895 6.32 33.065 6.49 ;
      RECT 32.895 7.8 33.065 7.97 ;
      RECT 32.545 0.1 32.715 0.27 ;
      RECT 32.525 2.76 32.695 2.93 ;
      RECT 32.525 5.95 32.695 6.12 ;
      RECT 31.845 0.105 32.015 0.275 ;
      RECT 31.535 2.025 31.705 2.195 ;
      RECT 31.535 6.685 31.705 6.855 ;
      RECT 31.165 0.105 31.335 0.275 ;
      RECT 31.105 0.915 31.275 1.085 ;
      RECT 31.105 1.655 31.275 1.825 ;
      RECT 31.105 7.055 31.275 7.225 ;
      RECT 31.105 7.795 31.275 7.965 ;
      RECT 30.73 2.395 30.9 2.565 ;
      RECT 30.73 6.315 30.9 6.485 ;
      RECT 30.485 0.105 30.655 0.275 ;
      RECT 29.805 0.105 29.975 0.275 ;
      RECT 28.18 1.415 28.35 1.585 ;
      RECT 27.81 2.875 27.98 3.045 ;
      RECT 27.72 1.415 27.89 1.585 ;
      RECT 27.49 2.045 27.66 2.215 ;
      RECT 27.345 2.485 27.515 2.655 ;
      RECT 27.26 1.415 27.43 1.585 ;
      RECT 26.8 1.415 26.97 1.585 ;
      RECT 26.755 6.685 26.925 6.855 ;
      RECT 26.735 2.525 26.905 2.695 ;
      RECT 26.39 2.16 26.56 2.33 ;
      RECT 26.38 3.52 26.55 3.69 ;
      RECT 26.34 1.415 26.51 1.585 ;
      RECT 26.325 7.055 26.495 7.225 ;
      RECT 26.325 7.795 26.495 7.965 ;
      RECT 25.965 2.76 26.135 2.93 ;
      RECT 25.88 1.415 26.05 1.585 ;
      RECT 25.615 2.235 25.785 2.405 ;
      RECT 25.435 3.55 25.605 3.72 ;
      RECT 25.42 1.415 25.59 1.585 ;
      RECT 25.155 2.865 25.325 3.035 ;
      RECT 24.96 1.415 25.13 1.585 ;
      RECT 24.835 2.49 25.005 2.66 ;
      RECT 24.5 1.415 24.67 1.585 ;
      RECT 24.145 1.97 24.315 2.14 ;
      RECT 24.07 2.44 24.24 2.61 ;
      RECT 24.04 1.415 24.21 1.585 ;
      RECT 23.58 1.415 23.75 1.585 ;
      RECT 23.22 2.165 23.39 2.335 ;
      RECT 23.12 1.415 23.29 1.585 ;
      RECT 22.88 3.36 23.05 3.53 ;
      RECT 22.845 2.695 23.015 2.865 ;
      RECT 22.66 1.415 22.83 1.585 ;
      RECT 22.235 2.55 22.405 2.72 ;
      RECT 22.2 1.415 22.37 1.585 ;
      RECT 22.165 3.25 22.335 3.42 ;
      RECT 22.105 2.085 22.275 2.255 ;
      RECT 21.74 1.415 21.91 1.585 ;
      RECT 21.465 3 21.635 3.17 ;
      RECT 21.28 1.415 21.45 1.585 ;
      RECT 20.96 2.505 21.13 2.675 ;
      RECT 20.82 1.415 20.99 1.585 ;
      RECT 20.74 3.25 20.91 3.42 ;
      RECT 20.535 2.13 20.705 2.3 ;
      RECT 20.36 1.415 20.53 1.585 ;
      RECT 20.265 3 20.435 3.17 ;
      RECT 20.225 2.43 20.395 2.6 ;
      RECT 19.9 1.415 20.07 1.585 ;
      RECT 19.68 3.475 19.85 3.645 ;
      RECT 19.54 2.095 19.71 2.265 ;
      RECT 19.44 1.415 19.61 1.585 ;
      RECT 18.98 1.415 19.15 1.585 ;
      RECT 18.97 3.015 19.14 3.185 ;
      RECT 18.105 7.8 18.275 7.97 ;
      RECT 17.755 0.1 17.925 0.27 ;
      RECT 17.735 2.76 17.905 2.93 ;
      RECT 17.735 5.95 17.905 6.12 ;
      RECT 17.115 0.91 17.285 1.08 ;
      RECT 17.115 2.39 17.285 2.56 ;
      RECT 17.115 6.32 17.285 6.49 ;
      RECT 17.115 7.8 17.285 7.97 ;
      RECT 16.765 0.1 16.935 0.27 ;
      RECT 16.745 2.76 16.915 2.93 ;
      RECT 16.745 5.95 16.915 6.12 ;
      RECT 16.065 0.105 16.235 0.275 ;
      RECT 15.755 2.025 15.925 2.195 ;
      RECT 15.755 6.685 15.925 6.855 ;
      RECT 15.385 0.105 15.555 0.275 ;
      RECT 15.325 0.915 15.495 1.085 ;
      RECT 15.325 1.655 15.495 1.825 ;
      RECT 15.325 7.055 15.495 7.225 ;
      RECT 15.325 7.795 15.495 7.965 ;
      RECT 14.95 2.395 15.12 2.565 ;
      RECT 14.95 6.315 15.12 6.485 ;
      RECT 14.705 0.105 14.875 0.275 ;
      RECT 14.025 0.105 14.195 0.275 ;
      RECT 12.4 1.415 12.57 1.585 ;
      RECT 12.03 2.875 12.2 3.045 ;
      RECT 11.94 1.415 12.11 1.585 ;
      RECT 11.71 2.045 11.88 2.215 ;
      RECT 11.565 2.485 11.735 2.655 ;
      RECT 11.48 1.415 11.65 1.585 ;
      RECT 11.02 1.415 11.19 1.585 ;
      RECT 10.975 6.685 11.145 6.855 ;
      RECT 10.955 2.525 11.125 2.695 ;
      RECT 10.61 2.16 10.78 2.33 ;
      RECT 10.6 3.52 10.77 3.69 ;
      RECT 10.56 1.415 10.73 1.585 ;
      RECT 10.545 7.055 10.715 7.225 ;
      RECT 10.545 7.795 10.715 7.965 ;
      RECT 10.185 2.76 10.355 2.93 ;
      RECT 10.1 1.415 10.27 1.585 ;
      RECT 9.835 2.235 10.005 2.405 ;
      RECT 9.655 3.55 9.825 3.72 ;
      RECT 9.64 1.415 9.81 1.585 ;
      RECT 9.375 2.865 9.545 3.035 ;
      RECT 9.18 1.415 9.35 1.585 ;
      RECT 9.055 2.49 9.225 2.66 ;
      RECT 8.72 1.415 8.89 1.585 ;
      RECT 8.365 1.97 8.535 2.14 ;
      RECT 8.29 2.44 8.46 2.61 ;
      RECT 8.26 1.415 8.43 1.585 ;
      RECT 7.8 1.415 7.97 1.585 ;
      RECT 7.44 2.165 7.61 2.335 ;
      RECT 7.34 1.415 7.51 1.585 ;
      RECT 7.1 3.36 7.27 3.53 ;
      RECT 7.065 2.695 7.235 2.865 ;
      RECT 6.88 1.415 7.05 1.585 ;
      RECT 6.455 2.55 6.625 2.72 ;
      RECT 6.42 1.415 6.59 1.585 ;
      RECT 6.385 3.25 6.555 3.42 ;
      RECT 6.325 2.085 6.495 2.255 ;
      RECT 5.96 1.415 6.13 1.585 ;
      RECT 5.685 3 5.855 3.17 ;
      RECT 5.5 1.415 5.67 1.585 ;
      RECT 5.18 2.505 5.35 2.675 ;
      RECT 5.04 1.415 5.21 1.585 ;
      RECT 4.96 3.25 5.13 3.42 ;
      RECT 4.755 2.13 4.925 2.3 ;
      RECT 4.58 1.415 4.75 1.585 ;
      RECT 4.485 3 4.655 3.17 ;
      RECT 4.445 2.43 4.615 2.6 ;
      RECT 4.12 1.415 4.29 1.585 ;
      RECT 3.9 3.475 4.07 3.645 ;
      RECT 3.76 2.095 3.93 2.265 ;
      RECT 3.66 1.415 3.83 1.585 ;
      RECT 3.2 1.415 3.37 1.585 ;
      RECT 3.19 3.015 3.36 3.185 ;
      RECT 1.61 7.055 1.78 7.225 ;
      RECT 1.61 7.795 1.78 7.965 ;
      RECT 1.235 6.315 1.405 6.485 ;
    LAYER li1 ;
      RECT 74.31 0 74.48 2.085 ;
      RECT 72.35 0 72.52 2.085 ;
      RECT 69.91 0 70.08 2.085 ;
      RECT 68.95 0 69.12 2.085 ;
      RECT 68.43 0 68.6 2.085 ;
      RECT 67.47 0 67.64 2.085 ;
      RECT 66.51 0 66.68 2.085 ;
      RECT 58.525 0 58.695 2.085 ;
      RECT 56.565 0 56.735 2.085 ;
      RECT 54.125 0 54.295 2.085 ;
      RECT 53.165 0 53.335 2.085 ;
      RECT 52.645 0 52.815 2.085 ;
      RECT 51.685 0 51.855 2.085 ;
      RECT 50.725 0 50.895 2.085 ;
      RECT 42.74 0 42.91 2.085 ;
      RECT 40.78 0 40.95 2.085 ;
      RECT 38.34 0 38.51 2.085 ;
      RECT 37.38 0 37.55 2.085 ;
      RECT 36.86 0 37.03 2.085 ;
      RECT 35.9 0 36.07 2.085 ;
      RECT 34.94 0 35.11 2.085 ;
      RECT 26.965 0 27.135 2.085 ;
      RECT 25.005 0 25.175 2.085 ;
      RECT 22.565 0 22.735 2.085 ;
      RECT 21.605 0 21.775 2.085 ;
      RECT 21.085 0 21.255 2.085 ;
      RECT 20.125 0 20.295 2.085 ;
      RECT 19.165 0 19.335 2.085 ;
      RECT 11.185 0 11.355 2.085 ;
      RECT 9.225 0 9.395 2.085 ;
      RECT 6.785 0 6.955 2.085 ;
      RECT 5.825 0 5.995 2.085 ;
      RECT 5.305 0 5.475 2.085 ;
      RECT 4.345 0 4.515 2.085 ;
      RECT 3.385 0 3.555 2.085 ;
      RECT 66.295 0 75.895 1.59 ;
      RECT 50.51 0 60.11 1.59 ;
      RECT 34.725 0 44.325 1.59 ;
      RECT 18.95 0 28.55 1.59 ;
      RECT 3.17 0 12.77 1.59 ;
      RECT 66.18 1.415 76.01 1.585 ;
      RECT 66.295 0 76.01 1.585 ;
      RECT 50.395 1.415 60.225 1.585 ;
      RECT 50.51 0 60.225 1.585 ;
      RECT 34.61 1.415 44.44 1.585 ;
      RECT 34.725 0 44.44 1.585 ;
      RECT 18.835 1.415 28.665 1.585 ;
      RECT 18.95 0 28.665 1.585 ;
      RECT 3.055 1.415 12.885 1.585 ;
      RECT 3.17 0 12.885 1.585 ;
      RECT 77.07 0 77.24 0.935 ;
      RECT 61.285 0 61.455 0.935 ;
      RECT 45.5 0 45.67 0.935 ;
      RECT 29.725 0 29.895 0.935 ;
      RECT 13.945 0 14.115 0.935 ;
      RECT 80.8 0 80.97 0.93 ;
      RECT 79.81 0 79.98 0.93 ;
      RECT 65.015 0 65.185 0.93 ;
      RECT 64.025 0 64.195 0.93 ;
      RECT 49.23 0 49.4 0.93 ;
      RECT 48.24 0 48.41 0.93 ;
      RECT 33.455 0 33.625 0.93 ;
      RECT 32.465 0 32.635 0.93 ;
      RECT 17.675 0 17.845 0.93 ;
      RECT 16.685 0 16.855 0.93 ;
      RECT 81.595 0 81.775 0.305 ;
      RECT 65.81 0 79.645 0.305 ;
      RECT 50.025 0 63.86 0.305 ;
      RECT 34.25 0 48.075 0.305 ;
      RECT 18.47 0 32.3 0.305 ;
      RECT 0 0 16.52 0.305 ;
      RECT 0 0 81.775 0.3 ;
      RECT 81.23 5.02 81.4 6.49 ;
      RECT 81.23 6.315 81.405 6.485 ;
      RECT 80.86 1.74 81.03 2.93 ;
      RECT 80.86 1.74 81.33 1.91 ;
      RECT 80.86 6.97 81.33 7.14 ;
      RECT 80.86 5.95 81.03 7.14 ;
      RECT 79.87 1.74 80.04 2.93 ;
      RECT 79.87 1.74 80.34 1.91 ;
      RECT 79.87 6.97 80.34 7.14 ;
      RECT 79.87 5.95 80.04 7.14 ;
      RECT 78.02 2.635 78.19 3.865 ;
      RECT 78.075 0.855 78.245 2.805 ;
      RECT 78.02 0.575 78.19 1.025 ;
      RECT 78.02 7.855 78.19 8.305 ;
      RECT 78.075 6.075 78.245 8.025 ;
      RECT 78.02 5.015 78.19 6.245 ;
      RECT 77.5 0.575 77.67 3.865 ;
      RECT 77.5 2.075 77.905 2.405 ;
      RECT 77.5 1.235 77.905 1.565 ;
      RECT 77.5 5.015 77.67 8.305 ;
      RECT 77.5 7.315 77.905 7.645 ;
      RECT 77.5 6.475 77.905 6.805 ;
      RECT 74.835 1.975 75.565 2.215 ;
      RECT 75.377 1.77 75.565 2.215 ;
      RECT 75.205 1.782 75.58 2.209 ;
      RECT 75.12 1.797 75.6 2.194 ;
      RECT 75.12 1.812 75.605 2.184 ;
      RECT 75.075 1.832 75.62 2.176 ;
      RECT 75.052 1.867 75.635 2.13 ;
      RECT 74.966 1.89 75.64 2.09 ;
      RECT 74.966 1.908 75.65 2.06 ;
      RECT 74.835 1.977 75.655 2.023 ;
      RECT 74.88 1.92 75.65 2.06 ;
      RECT 74.966 1.872 75.635 2.13 ;
      RECT 75.052 1.841 75.62 2.176 ;
      RECT 75.075 1.822 75.605 2.184 ;
      RECT 75.12 1.795 75.58 2.209 ;
      RECT 75.205 1.777 75.565 2.215 ;
      RECT 75.291 1.771 75.565 2.215 ;
      RECT 75.377 1.766 75.51 2.215 ;
      RECT 75.463 1.761 75.51 2.215 ;
      RECT 75.155 2.659 75.325 3.045 ;
      RECT 75.15 2.659 75.325 3.04 ;
      RECT 75.125 2.659 75.325 3.005 ;
      RECT 75.125 2.687 75.335 2.995 ;
      RECT 75.105 2.687 75.335 2.955 ;
      RECT 75.1 2.687 75.335 2.928 ;
      RECT 75.1 2.705 75.34 2.92 ;
      RECT 75.045 2.705 75.34 2.855 ;
      RECT 75.045 2.722 75.35 2.838 ;
      RECT 75.035 2.722 75.35 2.778 ;
      RECT 75.035 2.739 75.355 2.775 ;
      RECT 75.03 2.575 75.2 2.753 ;
      RECT 75.03 2.609 75.286 2.753 ;
      RECT 75.025 3.375 75.03 3.388 ;
      RECT 75.02 3.27 75.025 3.393 ;
      RECT 74.995 3.13 75.02 3.408 ;
      RECT 74.96 3.081 74.995 3.44 ;
      RECT 74.955 3.049 74.96 3.46 ;
      RECT 74.95 3.04 74.955 3.46 ;
      RECT 74.87 3.005 74.95 3.46 ;
      RECT 74.807 2.975 74.87 3.46 ;
      RECT 74.721 2.963 74.807 3.46 ;
      RECT 74.635 2.949 74.721 3.46 ;
      RECT 74.555 2.936 74.635 3.446 ;
      RECT 74.52 2.928 74.555 3.426 ;
      RECT 74.51 2.925 74.52 3.417 ;
      RECT 74.48 2.92 74.51 3.404 ;
      RECT 74.43 2.895 74.48 3.38 ;
      RECT 74.416 2.869 74.43 3.362 ;
      RECT 74.33 2.829 74.416 3.338 ;
      RECT 74.285 2.777 74.33 3.307 ;
      RECT 74.275 2.752 74.285 3.294 ;
      RECT 74.27 2.533 74.275 2.555 ;
      RECT 74.265 2.735 74.275 3.29 ;
      RECT 74.265 2.531 74.27 2.645 ;
      RECT 74.255 2.527 74.265 3.286 ;
      RECT 74.211 2.525 74.255 3.274 ;
      RECT 74.125 2.525 74.211 3.245 ;
      RECT 74.095 2.525 74.125 3.218 ;
      RECT 74.08 2.525 74.095 3.206 ;
      RECT 74.04 2.537 74.08 3.191 ;
      RECT 74.02 2.556 74.04 3.17 ;
      RECT 74.01 2.566 74.02 3.154 ;
      RECT 74 2.572 74.01 3.143 ;
      RECT 73.98 2.582 74 3.126 ;
      RECT 73.975 2.591 73.98 3.113 ;
      RECT 73.97 2.595 73.975 3.063 ;
      RECT 73.96 2.601 73.97 2.98 ;
      RECT 73.955 2.605 73.96 2.894 ;
      RECT 73.95 2.625 73.955 2.831 ;
      RECT 73.945 2.648 73.95 2.778 ;
      RECT 73.94 2.666 73.945 2.723 ;
      RECT 74.55 2.485 74.72 2.745 ;
      RECT 74.72 2.45 74.765 2.731 ;
      RECT 74.681 2.452 74.77 2.714 ;
      RECT 74.57 2.469 74.856 2.685 ;
      RECT 74.57 2.484 74.86 2.657 ;
      RECT 74.57 2.465 74.77 2.714 ;
      RECT 74.595 2.453 74.72 2.745 ;
      RECT 74.681 2.451 74.765 2.731 ;
      RECT 73.735 1.84 73.905 2.33 ;
      RECT 73.735 1.84 73.94 2.31 ;
      RECT 73.87 1.76 73.98 2.27 ;
      RECT 73.851 1.764 74 2.24 ;
      RECT 73.765 1.772 74.02 2.223 ;
      RECT 73.765 1.778 74.025 2.213 ;
      RECT 73.765 1.787 74.045 2.201 ;
      RECT 73.74 1.812 74.075 2.179 ;
      RECT 73.74 1.832 74.08 2.159 ;
      RECT 73.735 1.845 74.09 2.139 ;
      RECT 73.735 1.912 74.095 2.12 ;
      RECT 73.735 2.045 74.1 2.107 ;
      RECT 73.73 1.85 74.09 1.94 ;
      RECT 73.74 1.807 74.045 2.201 ;
      RECT 73.851 1.762 73.98 2.27 ;
      RECT 73.725 3.515 74.025 3.77 ;
      RECT 73.81 3.481 74.025 3.77 ;
      RECT 73.81 3.484 74.03 3.63 ;
      RECT 73.745 3.505 74.03 3.63 ;
      RECT 73.78 3.495 74.025 3.77 ;
      RECT 73.775 3.5 74.03 3.63 ;
      RECT 73.81 3.479 74.011 3.77 ;
      RECT 73.896 3.47 74.011 3.77 ;
      RECT 73.896 3.464 73.925 3.77 ;
      RECT 73.385 3.105 73.395 3.595 ;
      RECT 73.045 3.04 73.055 3.34 ;
      RECT 73.56 3.212 73.565 3.431 ;
      RECT 73.55 3.192 73.56 3.448 ;
      RECT 73.54 3.172 73.55 3.478 ;
      RECT 73.535 3.162 73.54 3.493 ;
      RECT 73.53 3.158 73.535 3.498 ;
      RECT 73.515 3.15 73.53 3.505 ;
      RECT 73.475 3.13 73.515 3.53 ;
      RECT 73.45 3.112 73.475 3.563 ;
      RECT 73.445 3.11 73.45 3.576 ;
      RECT 73.425 3.107 73.445 3.58 ;
      RECT 73.395 3.105 73.425 3.59 ;
      RECT 73.325 3.107 73.385 3.591 ;
      RECT 73.305 3.107 73.325 3.585 ;
      RECT 73.28 3.105 73.305 3.582 ;
      RECT 73.245 3.1 73.28 3.578 ;
      RECT 73.225 3.094 73.245 3.565 ;
      RECT 73.215 3.091 73.225 3.553 ;
      RECT 73.195 3.088 73.215 3.538 ;
      RECT 73.175 3.084 73.195 3.52 ;
      RECT 73.17 3.081 73.175 3.51 ;
      RECT 73.165 3.08 73.17 3.508 ;
      RECT 73.155 3.077 73.165 3.5 ;
      RECT 73.145 3.071 73.155 3.483 ;
      RECT 73.135 3.065 73.145 3.465 ;
      RECT 73.125 3.059 73.135 3.453 ;
      RECT 73.115 3.053 73.125 3.433 ;
      RECT 73.11 3.049 73.115 3.418 ;
      RECT 73.105 3.047 73.11 3.41 ;
      RECT 73.1 3.045 73.105 3.403 ;
      RECT 73.095 3.043 73.1 3.393 ;
      RECT 73.09 3.041 73.095 3.387 ;
      RECT 73.08 3.04 73.09 3.377 ;
      RECT 73.07 3.04 73.08 3.368 ;
      RECT 73.055 3.04 73.07 3.353 ;
      RECT 73.015 3.04 73.045 3.337 ;
      RECT 72.995 3.042 73.015 3.332 ;
      RECT 72.99 3.047 72.995 3.33 ;
      RECT 72.96 3.055 72.99 3.328 ;
      RECT 72.93 3.07 72.96 3.327 ;
      RECT 72.885 3.092 72.93 3.332 ;
      RECT 72.88 3.107 72.885 3.336 ;
      RECT 72.865 3.112 72.88 3.338 ;
      RECT 72.86 3.116 72.865 3.34 ;
      RECT 72.8 3.139 72.86 3.349 ;
      RECT 72.78 3.165 72.8 3.362 ;
      RECT 72.77 3.172 72.78 3.366 ;
      RECT 72.755 3.179 72.77 3.369 ;
      RECT 72.735 3.189 72.755 3.372 ;
      RECT 72.73 3.197 72.735 3.375 ;
      RECT 72.685 3.202 72.73 3.382 ;
      RECT 72.675 3.205 72.685 3.389 ;
      RECT 72.665 3.205 72.675 3.393 ;
      RECT 72.63 3.207 72.665 3.405 ;
      RECT 72.61 3.21 72.63 3.418 ;
      RECT 72.57 3.213 72.61 3.429 ;
      RECT 72.555 3.215 72.57 3.442 ;
      RECT 72.545 3.215 72.555 3.447 ;
      RECT 72.52 3.216 72.545 3.455 ;
      RECT 72.51 3.218 72.52 3.46 ;
      RECT 72.505 3.219 72.51 3.463 ;
      RECT 72.48 3.217 72.505 3.466 ;
      RECT 72.465 3.215 72.48 3.467 ;
      RECT 72.445 3.212 72.465 3.469 ;
      RECT 72.425 3.207 72.445 3.469 ;
      RECT 72.365 3.202 72.425 3.466 ;
      RECT 72.33 3.177 72.365 3.462 ;
      RECT 72.32 3.154 72.33 3.46 ;
      RECT 72.29 3.131 72.32 3.46 ;
      RECT 72.28 3.11 72.29 3.46 ;
      RECT 72.255 3.092 72.28 3.458 ;
      RECT 72.24 3.07 72.255 3.455 ;
      RECT 72.225 3.052 72.24 3.453 ;
      RECT 72.205 3.042 72.225 3.451 ;
      RECT 72.19 3.037 72.205 3.45 ;
      RECT 72.175 3.035 72.19 3.449 ;
      RECT 72.145 3.036 72.175 3.447 ;
      RECT 72.125 3.039 72.145 3.445 ;
      RECT 72.068 3.043 72.125 3.445 ;
      RECT 71.982 3.052 72.068 3.445 ;
      RECT 71.896 3.063 71.982 3.445 ;
      RECT 71.81 3.074 71.896 3.445 ;
      RECT 71.79 3.081 71.81 3.453 ;
      RECT 71.78 3.084 71.79 3.46 ;
      RECT 71.715 3.089 71.78 3.478 ;
      RECT 71.685 3.096 71.715 3.503 ;
      RECT 71.675 3.099 71.685 3.51 ;
      RECT 71.63 3.103 71.675 3.515 ;
      RECT 71.6 3.108 71.63 3.52 ;
      RECT 71.599 3.11 71.6 3.52 ;
      RECT 71.513 3.116 71.599 3.52 ;
      RECT 71.427 3.127 71.513 3.52 ;
      RECT 71.341 3.139 71.427 3.52 ;
      RECT 71.255 3.15 71.341 3.52 ;
      RECT 71.24 3.157 71.255 3.515 ;
      RECT 71.235 3.159 71.24 3.509 ;
      RECT 71.215 3.17 71.235 3.504 ;
      RECT 71.205 3.188 71.215 3.498 ;
      RECT 71.2 3.2 71.205 3.298 ;
      RECT 73.495 1.953 73.515 2.04 ;
      RECT 73.49 1.888 73.495 2.072 ;
      RECT 73.48 1.855 73.49 2.077 ;
      RECT 73.475 1.835 73.48 2.083 ;
      RECT 73.445 1.835 73.475 2.1 ;
      RECT 73.396 1.835 73.445 2.136 ;
      RECT 73.31 1.835 73.396 2.194 ;
      RECT 73.281 1.845 73.31 2.243 ;
      RECT 73.195 1.887 73.281 2.296 ;
      RECT 73.175 1.925 73.195 2.343 ;
      RECT 73.15 1.942 73.175 2.363 ;
      RECT 73.14 1.956 73.15 2.383 ;
      RECT 73.135 1.962 73.14 2.393 ;
      RECT 73.13 1.966 73.135 2.4 ;
      RECT 73.08 1.986 73.13 2.405 ;
      RECT 73.015 2.03 73.08 2.405 ;
      RECT 72.99 2.08 73.015 2.405 ;
      RECT 72.98 2.11 72.99 2.405 ;
      RECT 72.975 2.137 72.98 2.405 ;
      RECT 72.97 2.155 72.975 2.405 ;
      RECT 72.96 2.197 72.97 2.405 ;
      RECT 73.31 2.755 73.48 2.93 ;
      RECT 73.25 2.583 73.31 2.918 ;
      RECT 73.24 2.576 73.25 2.901 ;
      RECT 73.195 2.755 73.48 2.881 ;
      RECT 73.176 2.755 73.48 2.859 ;
      RECT 73.09 2.755 73.48 2.824 ;
      RECT 73.07 2.575 73.24 2.78 ;
      RECT 73.07 2.722 73.475 2.78 ;
      RECT 73.07 2.67 73.45 2.78 ;
      RECT 73.07 2.625 73.415 2.78 ;
      RECT 73.07 2.607 73.38 2.78 ;
      RECT 73.07 2.597 73.375 2.78 ;
      RECT 72.72 5.015 72.89 8.305 ;
      RECT 72.72 7.315 73.125 7.645 ;
      RECT 72.72 6.475 73.125 6.805 ;
      RECT 72.79 3.555 72.98 3.78 ;
      RECT 72.78 3.556 72.985 3.775 ;
      RECT 72.78 3.558 72.995 3.755 ;
      RECT 72.78 3.562 73 3.74 ;
      RECT 72.78 3.549 72.95 3.775 ;
      RECT 72.78 3.552 72.975 3.775 ;
      RECT 72.79 3.548 72.95 3.78 ;
      RECT 72.876 3.546 72.95 3.78 ;
      RECT 72.5 2.797 72.67 3.035 ;
      RECT 72.5 2.797 72.756 2.949 ;
      RECT 72.5 2.797 72.76 2.859 ;
      RECT 72.55 2.57 72.77 2.838 ;
      RECT 72.545 2.587 72.775 2.811 ;
      RECT 72.51 2.745 72.775 2.811 ;
      RECT 72.53 2.595 72.67 3.035 ;
      RECT 72.52 2.677 72.78 2.794 ;
      RECT 72.515 2.725 72.78 2.794 ;
      RECT 72.52 2.635 72.775 2.811 ;
      RECT 72.545 2.572 72.77 2.838 ;
      RECT 72.11 2.547 72.28 2.745 ;
      RECT 72.11 2.547 72.325 2.72 ;
      RECT 72.18 2.49 72.35 2.678 ;
      RECT 72.155 2.505 72.35 2.678 ;
      RECT 71.77 2.551 71.8 2.745 ;
      RECT 71.765 2.523 71.77 2.745 ;
      RECT 71.735 2.497 71.765 2.747 ;
      RECT 71.71 2.455 71.735 2.75 ;
      RECT 71.7 2.427 71.71 2.752 ;
      RECT 71.665 2.407 71.7 2.754 ;
      RECT 71.6 2.392 71.665 2.76 ;
      RECT 71.55 2.39 71.6 2.766 ;
      RECT 71.527 2.392 71.55 2.771 ;
      RECT 71.441 2.403 71.527 2.777 ;
      RECT 71.355 2.421 71.441 2.787 ;
      RECT 71.34 2.432 71.355 2.793 ;
      RECT 71.27 2.455 71.34 2.799 ;
      RECT 71.215 2.487 71.27 2.807 ;
      RECT 71.175 2.51 71.215 2.813 ;
      RECT 71.161 2.523 71.175 2.816 ;
      RECT 71.075 2.545 71.161 2.822 ;
      RECT 71.06 2.57 71.075 2.828 ;
      RECT 71.02 2.585 71.06 2.832 ;
      RECT 70.97 2.6 71.02 2.837 ;
      RECT 70.945 2.607 70.97 2.841 ;
      RECT 70.885 2.602 70.945 2.845 ;
      RECT 70.87 2.593 70.885 2.849 ;
      RECT 70.8 2.583 70.87 2.845 ;
      RECT 70.775 2.575 70.795 2.835 ;
      RECT 70.716 2.575 70.775 2.813 ;
      RECT 70.63 2.575 70.716 2.77 ;
      RECT 70.795 2.575 70.8 2.84 ;
      RECT 71.49 1.806 71.66 2.14 ;
      RECT 71.46 1.806 71.66 2.135 ;
      RECT 71.4 1.773 71.46 2.123 ;
      RECT 71.4 1.829 71.67 2.118 ;
      RECT 71.375 1.829 71.67 2.112 ;
      RECT 71.37 1.77 71.4 2.109 ;
      RECT 71.355 1.776 71.49 2.107 ;
      RECT 71.35 1.784 71.575 2.095 ;
      RECT 71.35 1.836 71.685 2.048 ;
      RECT 71.335 1.792 71.575 2.043 ;
      RECT 71.335 1.862 71.695 1.984 ;
      RECT 71.305 1.812 71.66 1.945 ;
      RECT 71.305 1.902 71.705 1.941 ;
      RECT 71.355 1.781 71.575 2.107 ;
      RECT 70.695 2.111 70.75 2.375 ;
      RECT 70.695 2.111 70.815 2.374 ;
      RECT 70.695 2.111 70.84 2.373 ;
      RECT 70.695 2.111 70.905 2.372 ;
      RECT 70.84 2.077 70.92 2.371 ;
      RECT 70.655 2.121 71.065 2.37 ;
      RECT 70.695 2.118 71.065 2.37 ;
      RECT 70.655 2.126 71.07 2.363 ;
      RECT 70.64 2.128 71.07 2.362 ;
      RECT 70.64 2.135 71.075 2.358 ;
      RECT 70.62 2.134 71.07 2.354 ;
      RECT 70.62 2.142 71.08 2.353 ;
      RECT 70.615 2.139 71.075 2.349 ;
      RECT 70.615 2.152 71.09 2.348 ;
      RECT 70.6 2.142 71.08 2.347 ;
      RECT 70.565 2.155 71.09 2.34 ;
      RECT 70.75 2.11 71.06 2.37 ;
      RECT 70.75 2.095 71.01 2.37 ;
      RECT 70.815 2.082 70.945 2.37 ;
      RECT 70.36 3.171 70.375 3.564 ;
      RECT 70.325 3.176 70.375 3.563 ;
      RECT 70.36 3.175 70.42 3.562 ;
      RECT 70.305 3.186 70.42 3.561 ;
      RECT 70.32 3.182 70.42 3.561 ;
      RECT 70.285 3.192 70.495 3.558 ;
      RECT 70.285 3.211 70.54 3.556 ;
      RECT 70.285 3.218 70.545 3.553 ;
      RECT 70.27 3.195 70.495 3.55 ;
      RECT 70.25 3.2 70.495 3.543 ;
      RECT 70.245 3.204 70.495 3.539 ;
      RECT 70.245 3.221 70.555 3.538 ;
      RECT 70.225 3.215 70.54 3.534 ;
      RECT 70.225 3.224 70.56 3.528 ;
      RECT 70.22 3.23 70.56 3.3 ;
      RECT 70.285 3.19 70.42 3.558 ;
      RECT 70.16 2.553 70.36 2.865 ;
      RECT 70.235 2.531 70.36 2.865 ;
      RECT 70.175 2.55 70.365 2.85 ;
      RECT 70.145 2.561 70.365 2.848 ;
      RECT 70.16 2.556 70.37 2.814 ;
      RECT 70.145 2.66 70.375 2.781 ;
      RECT 70.175 2.532 70.36 2.865 ;
      RECT 70.235 2.51 70.335 2.865 ;
      RECT 70.26 2.507 70.335 2.865 ;
      RECT 70.26 2.502 70.28 2.865 ;
      RECT 69.665 2.57 69.84 2.745 ;
      RECT 69.66 2.57 69.84 2.743 ;
      RECT 69.635 2.57 69.84 2.738 ;
      RECT 69.58 2.55 69.75 2.728 ;
      RECT 69.58 2.557 69.815 2.728 ;
      RECT 69.665 3.237 69.68 3.42 ;
      RECT 69.655 3.215 69.665 3.42 ;
      RECT 69.64 3.195 69.655 3.42 ;
      RECT 69.63 3.17 69.64 3.42 ;
      RECT 69.6 3.135 69.63 3.42 ;
      RECT 69.565 3.075 69.6 3.42 ;
      RECT 69.56 3.037 69.565 3.42 ;
      RECT 69.51 2.988 69.56 3.42 ;
      RECT 69.5 2.938 69.51 3.408 ;
      RECT 69.485 2.917 69.5 3.368 ;
      RECT 69.465 2.885 69.485 3.318 ;
      RECT 69.44 2.841 69.465 3.258 ;
      RECT 69.435 2.813 69.44 3.213 ;
      RECT 69.43 2.804 69.435 3.199 ;
      RECT 69.425 2.797 69.43 3.186 ;
      RECT 69.42 2.792 69.425 3.175 ;
      RECT 69.415 2.777 69.42 3.165 ;
      RECT 69.41 2.755 69.415 3.152 ;
      RECT 69.4 2.715 69.41 3.127 ;
      RECT 69.375 2.645 69.4 3.083 ;
      RECT 69.37 2.585 69.375 3.048 ;
      RECT 69.355 2.565 69.37 3.015 ;
      RECT 69.35 2.565 69.355 2.99 ;
      RECT 69.32 2.565 69.35 2.945 ;
      RECT 69.275 2.565 69.32 2.885 ;
      RECT 69.2 2.565 69.275 2.833 ;
      RECT 69.195 2.565 69.2 2.798 ;
      RECT 69.19 2.565 69.195 2.788 ;
      RECT 69.185 2.565 69.19 2.768 ;
      RECT 69.45 1.785 69.62 2.255 ;
      RECT 69.395 1.778 69.59 2.239 ;
      RECT 69.395 1.792 69.625 2.238 ;
      RECT 69.38 1.793 69.625 2.219 ;
      RECT 69.375 1.811 69.625 2.205 ;
      RECT 69.38 1.794 69.63 2.203 ;
      RECT 69.365 1.825 69.63 2.188 ;
      RECT 69.38 1.8 69.635 2.173 ;
      RECT 69.36 1.84 69.635 2.17 ;
      RECT 69.375 1.812 69.64 2.155 ;
      RECT 69.375 1.824 69.645 2.135 ;
      RECT 69.36 1.84 69.65 2.118 ;
      RECT 69.36 1.85 69.655 1.973 ;
      RECT 69.355 1.85 69.655 1.93 ;
      RECT 69.355 1.865 69.66 1.908 ;
      RECT 69.45 1.775 69.59 2.255 ;
      RECT 69.45 1.773 69.56 2.255 ;
      RECT 69.536 1.77 69.56 2.255 ;
      RECT 69.195 3.437 69.2 3.483 ;
      RECT 69.185 3.285 69.195 3.507 ;
      RECT 69.18 3.13 69.185 3.532 ;
      RECT 69.165 3.092 69.18 3.543 ;
      RECT 69.16 3.075 69.165 3.55 ;
      RECT 69.15 3.063 69.16 3.557 ;
      RECT 69.145 3.054 69.15 3.559 ;
      RECT 69.14 3.052 69.145 3.563 ;
      RECT 69.095 3.043 69.14 3.578 ;
      RECT 69.09 3.035 69.095 3.592 ;
      RECT 69.085 3.032 69.09 3.596 ;
      RECT 69.07 3.027 69.085 3.604 ;
      RECT 69.015 3.017 69.07 3.615 ;
      RECT 68.98 3.005 69.015 3.616 ;
      RECT 68.971 3 68.98 3.61 ;
      RECT 68.885 3 68.971 3.6 ;
      RECT 68.855 3 68.885 3.578 ;
      RECT 68.845 3 68.85 3.558 ;
      RECT 68.84 3 68.845 3.52 ;
      RECT 68.835 3 68.84 3.478 ;
      RECT 68.83 3 68.835 3.438 ;
      RECT 68.825 3 68.83 3.368 ;
      RECT 68.815 3 68.825 3.29 ;
      RECT 68.81 3 68.815 3.19 ;
      RECT 68.85 3 68.855 3.56 ;
      RECT 68.345 3.082 68.435 3.56 ;
      RECT 68.33 3.085 68.45 3.558 ;
      RECT 68.345 3.084 68.45 3.558 ;
      RECT 68.31 3.091 68.475 3.548 ;
      RECT 68.33 3.085 68.475 3.548 ;
      RECT 68.295 3.097 68.475 3.536 ;
      RECT 68.33 3.088 68.525 3.529 ;
      RECT 68.281 3.105 68.525 3.527 ;
      RECT 68.31 3.095 68.535 3.515 ;
      RECT 68.281 3.116 68.565 3.506 ;
      RECT 68.195 3.14 68.565 3.5 ;
      RECT 68.195 3.153 68.605 3.483 ;
      RECT 68.19 3.175 68.605 3.476 ;
      RECT 68.16 3.19 68.605 3.466 ;
      RECT 68.155 3.201 68.605 3.456 ;
      RECT 68.125 3.214 68.605 3.447 ;
      RECT 68.11 3.232 68.605 3.436 ;
      RECT 68.085 3.245 68.605 3.426 ;
      RECT 68.345 3.081 68.355 3.56 ;
      RECT 68.391 2.505 68.43 2.75 ;
      RECT 68.305 2.505 68.44 2.748 ;
      RECT 68.19 2.53 68.44 2.745 ;
      RECT 68.19 2.53 68.445 2.743 ;
      RECT 68.19 2.53 68.46 2.738 ;
      RECT 68.296 2.505 68.475 2.718 ;
      RECT 68.21 2.513 68.475 2.718 ;
      RECT 67.88 1.865 68.05 2.3 ;
      RECT 67.87 1.899 68.05 2.283 ;
      RECT 67.95 1.835 68.12 2.27 ;
      RECT 67.855 1.91 68.12 2.248 ;
      RECT 67.95 1.845 68.125 2.238 ;
      RECT 67.88 1.897 68.155 2.223 ;
      RECT 67.84 1.923 68.155 2.208 ;
      RECT 67.84 1.965 68.165 2.188 ;
      RECT 67.835 1.99 68.17 2.17 ;
      RECT 67.835 2 68.175 2.155 ;
      RECT 67.83 1.937 68.155 2.153 ;
      RECT 67.83 2.01 68.18 2.138 ;
      RECT 67.825 1.947 68.155 2.135 ;
      RECT 67.82 2.031 68.185 2.118 ;
      RECT 67.82 2.063 68.19 2.098 ;
      RECT 67.815 1.977 68.165 2.09 ;
      RECT 67.82 1.962 68.155 2.118 ;
      RECT 67.835 1.932 68.155 2.17 ;
      RECT 67.68 2.519 67.905 2.775 ;
      RECT 67.68 2.552 67.925 2.765 ;
      RECT 67.645 2.552 67.925 2.763 ;
      RECT 67.645 2.565 67.93 2.753 ;
      RECT 67.645 2.585 67.94 2.745 ;
      RECT 67.645 2.682 67.945 2.738 ;
      RECT 67.625 2.43 67.755 2.728 ;
      RECT 67.58 2.585 67.94 2.67 ;
      RECT 67.57 2.43 67.755 2.615 ;
      RECT 67.57 2.462 67.841 2.615 ;
      RECT 67.535 2.992 67.555 3.17 ;
      RECT 67.5 2.945 67.535 3.17 ;
      RECT 67.485 2.885 67.5 3.17 ;
      RECT 67.46 2.832 67.485 3.17 ;
      RECT 67.445 2.785 67.46 3.17 ;
      RECT 67.425 2.762 67.445 3.17 ;
      RECT 67.4 2.727 67.425 3.17 ;
      RECT 67.39 2.573 67.4 3.17 ;
      RECT 67.36 2.568 67.39 3.161 ;
      RECT 67.355 2.565 67.36 3.151 ;
      RECT 67.34 2.565 67.355 3.125 ;
      RECT 67.335 2.565 67.34 3.088 ;
      RECT 67.31 2.565 67.335 3.04 ;
      RECT 67.29 2.565 67.31 2.965 ;
      RECT 67.28 2.565 67.29 2.925 ;
      RECT 67.275 2.565 67.28 2.9 ;
      RECT 67.27 2.565 67.275 2.883 ;
      RECT 67.265 2.565 67.27 2.865 ;
      RECT 67.26 2.566 67.265 2.855 ;
      RECT 67.25 2.568 67.26 2.823 ;
      RECT 67.24 2.57 67.25 2.79 ;
      RECT 67.23 2.573 67.24 2.763 ;
      RECT 67.555 3 67.78 3.17 ;
      RECT 66.885 1.812 67.055 2.265 ;
      RECT 66.885 1.812 67.145 2.231 ;
      RECT 66.885 1.812 67.175 2.215 ;
      RECT 66.885 1.812 67.205 2.188 ;
      RECT 67.141 1.79 67.22 2.17 ;
      RECT 66.92 1.797 67.225 2.155 ;
      RECT 66.92 1.805 67.235 2.118 ;
      RECT 66.88 1.832 67.235 2.09 ;
      RECT 66.865 1.845 67.235 2.055 ;
      RECT 66.885 1.82 67.255 2.045 ;
      RECT 66.86 1.885 67.255 2.015 ;
      RECT 66.86 1.915 67.26 1.998 ;
      RECT 66.855 1.945 67.26 1.985 ;
      RECT 66.92 1.794 67.22 2.17 ;
      RECT 67.055 1.791 67.141 2.249 ;
      RECT 67.006 1.792 67.22 2.17 ;
      RECT 67.15 3.452 67.195 3.645 ;
      RECT 67.14 3.422 67.15 3.645 ;
      RECT 67.135 3.407 67.14 3.645 ;
      RECT 67.095 3.317 67.135 3.645 ;
      RECT 67.09 3.23 67.095 3.645 ;
      RECT 67.08 3.2 67.09 3.645 ;
      RECT 67.075 3.16 67.08 3.645 ;
      RECT 67.065 3.122 67.075 3.645 ;
      RECT 67.06 3.087 67.065 3.645 ;
      RECT 67.04 3.04 67.06 3.645 ;
      RECT 67.025 2.965 67.04 3.645 ;
      RECT 67.02 2.92 67.025 3.64 ;
      RECT 67.015 2.9 67.02 3.613 ;
      RECT 67.01 2.88 67.015 3.598 ;
      RECT 67.005 2.855 67.01 3.578 ;
      RECT 67 2.833 67.005 3.563 ;
      RECT 66.995 2.811 67 3.545 ;
      RECT 66.99 2.79 66.995 3.535 ;
      RECT 66.98 2.762 66.99 3.505 ;
      RECT 66.97 2.725 66.98 3.473 ;
      RECT 66.96 2.685 66.97 3.44 ;
      RECT 66.95 2.663 66.96 3.41 ;
      RECT 66.92 2.615 66.95 3.342 ;
      RECT 66.905 2.575 66.92 3.269 ;
      RECT 66.895 2.575 66.905 3.235 ;
      RECT 66.89 2.575 66.895 3.21 ;
      RECT 66.885 2.575 66.89 3.195 ;
      RECT 66.88 2.575 66.885 3.173 ;
      RECT 66.875 2.575 66.88 3.16 ;
      RECT 66.86 2.575 66.875 3.125 ;
      RECT 66.84 2.575 66.86 3.065 ;
      RECT 66.83 2.575 66.84 3.015 ;
      RECT 66.81 2.575 66.83 2.963 ;
      RECT 66.79 2.575 66.81 2.92 ;
      RECT 66.78 2.575 66.79 2.908 ;
      RECT 66.75 2.575 66.78 2.895 ;
      RECT 66.72 2.596 66.75 2.875 ;
      RECT 66.71 2.624 66.72 2.855 ;
      RECT 66.695 2.641 66.71 2.823 ;
      RECT 66.69 2.655 66.695 2.79 ;
      RECT 66.685 2.663 66.69 2.763 ;
      RECT 66.68 2.671 66.685 2.725 ;
      RECT 66.685 3.195 66.69 3.53 ;
      RECT 66.65 3.182 66.685 3.529 ;
      RECT 66.58 3.122 66.65 3.528 ;
      RECT 66.5 3.065 66.58 3.527 ;
      RECT 66.365 3.025 66.5 3.526 ;
      RECT 66.365 3.212 66.7 3.515 ;
      RECT 66.325 3.212 66.7 3.505 ;
      RECT 66.325 3.23 66.705 3.5 ;
      RECT 66.325 3.32 66.71 3.49 ;
      RECT 66.32 3.015 66.485 3.47 ;
      RECT 66.315 3.015 66.485 3.213 ;
      RECT 66.315 3.172 66.68 3.213 ;
      RECT 66.315 3.16 66.675 3.213 ;
      RECT 65.445 5.02 65.615 6.49 ;
      RECT 65.445 6.315 65.62 6.485 ;
      RECT 65.075 1.74 65.245 2.93 ;
      RECT 65.075 1.74 65.545 1.91 ;
      RECT 65.075 6.97 65.545 7.14 ;
      RECT 65.075 5.95 65.245 7.14 ;
      RECT 64.085 1.74 64.255 2.93 ;
      RECT 64.085 1.74 64.555 1.91 ;
      RECT 64.085 6.97 64.555 7.14 ;
      RECT 64.085 5.95 64.255 7.14 ;
      RECT 62.235 2.635 62.405 3.865 ;
      RECT 62.29 0.855 62.46 2.805 ;
      RECT 62.235 0.575 62.405 1.025 ;
      RECT 62.235 7.855 62.405 8.305 ;
      RECT 62.29 6.075 62.46 8.025 ;
      RECT 62.235 5.015 62.405 6.245 ;
      RECT 61.715 0.575 61.885 3.865 ;
      RECT 61.715 2.075 62.12 2.405 ;
      RECT 61.715 1.235 62.12 1.565 ;
      RECT 61.715 5.015 61.885 8.305 ;
      RECT 61.715 7.315 62.12 7.645 ;
      RECT 61.715 6.475 62.12 6.805 ;
      RECT 59.05 1.975 59.78 2.215 ;
      RECT 59.592 1.77 59.78 2.215 ;
      RECT 59.42 1.782 59.795 2.209 ;
      RECT 59.335 1.797 59.815 2.194 ;
      RECT 59.335 1.812 59.82 2.184 ;
      RECT 59.29 1.832 59.835 2.176 ;
      RECT 59.267 1.867 59.85 2.13 ;
      RECT 59.181 1.89 59.855 2.09 ;
      RECT 59.181 1.908 59.865 2.06 ;
      RECT 59.05 1.977 59.87 2.023 ;
      RECT 59.095 1.92 59.865 2.06 ;
      RECT 59.181 1.872 59.85 2.13 ;
      RECT 59.267 1.841 59.835 2.176 ;
      RECT 59.29 1.822 59.82 2.184 ;
      RECT 59.335 1.795 59.795 2.209 ;
      RECT 59.42 1.777 59.78 2.215 ;
      RECT 59.506 1.771 59.78 2.215 ;
      RECT 59.592 1.766 59.725 2.215 ;
      RECT 59.678 1.761 59.725 2.215 ;
      RECT 59.37 2.659 59.54 3.045 ;
      RECT 59.365 2.659 59.54 3.04 ;
      RECT 59.34 2.659 59.54 3.005 ;
      RECT 59.34 2.687 59.55 2.995 ;
      RECT 59.32 2.687 59.55 2.955 ;
      RECT 59.315 2.687 59.55 2.928 ;
      RECT 59.315 2.705 59.555 2.92 ;
      RECT 59.26 2.705 59.555 2.855 ;
      RECT 59.26 2.722 59.565 2.838 ;
      RECT 59.25 2.722 59.565 2.778 ;
      RECT 59.25 2.739 59.57 2.775 ;
      RECT 59.245 2.575 59.415 2.753 ;
      RECT 59.245 2.609 59.501 2.753 ;
      RECT 59.24 3.375 59.245 3.388 ;
      RECT 59.235 3.27 59.24 3.393 ;
      RECT 59.21 3.13 59.235 3.408 ;
      RECT 59.175 3.081 59.21 3.44 ;
      RECT 59.17 3.049 59.175 3.46 ;
      RECT 59.165 3.04 59.17 3.46 ;
      RECT 59.085 3.005 59.165 3.46 ;
      RECT 59.022 2.975 59.085 3.46 ;
      RECT 58.936 2.963 59.022 3.46 ;
      RECT 58.85 2.949 58.936 3.46 ;
      RECT 58.77 2.936 58.85 3.446 ;
      RECT 58.735 2.928 58.77 3.426 ;
      RECT 58.725 2.925 58.735 3.417 ;
      RECT 58.695 2.92 58.725 3.404 ;
      RECT 58.645 2.895 58.695 3.38 ;
      RECT 58.631 2.869 58.645 3.362 ;
      RECT 58.545 2.829 58.631 3.338 ;
      RECT 58.5 2.777 58.545 3.307 ;
      RECT 58.49 2.752 58.5 3.294 ;
      RECT 58.485 2.533 58.49 2.555 ;
      RECT 58.48 2.735 58.49 3.29 ;
      RECT 58.48 2.531 58.485 2.645 ;
      RECT 58.47 2.527 58.48 3.286 ;
      RECT 58.426 2.525 58.47 3.274 ;
      RECT 58.34 2.525 58.426 3.245 ;
      RECT 58.31 2.525 58.34 3.218 ;
      RECT 58.295 2.525 58.31 3.206 ;
      RECT 58.255 2.537 58.295 3.191 ;
      RECT 58.235 2.556 58.255 3.17 ;
      RECT 58.225 2.566 58.235 3.154 ;
      RECT 58.215 2.572 58.225 3.143 ;
      RECT 58.195 2.582 58.215 3.126 ;
      RECT 58.19 2.591 58.195 3.113 ;
      RECT 58.185 2.595 58.19 3.063 ;
      RECT 58.175 2.601 58.185 2.98 ;
      RECT 58.17 2.605 58.175 2.894 ;
      RECT 58.165 2.625 58.17 2.831 ;
      RECT 58.16 2.648 58.165 2.778 ;
      RECT 58.155 2.666 58.16 2.723 ;
      RECT 58.765 2.485 58.935 2.745 ;
      RECT 58.935 2.45 58.98 2.731 ;
      RECT 58.896 2.452 58.985 2.714 ;
      RECT 58.785 2.469 59.071 2.685 ;
      RECT 58.785 2.484 59.075 2.657 ;
      RECT 58.785 2.465 58.985 2.714 ;
      RECT 58.81 2.453 58.935 2.745 ;
      RECT 58.896 2.451 58.98 2.731 ;
      RECT 57.95 1.84 58.12 2.33 ;
      RECT 57.95 1.84 58.155 2.31 ;
      RECT 58.085 1.76 58.195 2.27 ;
      RECT 58.066 1.764 58.215 2.24 ;
      RECT 57.98 1.772 58.235 2.223 ;
      RECT 57.98 1.778 58.24 2.213 ;
      RECT 57.98 1.787 58.26 2.201 ;
      RECT 57.955 1.812 58.29 2.179 ;
      RECT 57.955 1.832 58.295 2.159 ;
      RECT 57.95 1.845 58.305 2.139 ;
      RECT 57.95 1.912 58.31 2.12 ;
      RECT 57.95 2.045 58.315 2.107 ;
      RECT 57.945 1.85 58.305 1.94 ;
      RECT 57.955 1.807 58.26 2.201 ;
      RECT 58.066 1.762 58.195 2.27 ;
      RECT 57.94 3.515 58.24 3.77 ;
      RECT 58.025 3.481 58.24 3.77 ;
      RECT 58.025 3.484 58.245 3.63 ;
      RECT 57.96 3.505 58.245 3.63 ;
      RECT 57.995 3.495 58.24 3.77 ;
      RECT 57.99 3.5 58.245 3.63 ;
      RECT 58.025 3.479 58.226 3.77 ;
      RECT 58.111 3.47 58.226 3.77 ;
      RECT 58.111 3.464 58.14 3.77 ;
      RECT 57.6 3.105 57.61 3.595 ;
      RECT 57.26 3.04 57.27 3.34 ;
      RECT 57.775 3.212 57.78 3.431 ;
      RECT 57.765 3.192 57.775 3.448 ;
      RECT 57.755 3.172 57.765 3.478 ;
      RECT 57.75 3.162 57.755 3.493 ;
      RECT 57.745 3.158 57.75 3.498 ;
      RECT 57.73 3.15 57.745 3.505 ;
      RECT 57.69 3.13 57.73 3.53 ;
      RECT 57.665 3.112 57.69 3.563 ;
      RECT 57.66 3.11 57.665 3.576 ;
      RECT 57.64 3.107 57.66 3.58 ;
      RECT 57.61 3.105 57.64 3.59 ;
      RECT 57.54 3.107 57.6 3.591 ;
      RECT 57.52 3.107 57.54 3.585 ;
      RECT 57.495 3.105 57.52 3.582 ;
      RECT 57.46 3.1 57.495 3.578 ;
      RECT 57.44 3.094 57.46 3.565 ;
      RECT 57.43 3.091 57.44 3.553 ;
      RECT 57.41 3.088 57.43 3.538 ;
      RECT 57.39 3.084 57.41 3.52 ;
      RECT 57.385 3.081 57.39 3.51 ;
      RECT 57.38 3.08 57.385 3.508 ;
      RECT 57.37 3.077 57.38 3.5 ;
      RECT 57.36 3.071 57.37 3.483 ;
      RECT 57.35 3.065 57.36 3.465 ;
      RECT 57.34 3.059 57.35 3.453 ;
      RECT 57.33 3.053 57.34 3.433 ;
      RECT 57.325 3.049 57.33 3.418 ;
      RECT 57.32 3.047 57.325 3.41 ;
      RECT 57.315 3.045 57.32 3.403 ;
      RECT 57.31 3.043 57.315 3.393 ;
      RECT 57.305 3.041 57.31 3.387 ;
      RECT 57.295 3.04 57.305 3.377 ;
      RECT 57.285 3.04 57.295 3.368 ;
      RECT 57.27 3.04 57.285 3.353 ;
      RECT 57.23 3.04 57.26 3.337 ;
      RECT 57.21 3.042 57.23 3.332 ;
      RECT 57.205 3.047 57.21 3.33 ;
      RECT 57.175 3.055 57.205 3.328 ;
      RECT 57.145 3.07 57.175 3.327 ;
      RECT 57.1 3.092 57.145 3.332 ;
      RECT 57.095 3.107 57.1 3.336 ;
      RECT 57.08 3.112 57.095 3.338 ;
      RECT 57.075 3.116 57.08 3.34 ;
      RECT 57.015 3.139 57.075 3.349 ;
      RECT 56.995 3.165 57.015 3.362 ;
      RECT 56.985 3.172 56.995 3.366 ;
      RECT 56.97 3.179 56.985 3.369 ;
      RECT 56.95 3.189 56.97 3.372 ;
      RECT 56.945 3.197 56.95 3.375 ;
      RECT 56.9 3.202 56.945 3.382 ;
      RECT 56.89 3.205 56.9 3.389 ;
      RECT 56.88 3.205 56.89 3.393 ;
      RECT 56.845 3.207 56.88 3.405 ;
      RECT 56.825 3.21 56.845 3.418 ;
      RECT 56.785 3.213 56.825 3.429 ;
      RECT 56.77 3.215 56.785 3.442 ;
      RECT 56.76 3.215 56.77 3.447 ;
      RECT 56.735 3.216 56.76 3.455 ;
      RECT 56.725 3.218 56.735 3.46 ;
      RECT 56.72 3.219 56.725 3.463 ;
      RECT 56.695 3.217 56.72 3.466 ;
      RECT 56.68 3.215 56.695 3.467 ;
      RECT 56.66 3.212 56.68 3.469 ;
      RECT 56.64 3.207 56.66 3.469 ;
      RECT 56.58 3.202 56.64 3.466 ;
      RECT 56.545 3.177 56.58 3.462 ;
      RECT 56.535 3.154 56.545 3.46 ;
      RECT 56.505 3.131 56.535 3.46 ;
      RECT 56.495 3.11 56.505 3.46 ;
      RECT 56.47 3.092 56.495 3.458 ;
      RECT 56.455 3.07 56.47 3.455 ;
      RECT 56.44 3.052 56.455 3.453 ;
      RECT 56.42 3.042 56.44 3.451 ;
      RECT 56.405 3.037 56.42 3.45 ;
      RECT 56.39 3.035 56.405 3.449 ;
      RECT 56.36 3.036 56.39 3.447 ;
      RECT 56.34 3.039 56.36 3.445 ;
      RECT 56.283 3.043 56.34 3.445 ;
      RECT 56.197 3.052 56.283 3.445 ;
      RECT 56.111 3.063 56.197 3.445 ;
      RECT 56.025 3.074 56.111 3.445 ;
      RECT 56.005 3.081 56.025 3.453 ;
      RECT 55.995 3.084 56.005 3.46 ;
      RECT 55.93 3.089 55.995 3.478 ;
      RECT 55.9 3.096 55.93 3.503 ;
      RECT 55.89 3.099 55.9 3.51 ;
      RECT 55.845 3.103 55.89 3.515 ;
      RECT 55.815 3.108 55.845 3.52 ;
      RECT 55.814 3.11 55.815 3.52 ;
      RECT 55.728 3.116 55.814 3.52 ;
      RECT 55.642 3.127 55.728 3.52 ;
      RECT 55.556 3.139 55.642 3.52 ;
      RECT 55.47 3.15 55.556 3.52 ;
      RECT 55.455 3.157 55.47 3.515 ;
      RECT 55.45 3.159 55.455 3.509 ;
      RECT 55.43 3.17 55.45 3.504 ;
      RECT 55.42 3.188 55.43 3.498 ;
      RECT 55.415 3.2 55.42 3.298 ;
      RECT 57.71 1.953 57.73 2.04 ;
      RECT 57.705 1.888 57.71 2.072 ;
      RECT 57.695 1.855 57.705 2.077 ;
      RECT 57.69 1.835 57.695 2.083 ;
      RECT 57.66 1.835 57.69 2.1 ;
      RECT 57.611 1.835 57.66 2.136 ;
      RECT 57.525 1.835 57.611 2.194 ;
      RECT 57.496 1.845 57.525 2.243 ;
      RECT 57.41 1.887 57.496 2.296 ;
      RECT 57.39 1.925 57.41 2.343 ;
      RECT 57.365 1.942 57.39 2.363 ;
      RECT 57.355 1.956 57.365 2.383 ;
      RECT 57.35 1.962 57.355 2.393 ;
      RECT 57.345 1.966 57.35 2.4 ;
      RECT 57.295 1.986 57.345 2.405 ;
      RECT 57.23 2.03 57.295 2.405 ;
      RECT 57.205 2.08 57.23 2.405 ;
      RECT 57.195 2.11 57.205 2.405 ;
      RECT 57.19 2.137 57.195 2.405 ;
      RECT 57.185 2.155 57.19 2.405 ;
      RECT 57.175 2.197 57.185 2.405 ;
      RECT 57.525 2.755 57.695 2.93 ;
      RECT 57.465 2.583 57.525 2.918 ;
      RECT 57.455 2.576 57.465 2.901 ;
      RECT 57.41 2.755 57.695 2.881 ;
      RECT 57.391 2.755 57.695 2.859 ;
      RECT 57.305 2.755 57.695 2.824 ;
      RECT 57.285 2.575 57.455 2.78 ;
      RECT 57.285 2.722 57.69 2.78 ;
      RECT 57.285 2.67 57.665 2.78 ;
      RECT 57.285 2.625 57.63 2.78 ;
      RECT 57.285 2.607 57.595 2.78 ;
      RECT 57.285 2.597 57.59 2.78 ;
      RECT 56.935 5.015 57.105 8.305 ;
      RECT 56.935 7.315 57.34 7.645 ;
      RECT 56.935 6.475 57.34 6.805 ;
      RECT 57.005 3.555 57.195 3.78 ;
      RECT 56.995 3.556 57.2 3.775 ;
      RECT 56.995 3.558 57.21 3.755 ;
      RECT 56.995 3.562 57.215 3.74 ;
      RECT 56.995 3.549 57.165 3.775 ;
      RECT 56.995 3.552 57.19 3.775 ;
      RECT 57.005 3.548 57.165 3.78 ;
      RECT 57.091 3.546 57.165 3.78 ;
      RECT 56.715 2.797 56.885 3.035 ;
      RECT 56.715 2.797 56.971 2.949 ;
      RECT 56.715 2.797 56.975 2.859 ;
      RECT 56.765 2.57 56.985 2.838 ;
      RECT 56.76 2.587 56.99 2.811 ;
      RECT 56.725 2.745 56.99 2.811 ;
      RECT 56.745 2.595 56.885 3.035 ;
      RECT 56.735 2.677 56.995 2.794 ;
      RECT 56.73 2.725 56.995 2.794 ;
      RECT 56.735 2.635 56.99 2.811 ;
      RECT 56.76 2.572 56.985 2.838 ;
      RECT 56.325 2.547 56.495 2.745 ;
      RECT 56.325 2.547 56.54 2.72 ;
      RECT 56.395 2.49 56.565 2.678 ;
      RECT 56.37 2.505 56.565 2.678 ;
      RECT 55.985 2.551 56.015 2.745 ;
      RECT 55.98 2.523 55.985 2.745 ;
      RECT 55.95 2.497 55.98 2.747 ;
      RECT 55.925 2.455 55.95 2.75 ;
      RECT 55.915 2.427 55.925 2.752 ;
      RECT 55.88 2.407 55.915 2.754 ;
      RECT 55.815 2.392 55.88 2.76 ;
      RECT 55.765 2.39 55.815 2.766 ;
      RECT 55.742 2.392 55.765 2.771 ;
      RECT 55.656 2.403 55.742 2.777 ;
      RECT 55.57 2.421 55.656 2.787 ;
      RECT 55.555 2.432 55.57 2.793 ;
      RECT 55.485 2.455 55.555 2.799 ;
      RECT 55.43 2.487 55.485 2.807 ;
      RECT 55.39 2.51 55.43 2.813 ;
      RECT 55.376 2.523 55.39 2.816 ;
      RECT 55.29 2.545 55.376 2.822 ;
      RECT 55.275 2.57 55.29 2.828 ;
      RECT 55.235 2.585 55.275 2.832 ;
      RECT 55.185 2.6 55.235 2.837 ;
      RECT 55.16 2.607 55.185 2.841 ;
      RECT 55.1 2.602 55.16 2.845 ;
      RECT 55.085 2.593 55.1 2.849 ;
      RECT 55.015 2.583 55.085 2.845 ;
      RECT 54.99 2.575 55.01 2.835 ;
      RECT 54.931 2.575 54.99 2.813 ;
      RECT 54.845 2.575 54.931 2.77 ;
      RECT 55.01 2.575 55.015 2.84 ;
      RECT 55.705 1.806 55.875 2.14 ;
      RECT 55.675 1.806 55.875 2.135 ;
      RECT 55.615 1.773 55.675 2.123 ;
      RECT 55.615 1.829 55.885 2.118 ;
      RECT 55.59 1.829 55.885 2.112 ;
      RECT 55.585 1.77 55.615 2.109 ;
      RECT 55.57 1.776 55.705 2.107 ;
      RECT 55.565 1.784 55.79 2.095 ;
      RECT 55.565 1.836 55.9 2.048 ;
      RECT 55.55 1.792 55.79 2.043 ;
      RECT 55.55 1.862 55.91 1.984 ;
      RECT 55.52 1.812 55.875 1.945 ;
      RECT 55.52 1.902 55.92 1.941 ;
      RECT 55.57 1.781 55.79 2.107 ;
      RECT 54.91 2.111 54.965 2.375 ;
      RECT 54.91 2.111 55.03 2.374 ;
      RECT 54.91 2.111 55.055 2.373 ;
      RECT 54.91 2.111 55.12 2.372 ;
      RECT 55.055 2.077 55.135 2.371 ;
      RECT 54.87 2.121 55.28 2.37 ;
      RECT 54.91 2.118 55.28 2.37 ;
      RECT 54.87 2.126 55.285 2.363 ;
      RECT 54.855 2.128 55.285 2.362 ;
      RECT 54.855 2.135 55.29 2.358 ;
      RECT 54.835 2.134 55.285 2.354 ;
      RECT 54.835 2.142 55.295 2.353 ;
      RECT 54.83 2.139 55.29 2.349 ;
      RECT 54.83 2.152 55.305 2.348 ;
      RECT 54.815 2.142 55.295 2.347 ;
      RECT 54.78 2.155 55.305 2.34 ;
      RECT 54.965 2.11 55.275 2.37 ;
      RECT 54.965 2.095 55.225 2.37 ;
      RECT 55.03 2.082 55.16 2.37 ;
      RECT 54.575 3.171 54.59 3.564 ;
      RECT 54.54 3.176 54.59 3.563 ;
      RECT 54.575 3.175 54.635 3.562 ;
      RECT 54.52 3.186 54.635 3.561 ;
      RECT 54.535 3.182 54.635 3.561 ;
      RECT 54.5 3.192 54.71 3.558 ;
      RECT 54.5 3.211 54.755 3.556 ;
      RECT 54.5 3.218 54.76 3.553 ;
      RECT 54.485 3.195 54.71 3.55 ;
      RECT 54.465 3.2 54.71 3.543 ;
      RECT 54.46 3.204 54.71 3.539 ;
      RECT 54.46 3.221 54.77 3.538 ;
      RECT 54.44 3.215 54.755 3.534 ;
      RECT 54.44 3.224 54.775 3.528 ;
      RECT 54.435 3.23 54.775 3.3 ;
      RECT 54.5 3.19 54.635 3.558 ;
      RECT 54.375 2.553 54.575 2.865 ;
      RECT 54.45 2.531 54.575 2.865 ;
      RECT 54.39 2.55 54.58 2.85 ;
      RECT 54.36 2.561 54.58 2.848 ;
      RECT 54.375 2.556 54.585 2.814 ;
      RECT 54.36 2.66 54.59 2.781 ;
      RECT 54.39 2.532 54.575 2.865 ;
      RECT 54.45 2.51 54.55 2.865 ;
      RECT 54.475 2.507 54.55 2.865 ;
      RECT 54.475 2.502 54.495 2.865 ;
      RECT 53.88 2.57 54.055 2.745 ;
      RECT 53.875 2.57 54.055 2.743 ;
      RECT 53.85 2.57 54.055 2.738 ;
      RECT 53.795 2.55 53.965 2.728 ;
      RECT 53.795 2.557 54.03 2.728 ;
      RECT 53.88 3.237 53.895 3.42 ;
      RECT 53.87 3.215 53.88 3.42 ;
      RECT 53.855 3.195 53.87 3.42 ;
      RECT 53.845 3.17 53.855 3.42 ;
      RECT 53.815 3.135 53.845 3.42 ;
      RECT 53.78 3.075 53.815 3.42 ;
      RECT 53.775 3.037 53.78 3.42 ;
      RECT 53.725 2.988 53.775 3.42 ;
      RECT 53.715 2.938 53.725 3.408 ;
      RECT 53.7 2.917 53.715 3.368 ;
      RECT 53.68 2.885 53.7 3.318 ;
      RECT 53.655 2.841 53.68 3.258 ;
      RECT 53.65 2.813 53.655 3.213 ;
      RECT 53.645 2.804 53.65 3.199 ;
      RECT 53.64 2.797 53.645 3.186 ;
      RECT 53.635 2.792 53.64 3.175 ;
      RECT 53.63 2.777 53.635 3.165 ;
      RECT 53.625 2.755 53.63 3.152 ;
      RECT 53.615 2.715 53.625 3.127 ;
      RECT 53.59 2.645 53.615 3.083 ;
      RECT 53.585 2.585 53.59 3.048 ;
      RECT 53.57 2.565 53.585 3.015 ;
      RECT 53.565 2.565 53.57 2.99 ;
      RECT 53.535 2.565 53.565 2.945 ;
      RECT 53.49 2.565 53.535 2.885 ;
      RECT 53.415 2.565 53.49 2.833 ;
      RECT 53.41 2.565 53.415 2.798 ;
      RECT 53.405 2.565 53.41 2.788 ;
      RECT 53.4 2.565 53.405 2.768 ;
      RECT 53.665 1.785 53.835 2.255 ;
      RECT 53.61 1.778 53.805 2.239 ;
      RECT 53.61 1.792 53.84 2.238 ;
      RECT 53.595 1.793 53.84 2.219 ;
      RECT 53.59 1.811 53.84 2.205 ;
      RECT 53.595 1.794 53.845 2.203 ;
      RECT 53.58 1.825 53.845 2.188 ;
      RECT 53.595 1.8 53.85 2.173 ;
      RECT 53.575 1.84 53.85 2.17 ;
      RECT 53.59 1.812 53.855 2.155 ;
      RECT 53.59 1.824 53.86 2.135 ;
      RECT 53.575 1.84 53.865 2.118 ;
      RECT 53.575 1.85 53.87 1.973 ;
      RECT 53.57 1.85 53.87 1.93 ;
      RECT 53.57 1.865 53.875 1.908 ;
      RECT 53.665 1.775 53.805 2.255 ;
      RECT 53.665 1.773 53.775 2.255 ;
      RECT 53.751 1.77 53.775 2.255 ;
      RECT 53.41 3.437 53.415 3.483 ;
      RECT 53.4 3.285 53.41 3.507 ;
      RECT 53.395 3.13 53.4 3.532 ;
      RECT 53.38 3.092 53.395 3.543 ;
      RECT 53.375 3.075 53.38 3.55 ;
      RECT 53.365 3.063 53.375 3.557 ;
      RECT 53.36 3.054 53.365 3.559 ;
      RECT 53.355 3.052 53.36 3.563 ;
      RECT 53.31 3.043 53.355 3.578 ;
      RECT 53.305 3.035 53.31 3.592 ;
      RECT 53.3 3.032 53.305 3.596 ;
      RECT 53.285 3.027 53.3 3.604 ;
      RECT 53.23 3.017 53.285 3.615 ;
      RECT 53.195 3.005 53.23 3.616 ;
      RECT 53.186 3 53.195 3.61 ;
      RECT 53.1 3 53.186 3.6 ;
      RECT 53.07 3 53.1 3.578 ;
      RECT 53.06 3 53.065 3.558 ;
      RECT 53.055 3 53.06 3.52 ;
      RECT 53.05 3 53.055 3.478 ;
      RECT 53.045 3 53.05 3.438 ;
      RECT 53.04 3 53.045 3.368 ;
      RECT 53.03 3 53.04 3.29 ;
      RECT 53.025 3 53.03 3.19 ;
      RECT 53.065 3 53.07 3.56 ;
      RECT 52.56 3.082 52.65 3.56 ;
      RECT 52.545 3.085 52.665 3.558 ;
      RECT 52.56 3.084 52.665 3.558 ;
      RECT 52.525 3.091 52.69 3.548 ;
      RECT 52.545 3.085 52.69 3.548 ;
      RECT 52.51 3.097 52.69 3.536 ;
      RECT 52.545 3.088 52.74 3.529 ;
      RECT 52.496 3.105 52.74 3.527 ;
      RECT 52.525 3.095 52.75 3.515 ;
      RECT 52.496 3.116 52.78 3.506 ;
      RECT 52.41 3.14 52.78 3.5 ;
      RECT 52.41 3.153 52.82 3.483 ;
      RECT 52.405 3.175 52.82 3.476 ;
      RECT 52.375 3.19 52.82 3.466 ;
      RECT 52.37 3.201 52.82 3.456 ;
      RECT 52.34 3.214 52.82 3.447 ;
      RECT 52.325 3.232 52.82 3.436 ;
      RECT 52.3 3.245 52.82 3.426 ;
      RECT 52.56 3.081 52.57 3.56 ;
      RECT 52.606 2.505 52.645 2.75 ;
      RECT 52.52 2.505 52.655 2.748 ;
      RECT 52.405 2.53 52.655 2.745 ;
      RECT 52.405 2.53 52.66 2.743 ;
      RECT 52.405 2.53 52.675 2.738 ;
      RECT 52.511 2.505 52.69 2.718 ;
      RECT 52.425 2.513 52.69 2.718 ;
      RECT 52.095 1.865 52.265 2.3 ;
      RECT 52.085 1.899 52.265 2.283 ;
      RECT 52.165 1.835 52.335 2.27 ;
      RECT 52.07 1.91 52.335 2.248 ;
      RECT 52.165 1.845 52.34 2.238 ;
      RECT 52.095 1.897 52.37 2.223 ;
      RECT 52.055 1.923 52.37 2.208 ;
      RECT 52.055 1.965 52.38 2.188 ;
      RECT 52.05 1.99 52.385 2.17 ;
      RECT 52.05 2 52.39 2.155 ;
      RECT 52.045 1.937 52.37 2.153 ;
      RECT 52.045 2.01 52.395 2.138 ;
      RECT 52.04 1.947 52.37 2.135 ;
      RECT 52.035 2.031 52.4 2.118 ;
      RECT 52.035 2.063 52.405 2.098 ;
      RECT 52.03 1.977 52.38 2.09 ;
      RECT 52.035 1.962 52.37 2.118 ;
      RECT 52.05 1.932 52.37 2.17 ;
      RECT 51.895 2.519 52.12 2.775 ;
      RECT 51.895 2.552 52.14 2.765 ;
      RECT 51.86 2.552 52.14 2.763 ;
      RECT 51.86 2.565 52.145 2.753 ;
      RECT 51.86 2.585 52.155 2.745 ;
      RECT 51.86 2.682 52.16 2.738 ;
      RECT 51.84 2.43 51.97 2.728 ;
      RECT 51.795 2.585 52.155 2.67 ;
      RECT 51.785 2.43 51.97 2.615 ;
      RECT 51.785 2.462 52.056 2.615 ;
      RECT 51.75 2.992 51.77 3.17 ;
      RECT 51.715 2.945 51.75 3.17 ;
      RECT 51.7 2.885 51.715 3.17 ;
      RECT 51.675 2.832 51.7 3.17 ;
      RECT 51.66 2.785 51.675 3.17 ;
      RECT 51.64 2.762 51.66 3.17 ;
      RECT 51.615 2.727 51.64 3.17 ;
      RECT 51.605 2.573 51.615 3.17 ;
      RECT 51.575 2.568 51.605 3.161 ;
      RECT 51.57 2.565 51.575 3.151 ;
      RECT 51.555 2.565 51.57 3.125 ;
      RECT 51.55 2.565 51.555 3.088 ;
      RECT 51.525 2.565 51.55 3.04 ;
      RECT 51.505 2.565 51.525 2.965 ;
      RECT 51.495 2.565 51.505 2.925 ;
      RECT 51.49 2.565 51.495 2.9 ;
      RECT 51.485 2.565 51.49 2.883 ;
      RECT 51.48 2.565 51.485 2.865 ;
      RECT 51.475 2.566 51.48 2.855 ;
      RECT 51.465 2.568 51.475 2.823 ;
      RECT 51.455 2.57 51.465 2.79 ;
      RECT 51.445 2.573 51.455 2.763 ;
      RECT 51.77 3 51.995 3.17 ;
      RECT 51.1 1.812 51.27 2.265 ;
      RECT 51.1 1.812 51.36 2.231 ;
      RECT 51.1 1.812 51.39 2.215 ;
      RECT 51.1 1.812 51.42 2.188 ;
      RECT 51.356 1.79 51.435 2.17 ;
      RECT 51.135 1.797 51.44 2.155 ;
      RECT 51.135 1.805 51.45 2.118 ;
      RECT 51.095 1.832 51.45 2.09 ;
      RECT 51.08 1.845 51.45 2.055 ;
      RECT 51.1 1.82 51.47 2.045 ;
      RECT 51.075 1.885 51.47 2.015 ;
      RECT 51.075 1.915 51.475 1.998 ;
      RECT 51.07 1.945 51.475 1.985 ;
      RECT 51.135 1.794 51.435 2.17 ;
      RECT 51.27 1.791 51.356 2.249 ;
      RECT 51.221 1.792 51.435 2.17 ;
      RECT 51.365 3.452 51.41 3.645 ;
      RECT 51.355 3.422 51.365 3.645 ;
      RECT 51.35 3.407 51.355 3.645 ;
      RECT 51.31 3.317 51.35 3.645 ;
      RECT 51.305 3.23 51.31 3.645 ;
      RECT 51.295 3.2 51.305 3.645 ;
      RECT 51.29 3.16 51.295 3.645 ;
      RECT 51.28 3.122 51.29 3.645 ;
      RECT 51.275 3.087 51.28 3.645 ;
      RECT 51.255 3.04 51.275 3.645 ;
      RECT 51.24 2.965 51.255 3.645 ;
      RECT 51.235 2.92 51.24 3.64 ;
      RECT 51.23 2.9 51.235 3.613 ;
      RECT 51.225 2.88 51.23 3.598 ;
      RECT 51.22 2.855 51.225 3.578 ;
      RECT 51.215 2.833 51.22 3.563 ;
      RECT 51.21 2.811 51.215 3.545 ;
      RECT 51.205 2.79 51.21 3.535 ;
      RECT 51.195 2.762 51.205 3.505 ;
      RECT 51.185 2.725 51.195 3.473 ;
      RECT 51.175 2.685 51.185 3.44 ;
      RECT 51.165 2.663 51.175 3.41 ;
      RECT 51.135 2.615 51.165 3.342 ;
      RECT 51.12 2.575 51.135 3.269 ;
      RECT 51.11 2.575 51.12 3.235 ;
      RECT 51.105 2.575 51.11 3.21 ;
      RECT 51.1 2.575 51.105 3.195 ;
      RECT 51.095 2.575 51.1 3.173 ;
      RECT 51.09 2.575 51.095 3.16 ;
      RECT 51.075 2.575 51.09 3.125 ;
      RECT 51.055 2.575 51.075 3.065 ;
      RECT 51.045 2.575 51.055 3.015 ;
      RECT 51.025 2.575 51.045 2.963 ;
      RECT 51.005 2.575 51.025 2.92 ;
      RECT 50.995 2.575 51.005 2.908 ;
      RECT 50.965 2.575 50.995 2.895 ;
      RECT 50.935 2.596 50.965 2.875 ;
      RECT 50.925 2.624 50.935 2.855 ;
      RECT 50.91 2.641 50.925 2.823 ;
      RECT 50.905 2.655 50.91 2.79 ;
      RECT 50.9 2.663 50.905 2.763 ;
      RECT 50.895 2.671 50.9 2.725 ;
      RECT 50.9 3.195 50.905 3.53 ;
      RECT 50.865 3.182 50.9 3.529 ;
      RECT 50.795 3.122 50.865 3.528 ;
      RECT 50.715 3.065 50.795 3.527 ;
      RECT 50.58 3.025 50.715 3.526 ;
      RECT 50.58 3.212 50.915 3.515 ;
      RECT 50.54 3.212 50.915 3.505 ;
      RECT 50.54 3.23 50.92 3.5 ;
      RECT 50.54 3.32 50.925 3.49 ;
      RECT 50.535 3.015 50.7 3.47 ;
      RECT 50.53 3.015 50.7 3.213 ;
      RECT 50.53 3.172 50.895 3.213 ;
      RECT 50.53 3.16 50.89 3.213 ;
      RECT 49.66 5.02 49.83 6.49 ;
      RECT 49.66 6.315 49.835 6.485 ;
      RECT 49.29 1.74 49.46 2.93 ;
      RECT 49.29 1.74 49.76 1.91 ;
      RECT 49.29 6.97 49.76 7.14 ;
      RECT 49.29 5.95 49.46 7.14 ;
      RECT 48.3 1.74 48.47 2.93 ;
      RECT 48.3 1.74 48.77 1.91 ;
      RECT 48.3 6.97 48.77 7.14 ;
      RECT 48.3 5.95 48.47 7.14 ;
      RECT 46.45 2.635 46.62 3.865 ;
      RECT 46.505 0.855 46.675 2.805 ;
      RECT 46.45 0.575 46.62 1.025 ;
      RECT 46.45 7.855 46.62 8.305 ;
      RECT 46.505 6.075 46.675 8.025 ;
      RECT 46.45 5.015 46.62 6.245 ;
      RECT 45.93 0.575 46.1 3.865 ;
      RECT 45.93 2.075 46.335 2.405 ;
      RECT 45.93 1.235 46.335 1.565 ;
      RECT 45.93 5.015 46.1 8.305 ;
      RECT 45.93 7.315 46.335 7.645 ;
      RECT 45.93 6.475 46.335 6.805 ;
      RECT 43.265 1.975 43.995 2.215 ;
      RECT 43.807 1.77 43.995 2.215 ;
      RECT 43.635 1.782 44.01 2.209 ;
      RECT 43.55 1.797 44.03 2.194 ;
      RECT 43.55 1.812 44.035 2.184 ;
      RECT 43.505 1.832 44.05 2.176 ;
      RECT 43.482 1.867 44.065 2.13 ;
      RECT 43.396 1.89 44.07 2.09 ;
      RECT 43.396 1.908 44.08 2.06 ;
      RECT 43.265 1.977 44.085 2.023 ;
      RECT 43.31 1.92 44.08 2.06 ;
      RECT 43.396 1.872 44.065 2.13 ;
      RECT 43.482 1.841 44.05 2.176 ;
      RECT 43.505 1.822 44.035 2.184 ;
      RECT 43.55 1.795 44.01 2.209 ;
      RECT 43.635 1.777 43.995 2.215 ;
      RECT 43.721 1.771 43.995 2.215 ;
      RECT 43.807 1.766 43.94 2.215 ;
      RECT 43.893 1.761 43.94 2.215 ;
      RECT 43.585 2.659 43.755 3.045 ;
      RECT 43.58 2.659 43.755 3.04 ;
      RECT 43.555 2.659 43.755 3.005 ;
      RECT 43.555 2.687 43.765 2.995 ;
      RECT 43.535 2.687 43.765 2.955 ;
      RECT 43.53 2.687 43.765 2.928 ;
      RECT 43.53 2.705 43.77 2.92 ;
      RECT 43.475 2.705 43.77 2.855 ;
      RECT 43.475 2.722 43.78 2.838 ;
      RECT 43.465 2.722 43.78 2.778 ;
      RECT 43.465 2.739 43.785 2.775 ;
      RECT 43.46 2.575 43.63 2.753 ;
      RECT 43.46 2.609 43.716 2.753 ;
      RECT 43.455 3.375 43.46 3.388 ;
      RECT 43.45 3.27 43.455 3.393 ;
      RECT 43.425 3.13 43.45 3.408 ;
      RECT 43.39 3.081 43.425 3.44 ;
      RECT 43.385 3.049 43.39 3.46 ;
      RECT 43.38 3.04 43.385 3.46 ;
      RECT 43.3 3.005 43.38 3.46 ;
      RECT 43.237 2.975 43.3 3.46 ;
      RECT 43.151 2.963 43.237 3.46 ;
      RECT 43.065 2.949 43.151 3.46 ;
      RECT 42.985 2.936 43.065 3.446 ;
      RECT 42.95 2.928 42.985 3.426 ;
      RECT 42.94 2.925 42.95 3.417 ;
      RECT 42.91 2.92 42.94 3.404 ;
      RECT 42.86 2.895 42.91 3.38 ;
      RECT 42.846 2.869 42.86 3.362 ;
      RECT 42.76 2.829 42.846 3.338 ;
      RECT 42.715 2.777 42.76 3.307 ;
      RECT 42.705 2.752 42.715 3.294 ;
      RECT 42.7 2.533 42.705 2.555 ;
      RECT 42.695 2.735 42.705 3.29 ;
      RECT 42.695 2.531 42.7 2.645 ;
      RECT 42.685 2.527 42.695 3.286 ;
      RECT 42.641 2.525 42.685 3.274 ;
      RECT 42.555 2.525 42.641 3.245 ;
      RECT 42.525 2.525 42.555 3.218 ;
      RECT 42.51 2.525 42.525 3.206 ;
      RECT 42.47 2.537 42.51 3.191 ;
      RECT 42.45 2.556 42.47 3.17 ;
      RECT 42.44 2.566 42.45 3.154 ;
      RECT 42.43 2.572 42.44 3.143 ;
      RECT 42.41 2.582 42.43 3.126 ;
      RECT 42.405 2.591 42.41 3.113 ;
      RECT 42.4 2.595 42.405 3.063 ;
      RECT 42.39 2.601 42.4 2.98 ;
      RECT 42.385 2.605 42.39 2.894 ;
      RECT 42.38 2.625 42.385 2.831 ;
      RECT 42.375 2.648 42.38 2.778 ;
      RECT 42.37 2.666 42.375 2.723 ;
      RECT 42.98 2.485 43.15 2.745 ;
      RECT 43.15 2.45 43.195 2.731 ;
      RECT 43.111 2.452 43.2 2.714 ;
      RECT 43 2.469 43.286 2.685 ;
      RECT 43 2.484 43.29 2.657 ;
      RECT 43 2.465 43.2 2.714 ;
      RECT 43.025 2.453 43.15 2.745 ;
      RECT 43.111 2.451 43.195 2.731 ;
      RECT 42.165 1.84 42.335 2.33 ;
      RECT 42.165 1.84 42.37 2.31 ;
      RECT 42.3 1.76 42.41 2.27 ;
      RECT 42.281 1.764 42.43 2.24 ;
      RECT 42.195 1.772 42.45 2.223 ;
      RECT 42.195 1.778 42.455 2.213 ;
      RECT 42.195 1.787 42.475 2.201 ;
      RECT 42.17 1.812 42.505 2.179 ;
      RECT 42.17 1.832 42.51 2.159 ;
      RECT 42.165 1.845 42.52 2.139 ;
      RECT 42.165 1.912 42.525 2.12 ;
      RECT 42.165 2.045 42.53 2.107 ;
      RECT 42.16 1.85 42.52 1.94 ;
      RECT 42.17 1.807 42.475 2.201 ;
      RECT 42.281 1.762 42.41 2.27 ;
      RECT 42.155 3.515 42.455 3.77 ;
      RECT 42.24 3.481 42.455 3.77 ;
      RECT 42.24 3.484 42.46 3.63 ;
      RECT 42.175 3.505 42.46 3.63 ;
      RECT 42.21 3.495 42.455 3.77 ;
      RECT 42.205 3.5 42.46 3.63 ;
      RECT 42.24 3.479 42.441 3.77 ;
      RECT 42.326 3.47 42.441 3.77 ;
      RECT 42.326 3.464 42.355 3.77 ;
      RECT 41.815 3.105 41.825 3.595 ;
      RECT 41.475 3.04 41.485 3.34 ;
      RECT 41.99 3.212 41.995 3.431 ;
      RECT 41.98 3.192 41.99 3.448 ;
      RECT 41.97 3.172 41.98 3.478 ;
      RECT 41.965 3.162 41.97 3.493 ;
      RECT 41.96 3.158 41.965 3.498 ;
      RECT 41.945 3.15 41.96 3.505 ;
      RECT 41.905 3.13 41.945 3.53 ;
      RECT 41.88 3.112 41.905 3.563 ;
      RECT 41.875 3.11 41.88 3.576 ;
      RECT 41.855 3.107 41.875 3.58 ;
      RECT 41.825 3.105 41.855 3.59 ;
      RECT 41.755 3.107 41.815 3.591 ;
      RECT 41.735 3.107 41.755 3.585 ;
      RECT 41.71 3.105 41.735 3.582 ;
      RECT 41.675 3.1 41.71 3.578 ;
      RECT 41.655 3.094 41.675 3.565 ;
      RECT 41.645 3.091 41.655 3.553 ;
      RECT 41.625 3.088 41.645 3.538 ;
      RECT 41.605 3.084 41.625 3.52 ;
      RECT 41.6 3.081 41.605 3.51 ;
      RECT 41.595 3.08 41.6 3.508 ;
      RECT 41.585 3.077 41.595 3.5 ;
      RECT 41.575 3.071 41.585 3.483 ;
      RECT 41.565 3.065 41.575 3.465 ;
      RECT 41.555 3.059 41.565 3.453 ;
      RECT 41.545 3.053 41.555 3.433 ;
      RECT 41.54 3.049 41.545 3.418 ;
      RECT 41.535 3.047 41.54 3.41 ;
      RECT 41.53 3.045 41.535 3.403 ;
      RECT 41.525 3.043 41.53 3.393 ;
      RECT 41.52 3.041 41.525 3.387 ;
      RECT 41.51 3.04 41.52 3.377 ;
      RECT 41.5 3.04 41.51 3.368 ;
      RECT 41.485 3.04 41.5 3.353 ;
      RECT 41.445 3.04 41.475 3.337 ;
      RECT 41.425 3.042 41.445 3.332 ;
      RECT 41.42 3.047 41.425 3.33 ;
      RECT 41.39 3.055 41.42 3.328 ;
      RECT 41.36 3.07 41.39 3.327 ;
      RECT 41.315 3.092 41.36 3.332 ;
      RECT 41.31 3.107 41.315 3.336 ;
      RECT 41.295 3.112 41.31 3.338 ;
      RECT 41.29 3.116 41.295 3.34 ;
      RECT 41.23 3.139 41.29 3.349 ;
      RECT 41.21 3.165 41.23 3.362 ;
      RECT 41.2 3.172 41.21 3.366 ;
      RECT 41.185 3.179 41.2 3.369 ;
      RECT 41.165 3.189 41.185 3.372 ;
      RECT 41.16 3.197 41.165 3.375 ;
      RECT 41.115 3.202 41.16 3.382 ;
      RECT 41.105 3.205 41.115 3.389 ;
      RECT 41.095 3.205 41.105 3.393 ;
      RECT 41.06 3.207 41.095 3.405 ;
      RECT 41.04 3.21 41.06 3.418 ;
      RECT 41 3.213 41.04 3.429 ;
      RECT 40.985 3.215 41 3.442 ;
      RECT 40.975 3.215 40.985 3.447 ;
      RECT 40.95 3.216 40.975 3.455 ;
      RECT 40.94 3.218 40.95 3.46 ;
      RECT 40.935 3.219 40.94 3.463 ;
      RECT 40.91 3.217 40.935 3.466 ;
      RECT 40.895 3.215 40.91 3.467 ;
      RECT 40.875 3.212 40.895 3.469 ;
      RECT 40.855 3.207 40.875 3.469 ;
      RECT 40.795 3.202 40.855 3.466 ;
      RECT 40.76 3.177 40.795 3.462 ;
      RECT 40.75 3.154 40.76 3.46 ;
      RECT 40.72 3.131 40.75 3.46 ;
      RECT 40.71 3.11 40.72 3.46 ;
      RECT 40.685 3.092 40.71 3.458 ;
      RECT 40.67 3.07 40.685 3.455 ;
      RECT 40.655 3.052 40.67 3.453 ;
      RECT 40.635 3.042 40.655 3.451 ;
      RECT 40.62 3.037 40.635 3.45 ;
      RECT 40.605 3.035 40.62 3.449 ;
      RECT 40.575 3.036 40.605 3.447 ;
      RECT 40.555 3.039 40.575 3.445 ;
      RECT 40.498 3.043 40.555 3.445 ;
      RECT 40.412 3.052 40.498 3.445 ;
      RECT 40.326 3.063 40.412 3.445 ;
      RECT 40.24 3.074 40.326 3.445 ;
      RECT 40.22 3.081 40.24 3.453 ;
      RECT 40.21 3.084 40.22 3.46 ;
      RECT 40.145 3.089 40.21 3.478 ;
      RECT 40.115 3.096 40.145 3.503 ;
      RECT 40.105 3.099 40.115 3.51 ;
      RECT 40.06 3.103 40.105 3.515 ;
      RECT 40.03 3.108 40.06 3.52 ;
      RECT 40.029 3.11 40.03 3.52 ;
      RECT 39.943 3.116 40.029 3.52 ;
      RECT 39.857 3.127 39.943 3.52 ;
      RECT 39.771 3.139 39.857 3.52 ;
      RECT 39.685 3.15 39.771 3.52 ;
      RECT 39.67 3.157 39.685 3.515 ;
      RECT 39.665 3.159 39.67 3.509 ;
      RECT 39.645 3.17 39.665 3.504 ;
      RECT 39.635 3.188 39.645 3.498 ;
      RECT 39.63 3.2 39.635 3.298 ;
      RECT 41.925 1.953 41.945 2.04 ;
      RECT 41.92 1.888 41.925 2.072 ;
      RECT 41.91 1.855 41.92 2.077 ;
      RECT 41.905 1.835 41.91 2.083 ;
      RECT 41.875 1.835 41.905 2.1 ;
      RECT 41.826 1.835 41.875 2.136 ;
      RECT 41.74 1.835 41.826 2.194 ;
      RECT 41.711 1.845 41.74 2.243 ;
      RECT 41.625 1.887 41.711 2.296 ;
      RECT 41.605 1.925 41.625 2.343 ;
      RECT 41.58 1.942 41.605 2.363 ;
      RECT 41.57 1.956 41.58 2.383 ;
      RECT 41.565 1.962 41.57 2.393 ;
      RECT 41.56 1.966 41.565 2.4 ;
      RECT 41.51 1.986 41.56 2.405 ;
      RECT 41.445 2.03 41.51 2.405 ;
      RECT 41.42 2.08 41.445 2.405 ;
      RECT 41.41 2.11 41.42 2.405 ;
      RECT 41.405 2.137 41.41 2.405 ;
      RECT 41.4 2.155 41.405 2.405 ;
      RECT 41.39 2.197 41.4 2.405 ;
      RECT 41.74 2.755 41.91 2.93 ;
      RECT 41.68 2.583 41.74 2.918 ;
      RECT 41.67 2.576 41.68 2.901 ;
      RECT 41.625 2.755 41.91 2.881 ;
      RECT 41.606 2.755 41.91 2.859 ;
      RECT 41.52 2.755 41.91 2.824 ;
      RECT 41.5 2.575 41.67 2.78 ;
      RECT 41.5 2.722 41.905 2.78 ;
      RECT 41.5 2.67 41.88 2.78 ;
      RECT 41.5 2.625 41.845 2.78 ;
      RECT 41.5 2.607 41.81 2.78 ;
      RECT 41.5 2.597 41.805 2.78 ;
      RECT 41.15 5.015 41.32 8.305 ;
      RECT 41.15 7.315 41.555 7.645 ;
      RECT 41.15 6.475 41.555 6.805 ;
      RECT 41.22 3.555 41.41 3.78 ;
      RECT 41.21 3.556 41.415 3.775 ;
      RECT 41.21 3.558 41.425 3.755 ;
      RECT 41.21 3.562 41.43 3.74 ;
      RECT 41.21 3.549 41.38 3.775 ;
      RECT 41.21 3.552 41.405 3.775 ;
      RECT 41.22 3.548 41.38 3.78 ;
      RECT 41.306 3.546 41.38 3.78 ;
      RECT 40.93 2.797 41.1 3.035 ;
      RECT 40.93 2.797 41.186 2.949 ;
      RECT 40.93 2.797 41.19 2.859 ;
      RECT 40.98 2.57 41.2 2.838 ;
      RECT 40.975 2.587 41.205 2.811 ;
      RECT 40.94 2.745 41.205 2.811 ;
      RECT 40.96 2.595 41.1 3.035 ;
      RECT 40.95 2.677 41.21 2.794 ;
      RECT 40.945 2.725 41.21 2.794 ;
      RECT 40.95 2.635 41.205 2.811 ;
      RECT 40.975 2.572 41.2 2.838 ;
      RECT 40.54 2.547 40.71 2.745 ;
      RECT 40.54 2.547 40.755 2.72 ;
      RECT 40.61 2.49 40.78 2.678 ;
      RECT 40.585 2.505 40.78 2.678 ;
      RECT 40.2 2.551 40.23 2.745 ;
      RECT 40.195 2.523 40.2 2.745 ;
      RECT 40.165 2.497 40.195 2.747 ;
      RECT 40.14 2.455 40.165 2.75 ;
      RECT 40.13 2.427 40.14 2.752 ;
      RECT 40.095 2.407 40.13 2.754 ;
      RECT 40.03 2.392 40.095 2.76 ;
      RECT 39.98 2.39 40.03 2.766 ;
      RECT 39.957 2.392 39.98 2.771 ;
      RECT 39.871 2.403 39.957 2.777 ;
      RECT 39.785 2.421 39.871 2.787 ;
      RECT 39.77 2.432 39.785 2.793 ;
      RECT 39.7 2.455 39.77 2.799 ;
      RECT 39.645 2.487 39.7 2.807 ;
      RECT 39.605 2.51 39.645 2.813 ;
      RECT 39.591 2.523 39.605 2.816 ;
      RECT 39.505 2.545 39.591 2.822 ;
      RECT 39.49 2.57 39.505 2.828 ;
      RECT 39.45 2.585 39.49 2.832 ;
      RECT 39.4 2.6 39.45 2.837 ;
      RECT 39.375 2.607 39.4 2.841 ;
      RECT 39.315 2.602 39.375 2.845 ;
      RECT 39.3 2.593 39.315 2.849 ;
      RECT 39.23 2.583 39.3 2.845 ;
      RECT 39.205 2.575 39.225 2.835 ;
      RECT 39.146 2.575 39.205 2.813 ;
      RECT 39.06 2.575 39.146 2.77 ;
      RECT 39.225 2.575 39.23 2.84 ;
      RECT 39.92 1.806 40.09 2.14 ;
      RECT 39.89 1.806 40.09 2.135 ;
      RECT 39.83 1.773 39.89 2.123 ;
      RECT 39.83 1.829 40.1 2.118 ;
      RECT 39.805 1.829 40.1 2.112 ;
      RECT 39.8 1.77 39.83 2.109 ;
      RECT 39.785 1.776 39.92 2.107 ;
      RECT 39.78 1.784 40.005 2.095 ;
      RECT 39.78 1.836 40.115 2.048 ;
      RECT 39.765 1.792 40.005 2.043 ;
      RECT 39.765 1.862 40.125 1.984 ;
      RECT 39.735 1.812 40.09 1.945 ;
      RECT 39.735 1.902 40.135 1.941 ;
      RECT 39.785 1.781 40.005 2.107 ;
      RECT 39.125 2.111 39.18 2.375 ;
      RECT 39.125 2.111 39.245 2.374 ;
      RECT 39.125 2.111 39.27 2.373 ;
      RECT 39.125 2.111 39.335 2.372 ;
      RECT 39.27 2.077 39.35 2.371 ;
      RECT 39.085 2.121 39.495 2.37 ;
      RECT 39.125 2.118 39.495 2.37 ;
      RECT 39.085 2.126 39.5 2.363 ;
      RECT 39.07 2.128 39.5 2.362 ;
      RECT 39.07 2.135 39.505 2.358 ;
      RECT 39.05 2.134 39.5 2.354 ;
      RECT 39.05 2.142 39.51 2.353 ;
      RECT 39.045 2.139 39.505 2.349 ;
      RECT 39.045 2.152 39.52 2.348 ;
      RECT 39.03 2.142 39.51 2.347 ;
      RECT 38.995 2.155 39.52 2.34 ;
      RECT 39.18 2.11 39.49 2.37 ;
      RECT 39.18 2.095 39.44 2.37 ;
      RECT 39.245 2.082 39.375 2.37 ;
      RECT 38.79 3.171 38.805 3.564 ;
      RECT 38.755 3.176 38.805 3.563 ;
      RECT 38.79 3.175 38.85 3.562 ;
      RECT 38.735 3.186 38.85 3.561 ;
      RECT 38.75 3.182 38.85 3.561 ;
      RECT 38.715 3.192 38.925 3.558 ;
      RECT 38.715 3.211 38.97 3.556 ;
      RECT 38.715 3.218 38.975 3.553 ;
      RECT 38.7 3.195 38.925 3.55 ;
      RECT 38.68 3.2 38.925 3.543 ;
      RECT 38.675 3.204 38.925 3.539 ;
      RECT 38.675 3.221 38.985 3.538 ;
      RECT 38.655 3.215 38.97 3.534 ;
      RECT 38.655 3.224 38.99 3.528 ;
      RECT 38.65 3.23 38.99 3.3 ;
      RECT 38.715 3.19 38.85 3.558 ;
      RECT 38.59 2.553 38.79 2.865 ;
      RECT 38.665 2.531 38.79 2.865 ;
      RECT 38.605 2.55 38.795 2.85 ;
      RECT 38.575 2.561 38.795 2.848 ;
      RECT 38.59 2.556 38.8 2.814 ;
      RECT 38.575 2.66 38.805 2.781 ;
      RECT 38.605 2.532 38.79 2.865 ;
      RECT 38.665 2.51 38.765 2.865 ;
      RECT 38.69 2.507 38.765 2.865 ;
      RECT 38.69 2.502 38.71 2.865 ;
      RECT 38.095 2.57 38.27 2.745 ;
      RECT 38.09 2.57 38.27 2.743 ;
      RECT 38.065 2.57 38.27 2.738 ;
      RECT 38.01 2.55 38.18 2.728 ;
      RECT 38.01 2.557 38.245 2.728 ;
      RECT 38.095 3.237 38.11 3.42 ;
      RECT 38.085 3.215 38.095 3.42 ;
      RECT 38.07 3.195 38.085 3.42 ;
      RECT 38.06 3.17 38.07 3.42 ;
      RECT 38.03 3.135 38.06 3.42 ;
      RECT 37.995 3.075 38.03 3.42 ;
      RECT 37.99 3.037 37.995 3.42 ;
      RECT 37.94 2.988 37.99 3.42 ;
      RECT 37.93 2.938 37.94 3.408 ;
      RECT 37.915 2.917 37.93 3.368 ;
      RECT 37.895 2.885 37.915 3.318 ;
      RECT 37.87 2.841 37.895 3.258 ;
      RECT 37.865 2.813 37.87 3.213 ;
      RECT 37.86 2.804 37.865 3.199 ;
      RECT 37.855 2.797 37.86 3.186 ;
      RECT 37.85 2.792 37.855 3.175 ;
      RECT 37.845 2.777 37.85 3.165 ;
      RECT 37.84 2.755 37.845 3.152 ;
      RECT 37.83 2.715 37.84 3.127 ;
      RECT 37.805 2.645 37.83 3.083 ;
      RECT 37.8 2.585 37.805 3.048 ;
      RECT 37.785 2.565 37.8 3.015 ;
      RECT 37.78 2.565 37.785 2.99 ;
      RECT 37.75 2.565 37.78 2.945 ;
      RECT 37.705 2.565 37.75 2.885 ;
      RECT 37.63 2.565 37.705 2.833 ;
      RECT 37.625 2.565 37.63 2.798 ;
      RECT 37.62 2.565 37.625 2.788 ;
      RECT 37.615 2.565 37.62 2.768 ;
      RECT 37.88 1.785 38.05 2.255 ;
      RECT 37.825 1.778 38.02 2.239 ;
      RECT 37.825 1.792 38.055 2.238 ;
      RECT 37.81 1.793 38.055 2.219 ;
      RECT 37.805 1.811 38.055 2.205 ;
      RECT 37.81 1.794 38.06 2.203 ;
      RECT 37.795 1.825 38.06 2.188 ;
      RECT 37.81 1.8 38.065 2.173 ;
      RECT 37.79 1.84 38.065 2.17 ;
      RECT 37.805 1.812 38.07 2.155 ;
      RECT 37.805 1.824 38.075 2.135 ;
      RECT 37.79 1.84 38.08 2.118 ;
      RECT 37.79 1.85 38.085 1.973 ;
      RECT 37.785 1.85 38.085 1.93 ;
      RECT 37.785 1.865 38.09 1.908 ;
      RECT 37.88 1.775 38.02 2.255 ;
      RECT 37.88 1.773 37.99 2.255 ;
      RECT 37.966 1.77 37.99 2.255 ;
      RECT 37.625 3.437 37.63 3.483 ;
      RECT 37.615 3.285 37.625 3.507 ;
      RECT 37.61 3.13 37.615 3.532 ;
      RECT 37.595 3.092 37.61 3.543 ;
      RECT 37.59 3.075 37.595 3.55 ;
      RECT 37.58 3.063 37.59 3.557 ;
      RECT 37.575 3.054 37.58 3.559 ;
      RECT 37.57 3.052 37.575 3.563 ;
      RECT 37.525 3.043 37.57 3.578 ;
      RECT 37.52 3.035 37.525 3.592 ;
      RECT 37.515 3.032 37.52 3.596 ;
      RECT 37.5 3.027 37.515 3.604 ;
      RECT 37.445 3.017 37.5 3.615 ;
      RECT 37.41 3.005 37.445 3.616 ;
      RECT 37.401 3 37.41 3.61 ;
      RECT 37.315 3 37.401 3.6 ;
      RECT 37.285 3 37.315 3.578 ;
      RECT 37.275 3 37.28 3.558 ;
      RECT 37.27 3 37.275 3.52 ;
      RECT 37.265 3 37.27 3.478 ;
      RECT 37.26 3 37.265 3.438 ;
      RECT 37.255 3 37.26 3.368 ;
      RECT 37.245 3 37.255 3.29 ;
      RECT 37.24 3 37.245 3.19 ;
      RECT 37.28 3 37.285 3.56 ;
      RECT 36.775 3.082 36.865 3.56 ;
      RECT 36.76 3.085 36.88 3.558 ;
      RECT 36.775 3.084 36.88 3.558 ;
      RECT 36.74 3.091 36.905 3.548 ;
      RECT 36.76 3.085 36.905 3.548 ;
      RECT 36.725 3.097 36.905 3.536 ;
      RECT 36.76 3.088 36.955 3.529 ;
      RECT 36.711 3.105 36.955 3.527 ;
      RECT 36.74 3.095 36.965 3.515 ;
      RECT 36.711 3.116 36.995 3.506 ;
      RECT 36.625 3.14 36.995 3.5 ;
      RECT 36.625 3.153 37.035 3.483 ;
      RECT 36.62 3.175 37.035 3.476 ;
      RECT 36.59 3.19 37.035 3.466 ;
      RECT 36.585 3.201 37.035 3.456 ;
      RECT 36.555 3.214 37.035 3.447 ;
      RECT 36.54 3.232 37.035 3.436 ;
      RECT 36.515 3.245 37.035 3.426 ;
      RECT 36.775 3.081 36.785 3.56 ;
      RECT 36.821 2.505 36.86 2.75 ;
      RECT 36.735 2.505 36.87 2.748 ;
      RECT 36.62 2.53 36.87 2.745 ;
      RECT 36.62 2.53 36.875 2.743 ;
      RECT 36.62 2.53 36.89 2.738 ;
      RECT 36.726 2.505 36.905 2.718 ;
      RECT 36.64 2.513 36.905 2.718 ;
      RECT 36.31 1.865 36.48 2.3 ;
      RECT 36.3 1.899 36.48 2.283 ;
      RECT 36.38 1.835 36.55 2.27 ;
      RECT 36.285 1.91 36.55 2.248 ;
      RECT 36.38 1.845 36.555 2.238 ;
      RECT 36.31 1.897 36.585 2.223 ;
      RECT 36.27 1.923 36.585 2.208 ;
      RECT 36.27 1.965 36.595 2.188 ;
      RECT 36.265 1.99 36.6 2.17 ;
      RECT 36.265 2 36.605 2.155 ;
      RECT 36.26 1.937 36.585 2.153 ;
      RECT 36.26 2.01 36.61 2.138 ;
      RECT 36.255 1.947 36.585 2.135 ;
      RECT 36.25 2.031 36.615 2.118 ;
      RECT 36.25 2.063 36.62 2.098 ;
      RECT 36.245 1.977 36.595 2.09 ;
      RECT 36.25 1.962 36.585 2.118 ;
      RECT 36.265 1.932 36.585 2.17 ;
      RECT 36.11 2.519 36.335 2.775 ;
      RECT 36.11 2.552 36.355 2.765 ;
      RECT 36.075 2.552 36.355 2.763 ;
      RECT 36.075 2.565 36.36 2.753 ;
      RECT 36.075 2.585 36.37 2.745 ;
      RECT 36.075 2.682 36.375 2.738 ;
      RECT 36.055 2.43 36.185 2.728 ;
      RECT 36.01 2.585 36.37 2.67 ;
      RECT 36 2.43 36.185 2.615 ;
      RECT 36 2.462 36.271 2.615 ;
      RECT 35.965 2.992 35.985 3.17 ;
      RECT 35.93 2.945 35.965 3.17 ;
      RECT 35.915 2.885 35.93 3.17 ;
      RECT 35.89 2.832 35.915 3.17 ;
      RECT 35.875 2.785 35.89 3.17 ;
      RECT 35.855 2.762 35.875 3.17 ;
      RECT 35.83 2.727 35.855 3.17 ;
      RECT 35.82 2.573 35.83 3.17 ;
      RECT 35.79 2.568 35.82 3.161 ;
      RECT 35.785 2.565 35.79 3.151 ;
      RECT 35.77 2.565 35.785 3.125 ;
      RECT 35.765 2.565 35.77 3.088 ;
      RECT 35.74 2.565 35.765 3.04 ;
      RECT 35.72 2.565 35.74 2.965 ;
      RECT 35.71 2.565 35.72 2.925 ;
      RECT 35.705 2.565 35.71 2.9 ;
      RECT 35.7 2.565 35.705 2.883 ;
      RECT 35.695 2.565 35.7 2.865 ;
      RECT 35.69 2.566 35.695 2.855 ;
      RECT 35.68 2.568 35.69 2.823 ;
      RECT 35.67 2.57 35.68 2.79 ;
      RECT 35.66 2.573 35.67 2.763 ;
      RECT 35.985 3 36.21 3.17 ;
      RECT 35.315 1.812 35.485 2.265 ;
      RECT 35.315 1.812 35.575 2.231 ;
      RECT 35.315 1.812 35.605 2.215 ;
      RECT 35.315 1.812 35.635 2.188 ;
      RECT 35.571 1.79 35.65 2.17 ;
      RECT 35.35 1.797 35.655 2.155 ;
      RECT 35.35 1.805 35.665 2.118 ;
      RECT 35.31 1.832 35.665 2.09 ;
      RECT 35.295 1.845 35.665 2.055 ;
      RECT 35.315 1.82 35.685 2.045 ;
      RECT 35.29 1.885 35.685 2.015 ;
      RECT 35.29 1.915 35.69 1.998 ;
      RECT 35.285 1.945 35.69 1.985 ;
      RECT 35.35 1.794 35.65 2.17 ;
      RECT 35.485 1.791 35.571 2.249 ;
      RECT 35.436 1.792 35.65 2.17 ;
      RECT 35.58 3.452 35.625 3.645 ;
      RECT 35.57 3.422 35.58 3.645 ;
      RECT 35.565 3.407 35.57 3.645 ;
      RECT 35.525 3.317 35.565 3.645 ;
      RECT 35.52 3.23 35.525 3.645 ;
      RECT 35.51 3.2 35.52 3.645 ;
      RECT 35.505 3.16 35.51 3.645 ;
      RECT 35.495 3.122 35.505 3.645 ;
      RECT 35.49 3.087 35.495 3.645 ;
      RECT 35.47 3.04 35.49 3.645 ;
      RECT 35.455 2.965 35.47 3.645 ;
      RECT 35.45 2.92 35.455 3.64 ;
      RECT 35.445 2.9 35.45 3.613 ;
      RECT 35.44 2.88 35.445 3.598 ;
      RECT 35.435 2.855 35.44 3.578 ;
      RECT 35.43 2.833 35.435 3.563 ;
      RECT 35.425 2.811 35.43 3.545 ;
      RECT 35.42 2.79 35.425 3.535 ;
      RECT 35.41 2.762 35.42 3.505 ;
      RECT 35.4 2.725 35.41 3.473 ;
      RECT 35.39 2.685 35.4 3.44 ;
      RECT 35.38 2.663 35.39 3.41 ;
      RECT 35.35 2.615 35.38 3.342 ;
      RECT 35.335 2.575 35.35 3.269 ;
      RECT 35.325 2.575 35.335 3.235 ;
      RECT 35.32 2.575 35.325 3.21 ;
      RECT 35.315 2.575 35.32 3.195 ;
      RECT 35.31 2.575 35.315 3.173 ;
      RECT 35.305 2.575 35.31 3.16 ;
      RECT 35.29 2.575 35.305 3.125 ;
      RECT 35.27 2.575 35.29 3.065 ;
      RECT 35.26 2.575 35.27 3.015 ;
      RECT 35.24 2.575 35.26 2.963 ;
      RECT 35.22 2.575 35.24 2.92 ;
      RECT 35.21 2.575 35.22 2.908 ;
      RECT 35.18 2.575 35.21 2.895 ;
      RECT 35.15 2.596 35.18 2.875 ;
      RECT 35.14 2.624 35.15 2.855 ;
      RECT 35.125 2.641 35.14 2.823 ;
      RECT 35.12 2.655 35.125 2.79 ;
      RECT 35.115 2.663 35.12 2.763 ;
      RECT 35.11 2.671 35.115 2.725 ;
      RECT 35.115 3.195 35.12 3.53 ;
      RECT 35.08 3.182 35.115 3.529 ;
      RECT 35.01 3.122 35.08 3.528 ;
      RECT 34.93 3.065 35.01 3.527 ;
      RECT 34.795 3.025 34.93 3.526 ;
      RECT 34.795 3.212 35.13 3.515 ;
      RECT 34.755 3.212 35.13 3.505 ;
      RECT 34.755 3.23 35.135 3.5 ;
      RECT 34.755 3.32 35.14 3.49 ;
      RECT 34.75 3.015 34.915 3.47 ;
      RECT 34.745 3.015 34.915 3.213 ;
      RECT 34.745 3.172 35.11 3.213 ;
      RECT 34.745 3.16 35.105 3.213 ;
      RECT 33.885 5.02 34.055 6.49 ;
      RECT 33.885 6.315 34.06 6.485 ;
      RECT 33.515 1.74 33.685 2.93 ;
      RECT 33.515 1.74 33.985 1.91 ;
      RECT 33.515 6.97 33.985 7.14 ;
      RECT 33.515 5.95 33.685 7.14 ;
      RECT 32.525 1.74 32.695 2.93 ;
      RECT 32.525 1.74 32.995 1.91 ;
      RECT 32.525 6.97 32.995 7.14 ;
      RECT 32.525 5.95 32.695 7.14 ;
      RECT 30.675 2.635 30.845 3.865 ;
      RECT 30.73 0.855 30.9 2.805 ;
      RECT 30.675 0.575 30.845 1.025 ;
      RECT 30.675 7.855 30.845 8.305 ;
      RECT 30.73 6.075 30.9 8.025 ;
      RECT 30.675 5.015 30.845 6.245 ;
      RECT 30.155 0.575 30.325 3.865 ;
      RECT 30.155 2.075 30.56 2.405 ;
      RECT 30.155 1.235 30.56 1.565 ;
      RECT 30.155 5.015 30.325 8.305 ;
      RECT 30.155 7.315 30.56 7.645 ;
      RECT 30.155 6.475 30.56 6.805 ;
      RECT 27.49 1.975 28.22 2.215 ;
      RECT 28.032 1.77 28.22 2.215 ;
      RECT 27.86 1.782 28.235 2.209 ;
      RECT 27.775 1.797 28.255 2.194 ;
      RECT 27.775 1.812 28.26 2.184 ;
      RECT 27.73 1.832 28.275 2.176 ;
      RECT 27.707 1.867 28.29 2.13 ;
      RECT 27.621 1.89 28.295 2.09 ;
      RECT 27.621 1.908 28.305 2.06 ;
      RECT 27.49 1.977 28.31 2.023 ;
      RECT 27.535 1.92 28.305 2.06 ;
      RECT 27.621 1.872 28.29 2.13 ;
      RECT 27.707 1.841 28.275 2.176 ;
      RECT 27.73 1.822 28.26 2.184 ;
      RECT 27.775 1.795 28.235 2.209 ;
      RECT 27.86 1.777 28.22 2.215 ;
      RECT 27.946 1.771 28.22 2.215 ;
      RECT 28.032 1.766 28.165 2.215 ;
      RECT 28.118 1.761 28.165 2.215 ;
      RECT 27.81 2.659 27.98 3.045 ;
      RECT 27.805 2.659 27.98 3.04 ;
      RECT 27.78 2.659 27.98 3.005 ;
      RECT 27.78 2.687 27.99 2.995 ;
      RECT 27.76 2.687 27.99 2.955 ;
      RECT 27.755 2.687 27.99 2.928 ;
      RECT 27.755 2.705 27.995 2.92 ;
      RECT 27.7 2.705 27.995 2.855 ;
      RECT 27.7 2.722 28.005 2.838 ;
      RECT 27.69 2.722 28.005 2.778 ;
      RECT 27.69 2.739 28.01 2.775 ;
      RECT 27.685 2.575 27.855 2.753 ;
      RECT 27.685 2.609 27.941 2.753 ;
      RECT 27.68 3.375 27.685 3.388 ;
      RECT 27.675 3.27 27.68 3.393 ;
      RECT 27.65 3.13 27.675 3.408 ;
      RECT 27.615 3.081 27.65 3.44 ;
      RECT 27.61 3.049 27.615 3.46 ;
      RECT 27.605 3.04 27.61 3.46 ;
      RECT 27.525 3.005 27.605 3.46 ;
      RECT 27.462 2.975 27.525 3.46 ;
      RECT 27.376 2.963 27.462 3.46 ;
      RECT 27.29 2.949 27.376 3.46 ;
      RECT 27.21 2.936 27.29 3.446 ;
      RECT 27.175 2.928 27.21 3.426 ;
      RECT 27.165 2.925 27.175 3.417 ;
      RECT 27.135 2.92 27.165 3.404 ;
      RECT 27.085 2.895 27.135 3.38 ;
      RECT 27.071 2.869 27.085 3.362 ;
      RECT 26.985 2.829 27.071 3.338 ;
      RECT 26.94 2.777 26.985 3.307 ;
      RECT 26.93 2.752 26.94 3.294 ;
      RECT 26.925 2.533 26.93 2.555 ;
      RECT 26.92 2.735 26.93 3.29 ;
      RECT 26.92 2.531 26.925 2.645 ;
      RECT 26.91 2.527 26.92 3.286 ;
      RECT 26.866 2.525 26.91 3.274 ;
      RECT 26.78 2.525 26.866 3.245 ;
      RECT 26.75 2.525 26.78 3.218 ;
      RECT 26.735 2.525 26.75 3.206 ;
      RECT 26.695 2.537 26.735 3.191 ;
      RECT 26.675 2.556 26.695 3.17 ;
      RECT 26.665 2.566 26.675 3.154 ;
      RECT 26.655 2.572 26.665 3.143 ;
      RECT 26.635 2.582 26.655 3.126 ;
      RECT 26.63 2.591 26.635 3.113 ;
      RECT 26.625 2.595 26.63 3.063 ;
      RECT 26.615 2.601 26.625 2.98 ;
      RECT 26.61 2.605 26.615 2.894 ;
      RECT 26.605 2.625 26.61 2.831 ;
      RECT 26.6 2.648 26.605 2.778 ;
      RECT 26.595 2.666 26.6 2.723 ;
      RECT 27.205 2.485 27.375 2.745 ;
      RECT 27.375 2.45 27.42 2.731 ;
      RECT 27.336 2.452 27.425 2.714 ;
      RECT 27.225 2.469 27.511 2.685 ;
      RECT 27.225 2.484 27.515 2.657 ;
      RECT 27.225 2.465 27.425 2.714 ;
      RECT 27.25 2.453 27.375 2.745 ;
      RECT 27.336 2.451 27.42 2.731 ;
      RECT 26.39 1.84 26.56 2.33 ;
      RECT 26.39 1.84 26.595 2.31 ;
      RECT 26.525 1.76 26.635 2.27 ;
      RECT 26.506 1.764 26.655 2.24 ;
      RECT 26.42 1.772 26.675 2.223 ;
      RECT 26.42 1.778 26.68 2.213 ;
      RECT 26.42 1.787 26.7 2.201 ;
      RECT 26.395 1.812 26.73 2.179 ;
      RECT 26.395 1.832 26.735 2.159 ;
      RECT 26.39 1.845 26.745 2.139 ;
      RECT 26.39 1.912 26.75 2.12 ;
      RECT 26.39 2.045 26.755 2.107 ;
      RECT 26.385 1.85 26.745 1.94 ;
      RECT 26.395 1.807 26.7 2.201 ;
      RECT 26.506 1.762 26.635 2.27 ;
      RECT 26.38 3.515 26.68 3.77 ;
      RECT 26.465 3.481 26.68 3.77 ;
      RECT 26.465 3.484 26.685 3.63 ;
      RECT 26.4 3.505 26.685 3.63 ;
      RECT 26.435 3.495 26.68 3.77 ;
      RECT 26.43 3.5 26.685 3.63 ;
      RECT 26.465 3.479 26.666 3.77 ;
      RECT 26.551 3.47 26.666 3.77 ;
      RECT 26.551 3.464 26.58 3.77 ;
      RECT 26.04 3.105 26.05 3.595 ;
      RECT 25.7 3.04 25.71 3.34 ;
      RECT 26.215 3.212 26.22 3.431 ;
      RECT 26.205 3.192 26.215 3.448 ;
      RECT 26.195 3.172 26.205 3.478 ;
      RECT 26.19 3.162 26.195 3.493 ;
      RECT 26.185 3.158 26.19 3.498 ;
      RECT 26.17 3.15 26.185 3.505 ;
      RECT 26.13 3.13 26.17 3.53 ;
      RECT 26.105 3.112 26.13 3.563 ;
      RECT 26.1 3.11 26.105 3.576 ;
      RECT 26.08 3.107 26.1 3.58 ;
      RECT 26.05 3.105 26.08 3.59 ;
      RECT 25.98 3.107 26.04 3.591 ;
      RECT 25.96 3.107 25.98 3.585 ;
      RECT 25.935 3.105 25.96 3.582 ;
      RECT 25.9 3.1 25.935 3.578 ;
      RECT 25.88 3.094 25.9 3.565 ;
      RECT 25.87 3.091 25.88 3.553 ;
      RECT 25.85 3.088 25.87 3.538 ;
      RECT 25.83 3.084 25.85 3.52 ;
      RECT 25.825 3.081 25.83 3.51 ;
      RECT 25.82 3.08 25.825 3.508 ;
      RECT 25.81 3.077 25.82 3.5 ;
      RECT 25.8 3.071 25.81 3.483 ;
      RECT 25.79 3.065 25.8 3.465 ;
      RECT 25.78 3.059 25.79 3.453 ;
      RECT 25.77 3.053 25.78 3.433 ;
      RECT 25.765 3.049 25.77 3.418 ;
      RECT 25.76 3.047 25.765 3.41 ;
      RECT 25.755 3.045 25.76 3.403 ;
      RECT 25.75 3.043 25.755 3.393 ;
      RECT 25.745 3.041 25.75 3.387 ;
      RECT 25.735 3.04 25.745 3.377 ;
      RECT 25.725 3.04 25.735 3.368 ;
      RECT 25.71 3.04 25.725 3.353 ;
      RECT 25.67 3.04 25.7 3.337 ;
      RECT 25.65 3.042 25.67 3.332 ;
      RECT 25.645 3.047 25.65 3.33 ;
      RECT 25.615 3.055 25.645 3.328 ;
      RECT 25.585 3.07 25.615 3.327 ;
      RECT 25.54 3.092 25.585 3.332 ;
      RECT 25.535 3.107 25.54 3.336 ;
      RECT 25.52 3.112 25.535 3.338 ;
      RECT 25.515 3.116 25.52 3.34 ;
      RECT 25.455 3.139 25.515 3.349 ;
      RECT 25.435 3.165 25.455 3.362 ;
      RECT 25.425 3.172 25.435 3.366 ;
      RECT 25.41 3.179 25.425 3.369 ;
      RECT 25.39 3.189 25.41 3.372 ;
      RECT 25.385 3.197 25.39 3.375 ;
      RECT 25.34 3.202 25.385 3.382 ;
      RECT 25.33 3.205 25.34 3.389 ;
      RECT 25.32 3.205 25.33 3.393 ;
      RECT 25.285 3.207 25.32 3.405 ;
      RECT 25.265 3.21 25.285 3.418 ;
      RECT 25.225 3.213 25.265 3.429 ;
      RECT 25.21 3.215 25.225 3.442 ;
      RECT 25.2 3.215 25.21 3.447 ;
      RECT 25.175 3.216 25.2 3.455 ;
      RECT 25.165 3.218 25.175 3.46 ;
      RECT 25.16 3.219 25.165 3.463 ;
      RECT 25.135 3.217 25.16 3.466 ;
      RECT 25.12 3.215 25.135 3.467 ;
      RECT 25.1 3.212 25.12 3.469 ;
      RECT 25.08 3.207 25.1 3.469 ;
      RECT 25.02 3.202 25.08 3.466 ;
      RECT 24.985 3.177 25.02 3.462 ;
      RECT 24.975 3.154 24.985 3.46 ;
      RECT 24.945 3.131 24.975 3.46 ;
      RECT 24.935 3.11 24.945 3.46 ;
      RECT 24.91 3.092 24.935 3.458 ;
      RECT 24.895 3.07 24.91 3.455 ;
      RECT 24.88 3.052 24.895 3.453 ;
      RECT 24.86 3.042 24.88 3.451 ;
      RECT 24.845 3.037 24.86 3.45 ;
      RECT 24.83 3.035 24.845 3.449 ;
      RECT 24.8 3.036 24.83 3.447 ;
      RECT 24.78 3.039 24.8 3.445 ;
      RECT 24.723 3.043 24.78 3.445 ;
      RECT 24.637 3.052 24.723 3.445 ;
      RECT 24.551 3.063 24.637 3.445 ;
      RECT 24.465 3.074 24.551 3.445 ;
      RECT 24.445 3.081 24.465 3.453 ;
      RECT 24.435 3.084 24.445 3.46 ;
      RECT 24.37 3.089 24.435 3.478 ;
      RECT 24.34 3.096 24.37 3.503 ;
      RECT 24.33 3.099 24.34 3.51 ;
      RECT 24.285 3.103 24.33 3.515 ;
      RECT 24.255 3.108 24.285 3.52 ;
      RECT 24.254 3.11 24.255 3.52 ;
      RECT 24.168 3.116 24.254 3.52 ;
      RECT 24.082 3.127 24.168 3.52 ;
      RECT 23.996 3.139 24.082 3.52 ;
      RECT 23.91 3.15 23.996 3.52 ;
      RECT 23.895 3.157 23.91 3.515 ;
      RECT 23.89 3.159 23.895 3.509 ;
      RECT 23.87 3.17 23.89 3.504 ;
      RECT 23.86 3.188 23.87 3.498 ;
      RECT 23.855 3.2 23.86 3.298 ;
      RECT 26.15 1.953 26.17 2.04 ;
      RECT 26.145 1.888 26.15 2.072 ;
      RECT 26.135 1.855 26.145 2.077 ;
      RECT 26.13 1.835 26.135 2.083 ;
      RECT 26.1 1.835 26.13 2.1 ;
      RECT 26.051 1.835 26.1 2.136 ;
      RECT 25.965 1.835 26.051 2.194 ;
      RECT 25.936 1.845 25.965 2.243 ;
      RECT 25.85 1.887 25.936 2.296 ;
      RECT 25.83 1.925 25.85 2.343 ;
      RECT 25.805 1.942 25.83 2.363 ;
      RECT 25.795 1.956 25.805 2.383 ;
      RECT 25.79 1.962 25.795 2.393 ;
      RECT 25.785 1.966 25.79 2.4 ;
      RECT 25.735 1.986 25.785 2.405 ;
      RECT 25.67 2.03 25.735 2.405 ;
      RECT 25.645 2.08 25.67 2.405 ;
      RECT 25.635 2.11 25.645 2.405 ;
      RECT 25.63 2.137 25.635 2.405 ;
      RECT 25.625 2.155 25.63 2.405 ;
      RECT 25.615 2.197 25.625 2.405 ;
      RECT 25.965 2.755 26.135 2.93 ;
      RECT 25.905 2.583 25.965 2.918 ;
      RECT 25.895 2.576 25.905 2.901 ;
      RECT 25.85 2.755 26.135 2.881 ;
      RECT 25.831 2.755 26.135 2.859 ;
      RECT 25.745 2.755 26.135 2.824 ;
      RECT 25.725 2.575 25.895 2.78 ;
      RECT 25.725 2.722 26.13 2.78 ;
      RECT 25.725 2.67 26.105 2.78 ;
      RECT 25.725 2.625 26.07 2.78 ;
      RECT 25.725 2.607 26.035 2.78 ;
      RECT 25.725 2.597 26.03 2.78 ;
      RECT 25.375 5.015 25.545 8.305 ;
      RECT 25.375 7.315 25.78 7.645 ;
      RECT 25.375 6.475 25.78 6.805 ;
      RECT 25.445 3.555 25.635 3.78 ;
      RECT 25.435 3.556 25.64 3.775 ;
      RECT 25.435 3.558 25.65 3.755 ;
      RECT 25.435 3.562 25.655 3.74 ;
      RECT 25.435 3.549 25.605 3.775 ;
      RECT 25.435 3.552 25.63 3.775 ;
      RECT 25.445 3.548 25.605 3.78 ;
      RECT 25.531 3.546 25.605 3.78 ;
      RECT 25.155 2.797 25.325 3.035 ;
      RECT 25.155 2.797 25.411 2.949 ;
      RECT 25.155 2.797 25.415 2.859 ;
      RECT 25.205 2.57 25.425 2.838 ;
      RECT 25.2 2.587 25.43 2.811 ;
      RECT 25.165 2.745 25.43 2.811 ;
      RECT 25.185 2.595 25.325 3.035 ;
      RECT 25.175 2.677 25.435 2.794 ;
      RECT 25.17 2.725 25.435 2.794 ;
      RECT 25.175 2.635 25.43 2.811 ;
      RECT 25.2 2.572 25.425 2.838 ;
      RECT 24.765 2.547 24.935 2.745 ;
      RECT 24.765 2.547 24.98 2.72 ;
      RECT 24.835 2.49 25.005 2.678 ;
      RECT 24.81 2.505 25.005 2.678 ;
      RECT 24.425 2.551 24.455 2.745 ;
      RECT 24.42 2.523 24.425 2.745 ;
      RECT 24.39 2.497 24.42 2.747 ;
      RECT 24.365 2.455 24.39 2.75 ;
      RECT 24.355 2.427 24.365 2.752 ;
      RECT 24.32 2.407 24.355 2.754 ;
      RECT 24.255 2.392 24.32 2.76 ;
      RECT 24.205 2.39 24.255 2.766 ;
      RECT 24.182 2.392 24.205 2.771 ;
      RECT 24.096 2.403 24.182 2.777 ;
      RECT 24.01 2.421 24.096 2.787 ;
      RECT 23.995 2.432 24.01 2.793 ;
      RECT 23.925 2.455 23.995 2.799 ;
      RECT 23.87 2.487 23.925 2.807 ;
      RECT 23.83 2.51 23.87 2.813 ;
      RECT 23.816 2.523 23.83 2.816 ;
      RECT 23.73 2.545 23.816 2.822 ;
      RECT 23.715 2.57 23.73 2.828 ;
      RECT 23.675 2.585 23.715 2.832 ;
      RECT 23.625 2.6 23.675 2.837 ;
      RECT 23.6 2.607 23.625 2.841 ;
      RECT 23.54 2.602 23.6 2.845 ;
      RECT 23.525 2.593 23.54 2.849 ;
      RECT 23.455 2.583 23.525 2.845 ;
      RECT 23.43 2.575 23.45 2.835 ;
      RECT 23.371 2.575 23.43 2.813 ;
      RECT 23.285 2.575 23.371 2.77 ;
      RECT 23.45 2.575 23.455 2.84 ;
      RECT 24.145 1.806 24.315 2.14 ;
      RECT 24.115 1.806 24.315 2.135 ;
      RECT 24.055 1.773 24.115 2.123 ;
      RECT 24.055 1.829 24.325 2.118 ;
      RECT 24.03 1.829 24.325 2.112 ;
      RECT 24.025 1.77 24.055 2.109 ;
      RECT 24.01 1.776 24.145 2.107 ;
      RECT 24.005 1.784 24.23 2.095 ;
      RECT 24.005 1.836 24.34 2.048 ;
      RECT 23.99 1.792 24.23 2.043 ;
      RECT 23.99 1.862 24.35 1.984 ;
      RECT 23.96 1.812 24.315 1.945 ;
      RECT 23.96 1.902 24.36 1.941 ;
      RECT 24.01 1.781 24.23 2.107 ;
      RECT 23.35 2.111 23.405 2.375 ;
      RECT 23.35 2.111 23.47 2.374 ;
      RECT 23.35 2.111 23.495 2.373 ;
      RECT 23.35 2.111 23.56 2.372 ;
      RECT 23.495 2.077 23.575 2.371 ;
      RECT 23.31 2.121 23.72 2.37 ;
      RECT 23.35 2.118 23.72 2.37 ;
      RECT 23.31 2.126 23.725 2.363 ;
      RECT 23.295 2.128 23.725 2.362 ;
      RECT 23.295 2.135 23.73 2.358 ;
      RECT 23.275 2.134 23.725 2.354 ;
      RECT 23.275 2.142 23.735 2.353 ;
      RECT 23.27 2.139 23.73 2.349 ;
      RECT 23.27 2.152 23.745 2.348 ;
      RECT 23.255 2.142 23.735 2.347 ;
      RECT 23.22 2.155 23.745 2.34 ;
      RECT 23.405 2.11 23.715 2.37 ;
      RECT 23.405 2.095 23.665 2.37 ;
      RECT 23.47 2.082 23.6 2.37 ;
      RECT 23.015 3.171 23.03 3.564 ;
      RECT 22.98 3.176 23.03 3.563 ;
      RECT 23.015 3.175 23.075 3.562 ;
      RECT 22.96 3.186 23.075 3.561 ;
      RECT 22.975 3.182 23.075 3.561 ;
      RECT 22.94 3.192 23.15 3.558 ;
      RECT 22.94 3.211 23.195 3.556 ;
      RECT 22.94 3.218 23.2 3.553 ;
      RECT 22.925 3.195 23.15 3.55 ;
      RECT 22.905 3.2 23.15 3.543 ;
      RECT 22.9 3.204 23.15 3.539 ;
      RECT 22.9 3.221 23.21 3.538 ;
      RECT 22.88 3.215 23.195 3.534 ;
      RECT 22.88 3.224 23.215 3.528 ;
      RECT 22.875 3.23 23.215 3.3 ;
      RECT 22.94 3.19 23.075 3.558 ;
      RECT 22.815 2.553 23.015 2.865 ;
      RECT 22.89 2.531 23.015 2.865 ;
      RECT 22.83 2.55 23.02 2.85 ;
      RECT 22.8 2.561 23.02 2.848 ;
      RECT 22.815 2.556 23.025 2.814 ;
      RECT 22.8 2.66 23.03 2.781 ;
      RECT 22.83 2.532 23.015 2.865 ;
      RECT 22.89 2.51 22.99 2.865 ;
      RECT 22.915 2.507 22.99 2.865 ;
      RECT 22.915 2.502 22.935 2.865 ;
      RECT 22.32 2.57 22.495 2.745 ;
      RECT 22.315 2.57 22.495 2.743 ;
      RECT 22.29 2.57 22.495 2.738 ;
      RECT 22.235 2.55 22.405 2.728 ;
      RECT 22.235 2.557 22.47 2.728 ;
      RECT 22.32 3.237 22.335 3.42 ;
      RECT 22.31 3.215 22.32 3.42 ;
      RECT 22.295 3.195 22.31 3.42 ;
      RECT 22.285 3.17 22.295 3.42 ;
      RECT 22.255 3.135 22.285 3.42 ;
      RECT 22.22 3.075 22.255 3.42 ;
      RECT 22.215 3.037 22.22 3.42 ;
      RECT 22.165 2.988 22.215 3.42 ;
      RECT 22.155 2.938 22.165 3.408 ;
      RECT 22.14 2.917 22.155 3.368 ;
      RECT 22.12 2.885 22.14 3.318 ;
      RECT 22.095 2.841 22.12 3.258 ;
      RECT 22.09 2.813 22.095 3.213 ;
      RECT 22.085 2.804 22.09 3.199 ;
      RECT 22.08 2.797 22.085 3.186 ;
      RECT 22.075 2.792 22.08 3.175 ;
      RECT 22.07 2.777 22.075 3.165 ;
      RECT 22.065 2.755 22.07 3.152 ;
      RECT 22.055 2.715 22.065 3.127 ;
      RECT 22.03 2.645 22.055 3.083 ;
      RECT 22.025 2.585 22.03 3.048 ;
      RECT 22.01 2.565 22.025 3.015 ;
      RECT 22.005 2.565 22.01 2.99 ;
      RECT 21.975 2.565 22.005 2.945 ;
      RECT 21.93 2.565 21.975 2.885 ;
      RECT 21.855 2.565 21.93 2.833 ;
      RECT 21.85 2.565 21.855 2.798 ;
      RECT 21.845 2.565 21.85 2.788 ;
      RECT 21.84 2.565 21.845 2.768 ;
      RECT 22.105 1.785 22.275 2.255 ;
      RECT 22.05 1.778 22.245 2.239 ;
      RECT 22.05 1.792 22.28 2.238 ;
      RECT 22.035 1.793 22.28 2.219 ;
      RECT 22.03 1.811 22.28 2.205 ;
      RECT 22.035 1.794 22.285 2.203 ;
      RECT 22.02 1.825 22.285 2.188 ;
      RECT 22.035 1.8 22.29 2.173 ;
      RECT 22.015 1.84 22.29 2.17 ;
      RECT 22.03 1.812 22.295 2.155 ;
      RECT 22.03 1.824 22.3 2.135 ;
      RECT 22.015 1.84 22.305 2.118 ;
      RECT 22.015 1.85 22.31 1.973 ;
      RECT 22.01 1.85 22.31 1.93 ;
      RECT 22.01 1.865 22.315 1.908 ;
      RECT 22.105 1.775 22.245 2.255 ;
      RECT 22.105 1.773 22.215 2.255 ;
      RECT 22.191 1.77 22.215 2.255 ;
      RECT 21.85 3.437 21.855 3.483 ;
      RECT 21.84 3.285 21.85 3.507 ;
      RECT 21.835 3.13 21.84 3.532 ;
      RECT 21.82 3.092 21.835 3.543 ;
      RECT 21.815 3.075 21.82 3.55 ;
      RECT 21.805 3.063 21.815 3.557 ;
      RECT 21.8 3.054 21.805 3.559 ;
      RECT 21.795 3.052 21.8 3.563 ;
      RECT 21.75 3.043 21.795 3.578 ;
      RECT 21.745 3.035 21.75 3.592 ;
      RECT 21.74 3.032 21.745 3.596 ;
      RECT 21.725 3.027 21.74 3.604 ;
      RECT 21.67 3.017 21.725 3.615 ;
      RECT 21.635 3.005 21.67 3.616 ;
      RECT 21.626 3 21.635 3.61 ;
      RECT 21.54 3 21.626 3.6 ;
      RECT 21.51 3 21.54 3.578 ;
      RECT 21.5 3 21.505 3.558 ;
      RECT 21.495 3 21.5 3.52 ;
      RECT 21.49 3 21.495 3.478 ;
      RECT 21.485 3 21.49 3.438 ;
      RECT 21.48 3 21.485 3.368 ;
      RECT 21.47 3 21.48 3.29 ;
      RECT 21.465 3 21.47 3.19 ;
      RECT 21.505 3 21.51 3.56 ;
      RECT 21 3.082 21.09 3.56 ;
      RECT 20.985 3.085 21.105 3.558 ;
      RECT 21 3.084 21.105 3.558 ;
      RECT 20.965 3.091 21.13 3.548 ;
      RECT 20.985 3.085 21.13 3.548 ;
      RECT 20.95 3.097 21.13 3.536 ;
      RECT 20.985 3.088 21.18 3.529 ;
      RECT 20.936 3.105 21.18 3.527 ;
      RECT 20.965 3.095 21.19 3.515 ;
      RECT 20.936 3.116 21.22 3.506 ;
      RECT 20.85 3.14 21.22 3.5 ;
      RECT 20.85 3.153 21.26 3.483 ;
      RECT 20.845 3.175 21.26 3.476 ;
      RECT 20.815 3.19 21.26 3.466 ;
      RECT 20.81 3.201 21.26 3.456 ;
      RECT 20.78 3.214 21.26 3.447 ;
      RECT 20.765 3.232 21.26 3.436 ;
      RECT 20.74 3.245 21.26 3.426 ;
      RECT 21 3.081 21.01 3.56 ;
      RECT 21.046 2.505 21.085 2.75 ;
      RECT 20.96 2.505 21.095 2.748 ;
      RECT 20.845 2.53 21.095 2.745 ;
      RECT 20.845 2.53 21.1 2.743 ;
      RECT 20.845 2.53 21.115 2.738 ;
      RECT 20.951 2.505 21.13 2.718 ;
      RECT 20.865 2.513 21.13 2.718 ;
      RECT 20.535 1.865 20.705 2.3 ;
      RECT 20.525 1.899 20.705 2.283 ;
      RECT 20.605 1.835 20.775 2.27 ;
      RECT 20.51 1.91 20.775 2.248 ;
      RECT 20.605 1.845 20.78 2.238 ;
      RECT 20.535 1.897 20.81 2.223 ;
      RECT 20.495 1.923 20.81 2.208 ;
      RECT 20.495 1.965 20.82 2.188 ;
      RECT 20.49 1.99 20.825 2.17 ;
      RECT 20.49 2 20.83 2.155 ;
      RECT 20.485 1.937 20.81 2.153 ;
      RECT 20.485 2.01 20.835 2.138 ;
      RECT 20.48 1.947 20.81 2.135 ;
      RECT 20.475 2.031 20.84 2.118 ;
      RECT 20.475 2.063 20.845 2.098 ;
      RECT 20.47 1.977 20.82 2.09 ;
      RECT 20.475 1.962 20.81 2.118 ;
      RECT 20.49 1.932 20.81 2.17 ;
      RECT 20.335 2.519 20.56 2.775 ;
      RECT 20.335 2.552 20.58 2.765 ;
      RECT 20.3 2.552 20.58 2.763 ;
      RECT 20.3 2.565 20.585 2.753 ;
      RECT 20.3 2.585 20.595 2.745 ;
      RECT 20.3 2.682 20.6 2.738 ;
      RECT 20.28 2.43 20.41 2.728 ;
      RECT 20.235 2.585 20.595 2.67 ;
      RECT 20.225 2.43 20.41 2.615 ;
      RECT 20.225 2.462 20.496 2.615 ;
      RECT 20.19 2.992 20.21 3.17 ;
      RECT 20.155 2.945 20.19 3.17 ;
      RECT 20.14 2.885 20.155 3.17 ;
      RECT 20.115 2.832 20.14 3.17 ;
      RECT 20.1 2.785 20.115 3.17 ;
      RECT 20.08 2.762 20.1 3.17 ;
      RECT 20.055 2.727 20.08 3.17 ;
      RECT 20.045 2.573 20.055 3.17 ;
      RECT 20.015 2.568 20.045 3.161 ;
      RECT 20.01 2.565 20.015 3.151 ;
      RECT 19.995 2.565 20.01 3.125 ;
      RECT 19.99 2.565 19.995 3.088 ;
      RECT 19.965 2.565 19.99 3.04 ;
      RECT 19.945 2.565 19.965 2.965 ;
      RECT 19.935 2.565 19.945 2.925 ;
      RECT 19.93 2.565 19.935 2.9 ;
      RECT 19.925 2.565 19.93 2.883 ;
      RECT 19.92 2.565 19.925 2.865 ;
      RECT 19.915 2.566 19.92 2.855 ;
      RECT 19.905 2.568 19.915 2.823 ;
      RECT 19.895 2.57 19.905 2.79 ;
      RECT 19.885 2.573 19.895 2.763 ;
      RECT 20.21 3 20.435 3.17 ;
      RECT 19.54 1.812 19.71 2.265 ;
      RECT 19.54 1.812 19.8 2.231 ;
      RECT 19.54 1.812 19.83 2.215 ;
      RECT 19.54 1.812 19.86 2.188 ;
      RECT 19.796 1.79 19.875 2.17 ;
      RECT 19.575 1.797 19.88 2.155 ;
      RECT 19.575 1.805 19.89 2.118 ;
      RECT 19.535 1.832 19.89 2.09 ;
      RECT 19.52 1.845 19.89 2.055 ;
      RECT 19.54 1.82 19.91 2.045 ;
      RECT 19.515 1.885 19.91 2.015 ;
      RECT 19.515 1.915 19.915 1.998 ;
      RECT 19.51 1.945 19.915 1.985 ;
      RECT 19.575 1.794 19.875 2.17 ;
      RECT 19.71 1.791 19.796 2.249 ;
      RECT 19.661 1.792 19.875 2.17 ;
      RECT 19.805 3.452 19.85 3.645 ;
      RECT 19.795 3.422 19.805 3.645 ;
      RECT 19.79 3.407 19.795 3.645 ;
      RECT 19.75 3.317 19.79 3.645 ;
      RECT 19.745 3.23 19.75 3.645 ;
      RECT 19.735 3.2 19.745 3.645 ;
      RECT 19.73 3.16 19.735 3.645 ;
      RECT 19.72 3.122 19.73 3.645 ;
      RECT 19.715 3.087 19.72 3.645 ;
      RECT 19.695 3.04 19.715 3.645 ;
      RECT 19.68 2.965 19.695 3.645 ;
      RECT 19.675 2.92 19.68 3.64 ;
      RECT 19.67 2.9 19.675 3.613 ;
      RECT 19.665 2.88 19.67 3.598 ;
      RECT 19.66 2.855 19.665 3.578 ;
      RECT 19.655 2.833 19.66 3.563 ;
      RECT 19.65 2.811 19.655 3.545 ;
      RECT 19.645 2.79 19.65 3.535 ;
      RECT 19.635 2.762 19.645 3.505 ;
      RECT 19.625 2.725 19.635 3.473 ;
      RECT 19.615 2.685 19.625 3.44 ;
      RECT 19.605 2.663 19.615 3.41 ;
      RECT 19.575 2.615 19.605 3.342 ;
      RECT 19.56 2.575 19.575 3.269 ;
      RECT 19.55 2.575 19.56 3.235 ;
      RECT 19.545 2.575 19.55 3.21 ;
      RECT 19.54 2.575 19.545 3.195 ;
      RECT 19.535 2.575 19.54 3.173 ;
      RECT 19.53 2.575 19.535 3.16 ;
      RECT 19.515 2.575 19.53 3.125 ;
      RECT 19.495 2.575 19.515 3.065 ;
      RECT 19.485 2.575 19.495 3.015 ;
      RECT 19.465 2.575 19.485 2.963 ;
      RECT 19.445 2.575 19.465 2.92 ;
      RECT 19.435 2.575 19.445 2.908 ;
      RECT 19.405 2.575 19.435 2.895 ;
      RECT 19.375 2.596 19.405 2.875 ;
      RECT 19.365 2.624 19.375 2.855 ;
      RECT 19.35 2.641 19.365 2.823 ;
      RECT 19.345 2.655 19.35 2.79 ;
      RECT 19.34 2.663 19.345 2.763 ;
      RECT 19.335 2.671 19.34 2.725 ;
      RECT 19.34 3.195 19.345 3.53 ;
      RECT 19.305 3.182 19.34 3.529 ;
      RECT 19.235 3.122 19.305 3.528 ;
      RECT 19.155 3.065 19.235 3.527 ;
      RECT 19.02 3.025 19.155 3.526 ;
      RECT 19.02 3.212 19.355 3.515 ;
      RECT 18.98 3.212 19.355 3.505 ;
      RECT 18.98 3.23 19.36 3.5 ;
      RECT 18.98 3.32 19.365 3.49 ;
      RECT 18.975 3.015 19.14 3.47 ;
      RECT 18.97 3.015 19.14 3.213 ;
      RECT 18.97 3.172 19.335 3.213 ;
      RECT 18.97 3.16 19.33 3.213 ;
      RECT 18.105 5.02 18.275 6.49 ;
      RECT 18.105 6.315 18.28 6.485 ;
      RECT 17.735 1.74 17.905 2.93 ;
      RECT 17.735 1.74 18.205 1.91 ;
      RECT 17.735 6.97 18.205 7.14 ;
      RECT 17.735 5.95 17.905 7.14 ;
      RECT 16.745 1.74 16.915 2.93 ;
      RECT 16.745 1.74 17.215 1.91 ;
      RECT 16.745 6.97 17.215 7.14 ;
      RECT 16.745 5.95 16.915 7.14 ;
      RECT 14.895 2.635 15.065 3.865 ;
      RECT 14.95 0.855 15.12 2.805 ;
      RECT 14.895 0.575 15.065 1.025 ;
      RECT 14.895 7.855 15.065 8.305 ;
      RECT 14.95 6.075 15.12 8.025 ;
      RECT 14.895 5.015 15.065 6.245 ;
      RECT 14.375 0.575 14.545 3.865 ;
      RECT 14.375 2.075 14.78 2.405 ;
      RECT 14.375 1.235 14.78 1.565 ;
      RECT 14.375 5.015 14.545 8.305 ;
      RECT 14.375 7.315 14.78 7.645 ;
      RECT 14.375 6.475 14.78 6.805 ;
      RECT 11.71 1.975 12.44 2.215 ;
      RECT 12.252 1.77 12.44 2.215 ;
      RECT 12.08 1.782 12.455 2.209 ;
      RECT 11.995 1.797 12.475 2.194 ;
      RECT 11.995 1.812 12.48 2.184 ;
      RECT 11.95 1.832 12.495 2.176 ;
      RECT 11.927 1.867 12.51 2.13 ;
      RECT 11.841 1.89 12.515 2.09 ;
      RECT 11.841 1.908 12.525 2.06 ;
      RECT 11.71 1.977 12.53 2.023 ;
      RECT 11.755 1.92 12.525 2.06 ;
      RECT 11.841 1.872 12.51 2.13 ;
      RECT 11.927 1.841 12.495 2.176 ;
      RECT 11.95 1.822 12.48 2.184 ;
      RECT 11.995 1.795 12.455 2.209 ;
      RECT 12.08 1.777 12.44 2.215 ;
      RECT 12.166 1.771 12.44 2.215 ;
      RECT 12.252 1.766 12.385 2.215 ;
      RECT 12.338 1.761 12.385 2.215 ;
      RECT 12.03 2.659 12.2 3.045 ;
      RECT 12.025 2.659 12.2 3.04 ;
      RECT 12 2.659 12.2 3.005 ;
      RECT 12 2.687 12.21 2.995 ;
      RECT 11.98 2.687 12.21 2.955 ;
      RECT 11.975 2.687 12.21 2.928 ;
      RECT 11.975 2.705 12.215 2.92 ;
      RECT 11.92 2.705 12.215 2.855 ;
      RECT 11.92 2.722 12.225 2.838 ;
      RECT 11.91 2.722 12.225 2.778 ;
      RECT 11.91 2.739 12.23 2.775 ;
      RECT 11.905 2.575 12.075 2.753 ;
      RECT 11.905 2.609 12.161 2.753 ;
      RECT 11.9 3.375 11.905 3.388 ;
      RECT 11.895 3.27 11.9 3.393 ;
      RECT 11.87 3.13 11.895 3.408 ;
      RECT 11.835 3.081 11.87 3.44 ;
      RECT 11.83 3.049 11.835 3.46 ;
      RECT 11.825 3.04 11.83 3.46 ;
      RECT 11.745 3.005 11.825 3.46 ;
      RECT 11.682 2.975 11.745 3.46 ;
      RECT 11.596 2.963 11.682 3.46 ;
      RECT 11.51 2.949 11.596 3.46 ;
      RECT 11.43 2.936 11.51 3.446 ;
      RECT 11.395 2.928 11.43 3.426 ;
      RECT 11.385 2.925 11.395 3.417 ;
      RECT 11.355 2.92 11.385 3.404 ;
      RECT 11.305 2.895 11.355 3.38 ;
      RECT 11.291 2.869 11.305 3.362 ;
      RECT 11.205 2.829 11.291 3.338 ;
      RECT 11.16 2.777 11.205 3.307 ;
      RECT 11.15 2.752 11.16 3.294 ;
      RECT 11.145 2.533 11.15 2.555 ;
      RECT 11.14 2.735 11.15 3.29 ;
      RECT 11.14 2.531 11.145 2.645 ;
      RECT 11.13 2.527 11.14 3.286 ;
      RECT 11.086 2.525 11.13 3.274 ;
      RECT 11 2.525 11.086 3.245 ;
      RECT 10.97 2.525 11 3.218 ;
      RECT 10.955 2.525 10.97 3.206 ;
      RECT 10.915 2.537 10.955 3.191 ;
      RECT 10.895 2.556 10.915 3.17 ;
      RECT 10.885 2.566 10.895 3.154 ;
      RECT 10.875 2.572 10.885 3.143 ;
      RECT 10.855 2.582 10.875 3.126 ;
      RECT 10.85 2.591 10.855 3.113 ;
      RECT 10.845 2.595 10.85 3.063 ;
      RECT 10.835 2.601 10.845 2.98 ;
      RECT 10.83 2.605 10.835 2.894 ;
      RECT 10.825 2.625 10.83 2.831 ;
      RECT 10.82 2.648 10.825 2.778 ;
      RECT 10.815 2.666 10.82 2.723 ;
      RECT 11.425 2.485 11.595 2.745 ;
      RECT 11.595 2.45 11.64 2.731 ;
      RECT 11.556 2.452 11.645 2.714 ;
      RECT 11.445 2.469 11.731 2.685 ;
      RECT 11.445 2.484 11.735 2.657 ;
      RECT 11.445 2.465 11.645 2.714 ;
      RECT 11.47 2.453 11.595 2.745 ;
      RECT 11.556 2.451 11.64 2.731 ;
      RECT 10.61 1.84 10.78 2.33 ;
      RECT 10.61 1.84 10.815 2.31 ;
      RECT 10.745 1.76 10.855 2.27 ;
      RECT 10.726 1.764 10.875 2.24 ;
      RECT 10.64 1.772 10.895 2.223 ;
      RECT 10.64 1.778 10.9 2.213 ;
      RECT 10.64 1.787 10.92 2.201 ;
      RECT 10.615 1.812 10.95 2.179 ;
      RECT 10.615 1.832 10.955 2.159 ;
      RECT 10.61 1.845 10.965 2.139 ;
      RECT 10.61 1.912 10.97 2.12 ;
      RECT 10.61 2.045 10.975 2.107 ;
      RECT 10.605 1.85 10.965 1.94 ;
      RECT 10.615 1.807 10.92 2.201 ;
      RECT 10.726 1.762 10.855 2.27 ;
      RECT 10.6 3.515 10.9 3.77 ;
      RECT 10.685 3.481 10.9 3.77 ;
      RECT 10.685 3.484 10.905 3.63 ;
      RECT 10.62 3.505 10.905 3.63 ;
      RECT 10.655 3.495 10.9 3.77 ;
      RECT 10.65 3.5 10.905 3.63 ;
      RECT 10.685 3.479 10.886 3.77 ;
      RECT 10.771 3.47 10.886 3.77 ;
      RECT 10.771 3.464 10.8 3.77 ;
      RECT 10.26 3.105 10.27 3.595 ;
      RECT 9.92 3.04 9.93 3.34 ;
      RECT 10.435 3.212 10.44 3.431 ;
      RECT 10.425 3.192 10.435 3.448 ;
      RECT 10.415 3.172 10.425 3.478 ;
      RECT 10.41 3.162 10.415 3.493 ;
      RECT 10.405 3.158 10.41 3.498 ;
      RECT 10.39 3.15 10.405 3.505 ;
      RECT 10.35 3.13 10.39 3.53 ;
      RECT 10.325 3.112 10.35 3.563 ;
      RECT 10.32 3.11 10.325 3.576 ;
      RECT 10.3 3.107 10.32 3.58 ;
      RECT 10.27 3.105 10.3 3.59 ;
      RECT 10.2 3.107 10.26 3.591 ;
      RECT 10.18 3.107 10.2 3.585 ;
      RECT 10.155 3.105 10.18 3.582 ;
      RECT 10.12 3.1 10.155 3.578 ;
      RECT 10.1 3.094 10.12 3.565 ;
      RECT 10.09 3.091 10.1 3.553 ;
      RECT 10.07 3.088 10.09 3.538 ;
      RECT 10.05 3.084 10.07 3.52 ;
      RECT 10.045 3.081 10.05 3.51 ;
      RECT 10.04 3.08 10.045 3.508 ;
      RECT 10.03 3.077 10.04 3.5 ;
      RECT 10.02 3.071 10.03 3.483 ;
      RECT 10.01 3.065 10.02 3.465 ;
      RECT 10 3.059 10.01 3.453 ;
      RECT 9.99 3.053 10 3.433 ;
      RECT 9.985 3.049 9.99 3.418 ;
      RECT 9.98 3.047 9.985 3.41 ;
      RECT 9.975 3.045 9.98 3.403 ;
      RECT 9.97 3.043 9.975 3.393 ;
      RECT 9.965 3.041 9.97 3.387 ;
      RECT 9.955 3.04 9.965 3.377 ;
      RECT 9.945 3.04 9.955 3.368 ;
      RECT 9.93 3.04 9.945 3.353 ;
      RECT 9.89 3.04 9.92 3.337 ;
      RECT 9.87 3.042 9.89 3.332 ;
      RECT 9.865 3.047 9.87 3.33 ;
      RECT 9.835 3.055 9.865 3.328 ;
      RECT 9.805 3.07 9.835 3.327 ;
      RECT 9.76 3.092 9.805 3.332 ;
      RECT 9.755 3.107 9.76 3.336 ;
      RECT 9.74 3.112 9.755 3.338 ;
      RECT 9.735 3.116 9.74 3.34 ;
      RECT 9.675 3.139 9.735 3.349 ;
      RECT 9.655 3.165 9.675 3.362 ;
      RECT 9.645 3.172 9.655 3.366 ;
      RECT 9.63 3.179 9.645 3.369 ;
      RECT 9.61 3.189 9.63 3.372 ;
      RECT 9.605 3.197 9.61 3.375 ;
      RECT 9.56 3.202 9.605 3.382 ;
      RECT 9.55 3.205 9.56 3.389 ;
      RECT 9.54 3.205 9.55 3.393 ;
      RECT 9.505 3.207 9.54 3.405 ;
      RECT 9.485 3.21 9.505 3.418 ;
      RECT 9.445 3.213 9.485 3.429 ;
      RECT 9.43 3.215 9.445 3.442 ;
      RECT 9.42 3.215 9.43 3.447 ;
      RECT 9.395 3.216 9.42 3.455 ;
      RECT 9.385 3.218 9.395 3.46 ;
      RECT 9.38 3.219 9.385 3.463 ;
      RECT 9.355 3.217 9.38 3.466 ;
      RECT 9.34 3.215 9.355 3.467 ;
      RECT 9.32 3.212 9.34 3.469 ;
      RECT 9.3 3.207 9.32 3.469 ;
      RECT 9.24 3.202 9.3 3.466 ;
      RECT 9.205 3.177 9.24 3.462 ;
      RECT 9.195 3.154 9.205 3.46 ;
      RECT 9.165 3.131 9.195 3.46 ;
      RECT 9.155 3.11 9.165 3.46 ;
      RECT 9.13 3.092 9.155 3.458 ;
      RECT 9.115 3.07 9.13 3.455 ;
      RECT 9.1 3.052 9.115 3.453 ;
      RECT 9.08 3.042 9.1 3.451 ;
      RECT 9.065 3.037 9.08 3.45 ;
      RECT 9.05 3.035 9.065 3.449 ;
      RECT 9.02 3.036 9.05 3.447 ;
      RECT 9 3.039 9.02 3.445 ;
      RECT 8.943 3.043 9 3.445 ;
      RECT 8.857 3.052 8.943 3.445 ;
      RECT 8.771 3.063 8.857 3.445 ;
      RECT 8.685 3.074 8.771 3.445 ;
      RECT 8.665 3.081 8.685 3.453 ;
      RECT 8.655 3.084 8.665 3.46 ;
      RECT 8.59 3.089 8.655 3.478 ;
      RECT 8.56 3.096 8.59 3.503 ;
      RECT 8.55 3.099 8.56 3.51 ;
      RECT 8.505 3.103 8.55 3.515 ;
      RECT 8.475 3.108 8.505 3.52 ;
      RECT 8.474 3.11 8.475 3.52 ;
      RECT 8.388 3.116 8.474 3.52 ;
      RECT 8.302 3.127 8.388 3.52 ;
      RECT 8.216 3.139 8.302 3.52 ;
      RECT 8.13 3.15 8.216 3.52 ;
      RECT 8.115 3.157 8.13 3.515 ;
      RECT 8.11 3.159 8.115 3.509 ;
      RECT 8.09 3.17 8.11 3.504 ;
      RECT 8.08 3.188 8.09 3.498 ;
      RECT 8.075 3.2 8.08 3.298 ;
      RECT 10.37 1.953 10.39 2.04 ;
      RECT 10.365 1.888 10.37 2.072 ;
      RECT 10.355 1.855 10.365 2.077 ;
      RECT 10.35 1.835 10.355 2.083 ;
      RECT 10.32 1.835 10.35 2.1 ;
      RECT 10.271 1.835 10.32 2.136 ;
      RECT 10.185 1.835 10.271 2.194 ;
      RECT 10.156 1.845 10.185 2.243 ;
      RECT 10.07 1.887 10.156 2.296 ;
      RECT 10.05 1.925 10.07 2.343 ;
      RECT 10.025 1.942 10.05 2.363 ;
      RECT 10.015 1.956 10.025 2.383 ;
      RECT 10.01 1.962 10.015 2.393 ;
      RECT 10.005 1.966 10.01 2.4 ;
      RECT 9.955 1.986 10.005 2.405 ;
      RECT 9.89 2.03 9.955 2.405 ;
      RECT 9.865 2.08 9.89 2.405 ;
      RECT 9.855 2.11 9.865 2.405 ;
      RECT 9.85 2.137 9.855 2.405 ;
      RECT 9.845 2.155 9.85 2.405 ;
      RECT 9.835 2.197 9.845 2.405 ;
      RECT 10.185 2.755 10.355 2.93 ;
      RECT 10.125 2.583 10.185 2.918 ;
      RECT 10.115 2.576 10.125 2.901 ;
      RECT 10.07 2.755 10.355 2.881 ;
      RECT 10.051 2.755 10.355 2.859 ;
      RECT 9.965 2.755 10.355 2.824 ;
      RECT 9.945 2.575 10.115 2.78 ;
      RECT 9.945 2.722 10.35 2.78 ;
      RECT 9.945 2.67 10.325 2.78 ;
      RECT 9.945 2.625 10.29 2.78 ;
      RECT 9.945 2.607 10.255 2.78 ;
      RECT 9.945 2.597 10.25 2.78 ;
      RECT 9.595 5.015 9.765 8.305 ;
      RECT 9.595 7.315 10 7.645 ;
      RECT 9.595 6.475 10 6.805 ;
      RECT 9.665 3.555 9.855 3.78 ;
      RECT 9.655 3.556 9.86 3.775 ;
      RECT 9.655 3.558 9.87 3.755 ;
      RECT 9.655 3.562 9.875 3.74 ;
      RECT 9.655 3.549 9.825 3.775 ;
      RECT 9.655 3.552 9.85 3.775 ;
      RECT 9.665 3.548 9.825 3.78 ;
      RECT 9.751 3.546 9.825 3.78 ;
      RECT 9.375 2.797 9.545 3.035 ;
      RECT 9.375 2.797 9.631 2.949 ;
      RECT 9.375 2.797 9.635 2.859 ;
      RECT 9.425 2.57 9.645 2.838 ;
      RECT 9.42 2.587 9.65 2.811 ;
      RECT 9.385 2.745 9.65 2.811 ;
      RECT 9.405 2.595 9.545 3.035 ;
      RECT 9.395 2.677 9.655 2.794 ;
      RECT 9.39 2.725 9.655 2.794 ;
      RECT 9.395 2.635 9.65 2.811 ;
      RECT 9.42 2.572 9.645 2.838 ;
      RECT 8.985 2.547 9.155 2.745 ;
      RECT 8.985 2.547 9.2 2.72 ;
      RECT 9.055 2.49 9.225 2.678 ;
      RECT 9.03 2.505 9.225 2.678 ;
      RECT 8.645 2.551 8.675 2.745 ;
      RECT 8.64 2.523 8.645 2.745 ;
      RECT 8.61 2.497 8.64 2.747 ;
      RECT 8.585 2.455 8.61 2.75 ;
      RECT 8.575 2.427 8.585 2.752 ;
      RECT 8.54 2.407 8.575 2.754 ;
      RECT 8.475 2.392 8.54 2.76 ;
      RECT 8.425 2.39 8.475 2.766 ;
      RECT 8.402 2.392 8.425 2.771 ;
      RECT 8.316 2.403 8.402 2.777 ;
      RECT 8.23 2.421 8.316 2.787 ;
      RECT 8.215 2.432 8.23 2.793 ;
      RECT 8.145 2.455 8.215 2.799 ;
      RECT 8.09 2.487 8.145 2.807 ;
      RECT 8.05 2.51 8.09 2.813 ;
      RECT 8.036 2.523 8.05 2.816 ;
      RECT 7.95 2.545 8.036 2.822 ;
      RECT 7.935 2.57 7.95 2.828 ;
      RECT 7.895 2.585 7.935 2.832 ;
      RECT 7.845 2.6 7.895 2.837 ;
      RECT 7.82 2.607 7.845 2.841 ;
      RECT 7.76 2.602 7.82 2.845 ;
      RECT 7.745 2.593 7.76 2.849 ;
      RECT 7.675 2.583 7.745 2.845 ;
      RECT 7.65 2.575 7.67 2.835 ;
      RECT 7.591 2.575 7.65 2.813 ;
      RECT 7.505 2.575 7.591 2.77 ;
      RECT 7.67 2.575 7.675 2.84 ;
      RECT 8.365 1.806 8.535 2.14 ;
      RECT 8.335 1.806 8.535 2.135 ;
      RECT 8.275 1.773 8.335 2.123 ;
      RECT 8.275 1.829 8.545 2.118 ;
      RECT 8.25 1.829 8.545 2.112 ;
      RECT 8.245 1.77 8.275 2.109 ;
      RECT 8.23 1.776 8.365 2.107 ;
      RECT 8.225 1.784 8.45 2.095 ;
      RECT 8.225 1.836 8.56 2.048 ;
      RECT 8.21 1.792 8.45 2.043 ;
      RECT 8.21 1.862 8.57 1.984 ;
      RECT 8.18 1.812 8.535 1.945 ;
      RECT 8.18 1.902 8.58 1.941 ;
      RECT 8.23 1.781 8.45 2.107 ;
      RECT 7.57 2.111 7.625 2.375 ;
      RECT 7.57 2.111 7.69 2.374 ;
      RECT 7.57 2.111 7.715 2.373 ;
      RECT 7.57 2.111 7.78 2.372 ;
      RECT 7.715 2.077 7.795 2.371 ;
      RECT 7.53 2.121 7.94 2.37 ;
      RECT 7.57 2.118 7.94 2.37 ;
      RECT 7.53 2.126 7.945 2.363 ;
      RECT 7.515 2.128 7.945 2.362 ;
      RECT 7.515 2.135 7.95 2.358 ;
      RECT 7.495 2.134 7.945 2.354 ;
      RECT 7.495 2.142 7.955 2.353 ;
      RECT 7.49 2.139 7.95 2.349 ;
      RECT 7.49 2.152 7.965 2.348 ;
      RECT 7.475 2.142 7.955 2.347 ;
      RECT 7.44 2.155 7.965 2.34 ;
      RECT 7.625 2.11 7.935 2.37 ;
      RECT 7.625 2.095 7.885 2.37 ;
      RECT 7.69 2.082 7.82 2.37 ;
      RECT 7.235 3.171 7.25 3.564 ;
      RECT 7.2 3.176 7.25 3.563 ;
      RECT 7.235 3.175 7.295 3.562 ;
      RECT 7.18 3.186 7.295 3.561 ;
      RECT 7.195 3.182 7.295 3.561 ;
      RECT 7.16 3.192 7.37 3.558 ;
      RECT 7.16 3.211 7.415 3.556 ;
      RECT 7.16 3.218 7.42 3.553 ;
      RECT 7.145 3.195 7.37 3.55 ;
      RECT 7.125 3.2 7.37 3.543 ;
      RECT 7.12 3.204 7.37 3.539 ;
      RECT 7.12 3.221 7.43 3.538 ;
      RECT 7.1 3.215 7.415 3.534 ;
      RECT 7.1 3.224 7.435 3.528 ;
      RECT 7.095 3.23 7.435 3.3 ;
      RECT 7.16 3.19 7.295 3.558 ;
      RECT 7.035 2.553 7.235 2.865 ;
      RECT 7.11 2.531 7.235 2.865 ;
      RECT 7.05 2.55 7.24 2.85 ;
      RECT 7.02 2.561 7.24 2.848 ;
      RECT 7.035 2.556 7.245 2.814 ;
      RECT 7.02 2.66 7.25 2.781 ;
      RECT 7.05 2.532 7.235 2.865 ;
      RECT 7.11 2.51 7.21 2.865 ;
      RECT 7.135 2.507 7.21 2.865 ;
      RECT 7.135 2.502 7.155 2.865 ;
      RECT 6.54 2.57 6.715 2.745 ;
      RECT 6.535 2.57 6.715 2.743 ;
      RECT 6.51 2.57 6.715 2.738 ;
      RECT 6.455 2.55 6.625 2.728 ;
      RECT 6.455 2.557 6.69 2.728 ;
      RECT 6.54 3.237 6.555 3.42 ;
      RECT 6.53 3.215 6.54 3.42 ;
      RECT 6.515 3.195 6.53 3.42 ;
      RECT 6.505 3.17 6.515 3.42 ;
      RECT 6.475 3.135 6.505 3.42 ;
      RECT 6.44 3.075 6.475 3.42 ;
      RECT 6.435 3.037 6.44 3.42 ;
      RECT 6.385 2.988 6.435 3.42 ;
      RECT 6.375 2.938 6.385 3.408 ;
      RECT 6.36 2.917 6.375 3.368 ;
      RECT 6.34 2.885 6.36 3.318 ;
      RECT 6.315 2.841 6.34 3.258 ;
      RECT 6.31 2.813 6.315 3.213 ;
      RECT 6.305 2.804 6.31 3.199 ;
      RECT 6.3 2.797 6.305 3.186 ;
      RECT 6.295 2.792 6.3 3.175 ;
      RECT 6.29 2.777 6.295 3.165 ;
      RECT 6.285 2.755 6.29 3.152 ;
      RECT 6.275 2.715 6.285 3.127 ;
      RECT 6.25 2.645 6.275 3.083 ;
      RECT 6.245 2.585 6.25 3.048 ;
      RECT 6.23 2.565 6.245 3.015 ;
      RECT 6.225 2.565 6.23 2.99 ;
      RECT 6.195 2.565 6.225 2.945 ;
      RECT 6.15 2.565 6.195 2.885 ;
      RECT 6.075 2.565 6.15 2.833 ;
      RECT 6.07 2.565 6.075 2.798 ;
      RECT 6.065 2.565 6.07 2.788 ;
      RECT 6.06 2.565 6.065 2.768 ;
      RECT 6.325 1.785 6.495 2.255 ;
      RECT 6.27 1.778 6.465 2.239 ;
      RECT 6.27 1.792 6.5 2.238 ;
      RECT 6.255 1.793 6.5 2.219 ;
      RECT 6.25 1.811 6.5 2.205 ;
      RECT 6.255 1.794 6.505 2.203 ;
      RECT 6.24 1.825 6.505 2.188 ;
      RECT 6.255 1.8 6.51 2.173 ;
      RECT 6.235 1.84 6.51 2.17 ;
      RECT 6.25 1.812 6.515 2.155 ;
      RECT 6.25 1.824 6.52 2.135 ;
      RECT 6.235 1.84 6.525 2.118 ;
      RECT 6.235 1.85 6.53 1.973 ;
      RECT 6.23 1.85 6.53 1.93 ;
      RECT 6.23 1.865 6.535 1.908 ;
      RECT 6.325 1.775 6.465 2.255 ;
      RECT 6.325 1.773 6.435 2.255 ;
      RECT 6.411 1.77 6.435 2.255 ;
      RECT 6.07 3.437 6.075 3.483 ;
      RECT 6.06 3.285 6.07 3.507 ;
      RECT 6.055 3.13 6.06 3.532 ;
      RECT 6.04 3.092 6.055 3.543 ;
      RECT 6.035 3.075 6.04 3.55 ;
      RECT 6.025 3.063 6.035 3.557 ;
      RECT 6.02 3.054 6.025 3.559 ;
      RECT 6.015 3.052 6.02 3.563 ;
      RECT 5.97 3.043 6.015 3.578 ;
      RECT 5.965 3.035 5.97 3.592 ;
      RECT 5.96 3.032 5.965 3.596 ;
      RECT 5.945 3.027 5.96 3.604 ;
      RECT 5.89 3.017 5.945 3.615 ;
      RECT 5.855 3.005 5.89 3.616 ;
      RECT 5.846 3 5.855 3.61 ;
      RECT 5.76 3 5.846 3.6 ;
      RECT 5.73 3 5.76 3.578 ;
      RECT 5.72 3 5.725 3.558 ;
      RECT 5.715 3 5.72 3.52 ;
      RECT 5.71 3 5.715 3.478 ;
      RECT 5.705 3 5.71 3.438 ;
      RECT 5.7 3 5.705 3.368 ;
      RECT 5.69 3 5.7 3.29 ;
      RECT 5.685 3 5.69 3.19 ;
      RECT 5.725 3 5.73 3.56 ;
      RECT 5.22 3.082 5.31 3.56 ;
      RECT 5.205 3.085 5.325 3.558 ;
      RECT 5.22 3.084 5.325 3.558 ;
      RECT 5.185 3.091 5.35 3.548 ;
      RECT 5.205 3.085 5.35 3.548 ;
      RECT 5.17 3.097 5.35 3.536 ;
      RECT 5.205 3.088 5.4 3.529 ;
      RECT 5.156 3.105 5.4 3.527 ;
      RECT 5.185 3.095 5.41 3.515 ;
      RECT 5.156 3.116 5.44 3.506 ;
      RECT 5.07 3.14 5.44 3.5 ;
      RECT 5.07 3.153 5.48 3.483 ;
      RECT 5.065 3.175 5.48 3.476 ;
      RECT 5.035 3.19 5.48 3.466 ;
      RECT 5.03 3.201 5.48 3.456 ;
      RECT 5 3.214 5.48 3.447 ;
      RECT 4.985 3.232 5.48 3.436 ;
      RECT 4.96 3.245 5.48 3.426 ;
      RECT 5.22 3.081 5.23 3.56 ;
      RECT 5.266 2.505 5.305 2.75 ;
      RECT 5.18 2.505 5.315 2.748 ;
      RECT 5.065 2.53 5.315 2.745 ;
      RECT 5.065 2.53 5.32 2.743 ;
      RECT 5.065 2.53 5.335 2.738 ;
      RECT 5.171 2.505 5.35 2.718 ;
      RECT 5.085 2.513 5.35 2.718 ;
      RECT 4.755 1.865 4.925 2.3 ;
      RECT 4.745 1.899 4.925 2.283 ;
      RECT 4.825 1.835 4.995 2.27 ;
      RECT 4.73 1.91 4.995 2.248 ;
      RECT 4.825 1.845 5 2.238 ;
      RECT 4.755 1.897 5.03 2.223 ;
      RECT 4.715 1.923 5.03 2.208 ;
      RECT 4.715 1.965 5.04 2.188 ;
      RECT 4.71 1.99 5.045 2.17 ;
      RECT 4.71 2 5.05 2.155 ;
      RECT 4.705 1.937 5.03 2.153 ;
      RECT 4.705 2.01 5.055 2.138 ;
      RECT 4.7 1.947 5.03 2.135 ;
      RECT 4.695 2.031 5.06 2.118 ;
      RECT 4.695 2.063 5.065 2.098 ;
      RECT 4.69 1.977 5.04 2.09 ;
      RECT 4.695 1.962 5.03 2.118 ;
      RECT 4.71 1.932 5.03 2.17 ;
      RECT 4.555 2.519 4.78 2.775 ;
      RECT 4.555 2.552 4.8 2.765 ;
      RECT 4.52 2.552 4.8 2.763 ;
      RECT 4.52 2.565 4.805 2.753 ;
      RECT 4.52 2.585 4.815 2.745 ;
      RECT 4.52 2.682 4.82 2.738 ;
      RECT 4.5 2.43 4.63 2.728 ;
      RECT 4.455 2.585 4.815 2.67 ;
      RECT 4.445 2.43 4.63 2.615 ;
      RECT 4.445 2.462 4.716 2.615 ;
      RECT 4.41 2.992 4.43 3.17 ;
      RECT 4.375 2.945 4.41 3.17 ;
      RECT 4.36 2.885 4.375 3.17 ;
      RECT 4.335 2.832 4.36 3.17 ;
      RECT 4.32 2.785 4.335 3.17 ;
      RECT 4.3 2.762 4.32 3.17 ;
      RECT 4.275 2.727 4.3 3.17 ;
      RECT 4.265 2.573 4.275 3.17 ;
      RECT 4.235 2.568 4.265 3.161 ;
      RECT 4.23 2.565 4.235 3.151 ;
      RECT 4.215 2.565 4.23 3.125 ;
      RECT 4.21 2.565 4.215 3.088 ;
      RECT 4.185 2.565 4.21 3.04 ;
      RECT 4.165 2.565 4.185 2.965 ;
      RECT 4.155 2.565 4.165 2.925 ;
      RECT 4.15 2.565 4.155 2.9 ;
      RECT 4.145 2.565 4.15 2.883 ;
      RECT 4.14 2.565 4.145 2.865 ;
      RECT 4.135 2.566 4.14 2.855 ;
      RECT 4.125 2.568 4.135 2.823 ;
      RECT 4.115 2.57 4.125 2.79 ;
      RECT 4.105 2.573 4.115 2.763 ;
      RECT 4.43 3 4.655 3.17 ;
      RECT 3.76 1.812 3.93 2.265 ;
      RECT 3.76 1.812 4.02 2.231 ;
      RECT 3.76 1.812 4.05 2.215 ;
      RECT 3.76 1.812 4.08 2.188 ;
      RECT 4.016 1.79 4.095 2.17 ;
      RECT 3.795 1.797 4.1 2.155 ;
      RECT 3.795 1.805 4.11 2.118 ;
      RECT 3.755 1.832 4.11 2.09 ;
      RECT 3.74 1.845 4.11 2.055 ;
      RECT 3.76 1.82 4.13 2.045 ;
      RECT 3.735 1.885 4.13 2.015 ;
      RECT 3.735 1.915 4.135 1.998 ;
      RECT 3.73 1.945 4.135 1.985 ;
      RECT 3.795 1.794 4.095 2.17 ;
      RECT 3.93 1.791 4.016 2.249 ;
      RECT 3.881 1.792 4.095 2.17 ;
      RECT 4.025 3.452 4.07 3.645 ;
      RECT 4.015 3.422 4.025 3.645 ;
      RECT 4.01 3.407 4.015 3.645 ;
      RECT 3.97 3.317 4.01 3.645 ;
      RECT 3.965 3.23 3.97 3.645 ;
      RECT 3.955 3.2 3.965 3.645 ;
      RECT 3.95 3.16 3.955 3.645 ;
      RECT 3.94 3.122 3.95 3.645 ;
      RECT 3.935 3.087 3.94 3.645 ;
      RECT 3.915 3.04 3.935 3.645 ;
      RECT 3.9 2.965 3.915 3.645 ;
      RECT 3.895 2.92 3.9 3.64 ;
      RECT 3.89 2.9 3.895 3.613 ;
      RECT 3.885 2.88 3.89 3.598 ;
      RECT 3.88 2.855 3.885 3.578 ;
      RECT 3.875 2.833 3.88 3.563 ;
      RECT 3.87 2.811 3.875 3.545 ;
      RECT 3.865 2.79 3.87 3.535 ;
      RECT 3.855 2.762 3.865 3.505 ;
      RECT 3.845 2.725 3.855 3.473 ;
      RECT 3.835 2.685 3.845 3.44 ;
      RECT 3.825 2.663 3.835 3.41 ;
      RECT 3.795 2.615 3.825 3.342 ;
      RECT 3.78 2.575 3.795 3.269 ;
      RECT 3.77 2.575 3.78 3.235 ;
      RECT 3.765 2.575 3.77 3.21 ;
      RECT 3.76 2.575 3.765 3.195 ;
      RECT 3.755 2.575 3.76 3.173 ;
      RECT 3.75 2.575 3.755 3.16 ;
      RECT 3.735 2.575 3.75 3.125 ;
      RECT 3.715 2.575 3.735 3.065 ;
      RECT 3.705 2.575 3.715 3.015 ;
      RECT 3.685 2.575 3.705 2.963 ;
      RECT 3.665 2.575 3.685 2.92 ;
      RECT 3.655 2.575 3.665 2.908 ;
      RECT 3.625 2.575 3.655 2.895 ;
      RECT 3.595 2.596 3.625 2.875 ;
      RECT 3.585 2.624 3.595 2.855 ;
      RECT 3.57 2.641 3.585 2.823 ;
      RECT 3.565 2.655 3.57 2.79 ;
      RECT 3.56 2.663 3.565 2.763 ;
      RECT 3.555 2.671 3.56 2.725 ;
      RECT 3.56 3.195 3.565 3.53 ;
      RECT 3.525 3.182 3.56 3.529 ;
      RECT 3.455 3.122 3.525 3.528 ;
      RECT 3.375 3.065 3.455 3.527 ;
      RECT 3.24 3.025 3.375 3.526 ;
      RECT 3.24 3.212 3.575 3.515 ;
      RECT 3.2 3.212 3.575 3.505 ;
      RECT 3.2 3.23 3.58 3.5 ;
      RECT 3.2 3.32 3.585 3.49 ;
      RECT 3.195 3.015 3.36 3.47 ;
      RECT 3.19 3.015 3.36 3.213 ;
      RECT 3.19 3.172 3.555 3.213 ;
      RECT 3.19 3.16 3.55 3.213 ;
      RECT 1.18 7.855 1.35 8.305 ;
      RECT 1.235 6.075 1.405 8.025 ;
      RECT 1.18 5.015 1.35 6.245 ;
      RECT 0.66 5.015 0.83 8.305 ;
      RECT 0.66 7.315 1.065 7.645 ;
      RECT 0.66 6.475 1.065 6.805 ;
      RECT 81.23 7.8 81.4 8.31 ;
      RECT 80.24 0.57 80.41 1.08 ;
      RECT 80.24 2.39 80.41 3.86 ;
      RECT 80.24 5.02 80.41 6.49 ;
      RECT 80.24 7.8 80.41 8.31 ;
      RECT 78.88 0.575 79.05 3.865 ;
      RECT 78.88 5.015 79.05 8.305 ;
      RECT 78.45 0.575 78.62 1.085 ;
      RECT 78.45 1.655 78.62 3.865 ;
      RECT 78.45 5.015 78.62 7.225 ;
      RECT 78.45 7.795 78.62 8.305 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 74.1 5.015 74.27 8.305 ;
      RECT 73.67 5.015 73.84 7.225 ;
      RECT 73.67 7.795 73.84 8.305 ;
      RECT 65.445 7.8 65.615 8.31 ;
      RECT 64.455 0.57 64.625 1.08 ;
      RECT 64.455 2.39 64.625 3.86 ;
      RECT 64.455 5.02 64.625 6.49 ;
      RECT 64.455 7.8 64.625 8.31 ;
      RECT 63.095 0.575 63.265 3.865 ;
      RECT 63.095 5.015 63.265 8.305 ;
      RECT 62.665 0.575 62.835 1.085 ;
      RECT 62.665 1.655 62.835 3.865 ;
      RECT 62.665 5.015 62.835 7.225 ;
      RECT 62.665 7.795 62.835 8.305 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 58.315 5.015 58.485 8.305 ;
      RECT 57.885 5.015 58.055 7.225 ;
      RECT 57.885 7.795 58.055 8.305 ;
      RECT 49.66 7.8 49.83 8.31 ;
      RECT 48.67 0.57 48.84 1.08 ;
      RECT 48.67 2.39 48.84 3.86 ;
      RECT 48.67 5.02 48.84 6.49 ;
      RECT 48.67 7.8 48.84 8.31 ;
      RECT 47.31 0.575 47.48 3.865 ;
      RECT 47.31 5.015 47.48 8.305 ;
      RECT 46.88 0.575 47.05 1.085 ;
      RECT 46.88 1.655 47.05 3.865 ;
      RECT 46.88 5.015 47.05 7.225 ;
      RECT 46.88 7.795 47.05 8.305 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 42.53 5.015 42.7 8.305 ;
      RECT 42.1 5.015 42.27 7.225 ;
      RECT 42.1 7.795 42.27 8.305 ;
      RECT 33.885 7.8 34.055 8.31 ;
      RECT 32.895 0.57 33.065 1.08 ;
      RECT 32.895 2.39 33.065 3.86 ;
      RECT 32.895 5.02 33.065 6.49 ;
      RECT 32.895 7.8 33.065 8.31 ;
      RECT 31.535 0.575 31.705 3.865 ;
      RECT 31.535 5.015 31.705 8.305 ;
      RECT 31.105 0.575 31.275 1.085 ;
      RECT 31.105 1.655 31.275 3.865 ;
      RECT 31.105 5.015 31.275 7.225 ;
      RECT 31.105 7.795 31.275 8.305 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 26.755 5.015 26.925 8.305 ;
      RECT 26.325 5.015 26.495 7.225 ;
      RECT 26.325 7.795 26.495 8.305 ;
      RECT 18.105 7.8 18.275 8.31 ;
      RECT 17.115 0.57 17.285 1.08 ;
      RECT 17.115 2.39 17.285 3.86 ;
      RECT 17.115 5.02 17.285 6.49 ;
      RECT 17.115 7.8 17.285 8.31 ;
      RECT 15.755 0.575 15.925 3.865 ;
      RECT 15.755 5.015 15.925 8.305 ;
      RECT 15.325 0.575 15.495 1.085 ;
      RECT 15.325 1.655 15.495 3.865 ;
      RECT 15.325 5.015 15.495 7.225 ;
      RECT 15.325 7.795 15.495 8.305 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 10.975 5.015 11.145 8.305 ;
      RECT 10.545 5.015 10.715 7.225 ;
      RECT 10.545 7.795 10.715 8.305 ;
      RECT 1.61 5.015 1.78 7.225 ;
      RECT 1.61 7.795 1.78 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r2 ;
  SIZE 81.765 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 18.1 0.915 18.27 1.085 ;
        RECT 18.095 0.91 18.265 1.08 ;
        RECT 18.095 2.39 18.265 2.56 ;
      LAYER li1 ;
        RECT 18.1 0.915 18.27 1.085 ;
        RECT 18.095 0.57 18.265 1.08 ;
        RECT 18.095 2.39 18.265 3.86 ;
      LAYER met1 ;
        RECT 18.035 2.36 18.325 2.59 ;
        RECT 18.035 0.88 18.325 1.11 ;
        RECT 18.095 0.88 18.265 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 33.88 0.915 34.05 1.085 ;
        RECT 33.875 0.91 34.045 1.08 ;
        RECT 33.875 2.39 34.045 2.56 ;
      LAYER li1 ;
        RECT 33.88 0.915 34.05 1.085 ;
        RECT 33.875 0.57 34.045 1.08 ;
        RECT 33.875 2.39 34.045 3.86 ;
      LAYER met1 ;
        RECT 33.815 2.36 34.105 2.59 ;
        RECT 33.815 0.88 34.105 1.11 ;
        RECT 33.875 0.88 34.045 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 49.655 0.915 49.825 1.085 ;
        RECT 49.65 0.91 49.82 1.08 ;
        RECT 49.65 2.39 49.82 2.56 ;
      LAYER li1 ;
        RECT 49.655 0.915 49.825 1.085 ;
        RECT 49.65 0.57 49.82 1.08 ;
        RECT 49.65 2.39 49.82 3.86 ;
      LAYER met1 ;
        RECT 49.59 2.36 49.88 2.59 ;
        RECT 49.59 0.88 49.88 1.11 ;
        RECT 49.65 0.88 49.82 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 65.44 0.915 65.61 1.085 ;
        RECT 65.435 0.91 65.605 1.08 ;
        RECT 65.435 2.39 65.605 2.56 ;
      LAYER li1 ;
        RECT 65.44 0.915 65.61 1.085 ;
        RECT 65.435 0.57 65.605 1.08 ;
        RECT 65.435 2.39 65.605 3.86 ;
      LAYER met1 ;
        RECT 65.375 2.36 65.665 2.59 ;
        RECT 65.375 0.88 65.665 1.11 ;
        RECT 65.435 0.88 65.605 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 81.225 0.915 81.395 1.085 ;
        RECT 81.22 0.91 81.39 1.08 ;
        RECT 81.22 2.39 81.39 2.56 ;
      LAYER li1 ;
        RECT 81.225 0.915 81.395 1.085 ;
        RECT 81.22 0.57 81.39 1.08 ;
        RECT 81.22 2.39 81.39 3.86 ;
      LAYER met1 ;
        RECT 81.16 2.36 81.45 2.59 ;
        RECT 81.16 0.88 81.45 1.11 ;
        RECT 81.22 0.88 81.39 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 13.86 5.855 14.21 6.205 ;
        RECT 13.855 2.705 14.205 3.055 ;
        RECT 13.93 2.705 14.105 6.205 ;
      LAYER li1 ;
        RECT 13.945 1.66 14.115 2.935 ;
        RECT 13.945 5.945 14.115 7.22 ;
        RECT 9.165 5.945 9.335 7.22 ;
      LAYER met1 ;
        RECT 13.855 2.765 14.345 2.935 ;
        RECT 13.855 2.705 14.205 3.055 ;
        RECT 9.105 5.945 14.345 6.115 ;
        RECT 13.86 5.855 14.21 6.205 ;
        RECT 9.105 5.915 9.395 6.145 ;
      LAYER mcon ;
        RECT 9.165 5.945 9.335 6.115 ;
        RECT 13.945 5.945 14.115 6.115 ;
        RECT 13.945 2.765 14.115 2.935 ;
      LAYER via1 ;
        RECT 13.955 2.805 14.105 2.955 ;
        RECT 13.96 5.955 14.11 6.105 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 29.64 5.855 29.99 6.205 ;
        RECT 29.635 2.705 29.985 3.055 ;
        RECT 29.71 2.705 29.885 6.205 ;
      LAYER li1 ;
        RECT 29.725 1.66 29.895 2.935 ;
        RECT 29.725 5.945 29.895 7.22 ;
        RECT 24.945 5.945 25.115 7.22 ;
      LAYER met1 ;
        RECT 29.635 2.765 30.125 2.935 ;
        RECT 29.635 2.705 29.985 3.055 ;
        RECT 24.885 5.945 30.125 6.115 ;
        RECT 29.64 5.855 29.99 6.205 ;
        RECT 24.885 5.915 25.175 6.145 ;
      LAYER mcon ;
        RECT 24.945 5.945 25.115 6.115 ;
        RECT 29.725 5.945 29.895 6.115 ;
        RECT 29.725 2.765 29.895 2.935 ;
      LAYER via1 ;
        RECT 29.735 2.805 29.885 2.955 ;
        RECT 29.74 5.955 29.89 6.105 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 45.415 5.855 45.765 6.205 ;
        RECT 45.41 2.705 45.76 3.055 ;
        RECT 45.485 2.705 45.66 6.205 ;
      LAYER li1 ;
        RECT 45.5 1.66 45.67 2.935 ;
        RECT 45.5 5.945 45.67 7.22 ;
        RECT 40.72 5.945 40.89 7.22 ;
      LAYER met1 ;
        RECT 45.41 2.765 45.9 2.935 ;
        RECT 45.41 2.705 45.76 3.055 ;
        RECT 40.66 5.945 45.9 6.115 ;
        RECT 45.415 5.855 45.765 6.205 ;
        RECT 40.66 5.915 40.95 6.145 ;
      LAYER mcon ;
        RECT 40.72 5.945 40.89 6.115 ;
        RECT 45.5 5.945 45.67 6.115 ;
        RECT 45.5 2.765 45.67 2.935 ;
      LAYER via1 ;
        RECT 45.51 2.805 45.66 2.955 ;
        RECT 45.515 5.955 45.665 6.105 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 61.2 5.855 61.55 6.205 ;
        RECT 61.195 2.705 61.545 3.055 ;
        RECT 61.27 2.705 61.445 6.205 ;
      LAYER li1 ;
        RECT 61.285 1.66 61.455 2.935 ;
        RECT 61.285 5.945 61.455 7.22 ;
        RECT 56.505 5.945 56.675 7.22 ;
      LAYER met1 ;
        RECT 61.195 2.765 61.685 2.935 ;
        RECT 61.195 2.705 61.545 3.055 ;
        RECT 56.445 5.945 61.685 6.115 ;
        RECT 61.2 5.855 61.55 6.205 ;
        RECT 56.445 5.915 56.735 6.145 ;
      LAYER mcon ;
        RECT 56.505 5.945 56.675 6.115 ;
        RECT 61.285 5.945 61.455 6.115 ;
        RECT 61.285 2.765 61.455 2.935 ;
      LAYER via1 ;
        RECT 61.295 2.805 61.445 2.955 ;
        RECT 61.3 5.955 61.45 6.105 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 76.985 5.855 77.335 6.205 ;
        RECT 76.98 2.705 77.33 3.055 ;
        RECT 77.055 2.705 77.23 6.205 ;
      LAYER li1 ;
        RECT 77.07 1.66 77.24 2.935 ;
        RECT 77.07 5.945 77.24 7.22 ;
        RECT 72.29 5.945 72.46 7.22 ;
      LAYER met1 ;
        RECT 76.98 2.765 77.47 2.935 ;
        RECT 76.98 2.705 77.33 3.055 ;
        RECT 72.23 5.945 77.47 6.115 ;
        RECT 76.985 5.855 77.335 6.205 ;
        RECT 72.23 5.915 72.52 6.145 ;
      LAYER mcon ;
        RECT 72.29 5.945 72.46 6.115 ;
        RECT 77.07 5.945 77.24 6.115 ;
        RECT 77.07 2.765 77.24 2.935 ;
      LAYER via1 ;
        RECT 77.08 2.805 77.23 2.955 ;
        RECT 77.085 5.955 77.235 6.105 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 5.945 0.4 7.22 ;
      LAYER met1 ;
        RECT 0.17 5.945 0.63 6.115 ;
        RECT 0.17 5.915 0.46 6.145 ;
      LAYER mcon ;
        RECT 0.23 5.945 0.4 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.295 4.24 2.1 4.62 ;
      LAYER met2 ;
        RECT 1.485 4.24 1.865 4.62 ;
      LAYER li1 ;
        RECT 0 4.44 81.765 4.745 ;
        RECT 1.76 4.135 81.765 4.745 ;
        RECT 79.63 4.13 81.61 4.75 ;
        RECT 80.79 3.4 80.96 5.48 ;
        RECT 79.8 3.4 79.97 5.48 ;
        RECT 77.06 3.405 77.23 5.475 ;
        RECT 75.26 3.635 75.43 4.745 ;
        RECT 74.3 3.635 74.47 4.745 ;
        RECT 72.28 4.135 72.45 5.475 ;
        RECT 71.86 3.635 72.03 4.745 ;
        RECT 70.86 3.635 71.03 4.745 ;
        RECT 69.9 3.635 70.07 4.745 ;
        RECT 67.46 3.635 67.63 4.745 ;
        RECT 63.845 4.13 65.825 4.75 ;
        RECT 65.005 3.4 65.175 5.48 ;
        RECT 64.015 3.4 64.185 5.48 ;
        RECT 61.275 3.405 61.445 5.475 ;
        RECT 59.475 3.635 59.645 4.745 ;
        RECT 58.515 3.635 58.685 4.745 ;
        RECT 56.495 4.135 56.665 5.475 ;
        RECT 56.075 3.635 56.245 4.745 ;
        RECT 55.075 3.635 55.245 4.745 ;
        RECT 54.115 3.635 54.285 4.745 ;
        RECT 51.675 3.635 51.845 4.745 ;
        RECT 48.06 4.13 50.04 4.75 ;
        RECT 49.22 3.4 49.39 5.48 ;
        RECT 48.23 3.4 48.4 5.48 ;
        RECT 45.49 3.405 45.66 5.475 ;
        RECT 43.69 3.635 43.86 4.745 ;
        RECT 42.73 3.635 42.9 4.745 ;
        RECT 40.71 4.135 40.88 5.475 ;
        RECT 40.29 3.635 40.46 4.745 ;
        RECT 39.29 3.635 39.46 4.745 ;
        RECT 38.33 3.635 38.5 4.745 ;
        RECT 35.89 3.635 36.06 4.745 ;
        RECT 32.285 4.13 34.265 4.75 ;
        RECT 33.445 3.4 33.615 5.48 ;
        RECT 32.455 3.4 32.625 5.48 ;
        RECT 29.715 3.405 29.885 5.475 ;
        RECT 27.915 3.635 28.085 4.745 ;
        RECT 26.955 3.635 27.125 4.745 ;
        RECT 24.935 4.135 25.105 5.475 ;
        RECT 24.515 3.635 24.685 4.745 ;
        RECT 23.515 3.635 23.685 4.745 ;
        RECT 22.555 3.635 22.725 4.745 ;
        RECT 20.115 3.635 20.285 4.745 ;
        RECT 16.505 4.13 18.485 4.75 ;
        RECT 17.665 3.4 17.835 5.48 ;
        RECT 16.675 3.4 16.845 5.48 ;
        RECT 13.935 3.405 14.105 5.475 ;
        RECT 12.135 3.635 12.305 4.745 ;
        RECT 11.175 3.635 11.345 4.745 ;
        RECT 9.155 4.135 9.325 5.475 ;
        RECT 8.735 3.635 8.905 4.745 ;
        RECT 7.735 3.635 7.905 4.745 ;
        RECT 6.775 3.635 6.945 4.745 ;
        RECT 4.335 3.635 4.505 4.745 ;
        RECT 2.03 4.135 2.2 8.305 ;
        RECT 0 4.135 81.765 4.315 ;
        RECT 0 4.135 1.59 4.745 ;
        RECT 0.22 4.135 0.39 5.475 ;
      LAYER met1 ;
        RECT 71.855 4.135 81.765 4.745 ;
        RECT 79.63 4.13 81.61 4.75 ;
        RECT 66.17 3.98 75.83 4.74 ;
        RECT 56.07 4.135 71.47 4.745 ;
        RECT 63.845 4.13 65.825 4.75 ;
        RECT 50.385 3.98 60.045 4.74 ;
        RECT 40.285 4.135 55.685 4.745 ;
        RECT 48.06 4.13 50.04 4.75 ;
        RECT 34.6 3.98 44.26 4.74 ;
        RECT 24.51 4.135 39.9 4.745 ;
        RECT 32.285 4.13 34.265 4.75 ;
        RECT 18.825 3.98 28.485 4.74 ;
        RECT 8.73 4.135 24.125 4.745 ;
        RECT 16.505 4.13 18.485 4.75 ;
        RECT 3.045 3.98 12.705 4.74 ;
        RECT 0 4.135 8.345 4.745 ;
        RECT 1.97 6.655 2.26 6.885 ;
        RECT 1.8 6.685 2.26 6.855 ;
      LAYER via2 ;
        RECT 1.575 4.33 1.775 4.53 ;
      LAYER mcon ;
        RECT 2.03 6.685 2.2 6.855 ;
        RECT 2.34 4.545 2.51 4.715 ;
        RECT 3.19 4.135 3.36 4.305 ;
        RECT 3.65 4.135 3.82 4.305 ;
        RECT 4.11 4.135 4.28 4.305 ;
        RECT 4.57 4.135 4.74 4.305 ;
        RECT 5.03 4.135 5.2 4.305 ;
        RECT 5.49 4.135 5.66 4.305 ;
        RECT 5.95 4.135 6.12 4.305 ;
        RECT 6.41 4.135 6.58 4.305 ;
        RECT 6.87 4.135 7.04 4.305 ;
        RECT 7.33 4.135 7.5 4.305 ;
        RECT 7.79 4.135 7.96 4.305 ;
        RECT 8.25 4.135 8.42 4.305 ;
        RECT 8.71 4.135 8.88 4.305 ;
        RECT 9.17 4.135 9.34 4.305 ;
        RECT 9.63 4.135 9.8 4.305 ;
        RECT 10.09 4.135 10.26 4.305 ;
        RECT 10.55 4.135 10.72 4.305 ;
        RECT 11.01 4.135 11.18 4.305 ;
        RECT 11.275 4.545 11.445 4.715 ;
        RECT 11.47 4.135 11.64 4.305 ;
        RECT 11.93 4.135 12.1 4.305 ;
        RECT 12.39 4.135 12.56 4.305 ;
        RECT 16.055 4.545 16.225 4.715 ;
        RECT 16.055 4.165 16.225 4.335 ;
        RECT 16.755 4.55 16.925 4.72 ;
        RECT 16.755 4.16 16.925 4.33 ;
        RECT 17.745 4.55 17.915 4.72 ;
        RECT 17.745 4.16 17.915 4.33 ;
        RECT 18.97 4.135 19.14 4.305 ;
        RECT 19.43 4.135 19.6 4.305 ;
        RECT 19.89 4.135 20.06 4.305 ;
        RECT 20.35 4.135 20.52 4.305 ;
        RECT 20.81 4.135 20.98 4.305 ;
        RECT 21.27 4.135 21.44 4.305 ;
        RECT 21.73 4.135 21.9 4.305 ;
        RECT 22.19 4.135 22.36 4.305 ;
        RECT 22.65 4.135 22.82 4.305 ;
        RECT 23.11 4.135 23.28 4.305 ;
        RECT 23.57 4.135 23.74 4.305 ;
        RECT 24.03 4.135 24.2 4.305 ;
        RECT 24.49 4.135 24.66 4.305 ;
        RECT 24.95 4.135 25.12 4.305 ;
        RECT 25.41 4.135 25.58 4.305 ;
        RECT 25.87 4.135 26.04 4.305 ;
        RECT 26.33 4.135 26.5 4.305 ;
        RECT 26.79 4.135 26.96 4.305 ;
        RECT 27.055 4.545 27.225 4.715 ;
        RECT 27.25 4.135 27.42 4.305 ;
        RECT 27.71 4.135 27.88 4.305 ;
        RECT 28.17 4.135 28.34 4.305 ;
        RECT 31.835 4.545 32.005 4.715 ;
        RECT 31.835 4.165 32.005 4.335 ;
        RECT 32.535 4.55 32.705 4.72 ;
        RECT 32.535 4.16 32.705 4.33 ;
        RECT 33.525 4.55 33.695 4.72 ;
        RECT 33.525 4.16 33.695 4.33 ;
        RECT 34.745 4.135 34.915 4.305 ;
        RECT 35.205 4.135 35.375 4.305 ;
        RECT 35.665 4.135 35.835 4.305 ;
        RECT 36.125 4.135 36.295 4.305 ;
        RECT 36.585 4.135 36.755 4.305 ;
        RECT 37.045 4.135 37.215 4.305 ;
        RECT 37.505 4.135 37.675 4.305 ;
        RECT 37.965 4.135 38.135 4.305 ;
        RECT 38.425 4.135 38.595 4.305 ;
        RECT 38.885 4.135 39.055 4.305 ;
        RECT 39.345 4.135 39.515 4.305 ;
        RECT 39.805 4.135 39.975 4.305 ;
        RECT 40.265 4.135 40.435 4.305 ;
        RECT 40.725 4.135 40.895 4.305 ;
        RECT 41.185 4.135 41.355 4.305 ;
        RECT 41.645 4.135 41.815 4.305 ;
        RECT 42.105 4.135 42.275 4.305 ;
        RECT 42.565 4.135 42.735 4.305 ;
        RECT 42.83 4.545 43 4.715 ;
        RECT 43.025 4.135 43.195 4.305 ;
        RECT 43.485 4.135 43.655 4.305 ;
        RECT 43.945 4.135 44.115 4.305 ;
        RECT 47.61 4.545 47.78 4.715 ;
        RECT 47.61 4.165 47.78 4.335 ;
        RECT 48.31 4.55 48.48 4.72 ;
        RECT 48.31 4.16 48.48 4.33 ;
        RECT 49.3 4.55 49.47 4.72 ;
        RECT 49.3 4.16 49.47 4.33 ;
        RECT 50.53 4.135 50.7 4.305 ;
        RECT 50.99 4.135 51.16 4.305 ;
        RECT 51.45 4.135 51.62 4.305 ;
        RECT 51.91 4.135 52.08 4.305 ;
        RECT 52.37 4.135 52.54 4.305 ;
        RECT 52.83 4.135 53 4.305 ;
        RECT 53.29 4.135 53.46 4.305 ;
        RECT 53.75 4.135 53.92 4.305 ;
        RECT 54.21 4.135 54.38 4.305 ;
        RECT 54.67 4.135 54.84 4.305 ;
        RECT 55.13 4.135 55.3 4.305 ;
        RECT 55.59 4.135 55.76 4.305 ;
        RECT 56.05 4.135 56.22 4.305 ;
        RECT 56.51 4.135 56.68 4.305 ;
        RECT 56.97 4.135 57.14 4.305 ;
        RECT 57.43 4.135 57.6 4.305 ;
        RECT 57.89 4.135 58.06 4.305 ;
        RECT 58.35 4.135 58.52 4.305 ;
        RECT 58.615 4.545 58.785 4.715 ;
        RECT 58.81 4.135 58.98 4.305 ;
        RECT 59.27 4.135 59.44 4.305 ;
        RECT 59.73 4.135 59.9 4.305 ;
        RECT 63.395 4.545 63.565 4.715 ;
        RECT 63.395 4.165 63.565 4.335 ;
        RECT 64.095 4.55 64.265 4.72 ;
        RECT 64.095 4.16 64.265 4.33 ;
        RECT 65.085 4.55 65.255 4.72 ;
        RECT 65.085 4.16 65.255 4.33 ;
        RECT 66.315 4.135 66.485 4.305 ;
        RECT 66.775 4.135 66.945 4.305 ;
        RECT 67.235 4.135 67.405 4.305 ;
        RECT 67.695 4.135 67.865 4.305 ;
        RECT 68.155 4.135 68.325 4.305 ;
        RECT 68.615 4.135 68.785 4.305 ;
        RECT 69.075 4.135 69.245 4.305 ;
        RECT 69.535 4.135 69.705 4.305 ;
        RECT 69.995 4.135 70.165 4.305 ;
        RECT 70.455 4.135 70.625 4.305 ;
        RECT 70.915 4.135 71.085 4.305 ;
        RECT 71.375 4.135 71.545 4.305 ;
        RECT 71.835 4.135 72.005 4.305 ;
        RECT 72.295 4.135 72.465 4.305 ;
        RECT 72.755 4.135 72.925 4.305 ;
        RECT 73.215 4.135 73.385 4.305 ;
        RECT 73.675 4.135 73.845 4.305 ;
        RECT 74.135 4.135 74.305 4.305 ;
        RECT 74.4 4.545 74.57 4.715 ;
        RECT 74.595 4.135 74.765 4.305 ;
        RECT 75.055 4.135 75.225 4.305 ;
        RECT 75.515 4.135 75.685 4.305 ;
        RECT 79.18 4.545 79.35 4.715 ;
        RECT 79.18 4.165 79.35 4.335 ;
        RECT 79.88 4.55 80.05 4.72 ;
        RECT 79.88 4.16 80.05 4.33 ;
        RECT 80.87 4.55 81.04 4.72 ;
        RECT 80.87 4.16 81.04 4.33 ;
      LAYER via1 ;
        RECT 1.6 4.355 1.75 4.505 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 73.56 7.04 73.93 7.41 ;
      RECT 73.6 6.72 73.93 7.41 ;
      RECT 73.6 6.72 76.39 7.025 ;
      RECT 76.085 2.85 76.39 7.025 ;
      RECT 76.05 2.85 76.42 3.22 ;
      RECT 75.31 0.815 75.615 4.02 ;
      RECT 75.06 2.975 75.615 3.705 ;
      RECT 75.27 0.815 75.64 1.185 ;
      RECT 71.42 1.85 71.75 2.745 ;
      RECT 70.54 2.015 70.87 2.745 ;
      RECT 71.415 1.85 71.785 2.65 ;
      RECT 74.58 1.85 74.91 2.58 ;
      RECT 74.54 1.735 74.72 2.385 ;
      RECT 70.55 1.85 74.91 2.22 ;
      RECT 71.04 3.535 71.37 3.865 ;
      RECT 69.835 3.55 71.37 3.85 ;
      RECT 69.835 2.43 70.135 3.85 ;
      RECT 69.58 2.415 69.91 2.745 ;
      RECT 57.775 7.04 58.145 7.41 ;
      RECT 57.815 6.72 58.145 7.41 ;
      RECT 57.815 6.72 60.605 7.025 ;
      RECT 60.3 2.85 60.605 7.025 ;
      RECT 60.265 2.85 60.635 3.22 ;
      RECT 59.525 0.815 59.83 4.02 ;
      RECT 59.275 2.975 59.83 3.705 ;
      RECT 59.485 0.815 59.855 1.185 ;
      RECT 55.635 1.85 55.965 2.745 ;
      RECT 54.755 2.015 55.085 2.745 ;
      RECT 55.63 1.85 56 2.65 ;
      RECT 58.795 1.85 59.125 2.58 ;
      RECT 58.755 1.735 58.935 2.385 ;
      RECT 54.765 1.85 59.125 2.22 ;
      RECT 55.255 3.535 55.585 3.865 ;
      RECT 54.05 3.55 55.585 3.85 ;
      RECT 54.05 2.43 54.35 3.85 ;
      RECT 53.795 2.415 54.125 2.745 ;
      RECT 41.99 7.04 42.36 7.41 ;
      RECT 42.03 6.72 42.36 7.41 ;
      RECT 42.03 6.72 44.82 7.025 ;
      RECT 44.515 2.85 44.82 7.025 ;
      RECT 44.48 2.85 44.85 3.22 ;
      RECT 43.74 0.815 44.045 4.02 ;
      RECT 43.49 2.975 44.045 3.705 ;
      RECT 43.7 0.815 44.07 1.185 ;
      RECT 39.85 1.85 40.18 2.745 ;
      RECT 38.97 2.015 39.3 2.745 ;
      RECT 39.845 1.85 40.215 2.65 ;
      RECT 43.01 1.85 43.34 2.58 ;
      RECT 42.97 1.735 43.15 2.385 ;
      RECT 38.98 1.85 43.34 2.22 ;
      RECT 39.47 3.535 39.8 3.865 ;
      RECT 38.265 3.55 39.8 3.85 ;
      RECT 38.265 2.43 38.565 3.85 ;
      RECT 38.01 2.415 38.34 2.745 ;
      RECT 26.215 7.04 26.585 7.41 ;
      RECT 26.255 6.72 26.585 7.41 ;
      RECT 26.255 6.72 29.045 7.025 ;
      RECT 28.74 2.85 29.045 7.025 ;
      RECT 28.705 2.85 29.075 3.22 ;
      RECT 27.965 0.815 28.27 4.02 ;
      RECT 27.715 2.975 28.27 3.705 ;
      RECT 27.925 0.815 28.295 1.185 ;
      RECT 24.075 1.85 24.405 2.745 ;
      RECT 23.195 2.015 23.525 2.745 ;
      RECT 24.07 1.85 24.44 2.65 ;
      RECT 27.235 1.85 27.565 2.58 ;
      RECT 27.195 1.735 27.375 2.385 ;
      RECT 23.205 1.85 27.565 2.22 ;
      RECT 23.695 3.535 24.025 3.865 ;
      RECT 22.49 3.55 24.025 3.85 ;
      RECT 22.49 2.43 22.79 3.85 ;
      RECT 22.235 2.415 22.565 2.745 ;
      RECT 10.435 7.04 10.805 7.41 ;
      RECT 10.475 6.72 10.805 7.41 ;
      RECT 10.475 6.72 13.265 7.025 ;
      RECT 12.96 2.85 13.265 7.025 ;
      RECT 12.925 2.85 13.295 3.22 ;
      RECT 12.185 0.815 12.49 4.02 ;
      RECT 11.935 2.975 12.49 3.705 ;
      RECT 12.145 0.815 12.515 1.185 ;
      RECT 8.295 1.85 8.625 2.745 ;
      RECT 7.415 2.015 7.745 2.745 ;
      RECT 8.29 1.85 8.66 2.65 ;
      RECT 11.455 1.85 11.785 2.58 ;
      RECT 11.415 1.735 11.595 2.385 ;
      RECT 7.425 1.85 11.785 2.22 ;
      RECT 7.915 3.535 8.245 3.865 ;
      RECT 6.71 3.55 8.245 3.85 ;
      RECT 6.71 2.43 7.01 3.85 ;
      RECT 6.455 2.415 6.785 2.745 ;
      RECT 72.98 2.575 73.31 3.305 ;
      RECT 68.86 2.415 69.19 3.145 ;
      RECT 67.86 1.855 68.19 2.585 ;
      RECT 66.42 2.575 66.75 3.305 ;
      RECT 57.195 2.575 57.525 3.305 ;
      RECT 53.075 2.415 53.405 3.145 ;
      RECT 52.075 1.855 52.405 2.585 ;
      RECT 50.635 2.575 50.965 3.305 ;
      RECT 41.41 2.575 41.74 3.305 ;
      RECT 37.29 2.415 37.62 3.145 ;
      RECT 36.29 1.855 36.62 2.585 ;
      RECT 34.85 2.575 35.18 3.305 ;
      RECT 25.635 2.575 25.965 3.305 ;
      RECT 21.515 2.415 21.845 3.145 ;
      RECT 20.515 1.855 20.845 2.585 ;
      RECT 19.075 2.575 19.405 3.305 ;
      RECT 9.855 2.575 10.185 3.305 ;
      RECT 5.735 2.415 6.065 3.145 ;
      RECT 4.735 1.855 5.065 2.585 ;
      RECT 3.295 2.575 3.625 3.305 ;
      RECT 0 0 0.805 0.38 ;
      RECT 0 8.5 0.805 8.88 ;
    LAYER via2 ;
      RECT 76.135 2.935 76.335 3.135 ;
      RECT 75.355 0.9 75.555 1.1 ;
      RECT 75.125 3.04 75.325 3.24 ;
      RECT 74.645 2.315 74.845 2.515 ;
      RECT 73.645 7.125 73.845 7.325 ;
      RECT 73.045 3.04 73.245 3.24 ;
      RECT 71.485 2.48 71.685 2.68 ;
      RECT 71.105 3.6 71.305 3.8 ;
      RECT 70.605 2.48 70.805 2.68 ;
      RECT 69.645 2.48 69.845 2.68 ;
      RECT 68.925 2.48 69.125 2.68 ;
      RECT 67.925 1.92 68.125 2.12 ;
      RECT 66.485 3.04 66.685 3.24 ;
      RECT 60.35 2.935 60.55 3.135 ;
      RECT 59.57 0.9 59.77 1.1 ;
      RECT 59.34 3.04 59.54 3.24 ;
      RECT 58.86 2.315 59.06 2.515 ;
      RECT 57.86 7.125 58.06 7.325 ;
      RECT 57.26 3.04 57.46 3.24 ;
      RECT 55.7 2.48 55.9 2.68 ;
      RECT 55.32 3.6 55.52 3.8 ;
      RECT 54.82 2.48 55.02 2.68 ;
      RECT 53.86 2.48 54.06 2.68 ;
      RECT 53.14 2.48 53.34 2.68 ;
      RECT 52.14 1.92 52.34 2.12 ;
      RECT 50.7 3.04 50.9 3.24 ;
      RECT 44.565 2.935 44.765 3.135 ;
      RECT 43.785 0.9 43.985 1.1 ;
      RECT 43.555 3.04 43.755 3.24 ;
      RECT 43.075 2.315 43.275 2.515 ;
      RECT 42.075 7.125 42.275 7.325 ;
      RECT 41.475 3.04 41.675 3.24 ;
      RECT 39.915 2.48 40.115 2.68 ;
      RECT 39.535 3.6 39.735 3.8 ;
      RECT 39.035 2.48 39.235 2.68 ;
      RECT 38.075 2.48 38.275 2.68 ;
      RECT 37.355 2.48 37.555 2.68 ;
      RECT 36.355 1.92 36.555 2.12 ;
      RECT 34.915 3.04 35.115 3.24 ;
      RECT 28.79 2.935 28.99 3.135 ;
      RECT 28.01 0.9 28.21 1.1 ;
      RECT 27.78 3.04 27.98 3.24 ;
      RECT 27.3 2.315 27.5 2.515 ;
      RECT 26.3 7.125 26.5 7.325 ;
      RECT 25.7 3.04 25.9 3.24 ;
      RECT 24.14 2.48 24.34 2.68 ;
      RECT 23.76 3.6 23.96 3.8 ;
      RECT 23.26 2.48 23.46 2.68 ;
      RECT 22.3 2.48 22.5 2.68 ;
      RECT 21.58 2.48 21.78 2.68 ;
      RECT 20.58 1.92 20.78 2.12 ;
      RECT 19.14 3.04 19.34 3.24 ;
      RECT 13.01 2.935 13.21 3.135 ;
      RECT 12.23 0.9 12.43 1.1 ;
      RECT 12 3.04 12.2 3.24 ;
      RECT 11.52 2.315 11.72 2.515 ;
      RECT 10.52 7.125 10.72 7.325 ;
      RECT 9.92 3.04 10.12 3.24 ;
      RECT 8.36 2.48 8.56 2.68 ;
      RECT 7.98 3.6 8.18 3.8 ;
      RECT 7.48 2.48 7.68 2.68 ;
      RECT 6.52 2.48 6.72 2.68 ;
      RECT 5.8 2.48 6 2.68 ;
      RECT 4.8 1.92 5 2.12 ;
      RECT 3.36 3.04 3.56 3.24 ;
      RECT 0.28 0.09 0.48 0.29 ;
      RECT 0.28 8.59 0.48 8.79 ;
    LAYER met2 ;
      RECT 1.225 8.4 81.395 8.57 ;
      RECT 81.225 7.275 81.395 8.57 ;
      RECT 1.225 6.255 1.395 8.57 ;
      RECT 81.195 7.275 81.545 7.625 ;
      RECT 1.165 6.255 1.455 6.605 ;
      RECT 78.035 6.22 78.355 6.545 ;
      RECT 78.065 5.695 78.235 6.545 ;
      RECT 78.065 5.695 78.24 6.045 ;
      RECT 78.065 5.695 79.04 5.87 ;
      RECT 78.865 1.965 79.04 5.87 ;
      RECT 78.81 1.965 79.16 2.315 ;
      RECT 78.835 6.655 79.16 6.98 ;
      RECT 77.72 6.745 79.16 6.915 ;
      RECT 77.72 2.395 77.88 6.915 ;
      RECT 78.035 2.365 78.355 2.685 ;
      RECT 77.72 2.395 78.355 2.565 ;
      RECT 66.445 3 66.725 3.28 ;
      RECT 66.415 3 66.725 3.265 ;
      RECT 66.41 3 66.725 3.263 ;
      RECT 66.405 1.33 66.575 3.257 ;
      RECT 66.4 2.967 66.67 3.25 ;
      RECT 66.395 3 66.725 3.243 ;
      RECT 66.365 2.97 66.67 3.23 ;
      RECT 66.365 2.997 66.69 3.23 ;
      RECT 66.365 2.987 66.685 3.23 ;
      RECT 66.365 2.972 66.68 3.23 ;
      RECT 66.405 2.962 66.67 3.257 ;
      RECT 66.405 2.957 66.66 3.257 ;
      RECT 66.405 2.956 66.645 3.257 ;
      RECT 76.375 1.34 76.725 1.69 ;
      RECT 76.37 1.34 76.725 1.595 ;
      RECT 66.405 1.33 76.615 1.5 ;
      RECT 76.05 2.85 76.42 3.22 ;
      RECT 76.135 2.235 76.305 3.22 ;
      RECT 72.155 2.455 72.39 2.715 ;
      RECT 75.3 2.235 75.465 2.495 ;
      RECT 75.205 2.225 75.22 2.495 ;
      RECT 75.3 2.235 76.305 2.415 ;
      RECT 73.805 1.795 73.845 1.935 ;
      RECT 75.22 2.23 75.3 2.495 ;
      RECT 75.165 2.225 75.205 2.461 ;
      RECT 75.151 2.225 75.165 2.461 ;
      RECT 75.065 2.23 75.151 2.463 ;
      RECT 75.02 2.237 75.065 2.465 ;
      RECT 74.99 2.237 75.02 2.467 ;
      RECT 74.965 2.232 74.99 2.469 ;
      RECT 74.935 2.228 74.965 2.478 ;
      RECT 74.925 2.225 74.935 2.49 ;
      RECT 74.92 2.225 74.925 2.498 ;
      RECT 74.915 2.225 74.92 2.503 ;
      RECT 74.905 2.224 74.915 2.513 ;
      RECT 74.9 2.223 74.905 2.523 ;
      RECT 74.885 2.222 74.9 2.528 ;
      RECT 74.857 2.219 74.885 2.555 ;
      RECT 74.771 2.211 74.857 2.555 ;
      RECT 74.685 2.2 74.771 2.555 ;
      RECT 74.645 2.185 74.685 2.555 ;
      RECT 74.605 2.159 74.645 2.555 ;
      RECT 74.6 2.141 74.605 2.367 ;
      RECT 74.59 2.137 74.6 2.357 ;
      RECT 74.575 2.127 74.59 2.344 ;
      RECT 74.555 2.111 74.575 2.329 ;
      RECT 74.54 2.096 74.555 2.314 ;
      RECT 74.53 2.085 74.54 2.304 ;
      RECT 74.505 2.069 74.53 2.293 ;
      RECT 74.5 2.056 74.505 2.283 ;
      RECT 74.495 2.052 74.5 2.278 ;
      RECT 74.44 2.038 74.495 2.256 ;
      RECT 74.401 2.019 74.44 2.22 ;
      RECT 74.315 1.993 74.401 2.173 ;
      RECT 74.311 1.975 74.315 2.139 ;
      RECT 74.225 1.956 74.311 2.117 ;
      RECT 74.22 1.938 74.225 2.095 ;
      RECT 74.215 1.936 74.22 2.093 ;
      RECT 74.205 1.935 74.215 2.088 ;
      RECT 74.145 1.922 74.205 2.074 ;
      RECT 74.1 1.9 74.145 2.053 ;
      RECT 74.04 1.877 74.1 2.032 ;
      RECT 73.976 1.852 74.04 2.007 ;
      RECT 73.89 1.822 73.976 1.976 ;
      RECT 73.875 1.802 73.89 1.955 ;
      RECT 73.845 1.797 73.875 1.946 ;
      RECT 73.792 1.795 73.805 1.935 ;
      RECT 73.706 1.795 73.792 1.937 ;
      RECT 73.62 1.795 73.706 1.939 ;
      RECT 73.6 1.795 73.62 1.943 ;
      RECT 73.555 1.797 73.6 1.954 ;
      RECT 73.515 1.807 73.555 1.97 ;
      RECT 73.511 1.816 73.515 1.978 ;
      RECT 73.425 1.836 73.511 1.994 ;
      RECT 73.415 1.855 73.425 2.012 ;
      RECT 73.41 1.857 73.415 2.015 ;
      RECT 73.4 1.861 73.41 2.018 ;
      RECT 73.38 1.866 73.4 2.028 ;
      RECT 73.35 1.876 73.38 2.048 ;
      RECT 73.345 1.883 73.35 2.062 ;
      RECT 73.335 1.887 73.345 2.069 ;
      RECT 73.32 1.895 73.335 2.08 ;
      RECT 73.31 1.905 73.32 2.091 ;
      RECT 73.3 1.912 73.31 2.099 ;
      RECT 73.275 1.925 73.3 2.114 ;
      RECT 73.211 1.961 73.275 2.153 ;
      RECT 73.125 2.024 73.211 2.217 ;
      RECT 73.09 2.075 73.125 2.27 ;
      RECT 73.085 2.092 73.09 2.287 ;
      RECT 73.07 2.101 73.085 2.294 ;
      RECT 73.05 2.116 73.07 2.308 ;
      RECT 73.045 2.127 73.05 2.318 ;
      RECT 73.025 2.14 73.045 2.328 ;
      RECT 73.02 2.15 73.025 2.338 ;
      RECT 73.005 2.155 73.02 2.347 ;
      RECT 72.995 2.165 73.005 2.358 ;
      RECT 72.965 2.182 72.995 2.375 ;
      RECT 72.955 2.2 72.965 2.393 ;
      RECT 72.94 2.211 72.955 2.404 ;
      RECT 72.9 2.235 72.94 2.42 ;
      RECT 72.865 2.269 72.9 2.437 ;
      RECT 72.835 2.292 72.865 2.449 ;
      RECT 72.82 2.302 72.835 2.458 ;
      RECT 72.78 2.312 72.82 2.469 ;
      RECT 72.76 2.323 72.78 2.481 ;
      RECT 72.755 2.327 72.76 2.488 ;
      RECT 72.74 2.331 72.755 2.493 ;
      RECT 72.73 2.336 72.74 2.498 ;
      RECT 72.725 2.339 72.73 2.501 ;
      RECT 72.695 2.345 72.725 2.508 ;
      RECT 72.66 2.355 72.695 2.522 ;
      RECT 72.6 2.37 72.66 2.542 ;
      RECT 72.545 2.39 72.6 2.566 ;
      RECT 72.516 2.405 72.545 2.584 ;
      RECT 72.43 2.425 72.516 2.609 ;
      RECT 72.425 2.44 72.43 2.629 ;
      RECT 72.415 2.443 72.425 2.63 ;
      RECT 72.39 2.45 72.415 2.715 ;
      RECT 75.085 2.943 75.365 3.28 ;
      RECT 75.085 2.953 75.37 3.238 ;
      RECT 75.085 2.962 75.375 3.135 ;
      RECT 75.085 2.977 75.38 3.003 ;
      RECT 75.085 2.805 75.345 3.28 ;
      RECT 65.385 6.655 65.735 7.005 ;
      RECT 74.21 6.61 74.56 6.96 ;
      RECT 65.385 6.685 74.56 6.885 ;
      RECT 72.805 3.685 72.815 3.875 ;
      RECT 71.065 3.56 71.345 3.84 ;
      RECT 74.11 2.5 74.115 2.985 ;
      RECT 74.005 2.5 74.065 2.76 ;
      RECT 74.33 3.47 74.335 3.545 ;
      RECT 74.32 3.337 74.33 3.58 ;
      RECT 74.31 3.172 74.32 3.601 ;
      RECT 74.305 3.042 74.31 3.617 ;
      RECT 74.295 2.932 74.305 3.633 ;
      RECT 74.29 2.831 74.295 3.65 ;
      RECT 74.285 2.813 74.29 3.66 ;
      RECT 74.28 2.795 74.285 3.67 ;
      RECT 74.27 2.77 74.28 3.685 ;
      RECT 74.265 2.75 74.27 3.7 ;
      RECT 74.245 2.5 74.265 3.725 ;
      RECT 74.23 2.5 74.245 3.758 ;
      RECT 74.2 2.5 74.23 3.78 ;
      RECT 74.18 2.5 74.2 3.794 ;
      RECT 74.16 2.5 74.18 3.31 ;
      RECT 74.175 3.377 74.18 3.799 ;
      RECT 74.17 3.407 74.175 3.801 ;
      RECT 74.165 3.42 74.17 3.804 ;
      RECT 74.16 3.43 74.165 3.808 ;
      RECT 74.155 2.5 74.16 3.228 ;
      RECT 74.155 3.44 74.16 3.81 ;
      RECT 74.15 2.5 74.155 3.205 ;
      RECT 74.14 3.462 74.155 3.81 ;
      RECT 74.135 2.5 74.15 3.15 ;
      RECT 74.13 3.487 74.14 3.81 ;
      RECT 74.13 2.5 74.135 3.095 ;
      RECT 74.12 2.5 74.13 3.043 ;
      RECT 74.125 3.5 74.13 3.811 ;
      RECT 74.12 3.512 74.125 3.812 ;
      RECT 74.115 2.5 74.12 3.003 ;
      RECT 74.115 3.525 74.12 3.813 ;
      RECT 74.1 3.54 74.115 3.814 ;
      RECT 74.105 2.5 74.11 2.965 ;
      RECT 74.1 2.5 74.105 2.93 ;
      RECT 74.095 2.5 74.1 2.905 ;
      RECT 74.09 3.567 74.1 3.816 ;
      RECT 74.085 2.5 74.095 2.863 ;
      RECT 74.085 3.585 74.09 3.817 ;
      RECT 74.08 2.5 74.085 2.823 ;
      RECT 74.08 3.592 74.085 3.818 ;
      RECT 74.075 2.5 74.08 2.795 ;
      RECT 74.07 3.61 74.08 3.819 ;
      RECT 74.065 2.5 74.075 2.775 ;
      RECT 74.06 3.63 74.07 3.821 ;
      RECT 74.05 3.647 74.06 3.822 ;
      RECT 74.015 3.67 74.05 3.825 ;
      RECT 73.96 3.688 74.015 3.831 ;
      RECT 73.874 3.696 73.96 3.84 ;
      RECT 73.788 3.707 73.874 3.851 ;
      RECT 73.702 3.717 73.788 3.862 ;
      RECT 73.616 3.727 73.702 3.874 ;
      RECT 73.53 3.737 73.616 3.885 ;
      RECT 73.51 3.743 73.53 3.891 ;
      RECT 73.43 3.745 73.51 3.895 ;
      RECT 73.425 3.744 73.43 3.9 ;
      RECT 73.417 3.743 73.425 3.9 ;
      RECT 73.331 3.739 73.417 3.898 ;
      RECT 73.245 3.731 73.331 3.895 ;
      RECT 73.159 3.722 73.245 3.891 ;
      RECT 73.073 3.714 73.159 3.888 ;
      RECT 72.987 3.706 73.073 3.884 ;
      RECT 72.901 3.697 72.987 3.881 ;
      RECT 72.815 3.689 72.901 3.877 ;
      RECT 72.76 3.682 72.805 3.875 ;
      RECT 72.675 3.675 72.76 3.873 ;
      RECT 72.601 3.667 72.675 3.869 ;
      RECT 72.515 3.659 72.601 3.866 ;
      RECT 72.512 3.655 72.515 3.864 ;
      RECT 72.426 3.651 72.512 3.863 ;
      RECT 72.34 3.643 72.426 3.86 ;
      RECT 72.255 3.638 72.34 3.857 ;
      RECT 72.169 3.635 72.255 3.854 ;
      RECT 72.083 3.633 72.169 3.851 ;
      RECT 71.997 3.63 72.083 3.848 ;
      RECT 71.911 3.627 71.997 3.845 ;
      RECT 71.825 3.624 71.911 3.842 ;
      RECT 71.749 3.622 71.825 3.839 ;
      RECT 71.663 3.619 71.749 3.836 ;
      RECT 71.577 3.616 71.663 3.834 ;
      RECT 71.491 3.614 71.577 3.831 ;
      RECT 71.405 3.611 71.491 3.828 ;
      RECT 71.345 3.602 71.405 3.826 ;
      RECT 73.855 3.22 73.93 3.48 ;
      RECT 73.835 3.2 73.84 3.48 ;
      RECT 73.155 2.985 73.26 3.28 ;
      RECT 67.6 2.96 67.67 3.22 ;
      RECT 73.495 2.835 73.5 3.206 ;
      RECT 73.485 2.89 73.49 3.206 ;
      RECT 73.79 2.06 73.85 2.32 ;
      RECT 73.845 3.215 73.855 3.48 ;
      RECT 73.84 3.205 73.845 3.48 ;
      RECT 73.76 3.152 73.835 3.48 ;
      RECT 73.785 2.06 73.79 2.34 ;
      RECT 73.775 2.06 73.785 2.36 ;
      RECT 73.76 2.06 73.775 2.39 ;
      RECT 73.745 2.06 73.76 2.433 ;
      RECT 73.74 3.095 73.76 3.48 ;
      RECT 73.73 2.06 73.745 2.47 ;
      RECT 73.725 3.075 73.74 3.48 ;
      RECT 73.725 2.06 73.73 2.493 ;
      RECT 73.715 2.06 73.725 2.518 ;
      RECT 73.685 3.042 73.725 3.48 ;
      RECT 73.69 2.06 73.715 2.568 ;
      RECT 73.685 2.06 73.69 2.623 ;
      RECT 73.68 2.06 73.685 2.665 ;
      RECT 73.67 3.005 73.685 3.48 ;
      RECT 73.675 2.06 73.68 2.708 ;
      RECT 73.67 2.06 73.675 2.773 ;
      RECT 73.665 2.06 73.67 2.795 ;
      RECT 73.665 2.993 73.67 3.345 ;
      RECT 73.66 2.06 73.665 2.863 ;
      RECT 73.66 2.985 73.665 3.328 ;
      RECT 73.655 2.06 73.66 2.908 ;
      RECT 73.65 2.967 73.66 3.305 ;
      RECT 73.65 2.06 73.655 2.945 ;
      RECT 73.64 2.06 73.65 3.285 ;
      RECT 73.635 2.06 73.64 3.268 ;
      RECT 73.63 2.06 73.635 3.253 ;
      RECT 73.625 2.06 73.63 3.238 ;
      RECT 73.605 2.06 73.625 3.228 ;
      RECT 73.6 2.06 73.605 3.218 ;
      RECT 73.59 2.06 73.6 3.214 ;
      RECT 73.585 2.337 73.59 3.213 ;
      RECT 73.58 2.36 73.585 3.212 ;
      RECT 73.575 2.39 73.58 3.211 ;
      RECT 73.57 2.417 73.575 3.21 ;
      RECT 73.565 2.445 73.57 3.21 ;
      RECT 73.56 2.472 73.565 3.21 ;
      RECT 73.555 2.492 73.56 3.21 ;
      RECT 73.55 2.52 73.555 3.21 ;
      RECT 73.54 2.562 73.55 3.21 ;
      RECT 73.53 2.607 73.54 3.209 ;
      RECT 73.525 2.66 73.53 3.208 ;
      RECT 73.52 2.692 73.525 3.207 ;
      RECT 73.515 2.712 73.52 3.206 ;
      RECT 73.51 2.75 73.515 3.206 ;
      RECT 73.505 2.772 73.51 3.206 ;
      RECT 73.5 2.797 73.505 3.206 ;
      RECT 73.49 2.862 73.495 3.206 ;
      RECT 73.475 2.922 73.485 3.206 ;
      RECT 73.46 2.932 73.475 3.206 ;
      RECT 73.44 2.942 73.46 3.206 ;
      RECT 73.41 2.947 73.44 3.203 ;
      RECT 73.35 2.957 73.41 3.2 ;
      RECT 73.33 2.966 73.35 3.205 ;
      RECT 73.305 2.972 73.33 3.218 ;
      RECT 73.285 2.977 73.305 3.233 ;
      RECT 73.26 2.982 73.285 3.28 ;
      RECT 73.131 2.984 73.155 3.28 ;
      RECT 73.045 2.979 73.131 3.28 ;
      RECT 73.005 2.976 73.045 3.28 ;
      RECT 72.955 2.978 73.005 3.26 ;
      RECT 72.925 2.982 72.955 3.26 ;
      RECT 72.846 2.992 72.925 3.26 ;
      RECT 72.76 3.007 72.846 3.261 ;
      RECT 72.71 3.017 72.76 3.262 ;
      RECT 72.702 3.02 72.71 3.262 ;
      RECT 72.616 3.022 72.702 3.263 ;
      RECT 72.53 3.026 72.616 3.263 ;
      RECT 72.444 3.03 72.53 3.264 ;
      RECT 72.358 3.033 72.444 3.265 ;
      RECT 72.272 3.037 72.358 3.265 ;
      RECT 72.186 3.041 72.272 3.266 ;
      RECT 72.1 3.044 72.186 3.267 ;
      RECT 72.014 3.048 72.1 3.267 ;
      RECT 71.928 3.052 72.014 3.268 ;
      RECT 71.842 3.056 71.928 3.269 ;
      RECT 71.756 3.059 71.842 3.269 ;
      RECT 71.67 3.063 71.756 3.27 ;
      RECT 71.64 3.065 71.67 3.27 ;
      RECT 71.554 3.068 71.64 3.271 ;
      RECT 71.468 3.072 71.554 3.272 ;
      RECT 71.382 3.076 71.468 3.273 ;
      RECT 71.296 3.079 71.382 3.273 ;
      RECT 71.21 3.083 71.296 3.274 ;
      RECT 71.175 3.088 71.21 3.275 ;
      RECT 71.12 3.098 71.175 3.282 ;
      RECT 71.095 3.11 71.12 3.292 ;
      RECT 71.06 3.123 71.095 3.3 ;
      RECT 71.02 3.14 71.06 3.323 ;
      RECT 71 3.153 71.02 3.35 ;
      RECT 70.97 3.165 71 3.378 ;
      RECT 70.965 3.173 70.97 3.398 ;
      RECT 70.96 3.176 70.965 3.408 ;
      RECT 70.91 3.188 70.96 3.442 ;
      RECT 70.9 3.203 70.91 3.475 ;
      RECT 70.89 3.209 70.9 3.488 ;
      RECT 70.88 3.216 70.89 3.5 ;
      RECT 70.855 3.229 70.88 3.518 ;
      RECT 70.84 3.244 70.855 3.54 ;
      RECT 70.83 3.252 70.84 3.556 ;
      RECT 70.815 3.261 70.83 3.571 ;
      RECT 70.805 3.271 70.815 3.585 ;
      RECT 70.786 3.284 70.805 3.602 ;
      RECT 70.7 3.329 70.786 3.667 ;
      RECT 70.685 3.374 70.7 3.725 ;
      RECT 70.68 3.383 70.685 3.738 ;
      RECT 70.67 3.39 70.68 3.743 ;
      RECT 70.665 3.395 70.67 3.747 ;
      RECT 70.645 3.405 70.665 3.754 ;
      RECT 70.62 3.425 70.645 3.768 ;
      RECT 70.585 3.45 70.62 3.788 ;
      RECT 70.57 3.473 70.585 3.803 ;
      RECT 70.56 3.483 70.57 3.808 ;
      RECT 70.55 3.491 70.56 3.815 ;
      RECT 70.54 3.5 70.55 3.821 ;
      RECT 70.52 3.512 70.54 3.823 ;
      RECT 70.51 3.525 70.52 3.825 ;
      RECT 70.485 3.54 70.51 3.828 ;
      RECT 70.465 3.557 70.485 3.832 ;
      RECT 70.425 3.585 70.465 3.838 ;
      RECT 70.36 3.632 70.425 3.847 ;
      RECT 70.345 3.665 70.36 3.855 ;
      RECT 70.34 3.672 70.345 3.857 ;
      RECT 70.29 3.697 70.34 3.862 ;
      RECT 70.275 3.721 70.29 3.869 ;
      RECT 70.225 3.726 70.275 3.87 ;
      RECT 70.139 3.73 70.225 3.87 ;
      RECT 70.053 3.73 70.139 3.87 ;
      RECT 69.967 3.73 70.053 3.871 ;
      RECT 69.881 3.73 69.967 3.871 ;
      RECT 69.795 3.73 69.881 3.871 ;
      RECT 69.729 3.73 69.795 3.871 ;
      RECT 69.643 3.73 69.729 3.872 ;
      RECT 69.557 3.73 69.643 3.872 ;
      RECT 69.471 3.731 69.557 3.873 ;
      RECT 69.385 3.731 69.471 3.873 ;
      RECT 69.299 3.731 69.385 3.873 ;
      RECT 69.213 3.731 69.299 3.874 ;
      RECT 69.127 3.731 69.213 3.874 ;
      RECT 69.041 3.732 69.127 3.875 ;
      RECT 68.955 3.732 69.041 3.875 ;
      RECT 68.935 3.732 68.955 3.875 ;
      RECT 68.849 3.732 68.935 3.875 ;
      RECT 68.763 3.732 68.849 3.875 ;
      RECT 68.677 3.733 68.763 3.875 ;
      RECT 68.591 3.733 68.677 3.875 ;
      RECT 68.505 3.733 68.591 3.875 ;
      RECT 68.419 3.734 68.505 3.875 ;
      RECT 68.333 3.734 68.419 3.875 ;
      RECT 68.247 3.734 68.333 3.875 ;
      RECT 68.161 3.734 68.247 3.875 ;
      RECT 68.075 3.735 68.161 3.875 ;
      RECT 68.025 3.732 68.075 3.875 ;
      RECT 68.015 3.73 68.025 3.874 ;
      RECT 68.011 3.73 68.015 3.873 ;
      RECT 67.925 3.725 68.011 3.868 ;
      RECT 67.903 3.718 67.925 3.862 ;
      RECT 67.817 3.709 67.903 3.856 ;
      RECT 67.731 3.696 67.817 3.847 ;
      RECT 67.645 3.682 67.731 3.837 ;
      RECT 67.6 3.672 67.645 3.83 ;
      RECT 67.58 2.96 67.6 3.238 ;
      RECT 67.58 3.665 67.6 3.826 ;
      RECT 67.55 2.96 67.58 3.26 ;
      RECT 67.54 3.632 67.58 3.823 ;
      RECT 67.535 2.96 67.55 3.28 ;
      RECT 67.535 3.597 67.54 3.821 ;
      RECT 67.53 2.96 67.535 3.405 ;
      RECT 67.53 3.557 67.535 3.821 ;
      RECT 67.52 2.96 67.53 3.821 ;
      RECT 67.445 2.96 67.52 3.815 ;
      RECT 67.415 2.96 67.445 3.805 ;
      RECT 67.41 2.96 67.415 3.797 ;
      RECT 67.405 3.002 67.41 3.79 ;
      RECT 67.395 3.071 67.405 3.781 ;
      RECT 67.39 3.141 67.395 3.733 ;
      RECT 67.385 3.205 67.39 3.63 ;
      RECT 67.38 3.24 67.385 3.585 ;
      RECT 67.378 3.277 67.38 3.477 ;
      RECT 67.375 3.285 67.378 3.47 ;
      RECT 67.37 3.35 67.375 3.413 ;
      RECT 71.445 2.44 71.725 2.72 ;
      RECT 71.435 2.44 71.725 2.583 ;
      RECT 71.39 2.305 71.65 2.565 ;
      RECT 71.39 2.42 71.705 2.565 ;
      RECT 71.39 2.39 71.7 2.565 ;
      RECT 71.39 2.377 71.69 2.565 ;
      RECT 71.39 2.367 71.685 2.565 ;
      RECT 67.365 2.35 67.625 2.61 ;
      RECT 71.135 1.9 71.395 2.16 ;
      RECT 71.125 1.925 71.395 2.12 ;
      RECT 71.12 1.925 71.125 2.119 ;
      RECT 71.05 1.92 71.12 2.111 ;
      RECT 70.965 1.907 71.05 2.094 ;
      RECT 70.961 1.899 70.965 2.084 ;
      RECT 70.875 1.892 70.961 2.074 ;
      RECT 70.866 1.884 70.875 2.064 ;
      RECT 70.78 1.877 70.866 2.052 ;
      RECT 70.76 1.868 70.78 2.038 ;
      RECT 70.705 1.863 70.76 2.03 ;
      RECT 70.695 1.857 70.705 2.024 ;
      RECT 70.675 1.855 70.695 2.02 ;
      RECT 70.667 1.854 70.675 2.016 ;
      RECT 70.581 1.846 70.667 2.005 ;
      RECT 70.495 1.832 70.581 1.985 ;
      RECT 70.435 1.82 70.495 1.97 ;
      RECT 70.425 1.815 70.435 1.965 ;
      RECT 70.375 1.815 70.425 1.967 ;
      RECT 70.328 1.817 70.375 1.971 ;
      RECT 70.242 1.824 70.328 1.976 ;
      RECT 70.156 1.832 70.242 1.982 ;
      RECT 70.07 1.841 70.156 1.988 ;
      RECT 70.011 1.847 70.07 1.993 ;
      RECT 69.925 1.852 70.011 1.999 ;
      RECT 69.85 1.857 69.925 2.005 ;
      RECT 69.811 1.859 69.85 2.01 ;
      RECT 69.725 1.856 69.811 2.015 ;
      RECT 69.64 1.854 69.725 2.022 ;
      RECT 69.608 1.853 69.64 2.025 ;
      RECT 69.522 1.852 69.608 2.026 ;
      RECT 69.436 1.851 69.522 2.027 ;
      RECT 69.35 1.85 69.436 2.027 ;
      RECT 69.264 1.849 69.35 2.028 ;
      RECT 69.178 1.848 69.264 2.029 ;
      RECT 69.092 1.847 69.178 2.03 ;
      RECT 69.006 1.846 69.092 2.03 ;
      RECT 68.92 1.845 69.006 2.031 ;
      RECT 68.87 1.845 68.92 2.032 ;
      RECT 68.856 1.846 68.87 2.032 ;
      RECT 68.77 1.853 68.856 2.033 ;
      RECT 68.696 1.864 68.77 2.034 ;
      RECT 68.61 1.873 68.696 2.035 ;
      RECT 68.575 1.88 68.61 2.05 ;
      RECT 68.55 1.883 68.575 2.08 ;
      RECT 68.525 1.892 68.55 2.109 ;
      RECT 68.515 1.903 68.525 2.129 ;
      RECT 68.505 1.911 68.515 2.143 ;
      RECT 68.5 1.917 68.505 2.153 ;
      RECT 68.475 1.934 68.5 2.17 ;
      RECT 68.46 1.956 68.475 2.198 ;
      RECT 68.43 1.982 68.46 2.228 ;
      RECT 68.41 2.011 68.43 2.258 ;
      RECT 68.405 2.026 68.41 2.275 ;
      RECT 68.385 2.041 68.405 2.29 ;
      RECT 68.375 2.059 68.385 2.308 ;
      RECT 68.365 2.07 68.375 2.323 ;
      RECT 68.315 2.102 68.365 2.349 ;
      RECT 68.31 2.132 68.315 2.369 ;
      RECT 68.3 2.145 68.31 2.375 ;
      RECT 68.291 2.155 68.3 2.383 ;
      RECT 68.28 2.166 68.291 2.391 ;
      RECT 68.275 2.176 68.28 2.397 ;
      RECT 68.26 2.197 68.275 2.404 ;
      RECT 68.245 2.227 68.26 2.412 ;
      RECT 68.21 2.257 68.245 2.418 ;
      RECT 68.185 2.275 68.21 2.425 ;
      RECT 68.135 2.283 68.185 2.434 ;
      RECT 68.11 2.288 68.135 2.443 ;
      RECT 68.055 2.294 68.11 2.453 ;
      RECT 68.05 2.299 68.055 2.461 ;
      RECT 68.036 2.302 68.05 2.463 ;
      RECT 67.95 2.314 68.036 2.475 ;
      RECT 67.94 2.326 67.95 2.488 ;
      RECT 67.855 2.339 67.94 2.5 ;
      RECT 67.811 2.356 67.855 2.514 ;
      RECT 67.725 2.373 67.811 2.53 ;
      RECT 67.695 2.387 67.725 2.544 ;
      RECT 67.685 2.392 67.695 2.549 ;
      RECT 67.625 2.395 67.685 2.558 ;
      RECT 70.515 2.665 70.775 2.925 ;
      RECT 70.515 2.665 70.795 2.778 ;
      RECT 70.515 2.665 70.82 2.745 ;
      RECT 70.515 2.665 70.825 2.725 ;
      RECT 70.565 2.44 70.845 2.72 ;
      RECT 70.12 3.175 70.38 3.435 ;
      RECT 70.11 3.032 70.305 3.373 ;
      RECT 70.105 3.14 70.32 3.365 ;
      RECT 70.1 3.19 70.38 3.355 ;
      RECT 70.09 3.267 70.38 3.34 ;
      RECT 70.11 3.115 70.32 3.373 ;
      RECT 70.12 2.99 70.305 3.435 ;
      RECT 70.12 2.885 70.285 3.435 ;
      RECT 70.13 2.872 70.285 3.435 ;
      RECT 70.13 2.83 70.275 3.435 ;
      RECT 70.135 2.755 70.275 3.435 ;
      RECT 70.165 2.405 70.275 3.435 ;
      RECT 70.17 2.135 70.295 2.758 ;
      RECT 70.14 2.71 70.295 2.758 ;
      RECT 70.155 2.512 70.275 3.435 ;
      RECT 70.145 2.622 70.295 2.758 ;
      RECT 70.17 2.135 70.31 2.615 ;
      RECT 70.17 2.135 70.33 2.49 ;
      RECT 70.135 2.135 70.395 2.395 ;
      RECT 69.605 2.44 69.885 2.72 ;
      RECT 69.59 2.44 69.885 2.7 ;
      RECT 67.645 3.305 67.905 3.565 ;
      RECT 69.43 3.16 69.69 3.42 ;
      RECT 69.41 3.18 69.69 3.395 ;
      RECT 69.367 3.18 69.41 3.394 ;
      RECT 69.281 3.181 69.367 3.391 ;
      RECT 69.195 3.182 69.281 3.387 ;
      RECT 69.12 3.184 69.195 3.384 ;
      RECT 69.097 3.185 69.12 3.382 ;
      RECT 69.011 3.186 69.097 3.38 ;
      RECT 68.925 3.187 69.011 3.377 ;
      RECT 68.901 3.188 68.925 3.375 ;
      RECT 68.815 3.19 68.901 3.372 ;
      RECT 68.73 3.192 68.815 3.373 ;
      RECT 68.673 3.193 68.73 3.379 ;
      RECT 68.587 3.195 68.673 3.389 ;
      RECT 68.501 3.198 68.587 3.402 ;
      RECT 68.415 3.2 68.501 3.414 ;
      RECT 68.401 3.201 68.415 3.421 ;
      RECT 68.315 3.202 68.401 3.429 ;
      RECT 68.275 3.204 68.315 3.438 ;
      RECT 68.266 3.205 68.275 3.441 ;
      RECT 68.18 3.213 68.266 3.447 ;
      RECT 68.16 3.222 68.18 3.455 ;
      RECT 68.075 3.237 68.16 3.463 ;
      RECT 68.015 3.26 68.075 3.474 ;
      RECT 68.005 3.272 68.015 3.479 ;
      RECT 67.965 3.282 68.005 3.483 ;
      RECT 67.91 3.299 67.965 3.491 ;
      RECT 67.905 3.309 67.91 3.495 ;
      RECT 68.971 2.44 69.03 2.837 ;
      RECT 68.885 2.44 69.09 2.828 ;
      RECT 68.88 2.47 69.09 2.823 ;
      RECT 68.846 2.47 69.09 2.821 ;
      RECT 68.76 2.47 69.09 2.815 ;
      RECT 68.715 2.47 69.11 2.793 ;
      RECT 68.715 2.47 69.13 2.748 ;
      RECT 68.675 2.47 69.13 2.738 ;
      RECT 68.885 2.44 69.165 2.72 ;
      RECT 68.62 2.44 68.88 2.7 ;
      RECT 67.805 1.92 68.065 2.18 ;
      RECT 67.885 1.88 68.165 2.16 ;
      RECT 62.25 6.22 62.57 6.545 ;
      RECT 62.28 5.695 62.45 6.545 ;
      RECT 62.28 5.695 62.455 6.045 ;
      RECT 62.28 5.695 63.255 5.87 ;
      RECT 63.08 1.965 63.255 5.87 ;
      RECT 63.025 1.965 63.375 2.315 ;
      RECT 63.05 6.655 63.375 6.98 ;
      RECT 61.935 6.745 63.375 6.915 ;
      RECT 61.935 2.395 62.095 6.915 ;
      RECT 62.25 2.365 62.57 2.685 ;
      RECT 61.935 2.395 62.57 2.565 ;
      RECT 50.66 3 50.94 3.28 ;
      RECT 50.63 3 50.94 3.265 ;
      RECT 50.625 3 50.94 3.263 ;
      RECT 50.62 1.33 50.79 3.257 ;
      RECT 50.615 2.967 50.885 3.25 ;
      RECT 50.61 3 50.94 3.243 ;
      RECT 50.58 2.97 50.885 3.23 ;
      RECT 50.58 2.997 50.905 3.23 ;
      RECT 50.58 2.987 50.9 3.23 ;
      RECT 50.58 2.972 50.895 3.23 ;
      RECT 50.62 2.962 50.885 3.257 ;
      RECT 50.62 2.957 50.875 3.257 ;
      RECT 50.62 2.956 50.86 3.257 ;
      RECT 60.59 1.34 60.94 1.69 ;
      RECT 60.585 1.34 60.94 1.595 ;
      RECT 50.62 1.33 60.83 1.5 ;
      RECT 60.265 2.85 60.635 3.22 ;
      RECT 60.35 2.235 60.52 3.22 ;
      RECT 56.37 2.455 56.605 2.715 ;
      RECT 59.515 2.235 59.68 2.495 ;
      RECT 59.42 2.225 59.435 2.495 ;
      RECT 59.515 2.235 60.52 2.415 ;
      RECT 58.02 1.795 58.06 1.935 ;
      RECT 59.435 2.23 59.515 2.495 ;
      RECT 59.38 2.225 59.42 2.461 ;
      RECT 59.366 2.225 59.38 2.461 ;
      RECT 59.28 2.23 59.366 2.463 ;
      RECT 59.235 2.237 59.28 2.465 ;
      RECT 59.205 2.237 59.235 2.467 ;
      RECT 59.18 2.232 59.205 2.469 ;
      RECT 59.15 2.228 59.18 2.478 ;
      RECT 59.14 2.225 59.15 2.49 ;
      RECT 59.135 2.225 59.14 2.498 ;
      RECT 59.13 2.225 59.135 2.503 ;
      RECT 59.12 2.224 59.13 2.513 ;
      RECT 59.115 2.223 59.12 2.523 ;
      RECT 59.1 2.222 59.115 2.528 ;
      RECT 59.072 2.219 59.1 2.555 ;
      RECT 58.986 2.211 59.072 2.555 ;
      RECT 58.9 2.2 58.986 2.555 ;
      RECT 58.86 2.185 58.9 2.555 ;
      RECT 58.82 2.159 58.86 2.555 ;
      RECT 58.815 2.141 58.82 2.367 ;
      RECT 58.805 2.137 58.815 2.357 ;
      RECT 58.79 2.127 58.805 2.344 ;
      RECT 58.77 2.111 58.79 2.329 ;
      RECT 58.755 2.096 58.77 2.314 ;
      RECT 58.745 2.085 58.755 2.304 ;
      RECT 58.72 2.069 58.745 2.293 ;
      RECT 58.715 2.056 58.72 2.283 ;
      RECT 58.71 2.052 58.715 2.278 ;
      RECT 58.655 2.038 58.71 2.256 ;
      RECT 58.616 2.019 58.655 2.22 ;
      RECT 58.53 1.993 58.616 2.173 ;
      RECT 58.526 1.975 58.53 2.139 ;
      RECT 58.44 1.956 58.526 2.117 ;
      RECT 58.435 1.938 58.44 2.095 ;
      RECT 58.43 1.936 58.435 2.093 ;
      RECT 58.42 1.935 58.43 2.088 ;
      RECT 58.36 1.922 58.42 2.074 ;
      RECT 58.315 1.9 58.36 2.053 ;
      RECT 58.255 1.877 58.315 2.032 ;
      RECT 58.191 1.852 58.255 2.007 ;
      RECT 58.105 1.822 58.191 1.976 ;
      RECT 58.09 1.802 58.105 1.955 ;
      RECT 58.06 1.797 58.09 1.946 ;
      RECT 58.007 1.795 58.02 1.935 ;
      RECT 57.921 1.795 58.007 1.937 ;
      RECT 57.835 1.795 57.921 1.939 ;
      RECT 57.815 1.795 57.835 1.943 ;
      RECT 57.77 1.797 57.815 1.954 ;
      RECT 57.73 1.807 57.77 1.97 ;
      RECT 57.726 1.816 57.73 1.978 ;
      RECT 57.64 1.836 57.726 1.994 ;
      RECT 57.63 1.855 57.64 2.012 ;
      RECT 57.625 1.857 57.63 2.015 ;
      RECT 57.615 1.861 57.625 2.018 ;
      RECT 57.595 1.866 57.615 2.028 ;
      RECT 57.565 1.876 57.595 2.048 ;
      RECT 57.56 1.883 57.565 2.062 ;
      RECT 57.55 1.887 57.56 2.069 ;
      RECT 57.535 1.895 57.55 2.08 ;
      RECT 57.525 1.905 57.535 2.091 ;
      RECT 57.515 1.912 57.525 2.099 ;
      RECT 57.49 1.925 57.515 2.114 ;
      RECT 57.426 1.961 57.49 2.153 ;
      RECT 57.34 2.024 57.426 2.217 ;
      RECT 57.305 2.075 57.34 2.27 ;
      RECT 57.3 2.092 57.305 2.287 ;
      RECT 57.285 2.101 57.3 2.294 ;
      RECT 57.265 2.116 57.285 2.308 ;
      RECT 57.26 2.127 57.265 2.318 ;
      RECT 57.24 2.14 57.26 2.328 ;
      RECT 57.235 2.15 57.24 2.338 ;
      RECT 57.22 2.155 57.235 2.347 ;
      RECT 57.21 2.165 57.22 2.358 ;
      RECT 57.18 2.182 57.21 2.375 ;
      RECT 57.17 2.2 57.18 2.393 ;
      RECT 57.155 2.211 57.17 2.404 ;
      RECT 57.115 2.235 57.155 2.42 ;
      RECT 57.08 2.269 57.115 2.437 ;
      RECT 57.05 2.292 57.08 2.449 ;
      RECT 57.035 2.302 57.05 2.458 ;
      RECT 56.995 2.312 57.035 2.469 ;
      RECT 56.975 2.323 56.995 2.481 ;
      RECT 56.97 2.327 56.975 2.488 ;
      RECT 56.955 2.331 56.97 2.493 ;
      RECT 56.945 2.336 56.955 2.498 ;
      RECT 56.94 2.339 56.945 2.501 ;
      RECT 56.91 2.345 56.94 2.508 ;
      RECT 56.875 2.355 56.91 2.522 ;
      RECT 56.815 2.37 56.875 2.542 ;
      RECT 56.76 2.39 56.815 2.566 ;
      RECT 56.731 2.405 56.76 2.584 ;
      RECT 56.645 2.425 56.731 2.609 ;
      RECT 56.64 2.44 56.645 2.629 ;
      RECT 56.63 2.443 56.64 2.63 ;
      RECT 56.605 2.45 56.63 2.715 ;
      RECT 59.3 2.943 59.58 3.28 ;
      RECT 59.3 2.953 59.585 3.238 ;
      RECT 59.3 2.962 59.59 3.135 ;
      RECT 59.3 2.977 59.595 3.003 ;
      RECT 59.3 2.805 59.56 3.28 ;
      RECT 49.6 6.655 49.95 7.005 ;
      RECT 58.425 6.61 58.775 6.96 ;
      RECT 49.6 6.685 58.775 6.885 ;
      RECT 57.02 3.685 57.03 3.875 ;
      RECT 55.28 3.56 55.56 3.84 ;
      RECT 58.325 2.5 58.33 2.985 ;
      RECT 58.22 2.5 58.28 2.76 ;
      RECT 58.545 3.47 58.55 3.545 ;
      RECT 58.535 3.337 58.545 3.58 ;
      RECT 58.525 3.172 58.535 3.601 ;
      RECT 58.52 3.042 58.525 3.617 ;
      RECT 58.51 2.932 58.52 3.633 ;
      RECT 58.505 2.831 58.51 3.65 ;
      RECT 58.5 2.813 58.505 3.66 ;
      RECT 58.495 2.795 58.5 3.67 ;
      RECT 58.485 2.77 58.495 3.685 ;
      RECT 58.48 2.75 58.485 3.7 ;
      RECT 58.46 2.5 58.48 3.725 ;
      RECT 58.445 2.5 58.46 3.758 ;
      RECT 58.415 2.5 58.445 3.78 ;
      RECT 58.395 2.5 58.415 3.794 ;
      RECT 58.375 2.5 58.395 3.31 ;
      RECT 58.39 3.377 58.395 3.799 ;
      RECT 58.385 3.407 58.39 3.801 ;
      RECT 58.38 3.42 58.385 3.804 ;
      RECT 58.375 3.43 58.38 3.808 ;
      RECT 58.37 2.5 58.375 3.228 ;
      RECT 58.37 3.44 58.375 3.81 ;
      RECT 58.365 2.5 58.37 3.205 ;
      RECT 58.355 3.462 58.37 3.81 ;
      RECT 58.35 2.5 58.365 3.15 ;
      RECT 58.345 3.487 58.355 3.81 ;
      RECT 58.345 2.5 58.35 3.095 ;
      RECT 58.335 2.5 58.345 3.043 ;
      RECT 58.34 3.5 58.345 3.811 ;
      RECT 58.335 3.512 58.34 3.812 ;
      RECT 58.33 2.5 58.335 3.003 ;
      RECT 58.33 3.525 58.335 3.813 ;
      RECT 58.315 3.54 58.33 3.814 ;
      RECT 58.32 2.5 58.325 2.965 ;
      RECT 58.315 2.5 58.32 2.93 ;
      RECT 58.31 2.5 58.315 2.905 ;
      RECT 58.305 3.567 58.315 3.816 ;
      RECT 58.3 2.5 58.31 2.863 ;
      RECT 58.3 3.585 58.305 3.817 ;
      RECT 58.295 2.5 58.3 2.823 ;
      RECT 58.295 3.592 58.3 3.818 ;
      RECT 58.29 2.5 58.295 2.795 ;
      RECT 58.285 3.61 58.295 3.819 ;
      RECT 58.28 2.5 58.29 2.775 ;
      RECT 58.275 3.63 58.285 3.821 ;
      RECT 58.265 3.647 58.275 3.822 ;
      RECT 58.23 3.67 58.265 3.825 ;
      RECT 58.175 3.688 58.23 3.831 ;
      RECT 58.089 3.696 58.175 3.84 ;
      RECT 58.003 3.707 58.089 3.851 ;
      RECT 57.917 3.717 58.003 3.862 ;
      RECT 57.831 3.727 57.917 3.874 ;
      RECT 57.745 3.737 57.831 3.885 ;
      RECT 57.725 3.743 57.745 3.891 ;
      RECT 57.645 3.745 57.725 3.895 ;
      RECT 57.64 3.744 57.645 3.9 ;
      RECT 57.632 3.743 57.64 3.9 ;
      RECT 57.546 3.739 57.632 3.898 ;
      RECT 57.46 3.731 57.546 3.895 ;
      RECT 57.374 3.722 57.46 3.891 ;
      RECT 57.288 3.714 57.374 3.888 ;
      RECT 57.202 3.706 57.288 3.884 ;
      RECT 57.116 3.697 57.202 3.881 ;
      RECT 57.03 3.689 57.116 3.877 ;
      RECT 56.975 3.682 57.02 3.875 ;
      RECT 56.89 3.675 56.975 3.873 ;
      RECT 56.816 3.667 56.89 3.869 ;
      RECT 56.73 3.659 56.816 3.866 ;
      RECT 56.727 3.655 56.73 3.864 ;
      RECT 56.641 3.651 56.727 3.863 ;
      RECT 56.555 3.643 56.641 3.86 ;
      RECT 56.47 3.638 56.555 3.857 ;
      RECT 56.384 3.635 56.47 3.854 ;
      RECT 56.298 3.633 56.384 3.851 ;
      RECT 56.212 3.63 56.298 3.848 ;
      RECT 56.126 3.627 56.212 3.845 ;
      RECT 56.04 3.624 56.126 3.842 ;
      RECT 55.964 3.622 56.04 3.839 ;
      RECT 55.878 3.619 55.964 3.836 ;
      RECT 55.792 3.616 55.878 3.834 ;
      RECT 55.706 3.614 55.792 3.831 ;
      RECT 55.62 3.611 55.706 3.828 ;
      RECT 55.56 3.602 55.62 3.826 ;
      RECT 58.07 3.22 58.145 3.48 ;
      RECT 58.05 3.2 58.055 3.48 ;
      RECT 57.37 2.985 57.475 3.28 ;
      RECT 51.815 2.96 51.885 3.22 ;
      RECT 57.71 2.835 57.715 3.206 ;
      RECT 57.7 2.89 57.705 3.206 ;
      RECT 58.005 2.06 58.065 2.32 ;
      RECT 58.06 3.215 58.07 3.48 ;
      RECT 58.055 3.205 58.06 3.48 ;
      RECT 57.975 3.152 58.05 3.48 ;
      RECT 58 2.06 58.005 2.34 ;
      RECT 57.99 2.06 58 2.36 ;
      RECT 57.975 2.06 57.99 2.39 ;
      RECT 57.96 2.06 57.975 2.433 ;
      RECT 57.955 3.095 57.975 3.48 ;
      RECT 57.945 2.06 57.96 2.47 ;
      RECT 57.94 3.075 57.955 3.48 ;
      RECT 57.94 2.06 57.945 2.493 ;
      RECT 57.93 2.06 57.94 2.518 ;
      RECT 57.9 3.042 57.94 3.48 ;
      RECT 57.905 2.06 57.93 2.568 ;
      RECT 57.9 2.06 57.905 2.623 ;
      RECT 57.895 2.06 57.9 2.665 ;
      RECT 57.885 3.005 57.9 3.48 ;
      RECT 57.89 2.06 57.895 2.708 ;
      RECT 57.885 2.06 57.89 2.773 ;
      RECT 57.88 2.06 57.885 2.795 ;
      RECT 57.88 2.993 57.885 3.345 ;
      RECT 57.875 2.06 57.88 2.863 ;
      RECT 57.875 2.985 57.88 3.328 ;
      RECT 57.87 2.06 57.875 2.908 ;
      RECT 57.865 2.967 57.875 3.305 ;
      RECT 57.865 2.06 57.87 2.945 ;
      RECT 57.855 2.06 57.865 3.285 ;
      RECT 57.85 2.06 57.855 3.268 ;
      RECT 57.845 2.06 57.85 3.253 ;
      RECT 57.84 2.06 57.845 3.238 ;
      RECT 57.82 2.06 57.84 3.228 ;
      RECT 57.815 2.06 57.82 3.218 ;
      RECT 57.805 2.06 57.815 3.214 ;
      RECT 57.8 2.337 57.805 3.213 ;
      RECT 57.795 2.36 57.8 3.212 ;
      RECT 57.79 2.39 57.795 3.211 ;
      RECT 57.785 2.417 57.79 3.21 ;
      RECT 57.78 2.445 57.785 3.21 ;
      RECT 57.775 2.472 57.78 3.21 ;
      RECT 57.77 2.492 57.775 3.21 ;
      RECT 57.765 2.52 57.77 3.21 ;
      RECT 57.755 2.562 57.765 3.21 ;
      RECT 57.745 2.607 57.755 3.209 ;
      RECT 57.74 2.66 57.745 3.208 ;
      RECT 57.735 2.692 57.74 3.207 ;
      RECT 57.73 2.712 57.735 3.206 ;
      RECT 57.725 2.75 57.73 3.206 ;
      RECT 57.72 2.772 57.725 3.206 ;
      RECT 57.715 2.797 57.72 3.206 ;
      RECT 57.705 2.862 57.71 3.206 ;
      RECT 57.69 2.922 57.7 3.206 ;
      RECT 57.675 2.932 57.69 3.206 ;
      RECT 57.655 2.942 57.675 3.206 ;
      RECT 57.625 2.947 57.655 3.203 ;
      RECT 57.565 2.957 57.625 3.2 ;
      RECT 57.545 2.966 57.565 3.205 ;
      RECT 57.52 2.972 57.545 3.218 ;
      RECT 57.5 2.977 57.52 3.233 ;
      RECT 57.475 2.982 57.5 3.28 ;
      RECT 57.346 2.984 57.37 3.28 ;
      RECT 57.26 2.979 57.346 3.28 ;
      RECT 57.22 2.976 57.26 3.28 ;
      RECT 57.17 2.978 57.22 3.26 ;
      RECT 57.14 2.982 57.17 3.26 ;
      RECT 57.061 2.992 57.14 3.26 ;
      RECT 56.975 3.007 57.061 3.261 ;
      RECT 56.925 3.017 56.975 3.262 ;
      RECT 56.917 3.02 56.925 3.262 ;
      RECT 56.831 3.022 56.917 3.263 ;
      RECT 56.745 3.026 56.831 3.263 ;
      RECT 56.659 3.03 56.745 3.264 ;
      RECT 56.573 3.033 56.659 3.265 ;
      RECT 56.487 3.037 56.573 3.265 ;
      RECT 56.401 3.041 56.487 3.266 ;
      RECT 56.315 3.044 56.401 3.267 ;
      RECT 56.229 3.048 56.315 3.267 ;
      RECT 56.143 3.052 56.229 3.268 ;
      RECT 56.057 3.056 56.143 3.269 ;
      RECT 55.971 3.059 56.057 3.269 ;
      RECT 55.885 3.063 55.971 3.27 ;
      RECT 55.855 3.065 55.885 3.27 ;
      RECT 55.769 3.068 55.855 3.271 ;
      RECT 55.683 3.072 55.769 3.272 ;
      RECT 55.597 3.076 55.683 3.273 ;
      RECT 55.511 3.079 55.597 3.273 ;
      RECT 55.425 3.083 55.511 3.274 ;
      RECT 55.39 3.088 55.425 3.275 ;
      RECT 55.335 3.098 55.39 3.282 ;
      RECT 55.31 3.11 55.335 3.292 ;
      RECT 55.275 3.123 55.31 3.3 ;
      RECT 55.235 3.14 55.275 3.323 ;
      RECT 55.215 3.153 55.235 3.35 ;
      RECT 55.185 3.165 55.215 3.378 ;
      RECT 55.18 3.173 55.185 3.398 ;
      RECT 55.175 3.176 55.18 3.408 ;
      RECT 55.125 3.188 55.175 3.442 ;
      RECT 55.115 3.203 55.125 3.475 ;
      RECT 55.105 3.209 55.115 3.488 ;
      RECT 55.095 3.216 55.105 3.5 ;
      RECT 55.07 3.229 55.095 3.518 ;
      RECT 55.055 3.244 55.07 3.54 ;
      RECT 55.045 3.252 55.055 3.556 ;
      RECT 55.03 3.261 55.045 3.571 ;
      RECT 55.02 3.271 55.03 3.585 ;
      RECT 55.001 3.284 55.02 3.602 ;
      RECT 54.915 3.329 55.001 3.667 ;
      RECT 54.9 3.374 54.915 3.725 ;
      RECT 54.895 3.383 54.9 3.738 ;
      RECT 54.885 3.39 54.895 3.743 ;
      RECT 54.88 3.395 54.885 3.747 ;
      RECT 54.86 3.405 54.88 3.754 ;
      RECT 54.835 3.425 54.86 3.768 ;
      RECT 54.8 3.45 54.835 3.788 ;
      RECT 54.785 3.473 54.8 3.803 ;
      RECT 54.775 3.483 54.785 3.808 ;
      RECT 54.765 3.491 54.775 3.815 ;
      RECT 54.755 3.5 54.765 3.821 ;
      RECT 54.735 3.512 54.755 3.823 ;
      RECT 54.725 3.525 54.735 3.825 ;
      RECT 54.7 3.54 54.725 3.828 ;
      RECT 54.68 3.557 54.7 3.832 ;
      RECT 54.64 3.585 54.68 3.838 ;
      RECT 54.575 3.632 54.64 3.847 ;
      RECT 54.56 3.665 54.575 3.855 ;
      RECT 54.555 3.672 54.56 3.857 ;
      RECT 54.505 3.697 54.555 3.862 ;
      RECT 54.49 3.721 54.505 3.869 ;
      RECT 54.44 3.726 54.49 3.87 ;
      RECT 54.354 3.73 54.44 3.87 ;
      RECT 54.268 3.73 54.354 3.87 ;
      RECT 54.182 3.73 54.268 3.871 ;
      RECT 54.096 3.73 54.182 3.871 ;
      RECT 54.01 3.73 54.096 3.871 ;
      RECT 53.944 3.73 54.01 3.871 ;
      RECT 53.858 3.73 53.944 3.872 ;
      RECT 53.772 3.73 53.858 3.872 ;
      RECT 53.686 3.731 53.772 3.873 ;
      RECT 53.6 3.731 53.686 3.873 ;
      RECT 53.514 3.731 53.6 3.873 ;
      RECT 53.428 3.731 53.514 3.874 ;
      RECT 53.342 3.731 53.428 3.874 ;
      RECT 53.256 3.732 53.342 3.875 ;
      RECT 53.17 3.732 53.256 3.875 ;
      RECT 53.15 3.732 53.17 3.875 ;
      RECT 53.064 3.732 53.15 3.875 ;
      RECT 52.978 3.732 53.064 3.875 ;
      RECT 52.892 3.733 52.978 3.875 ;
      RECT 52.806 3.733 52.892 3.875 ;
      RECT 52.72 3.733 52.806 3.875 ;
      RECT 52.634 3.734 52.72 3.875 ;
      RECT 52.548 3.734 52.634 3.875 ;
      RECT 52.462 3.734 52.548 3.875 ;
      RECT 52.376 3.734 52.462 3.875 ;
      RECT 52.29 3.735 52.376 3.875 ;
      RECT 52.24 3.732 52.29 3.875 ;
      RECT 52.23 3.73 52.24 3.874 ;
      RECT 52.226 3.73 52.23 3.873 ;
      RECT 52.14 3.725 52.226 3.868 ;
      RECT 52.118 3.718 52.14 3.862 ;
      RECT 52.032 3.709 52.118 3.856 ;
      RECT 51.946 3.696 52.032 3.847 ;
      RECT 51.86 3.682 51.946 3.837 ;
      RECT 51.815 3.672 51.86 3.83 ;
      RECT 51.795 2.96 51.815 3.238 ;
      RECT 51.795 3.665 51.815 3.826 ;
      RECT 51.765 2.96 51.795 3.26 ;
      RECT 51.755 3.632 51.795 3.823 ;
      RECT 51.75 2.96 51.765 3.28 ;
      RECT 51.75 3.597 51.755 3.821 ;
      RECT 51.745 2.96 51.75 3.405 ;
      RECT 51.745 3.557 51.75 3.821 ;
      RECT 51.735 2.96 51.745 3.821 ;
      RECT 51.66 2.96 51.735 3.815 ;
      RECT 51.63 2.96 51.66 3.805 ;
      RECT 51.625 2.96 51.63 3.797 ;
      RECT 51.62 3.002 51.625 3.79 ;
      RECT 51.61 3.071 51.62 3.781 ;
      RECT 51.605 3.141 51.61 3.733 ;
      RECT 51.6 3.205 51.605 3.63 ;
      RECT 51.595 3.24 51.6 3.585 ;
      RECT 51.593 3.277 51.595 3.477 ;
      RECT 51.59 3.285 51.593 3.47 ;
      RECT 51.585 3.35 51.59 3.413 ;
      RECT 55.66 2.44 55.94 2.72 ;
      RECT 55.65 2.44 55.94 2.583 ;
      RECT 55.605 2.305 55.865 2.565 ;
      RECT 55.605 2.42 55.92 2.565 ;
      RECT 55.605 2.39 55.915 2.565 ;
      RECT 55.605 2.377 55.905 2.565 ;
      RECT 55.605 2.367 55.9 2.565 ;
      RECT 51.58 2.35 51.84 2.61 ;
      RECT 55.35 1.9 55.61 2.16 ;
      RECT 55.34 1.925 55.61 2.12 ;
      RECT 55.335 1.925 55.34 2.119 ;
      RECT 55.265 1.92 55.335 2.111 ;
      RECT 55.18 1.907 55.265 2.094 ;
      RECT 55.176 1.899 55.18 2.084 ;
      RECT 55.09 1.892 55.176 2.074 ;
      RECT 55.081 1.884 55.09 2.064 ;
      RECT 54.995 1.877 55.081 2.052 ;
      RECT 54.975 1.868 54.995 2.038 ;
      RECT 54.92 1.863 54.975 2.03 ;
      RECT 54.91 1.857 54.92 2.024 ;
      RECT 54.89 1.855 54.91 2.02 ;
      RECT 54.882 1.854 54.89 2.016 ;
      RECT 54.796 1.846 54.882 2.005 ;
      RECT 54.71 1.832 54.796 1.985 ;
      RECT 54.65 1.82 54.71 1.97 ;
      RECT 54.64 1.815 54.65 1.965 ;
      RECT 54.59 1.815 54.64 1.967 ;
      RECT 54.543 1.817 54.59 1.971 ;
      RECT 54.457 1.824 54.543 1.976 ;
      RECT 54.371 1.832 54.457 1.982 ;
      RECT 54.285 1.841 54.371 1.988 ;
      RECT 54.226 1.847 54.285 1.993 ;
      RECT 54.14 1.852 54.226 1.999 ;
      RECT 54.065 1.857 54.14 2.005 ;
      RECT 54.026 1.859 54.065 2.01 ;
      RECT 53.94 1.856 54.026 2.015 ;
      RECT 53.855 1.854 53.94 2.022 ;
      RECT 53.823 1.853 53.855 2.025 ;
      RECT 53.737 1.852 53.823 2.026 ;
      RECT 53.651 1.851 53.737 2.027 ;
      RECT 53.565 1.85 53.651 2.027 ;
      RECT 53.479 1.849 53.565 2.028 ;
      RECT 53.393 1.848 53.479 2.029 ;
      RECT 53.307 1.847 53.393 2.03 ;
      RECT 53.221 1.846 53.307 2.03 ;
      RECT 53.135 1.845 53.221 2.031 ;
      RECT 53.085 1.845 53.135 2.032 ;
      RECT 53.071 1.846 53.085 2.032 ;
      RECT 52.985 1.853 53.071 2.033 ;
      RECT 52.911 1.864 52.985 2.034 ;
      RECT 52.825 1.873 52.911 2.035 ;
      RECT 52.79 1.88 52.825 2.05 ;
      RECT 52.765 1.883 52.79 2.08 ;
      RECT 52.74 1.892 52.765 2.109 ;
      RECT 52.73 1.903 52.74 2.129 ;
      RECT 52.72 1.911 52.73 2.143 ;
      RECT 52.715 1.917 52.72 2.153 ;
      RECT 52.69 1.934 52.715 2.17 ;
      RECT 52.675 1.956 52.69 2.198 ;
      RECT 52.645 1.982 52.675 2.228 ;
      RECT 52.625 2.011 52.645 2.258 ;
      RECT 52.62 2.026 52.625 2.275 ;
      RECT 52.6 2.041 52.62 2.29 ;
      RECT 52.59 2.059 52.6 2.308 ;
      RECT 52.58 2.07 52.59 2.323 ;
      RECT 52.53 2.102 52.58 2.349 ;
      RECT 52.525 2.132 52.53 2.369 ;
      RECT 52.515 2.145 52.525 2.375 ;
      RECT 52.506 2.155 52.515 2.383 ;
      RECT 52.495 2.166 52.506 2.391 ;
      RECT 52.49 2.176 52.495 2.397 ;
      RECT 52.475 2.197 52.49 2.404 ;
      RECT 52.46 2.227 52.475 2.412 ;
      RECT 52.425 2.257 52.46 2.418 ;
      RECT 52.4 2.275 52.425 2.425 ;
      RECT 52.35 2.283 52.4 2.434 ;
      RECT 52.325 2.288 52.35 2.443 ;
      RECT 52.27 2.294 52.325 2.453 ;
      RECT 52.265 2.299 52.27 2.461 ;
      RECT 52.251 2.302 52.265 2.463 ;
      RECT 52.165 2.314 52.251 2.475 ;
      RECT 52.155 2.326 52.165 2.488 ;
      RECT 52.07 2.339 52.155 2.5 ;
      RECT 52.026 2.356 52.07 2.514 ;
      RECT 51.94 2.373 52.026 2.53 ;
      RECT 51.91 2.387 51.94 2.544 ;
      RECT 51.9 2.392 51.91 2.549 ;
      RECT 51.84 2.395 51.9 2.558 ;
      RECT 54.73 2.665 54.99 2.925 ;
      RECT 54.73 2.665 55.01 2.778 ;
      RECT 54.73 2.665 55.035 2.745 ;
      RECT 54.73 2.665 55.04 2.725 ;
      RECT 54.78 2.44 55.06 2.72 ;
      RECT 54.335 3.175 54.595 3.435 ;
      RECT 54.325 3.032 54.52 3.373 ;
      RECT 54.32 3.14 54.535 3.365 ;
      RECT 54.315 3.19 54.595 3.355 ;
      RECT 54.305 3.267 54.595 3.34 ;
      RECT 54.325 3.115 54.535 3.373 ;
      RECT 54.335 2.99 54.52 3.435 ;
      RECT 54.335 2.885 54.5 3.435 ;
      RECT 54.345 2.872 54.5 3.435 ;
      RECT 54.345 2.83 54.49 3.435 ;
      RECT 54.35 2.755 54.49 3.435 ;
      RECT 54.38 2.405 54.49 3.435 ;
      RECT 54.385 2.135 54.51 2.758 ;
      RECT 54.355 2.71 54.51 2.758 ;
      RECT 54.37 2.512 54.49 3.435 ;
      RECT 54.36 2.622 54.51 2.758 ;
      RECT 54.385 2.135 54.525 2.615 ;
      RECT 54.385 2.135 54.545 2.49 ;
      RECT 54.35 2.135 54.61 2.395 ;
      RECT 53.82 2.44 54.1 2.72 ;
      RECT 53.805 2.44 54.1 2.7 ;
      RECT 51.86 3.305 52.12 3.565 ;
      RECT 53.645 3.16 53.905 3.42 ;
      RECT 53.625 3.18 53.905 3.395 ;
      RECT 53.582 3.18 53.625 3.394 ;
      RECT 53.496 3.181 53.582 3.391 ;
      RECT 53.41 3.182 53.496 3.387 ;
      RECT 53.335 3.184 53.41 3.384 ;
      RECT 53.312 3.185 53.335 3.382 ;
      RECT 53.226 3.186 53.312 3.38 ;
      RECT 53.14 3.187 53.226 3.377 ;
      RECT 53.116 3.188 53.14 3.375 ;
      RECT 53.03 3.19 53.116 3.372 ;
      RECT 52.945 3.192 53.03 3.373 ;
      RECT 52.888 3.193 52.945 3.379 ;
      RECT 52.802 3.195 52.888 3.389 ;
      RECT 52.716 3.198 52.802 3.402 ;
      RECT 52.63 3.2 52.716 3.414 ;
      RECT 52.616 3.201 52.63 3.421 ;
      RECT 52.53 3.202 52.616 3.429 ;
      RECT 52.49 3.204 52.53 3.438 ;
      RECT 52.481 3.205 52.49 3.441 ;
      RECT 52.395 3.213 52.481 3.447 ;
      RECT 52.375 3.222 52.395 3.455 ;
      RECT 52.29 3.237 52.375 3.463 ;
      RECT 52.23 3.26 52.29 3.474 ;
      RECT 52.22 3.272 52.23 3.479 ;
      RECT 52.18 3.282 52.22 3.483 ;
      RECT 52.125 3.299 52.18 3.491 ;
      RECT 52.12 3.309 52.125 3.495 ;
      RECT 53.186 2.44 53.245 2.837 ;
      RECT 53.1 2.44 53.305 2.828 ;
      RECT 53.095 2.47 53.305 2.823 ;
      RECT 53.061 2.47 53.305 2.821 ;
      RECT 52.975 2.47 53.305 2.815 ;
      RECT 52.93 2.47 53.325 2.793 ;
      RECT 52.93 2.47 53.345 2.748 ;
      RECT 52.89 2.47 53.345 2.738 ;
      RECT 53.1 2.44 53.38 2.72 ;
      RECT 52.835 2.44 53.095 2.7 ;
      RECT 52.02 1.92 52.28 2.18 ;
      RECT 52.1 1.88 52.38 2.16 ;
      RECT 46.465 6.22 46.785 6.545 ;
      RECT 46.495 5.695 46.665 6.545 ;
      RECT 46.495 5.695 46.67 6.045 ;
      RECT 46.495 5.695 47.47 5.87 ;
      RECT 47.295 1.965 47.47 5.87 ;
      RECT 47.24 1.965 47.59 2.315 ;
      RECT 47.265 6.655 47.59 6.98 ;
      RECT 46.15 6.745 47.59 6.915 ;
      RECT 46.15 2.395 46.31 6.915 ;
      RECT 46.465 2.365 46.785 2.685 ;
      RECT 46.15 2.395 46.785 2.565 ;
      RECT 34.875 3 35.155 3.28 ;
      RECT 34.845 3 35.155 3.265 ;
      RECT 34.84 3 35.155 3.263 ;
      RECT 34.835 1.33 35.005 3.257 ;
      RECT 34.83 2.967 35.1 3.25 ;
      RECT 34.825 3 35.155 3.243 ;
      RECT 34.795 2.97 35.1 3.23 ;
      RECT 34.795 2.997 35.12 3.23 ;
      RECT 34.795 2.987 35.115 3.23 ;
      RECT 34.795 2.972 35.11 3.23 ;
      RECT 34.835 2.962 35.1 3.257 ;
      RECT 34.835 2.957 35.09 3.257 ;
      RECT 34.835 2.956 35.075 3.257 ;
      RECT 44.805 1.34 45.155 1.69 ;
      RECT 44.8 1.34 45.155 1.595 ;
      RECT 34.835 1.33 45.045 1.5 ;
      RECT 44.48 2.85 44.85 3.22 ;
      RECT 44.565 2.235 44.735 3.22 ;
      RECT 40.585 2.455 40.82 2.715 ;
      RECT 43.73 2.235 43.895 2.495 ;
      RECT 43.635 2.225 43.65 2.495 ;
      RECT 43.73 2.235 44.735 2.415 ;
      RECT 42.235 1.795 42.275 1.935 ;
      RECT 43.65 2.23 43.73 2.495 ;
      RECT 43.595 2.225 43.635 2.461 ;
      RECT 43.581 2.225 43.595 2.461 ;
      RECT 43.495 2.23 43.581 2.463 ;
      RECT 43.45 2.237 43.495 2.465 ;
      RECT 43.42 2.237 43.45 2.467 ;
      RECT 43.395 2.232 43.42 2.469 ;
      RECT 43.365 2.228 43.395 2.478 ;
      RECT 43.355 2.225 43.365 2.49 ;
      RECT 43.35 2.225 43.355 2.498 ;
      RECT 43.345 2.225 43.35 2.503 ;
      RECT 43.335 2.224 43.345 2.513 ;
      RECT 43.33 2.223 43.335 2.523 ;
      RECT 43.315 2.222 43.33 2.528 ;
      RECT 43.287 2.219 43.315 2.555 ;
      RECT 43.201 2.211 43.287 2.555 ;
      RECT 43.115 2.2 43.201 2.555 ;
      RECT 43.075 2.185 43.115 2.555 ;
      RECT 43.035 2.159 43.075 2.555 ;
      RECT 43.03 2.141 43.035 2.367 ;
      RECT 43.02 2.137 43.03 2.357 ;
      RECT 43.005 2.127 43.02 2.344 ;
      RECT 42.985 2.111 43.005 2.329 ;
      RECT 42.97 2.096 42.985 2.314 ;
      RECT 42.96 2.085 42.97 2.304 ;
      RECT 42.935 2.069 42.96 2.293 ;
      RECT 42.93 2.056 42.935 2.283 ;
      RECT 42.925 2.052 42.93 2.278 ;
      RECT 42.87 2.038 42.925 2.256 ;
      RECT 42.831 2.019 42.87 2.22 ;
      RECT 42.745 1.993 42.831 2.173 ;
      RECT 42.741 1.975 42.745 2.139 ;
      RECT 42.655 1.956 42.741 2.117 ;
      RECT 42.65 1.938 42.655 2.095 ;
      RECT 42.645 1.936 42.65 2.093 ;
      RECT 42.635 1.935 42.645 2.088 ;
      RECT 42.575 1.922 42.635 2.074 ;
      RECT 42.53 1.9 42.575 2.053 ;
      RECT 42.47 1.877 42.53 2.032 ;
      RECT 42.406 1.852 42.47 2.007 ;
      RECT 42.32 1.822 42.406 1.976 ;
      RECT 42.305 1.802 42.32 1.955 ;
      RECT 42.275 1.797 42.305 1.946 ;
      RECT 42.222 1.795 42.235 1.935 ;
      RECT 42.136 1.795 42.222 1.937 ;
      RECT 42.05 1.795 42.136 1.939 ;
      RECT 42.03 1.795 42.05 1.943 ;
      RECT 41.985 1.797 42.03 1.954 ;
      RECT 41.945 1.807 41.985 1.97 ;
      RECT 41.941 1.816 41.945 1.978 ;
      RECT 41.855 1.836 41.941 1.994 ;
      RECT 41.845 1.855 41.855 2.012 ;
      RECT 41.84 1.857 41.845 2.015 ;
      RECT 41.83 1.861 41.84 2.018 ;
      RECT 41.81 1.866 41.83 2.028 ;
      RECT 41.78 1.876 41.81 2.048 ;
      RECT 41.775 1.883 41.78 2.062 ;
      RECT 41.765 1.887 41.775 2.069 ;
      RECT 41.75 1.895 41.765 2.08 ;
      RECT 41.74 1.905 41.75 2.091 ;
      RECT 41.73 1.912 41.74 2.099 ;
      RECT 41.705 1.925 41.73 2.114 ;
      RECT 41.641 1.961 41.705 2.153 ;
      RECT 41.555 2.024 41.641 2.217 ;
      RECT 41.52 2.075 41.555 2.27 ;
      RECT 41.515 2.092 41.52 2.287 ;
      RECT 41.5 2.101 41.515 2.294 ;
      RECT 41.48 2.116 41.5 2.308 ;
      RECT 41.475 2.127 41.48 2.318 ;
      RECT 41.455 2.14 41.475 2.328 ;
      RECT 41.45 2.15 41.455 2.338 ;
      RECT 41.435 2.155 41.45 2.347 ;
      RECT 41.425 2.165 41.435 2.358 ;
      RECT 41.395 2.182 41.425 2.375 ;
      RECT 41.385 2.2 41.395 2.393 ;
      RECT 41.37 2.211 41.385 2.404 ;
      RECT 41.33 2.235 41.37 2.42 ;
      RECT 41.295 2.269 41.33 2.437 ;
      RECT 41.265 2.292 41.295 2.449 ;
      RECT 41.25 2.302 41.265 2.458 ;
      RECT 41.21 2.312 41.25 2.469 ;
      RECT 41.19 2.323 41.21 2.481 ;
      RECT 41.185 2.327 41.19 2.488 ;
      RECT 41.17 2.331 41.185 2.493 ;
      RECT 41.16 2.336 41.17 2.498 ;
      RECT 41.155 2.339 41.16 2.501 ;
      RECT 41.125 2.345 41.155 2.508 ;
      RECT 41.09 2.355 41.125 2.522 ;
      RECT 41.03 2.37 41.09 2.542 ;
      RECT 40.975 2.39 41.03 2.566 ;
      RECT 40.946 2.405 40.975 2.584 ;
      RECT 40.86 2.425 40.946 2.609 ;
      RECT 40.855 2.44 40.86 2.629 ;
      RECT 40.845 2.443 40.855 2.63 ;
      RECT 40.82 2.45 40.845 2.715 ;
      RECT 43.515 2.943 43.795 3.28 ;
      RECT 43.515 2.953 43.8 3.238 ;
      RECT 43.515 2.962 43.805 3.135 ;
      RECT 43.515 2.977 43.81 3.003 ;
      RECT 43.515 2.805 43.775 3.28 ;
      RECT 33.87 6.66 34.22 7.01 ;
      RECT 42.695 6.615 43.045 6.965 ;
      RECT 33.87 6.69 43.045 6.89 ;
      RECT 41.235 3.685 41.245 3.875 ;
      RECT 39.495 3.56 39.775 3.84 ;
      RECT 42.54 2.5 42.545 2.985 ;
      RECT 42.435 2.5 42.495 2.76 ;
      RECT 42.76 3.47 42.765 3.545 ;
      RECT 42.75 3.337 42.76 3.58 ;
      RECT 42.74 3.172 42.75 3.601 ;
      RECT 42.735 3.042 42.74 3.617 ;
      RECT 42.725 2.932 42.735 3.633 ;
      RECT 42.72 2.831 42.725 3.65 ;
      RECT 42.715 2.813 42.72 3.66 ;
      RECT 42.71 2.795 42.715 3.67 ;
      RECT 42.7 2.77 42.71 3.685 ;
      RECT 42.695 2.75 42.7 3.7 ;
      RECT 42.675 2.5 42.695 3.725 ;
      RECT 42.66 2.5 42.675 3.758 ;
      RECT 42.63 2.5 42.66 3.78 ;
      RECT 42.61 2.5 42.63 3.794 ;
      RECT 42.59 2.5 42.61 3.31 ;
      RECT 42.605 3.377 42.61 3.799 ;
      RECT 42.6 3.407 42.605 3.801 ;
      RECT 42.595 3.42 42.6 3.804 ;
      RECT 42.59 3.43 42.595 3.808 ;
      RECT 42.585 2.5 42.59 3.228 ;
      RECT 42.585 3.44 42.59 3.81 ;
      RECT 42.58 2.5 42.585 3.205 ;
      RECT 42.57 3.462 42.585 3.81 ;
      RECT 42.565 2.5 42.58 3.15 ;
      RECT 42.56 3.487 42.57 3.81 ;
      RECT 42.56 2.5 42.565 3.095 ;
      RECT 42.55 2.5 42.56 3.043 ;
      RECT 42.555 3.5 42.56 3.811 ;
      RECT 42.55 3.512 42.555 3.812 ;
      RECT 42.545 2.5 42.55 3.003 ;
      RECT 42.545 3.525 42.55 3.813 ;
      RECT 42.53 3.54 42.545 3.814 ;
      RECT 42.535 2.5 42.54 2.965 ;
      RECT 42.53 2.5 42.535 2.93 ;
      RECT 42.525 2.5 42.53 2.905 ;
      RECT 42.52 3.567 42.53 3.816 ;
      RECT 42.515 2.5 42.525 2.863 ;
      RECT 42.515 3.585 42.52 3.817 ;
      RECT 42.51 2.5 42.515 2.823 ;
      RECT 42.51 3.592 42.515 3.818 ;
      RECT 42.505 2.5 42.51 2.795 ;
      RECT 42.5 3.61 42.51 3.819 ;
      RECT 42.495 2.5 42.505 2.775 ;
      RECT 42.49 3.63 42.5 3.821 ;
      RECT 42.48 3.647 42.49 3.822 ;
      RECT 42.445 3.67 42.48 3.825 ;
      RECT 42.39 3.688 42.445 3.831 ;
      RECT 42.304 3.696 42.39 3.84 ;
      RECT 42.218 3.707 42.304 3.851 ;
      RECT 42.132 3.717 42.218 3.862 ;
      RECT 42.046 3.727 42.132 3.874 ;
      RECT 41.96 3.737 42.046 3.885 ;
      RECT 41.94 3.743 41.96 3.891 ;
      RECT 41.86 3.745 41.94 3.895 ;
      RECT 41.855 3.744 41.86 3.9 ;
      RECT 41.847 3.743 41.855 3.9 ;
      RECT 41.761 3.739 41.847 3.898 ;
      RECT 41.675 3.731 41.761 3.895 ;
      RECT 41.589 3.722 41.675 3.891 ;
      RECT 41.503 3.714 41.589 3.888 ;
      RECT 41.417 3.706 41.503 3.884 ;
      RECT 41.331 3.697 41.417 3.881 ;
      RECT 41.245 3.689 41.331 3.877 ;
      RECT 41.19 3.682 41.235 3.875 ;
      RECT 41.105 3.675 41.19 3.873 ;
      RECT 41.031 3.667 41.105 3.869 ;
      RECT 40.945 3.659 41.031 3.866 ;
      RECT 40.942 3.655 40.945 3.864 ;
      RECT 40.856 3.651 40.942 3.863 ;
      RECT 40.77 3.643 40.856 3.86 ;
      RECT 40.685 3.638 40.77 3.857 ;
      RECT 40.599 3.635 40.685 3.854 ;
      RECT 40.513 3.633 40.599 3.851 ;
      RECT 40.427 3.63 40.513 3.848 ;
      RECT 40.341 3.627 40.427 3.845 ;
      RECT 40.255 3.624 40.341 3.842 ;
      RECT 40.179 3.622 40.255 3.839 ;
      RECT 40.093 3.619 40.179 3.836 ;
      RECT 40.007 3.616 40.093 3.834 ;
      RECT 39.921 3.614 40.007 3.831 ;
      RECT 39.835 3.611 39.921 3.828 ;
      RECT 39.775 3.602 39.835 3.826 ;
      RECT 42.285 3.22 42.36 3.48 ;
      RECT 42.265 3.2 42.27 3.48 ;
      RECT 41.585 2.985 41.69 3.28 ;
      RECT 36.03 2.96 36.1 3.22 ;
      RECT 41.925 2.835 41.93 3.206 ;
      RECT 41.915 2.89 41.92 3.206 ;
      RECT 42.22 2.06 42.28 2.32 ;
      RECT 42.275 3.215 42.285 3.48 ;
      RECT 42.27 3.205 42.275 3.48 ;
      RECT 42.19 3.152 42.265 3.48 ;
      RECT 42.215 2.06 42.22 2.34 ;
      RECT 42.205 2.06 42.215 2.36 ;
      RECT 42.19 2.06 42.205 2.39 ;
      RECT 42.175 2.06 42.19 2.433 ;
      RECT 42.17 3.095 42.19 3.48 ;
      RECT 42.16 2.06 42.175 2.47 ;
      RECT 42.155 3.075 42.17 3.48 ;
      RECT 42.155 2.06 42.16 2.493 ;
      RECT 42.145 2.06 42.155 2.518 ;
      RECT 42.115 3.042 42.155 3.48 ;
      RECT 42.12 2.06 42.145 2.568 ;
      RECT 42.115 2.06 42.12 2.623 ;
      RECT 42.11 2.06 42.115 2.665 ;
      RECT 42.1 3.005 42.115 3.48 ;
      RECT 42.105 2.06 42.11 2.708 ;
      RECT 42.1 2.06 42.105 2.773 ;
      RECT 42.095 2.06 42.1 2.795 ;
      RECT 42.095 2.993 42.1 3.345 ;
      RECT 42.09 2.06 42.095 2.863 ;
      RECT 42.09 2.985 42.095 3.328 ;
      RECT 42.085 2.06 42.09 2.908 ;
      RECT 42.08 2.967 42.09 3.305 ;
      RECT 42.08 2.06 42.085 2.945 ;
      RECT 42.07 2.06 42.08 3.285 ;
      RECT 42.065 2.06 42.07 3.268 ;
      RECT 42.06 2.06 42.065 3.253 ;
      RECT 42.055 2.06 42.06 3.238 ;
      RECT 42.035 2.06 42.055 3.228 ;
      RECT 42.03 2.06 42.035 3.218 ;
      RECT 42.02 2.06 42.03 3.214 ;
      RECT 42.015 2.337 42.02 3.213 ;
      RECT 42.01 2.36 42.015 3.212 ;
      RECT 42.005 2.39 42.01 3.211 ;
      RECT 42 2.417 42.005 3.21 ;
      RECT 41.995 2.445 42 3.21 ;
      RECT 41.99 2.472 41.995 3.21 ;
      RECT 41.985 2.492 41.99 3.21 ;
      RECT 41.98 2.52 41.985 3.21 ;
      RECT 41.97 2.562 41.98 3.21 ;
      RECT 41.96 2.607 41.97 3.209 ;
      RECT 41.955 2.66 41.96 3.208 ;
      RECT 41.95 2.692 41.955 3.207 ;
      RECT 41.945 2.712 41.95 3.206 ;
      RECT 41.94 2.75 41.945 3.206 ;
      RECT 41.935 2.772 41.94 3.206 ;
      RECT 41.93 2.797 41.935 3.206 ;
      RECT 41.92 2.862 41.925 3.206 ;
      RECT 41.905 2.922 41.915 3.206 ;
      RECT 41.89 2.932 41.905 3.206 ;
      RECT 41.87 2.942 41.89 3.206 ;
      RECT 41.84 2.947 41.87 3.203 ;
      RECT 41.78 2.957 41.84 3.2 ;
      RECT 41.76 2.966 41.78 3.205 ;
      RECT 41.735 2.972 41.76 3.218 ;
      RECT 41.715 2.977 41.735 3.233 ;
      RECT 41.69 2.982 41.715 3.28 ;
      RECT 41.561 2.984 41.585 3.28 ;
      RECT 41.475 2.979 41.561 3.28 ;
      RECT 41.435 2.976 41.475 3.28 ;
      RECT 41.385 2.978 41.435 3.26 ;
      RECT 41.355 2.982 41.385 3.26 ;
      RECT 41.276 2.992 41.355 3.26 ;
      RECT 41.19 3.007 41.276 3.261 ;
      RECT 41.14 3.017 41.19 3.262 ;
      RECT 41.132 3.02 41.14 3.262 ;
      RECT 41.046 3.022 41.132 3.263 ;
      RECT 40.96 3.026 41.046 3.263 ;
      RECT 40.874 3.03 40.96 3.264 ;
      RECT 40.788 3.033 40.874 3.265 ;
      RECT 40.702 3.037 40.788 3.265 ;
      RECT 40.616 3.041 40.702 3.266 ;
      RECT 40.53 3.044 40.616 3.267 ;
      RECT 40.444 3.048 40.53 3.267 ;
      RECT 40.358 3.052 40.444 3.268 ;
      RECT 40.272 3.056 40.358 3.269 ;
      RECT 40.186 3.059 40.272 3.269 ;
      RECT 40.1 3.063 40.186 3.27 ;
      RECT 40.07 3.065 40.1 3.27 ;
      RECT 39.984 3.068 40.07 3.271 ;
      RECT 39.898 3.072 39.984 3.272 ;
      RECT 39.812 3.076 39.898 3.273 ;
      RECT 39.726 3.079 39.812 3.273 ;
      RECT 39.64 3.083 39.726 3.274 ;
      RECT 39.605 3.088 39.64 3.275 ;
      RECT 39.55 3.098 39.605 3.282 ;
      RECT 39.525 3.11 39.55 3.292 ;
      RECT 39.49 3.123 39.525 3.3 ;
      RECT 39.45 3.14 39.49 3.323 ;
      RECT 39.43 3.153 39.45 3.35 ;
      RECT 39.4 3.165 39.43 3.378 ;
      RECT 39.395 3.173 39.4 3.398 ;
      RECT 39.39 3.176 39.395 3.408 ;
      RECT 39.34 3.188 39.39 3.442 ;
      RECT 39.33 3.203 39.34 3.475 ;
      RECT 39.32 3.209 39.33 3.488 ;
      RECT 39.31 3.216 39.32 3.5 ;
      RECT 39.285 3.229 39.31 3.518 ;
      RECT 39.27 3.244 39.285 3.54 ;
      RECT 39.26 3.252 39.27 3.556 ;
      RECT 39.245 3.261 39.26 3.571 ;
      RECT 39.235 3.271 39.245 3.585 ;
      RECT 39.216 3.284 39.235 3.602 ;
      RECT 39.13 3.329 39.216 3.667 ;
      RECT 39.115 3.374 39.13 3.725 ;
      RECT 39.11 3.383 39.115 3.738 ;
      RECT 39.1 3.39 39.11 3.743 ;
      RECT 39.095 3.395 39.1 3.747 ;
      RECT 39.075 3.405 39.095 3.754 ;
      RECT 39.05 3.425 39.075 3.768 ;
      RECT 39.015 3.45 39.05 3.788 ;
      RECT 39 3.473 39.015 3.803 ;
      RECT 38.99 3.483 39 3.808 ;
      RECT 38.98 3.491 38.99 3.815 ;
      RECT 38.97 3.5 38.98 3.821 ;
      RECT 38.95 3.512 38.97 3.823 ;
      RECT 38.94 3.525 38.95 3.825 ;
      RECT 38.915 3.54 38.94 3.828 ;
      RECT 38.895 3.557 38.915 3.832 ;
      RECT 38.855 3.585 38.895 3.838 ;
      RECT 38.79 3.632 38.855 3.847 ;
      RECT 38.775 3.665 38.79 3.855 ;
      RECT 38.77 3.672 38.775 3.857 ;
      RECT 38.72 3.697 38.77 3.862 ;
      RECT 38.705 3.721 38.72 3.869 ;
      RECT 38.655 3.726 38.705 3.87 ;
      RECT 38.569 3.73 38.655 3.87 ;
      RECT 38.483 3.73 38.569 3.87 ;
      RECT 38.397 3.73 38.483 3.871 ;
      RECT 38.311 3.73 38.397 3.871 ;
      RECT 38.225 3.73 38.311 3.871 ;
      RECT 38.159 3.73 38.225 3.871 ;
      RECT 38.073 3.73 38.159 3.872 ;
      RECT 37.987 3.73 38.073 3.872 ;
      RECT 37.901 3.731 37.987 3.873 ;
      RECT 37.815 3.731 37.901 3.873 ;
      RECT 37.729 3.731 37.815 3.873 ;
      RECT 37.643 3.731 37.729 3.874 ;
      RECT 37.557 3.731 37.643 3.874 ;
      RECT 37.471 3.732 37.557 3.875 ;
      RECT 37.385 3.732 37.471 3.875 ;
      RECT 37.365 3.732 37.385 3.875 ;
      RECT 37.279 3.732 37.365 3.875 ;
      RECT 37.193 3.732 37.279 3.875 ;
      RECT 37.107 3.733 37.193 3.875 ;
      RECT 37.021 3.733 37.107 3.875 ;
      RECT 36.935 3.733 37.021 3.875 ;
      RECT 36.849 3.734 36.935 3.875 ;
      RECT 36.763 3.734 36.849 3.875 ;
      RECT 36.677 3.734 36.763 3.875 ;
      RECT 36.591 3.734 36.677 3.875 ;
      RECT 36.505 3.735 36.591 3.875 ;
      RECT 36.455 3.732 36.505 3.875 ;
      RECT 36.445 3.73 36.455 3.874 ;
      RECT 36.441 3.73 36.445 3.873 ;
      RECT 36.355 3.725 36.441 3.868 ;
      RECT 36.333 3.718 36.355 3.862 ;
      RECT 36.247 3.709 36.333 3.856 ;
      RECT 36.161 3.696 36.247 3.847 ;
      RECT 36.075 3.682 36.161 3.837 ;
      RECT 36.03 3.672 36.075 3.83 ;
      RECT 36.01 2.96 36.03 3.238 ;
      RECT 36.01 3.665 36.03 3.826 ;
      RECT 35.98 2.96 36.01 3.26 ;
      RECT 35.97 3.632 36.01 3.823 ;
      RECT 35.965 2.96 35.98 3.28 ;
      RECT 35.965 3.597 35.97 3.821 ;
      RECT 35.96 2.96 35.965 3.405 ;
      RECT 35.96 3.557 35.965 3.821 ;
      RECT 35.95 2.96 35.96 3.821 ;
      RECT 35.875 2.96 35.95 3.815 ;
      RECT 35.845 2.96 35.875 3.805 ;
      RECT 35.84 2.96 35.845 3.797 ;
      RECT 35.835 3.002 35.84 3.79 ;
      RECT 35.825 3.071 35.835 3.781 ;
      RECT 35.82 3.141 35.825 3.733 ;
      RECT 35.815 3.205 35.82 3.63 ;
      RECT 35.81 3.24 35.815 3.585 ;
      RECT 35.808 3.277 35.81 3.477 ;
      RECT 35.805 3.285 35.808 3.47 ;
      RECT 35.8 3.35 35.805 3.413 ;
      RECT 39.875 2.44 40.155 2.72 ;
      RECT 39.865 2.44 40.155 2.583 ;
      RECT 39.82 2.305 40.08 2.565 ;
      RECT 39.82 2.42 40.135 2.565 ;
      RECT 39.82 2.39 40.13 2.565 ;
      RECT 39.82 2.377 40.12 2.565 ;
      RECT 39.82 2.367 40.115 2.565 ;
      RECT 35.795 2.35 36.055 2.61 ;
      RECT 39.565 1.9 39.825 2.16 ;
      RECT 39.555 1.925 39.825 2.12 ;
      RECT 39.55 1.925 39.555 2.119 ;
      RECT 39.48 1.92 39.55 2.111 ;
      RECT 39.395 1.907 39.48 2.094 ;
      RECT 39.391 1.899 39.395 2.084 ;
      RECT 39.305 1.892 39.391 2.074 ;
      RECT 39.296 1.884 39.305 2.064 ;
      RECT 39.21 1.877 39.296 2.052 ;
      RECT 39.19 1.868 39.21 2.038 ;
      RECT 39.135 1.863 39.19 2.03 ;
      RECT 39.125 1.857 39.135 2.024 ;
      RECT 39.105 1.855 39.125 2.02 ;
      RECT 39.097 1.854 39.105 2.016 ;
      RECT 39.011 1.846 39.097 2.005 ;
      RECT 38.925 1.832 39.011 1.985 ;
      RECT 38.865 1.82 38.925 1.97 ;
      RECT 38.855 1.815 38.865 1.965 ;
      RECT 38.805 1.815 38.855 1.967 ;
      RECT 38.758 1.817 38.805 1.971 ;
      RECT 38.672 1.824 38.758 1.976 ;
      RECT 38.586 1.832 38.672 1.982 ;
      RECT 38.5 1.841 38.586 1.988 ;
      RECT 38.441 1.847 38.5 1.993 ;
      RECT 38.355 1.852 38.441 1.999 ;
      RECT 38.28 1.857 38.355 2.005 ;
      RECT 38.241 1.859 38.28 2.01 ;
      RECT 38.155 1.856 38.241 2.015 ;
      RECT 38.07 1.854 38.155 2.022 ;
      RECT 38.038 1.853 38.07 2.025 ;
      RECT 37.952 1.852 38.038 2.026 ;
      RECT 37.866 1.851 37.952 2.027 ;
      RECT 37.78 1.85 37.866 2.027 ;
      RECT 37.694 1.849 37.78 2.028 ;
      RECT 37.608 1.848 37.694 2.029 ;
      RECT 37.522 1.847 37.608 2.03 ;
      RECT 37.436 1.846 37.522 2.03 ;
      RECT 37.35 1.845 37.436 2.031 ;
      RECT 37.3 1.845 37.35 2.032 ;
      RECT 37.286 1.846 37.3 2.032 ;
      RECT 37.2 1.853 37.286 2.033 ;
      RECT 37.126 1.864 37.2 2.034 ;
      RECT 37.04 1.873 37.126 2.035 ;
      RECT 37.005 1.88 37.04 2.05 ;
      RECT 36.98 1.883 37.005 2.08 ;
      RECT 36.955 1.892 36.98 2.109 ;
      RECT 36.945 1.903 36.955 2.129 ;
      RECT 36.935 1.911 36.945 2.143 ;
      RECT 36.93 1.917 36.935 2.153 ;
      RECT 36.905 1.934 36.93 2.17 ;
      RECT 36.89 1.956 36.905 2.198 ;
      RECT 36.86 1.982 36.89 2.228 ;
      RECT 36.84 2.011 36.86 2.258 ;
      RECT 36.835 2.026 36.84 2.275 ;
      RECT 36.815 2.041 36.835 2.29 ;
      RECT 36.805 2.059 36.815 2.308 ;
      RECT 36.795 2.07 36.805 2.323 ;
      RECT 36.745 2.102 36.795 2.349 ;
      RECT 36.74 2.132 36.745 2.369 ;
      RECT 36.73 2.145 36.74 2.375 ;
      RECT 36.721 2.155 36.73 2.383 ;
      RECT 36.71 2.166 36.721 2.391 ;
      RECT 36.705 2.176 36.71 2.397 ;
      RECT 36.69 2.197 36.705 2.404 ;
      RECT 36.675 2.227 36.69 2.412 ;
      RECT 36.64 2.257 36.675 2.418 ;
      RECT 36.615 2.275 36.64 2.425 ;
      RECT 36.565 2.283 36.615 2.434 ;
      RECT 36.54 2.288 36.565 2.443 ;
      RECT 36.485 2.294 36.54 2.453 ;
      RECT 36.48 2.299 36.485 2.461 ;
      RECT 36.466 2.302 36.48 2.463 ;
      RECT 36.38 2.314 36.466 2.475 ;
      RECT 36.37 2.326 36.38 2.488 ;
      RECT 36.285 2.339 36.37 2.5 ;
      RECT 36.241 2.356 36.285 2.514 ;
      RECT 36.155 2.373 36.241 2.53 ;
      RECT 36.125 2.387 36.155 2.544 ;
      RECT 36.115 2.392 36.125 2.549 ;
      RECT 36.055 2.395 36.115 2.558 ;
      RECT 38.945 2.665 39.205 2.925 ;
      RECT 38.945 2.665 39.225 2.778 ;
      RECT 38.945 2.665 39.25 2.745 ;
      RECT 38.945 2.665 39.255 2.725 ;
      RECT 38.995 2.44 39.275 2.72 ;
      RECT 38.55 3.175 38.81 3.435 ;
      RECT 38.54 3.032 38.735 3.373 ;
      RECT 38.535 3.14 38.75 3.365 ;
      RECT 38.53 3.19 38.81 3.355 ;
      RECT 38.52 3.267 38.81 3.34 ;
      RECT 38.54 3.115 38.75 3.373 ;
      RECT 38.55 2.99 38.735 3.435 ;
      RECT 38.55 2.885 38.715 3.435 ;
      RECT 38.56 2.872 38.715 3.435 ;
      RECT 38.56 2.83 38.705 3.435 ;
      RECT 38.565 2.755 38.705 3.435 ;
      RECT 38.595 2.405 38.705 3.435 ;
      RECT 38.6 2.135 38.725 2.758 ;
      RECT 38.57 2.71 38.725 2.758 ;
      RECT 38.585 2.512 38.705 3.435 ;
      RECT 38.575 2.622 38.725 2.758 ;
      RECT 38.6 2.135 38.74 2.615 ;
      RECT 38.6 2.135 38.76 2.49 ;
      RECT 38.565 2.135 38.825 2.395 ;
      RECT 38.035 2.44 38.315 2.72 ;
      RECT 38.02 2.44 38.315 2.7 ;
      RECT 36.075 3.305 36.335 3.565 ;
      RECT 37.86 3.16 38.12 3.42 ;
      RECT 37.84 3.18 38.12 3.395 ;
      RECT 37.797 3.18 37.84 3.394 ;
      RECT 37.711 3.181 37.797 3.391 ;
      RECT 37.625 3.182 37.711 3.387 ;
      RECT 37.55 3.184 37.625 3.384 ;
      RECT 37.527 3.185 37.55 3.382 ;
      RECT 37.441 3.186 37.527 3.38 ;
      RECT 37.355 3.187 37.441 3.377 ;
      RECT 37.331 3.188 37.355 3.375 ;
      RECT 37.245 3.19 37.331 3.372 ;
      RECT 37.16 3.192 37.245 3.373 ;
      RECT 37.103 3.193 37.16 3.379 ;
      RECT 37.017 3.195 37.103 3.389 ;
      RECT 36.931 3.198 37.017 3.402 ;
      RECT 36.845 3.2 36.931 3.414 ;
      RECT 36.831 3.201 36.845 3.421 ;
      RECT 36.745 3.202 36.831 3.429 ;
      RECT 36.705 3.204 36.745 3.438 ;
      RECT 36.696 3.205 36.705 3.441 ;
      RECT 36.61 3.213 36.696 3.447 ;
      RECT 36.59 3.222 36.61 3.455 ;
      RECT 36.505 3.237 36.59 3.463 ;
      RECT 36.445 3.26 36.505 3.474 ;
      RECT 36.435 3.272 36.445 3.479 ;
      RECT 36.395 3.282 36.435 3.483 ;
      RECT 36.34 3.299 36.395 3.491 ;
      RECT 36.335 3.309 36.34 3.495 ;
      RECT 37.401 2.44 37.46 2.837 ;
      RECT 37.315 2.44 37.52 2.828 ;
      RECT 37.31 2.47 37.52 2.823 ;
      RECT 37.276 2.47 37.52 2.821 ;
      RECT 37.19 2.47 37.52 2.815 ;
      RECT 37.145 2.47 37.54 2.793 ;
      RECT 37.145 2.47 37.56 2.748 ;
      RECT 37.105 2.47 37.56 2.738 ;
      RECT 37.315 2.44 37.595 2.72 ;
      RECT 37.05 2.44 37.31 2.7 ;
      RECT 36.235 1.92 36.495 2.18 ;
      RECT 36.315 1.88 36.595 2.16 ;
      RECT 30.69 6.22 31.01 6.545 ;
      RECT 30.72 5.695 30.89 6.545 ;
      RECT 30.72 5.695 30.895 6.045 ;
      RECT 30.72 5.695 31.695 5.87 ;
      RECT 31.52 1.965 31.695 5.87 ;
      RECT 31.465 1.965 31.815 2.315 ;
      RECT 31.49 6.655 31.815 6.98 ;
      RECT 30.375 6.745 31.815 6.915 ;
      RECT 30.375 2.395 30.535 6.915 ;
      RECT 30.69 2.365 31.01 2.685 ;
      RECT 30.375 2.395 31.01 2.565 ;
      RECT 19.1 3 19.38 3.28 ;
      RECT 19.07 3 19.38 3.265 ;
      RECT 19.065 3 19.38 3.263 ;
      RECT 19.06 1.33 19.23 3.257 ;
      RECT 19.055 2.967 19.325 3.25 ;
      RECT 19.05 3 19.38 3.243 ;
      RECT 19.02 2.97 19.325 3.23 ;
      RECT 19.02 2.997 19.345 3.23 ;
      RECT 19.02 2.987 19.34 3.23 ;
      RECT 19.02 2.972 19.335 3.23 ;
      RECT 19.06 2.962 19.325 3.257 ;
      RECT 19.06 2.957 19.315 3.257 ;
      RECT 19.06 2.956 19.3 3.257 ;
      RECT 29.03 1.34 29.38 1.69 ;
      RECT 29.025 1.34 29.38 1.595 ;
      RECT 19.06 1.33 29.27 1.5 ;
      RECT 28.705 2.85 29.075 3.22 ;
      RECT 28.79 2.235 28.96 3.22 ;
      RECT 24.81 2.455 25.045 2.715 ;
      RECT 27.955 2.235 28.12 2.495 ;
      RECT 27.86 2.225 27.875 2.495 ;
      RECT 27.955 2.235 28.96 2.415 ;
      RECT 26.46 1.795 26.5 1.935 ;
      RECT 27.875 2.23 27.955 2.495 ;
      RECT 27.82 2.225 27.86 2.461 ;
      RECT 27.806 2.225 27.82 2.461 ;
      RECT 27.72 2.23 27.806 2.463 ;
      RECT 27.675 2.237 27.72 2.465 ;
      RECT 27.645 2.237 27.675 2.467 ;
      RECT 27.62 2.232 27.645 2.469 ;
      RECT 27.59 2.228 27.62 2.478 ;
      RECT 27.58 2.225 27.59 2.49 ;
      RECT 27.575 2.225 27.58 2.498 ;
      RECT 27.57 2.225 27.575 2.503 ;
      RECT 27.56 2.224 27.57 2.513 ;
      RECT 27.555 2.223 27.56 2.523 ;
      RECT 27.54 2.222 27.555 2.528 ;
      RECT 27.512 2.219 27.54 2.555 ;
      RECT 27.426 2.211 27.512 2.555 ;
      RECT 27.34 2.2 27.426 2.555 ;
      RECT 27.3 2.185 27.34 2.555 ;
      RECT 27.26 2.159 27.3 2.555 ;
      RECT 27.255 2.141 27.26 2.367 ;
      RECT 27.245 2.137 27.255 2.357 ;
      RECT 27.23 2.127 27.245 2.344 ;
      RECT 27.21 2.111 27.23 2.329 ;
      RECT 27.195 2.096 27.21 2.314 ;
      RECT 27.185 2.085 27.195 2.304 ;
      RECT 27.16 2.069 27.185 2.293 ;
      RECT 27.155 2.056 27.16 2.283 ;
      RECT 27.15 2.052 27.155 2.278 ;
      RECT 27.095 2.038 27.15 2.256 ;
      RECT 27.056 2.019 27.095 2.22 ;
      RECT 26.97 1.993 27.056 2.173 ;
      RECT 26.966 1.975 26.97 2.139 ;
      RECT 26.88 1.956 26.966 2.117 ;
      RECT 26.875 1.938 26.88 2.095 ;
      RECT 26.87 1.936 26.875 2.093 ;
      RECT 26.86 1.935 26.87 2.088 ;
      RECT 26.8 1.922 26.86 2.074 ;
      RECT 26.755 1.9 26.8 2.053 ;
      RECT 26.695 1.877 26.755 2.032 ;
      RECT 26.631 1.852 26.695 2.007 ;
      RECT 26.545 1.822 26.631 1.976 ;
      RECT 26.53 1.802 26.545 1.955 ;
      RECT 26.5 1.797 26.53 1.946 ;
      RECT 26.447 1.795 26.46 1.935 ;
      RECT 26.361 1.795 26.447 1.937 ;
      RECT 26.275 1.795 26.361 1.939 ;
      RECT 26.255 1.795 26.275 1.943 ;
      RECT 26.21 1.797 26.255 1.954 ;
      RECT 26.17 1.807 26.21 1.97 ;
      RECT 26.166 1.816 26.17 1.978 ;
      RECT 26.08 1.836 26.166 1.994 ;
      RECT 26.07 1.855 26.08 2.012 ;
      RECT 26.065 1.857 26.07 2.015 ;
      RECT 26.055 1.861 26.065 2.018 ;
      RECT 26.035 1.866 26.055 2.028 ;
      RECT 26.005 1.876 26.035 2.048 ;
      RECT 26 1.883 26.005 2.062 ;
      RECT 25.99 1.887 26 2.069 ;
      RECT 25.975 1.895 25.99 2.08 ;
      RECT 25.965 1.905 25.975 2.091 ;
      RECT 25.955 1.912 25.965 2.099 ;
      RECT 25.93 1.925 25.955 2.114 ;
      RECT 25.866 1.961 25.93 2.153 ;
      RECT 25.78 2.024 25.866 2.217 ;
      RECT 25.745 2.075 25.78 2.27 ;
      RECT 25.74 2.092 25.745 2.287 ;
      RECT 25.725 2.101 25.74 2.294 ;
      RECT 25.705 2.116 25.725 2.308 ;
      RECT 25.7 2.127 25.705 2.318 ;
      RECT 25.68 2.14 25.7 2.328 ;
      RECT 25.675 2.15 25.68 2.338 ;
      RECT 25.66 2.155 25.675 2.347 ;
      RECT 25.65 2.165 25.66 2.358 ;
      RECT 25.62 2.182 25.65 2.375 ;
      RECT 25.61 2.2 25.62 2.393 ;
      RECT 25.595 2.211 25.61 2.404 ;
      RECT 25.555 2.235 25.595 2.42 ;
      RECT 25.52 2.269 25.555 2.437 ;
      RECT 25.49 2.292 25.52 2.449 ;
      RECT 25.475 2.302 25.49 2.458 ;
      RECT 25.435 2.312 25.475 2.469 ;
      RECT 25.415 2.323 25.435 2.481 ;
      RECT 25.41 2.327 25.415 2.488 ;
      RECT 25.395 2.331 25.41 2.493 ;
      RECT 25.385 2.336 25.395 2.498 ;
      RECT 25.38 2.339 25.385 2.501 ;
      RECT 25.35 2.345 25.38 2.508 ;
      RECT 25.315 2.355 25.35 2.522 ;
      RECT 25.255 2.37 25.315 2.542 ;
      RECT 25.2 2.39 25.255 2.566 ;
      RECT 25.171 2.405 25.2 2.584 ;
      RECT 25.085 2.425 25.171 2.609 ;
      RECT 25.08 2.44 25.085 2.629 ;
      RECT 25.07 2.443 25.08 2.63 ;
      RECT 25.045 2.45 25.07 2.715 ;
      RECT 27.74 2.943 28.02 3.28 ;
      RECT 27.74 2.953 28.025 3.238 ;
      RECT 27.74 2.962 28.03 3.135 ;
      RECT 27.74 2.977 28.035 3.003 ;
      RECT 27.74 2.805 28 3.28 ;
      RECT 18.09 6.655 18.44 7.005 ;
      RECT 26.915 6.61 27.265 6.96 ;
      RECT 18.09 6.685 27.265 6.885 ;
      RECT 25.46 3.685 25.47 3.875 ;
      RECT 23.72 3.56 24 3.84 ;
      RECT 26.765 2.5 26.77 2.985 ;
      RECT 26.66 2.5 26.72 2.76 ;
      RECT 26.985 3.47 26.99 3.545 ;
      RECT 26.975 3.337 26.985 3.58 ;
      RECT 26.965 3.172 26.975 3.601 ;
      RECT 26.96 3.042 26.965 3.617 ;
      RECT 26.95 2.932 26.96 3.633 ;
      RECT 26.945 2.831 26.95 3.65 ;
      RECT 26.94 2.813 26.945 3.66 ;
      RECT 26.935 2.795 26.94 3.67 ;
      RECT 26.925 2.77 26.935 3.685 ;
      RECT 26.92 2.75 26.925 3.7 ;
      RECT 26.9 2.5 26.92 3.725 ;
      RECT 26.885 2.5 26.9 3.758 ;
      RECT 26.855 2.5 26.885 3.78 ;
      RECT 26.835 2.5 26.855 3.794 ;
      RECT 26.815 2.5 26.835 3.31 ;
      RECT 26.83 3.377 26.835 3.799 ;
      RECT 26.825 3.407 26.83 3.801 ;
      RECT 26.82 3.42 26.825 3.804 ;
      RECT 26.815 3.43 26.82 3.808 ;
      RECT 26.81 2.5 26.815 3.228 ;
      RECT 26.81 3.44 26.815 3.81 ;
      RECT 26.805 2.5 26.81 3.205 ;
      RECT 26.795 3.462 26.81 3.81 ;
      RECT 26.79 2.5 26.805 3.15 ;
      RECT 26.785 3.487 26.795 3.81 ;
      RECT 26.785 2.5 26.79 3.095 ;
      RECT 26.775 2.5 26.785 3.043 ;
      RECT 26.78 3.5 26.785 3.811 ;
      RECT 26.775 3.512 26.78 3.812 ;
      RECT 26.77 2.5 26.775 3.003 ;
      RECT 26.77 3.525 26.775 3.813 ;
      RECT 26.755 3.54 26.77 3.814 ;
      RECT 26.76 2.5 26.765 2.965 ;
      RECT 26.755 2.5 26.76 2.93 ;
      RECT 26.75 2.5 26.755 2.905 ;
      RECT 26.745 3.567 26.755 3.816 ;
      RECT 26.74 2.5 26.75 2.863 ;
      RECT 26.74 3.585 26.745 3.817 ;
      RECT 26.735 2.5 26.74 2.823 ;
      RECT 26.735 3.592 26.74 3.818 ;
      RECT 26.73 2.5 26.735 2.795 ;
      RECT 26.725 3.61 26.735 3.819 ;
      RECT 26.72 2.5 26.73 2.775 ;
      RECT 26.715 3.63 26.725 3.821 ;
      RECT 26.705 3.647 26.715 3.822 ;
      RECT 26.67 3.67 26.705 3.825 ;
      RECT 26.615 3.688 26.67 3.831 ;
      RECT 26.529 3.696 26.615 3.84 ;
      RECT 26.443 3.707 26.529 3.851 ;
      RECT 26.357 3.717 26.443 3.862 ;
      RECT 26.271 3.727 26.357 3.874 ;
      RECT 26.185 3.737 26.271 3.885 ;
      RECT 26.165 3.743 26.185 3.891 ;
      RECT 26.085 3.745 26.165 3.895 ;
      RECT 26.08 3.744 26.085 3.9 ;
      RECT 26.072 3.743 26.08 3.9 ;
      RECT 25.986 3.739 26.072 3.898 ;
      RECT 25.9 3.731 25.986 3.895 ;
      RECT 25.814 3.722 25.9 3.891 ;
      RECT 25.728 3.714 25.814 3.888 ;
      RECT 25.642 3.706 25.728 3.884 ;
      RECT 25.556 3.697 25.642 3.881 ;
      RECT 25.47 3.689 25.556 3.877 ;
      RECT 25.415 3.682 25.46 3.875 ;
      RECT 25.33 3.675 25.415 3.873 ;
      RECT 25.256 3.667 25.33 3.869 ;
      RECT 25.17 3.659 25.256 3.866 ;
      RECT 25.167 3.655 25.17 3.864 ;
      RECT 25.081 3.651 25.167 3.863 ;
      RECT 24.995 3.643 25.081 3.86 ;
      RECT 24.91 3.638 24.995 3.857 ;
      RECT 24.824 3.635 24.91 3.854 ;
      RECT 24.738 3.633 24.824 3.851 ;
      RECT 24.652 3.63 24.738 3.848 ;
      RECT 24.566 3.627 24.652 3.845 ;
      RECT 24.48 3.624 24.566 3.842 ;
      RECT 24.404 3.622 24.48 3.839 ;
      RECT 24.318 3.619 24.404 3.836 ;
      RECT 24.232 3.616 24.318 3.834 ;
      RECT 24.146 3.614 24.232 3.831 ;
      RECT 24.06 3.611 24.146 3.828 ;
      RECT 24 3.602 24.06 3.826 ;
      RECT 26.51 3.22 26.585 3.48 ;
      RECT 26.49 3.2 26.495 3.48 ;
      RECT 25.81 2.985 25.915 3.28 ;
      RECT 20.255 2.96 20.325 3.22 ;
      RECT 26.15 2.835 26.155 3.206 ;
      RECT 26.14 2.89 26.145 3.206 ;
      RECT 26.445 2.06 26.505 2.32 ;
      RECT 26.5 3.215 26.51 3.48 ;
      RECT 26.495 3.205 26.5 3.48 ;
      RECT 26.415 3.152 26.49 3.48 ;
      RECT 26.44 2.06 26.445 2.34 ;
      RECT 26.43 2.06 26.44 2.36 ;
      RECT 26.415 2.06 26.43 2.39 ;
      RECT 26.4 2.06 26.415 2.433 ;
      RECT 26.395 3.095 26.415 3.48 ;
      RECT 26.385 2.06 26.4 2.47 ;
      RECT 26.38 3.075 26.395 3.48 ;
      RECT 26.38 2.06 26.385 2.493 ;
      RECT 26.37 2.06 26.38 2.518 ;
      RECT 26.34 3.042 26.38 3.48 ;
      RECT 26.345 2.06 26.37 2.568 ;
      RECT 26.34 2.06 26.345 2.623 ;
      RECT 26.335 2.06 26.34 2.665 ;
      RECT 26.325 3.005 26.34 3.48 ;
      RECT 26.33 2.06 26.335 2.708 ;
      RECT 26.325 2.06 26.33 2.773 ;
      RECT 26.32 2.06 26.325 2.795 ;
      RECT 26.32 2.993 26.325 3.345 ;
      RECT 26.315 2.06 26.32 2.863 ;
      RECT 26.315 2.985 26.32 3.328 ;
      RECT 26.31 2.06 26.315 2.908 ;
      RECT 26.305 2.967 26.315 3.305 ;
      RECT 26.305 2.06 26.31 2.945 ;
      RECT 26.295 2.06 26.305 3.285 ;
      RECT 26.29 2.06 26.295 3.268 ;
      RECT 26.285 2.06 26.29 3.253 ;
      RECT 26.28 2.06 26.285 3.238 ;
      RECT 26.26 2.06 26.28 3.228 ;
      RECT 26.255 2.06 26.26 3.218 ;
      RECT 26.245 2.06 26.255 3.214 ;
      RECT 26.24 2.337 26.245 3.213 ;
      RECT 26.235 2.36 26.24 3.212 ;
      RECT 26.23 2.39 26.235 3.211 ;
      RECT 26.225 2.417 26.23 3.21 ;
      RECT 26.22 2.445 26.225 3.21 ;
      RECT 26.215 2.472 26.22 3.21 ;
      RECT 26.21 2.492 26.215 3.21 ;
      RECT 26.205 2.52 26.21 3.21 ;
      RECT 26.195 2.562 26.205 3.21 ;
      RECT 26.185 2.607 26.195 3.209 ;
      RECT 26.18 2.66 26.185 3.208 ;
      RECT 26.175 2.692 26.18 3.207 ;
      RECT 26.17 2.712 26.175 3.206 ;
      RECT 26.165 2.75 26.17 3.206 ;
      RECT 26.16 2.772 26.165 3.206 ;
      RECT 26.155 2.797 26.16 3.206 ;
      RECT 26.145 2.862 26.15 3.206 ;
      RECT 26.13 2.922 26.14 3.206 ;
      RECT 26.115 2.932 26.13 3.206 ;
      RECT 26.095 2.942 26.115 3.206 ;
      RECT 26.065 2.947 26.095 3.203 ;
      RECT 26.005 2.957 26.065 3.2 ;
      RECT 25.985 2.966 26.005 3.205 ;
      RECT 25.96 2.972 25.985 3.218 ;
      RECT 25.94 2.977 25.96 3.233 ;
      RECT 25.915 2.982 25.94 3.28 ;
      RECT 25.786 2.984 25.81 3.28 ;
      RECT 25.7 2.979 25.786 3.28 ;
      RECT 25.66 2.976 25.7 3.28 ;
      RECT 25.61 2.978 25.66 3.26 ;
      RECT 25.58 2.982 25.61 3.26 ;
      RECT 25.501 2.992 25.58 3.26 ;
      RECT 25.415 3.007 25.501 3.261 ;
      RECT 25.365 3.017 25.415 3.262 ;
      RECT 25.357 3.02 25.365 3.262 ;
      RECT 25.271 3.022 25.357 3.263 ;
      RECT 25.185 3.026 25.271 3.263 ;
      RECT 25.099 3.03 25.185 3.264 ;
      RECT 25.013 3.033 25.099 3.265 ;
      RECT 24.927 3.037 25.013 3.265 ;
      RECT 24.841 3.041 24.927 3.266 ;
      RECT 24.755 3.044 24.841 3.267 ;
      RECT 24.669 3.048 24.755 3.267 ;
      RECT 24.583 3.052 24.669 3.268 ;
      RECT 24.497 3.056 24.583 3.269 ;
      RECT 24.411 3.059 24.497 3.269 ;
      RECT 24.325 3.063 24.411 3.27 ;
      RECT 24.295 3.065 24.325 3.27 ;
      RECT 24.209 3.068 24.295 3.271 ;
      RECT 24.123 3.072 24.209 3.272 ;
      RECT 24.037 3.076 24.123 3.273 ;
      RECT 23.951 3.079 24.037 3.273 ;
      RECT 23.865 3.083 23.951 3.274 ;
      RECT 23.83 3.088 23.865 3.275 ;
      RECT 23.775 3.098 23.83 3.282 ;
      RECT 23.75 3.11 23.775 3.292 ;
      RECT 23.715 3.123 23.75 3.3 ;
      RECT 23.675 3.14 23.715 3.323 ;
      RECT 23.655 3.153 23.675 3.35 ;
      RECT 23.625 3.165 23.655 3.378 ;
      RECT 23.62 3.173 23.625 3.398 ;
      RECT 23.615 3.176 23.62 3.408 ;
      RECT 23.565 3.188 23.615 3.442 ;
      RECT 23.555 3.203 23.565 3.475 ;
      RECT 23.545 3.209 23.555 3.488 ;
      RECT 23.535 3.216 23.545 3.5 ;
      RECT 23.51 3.229 23.535 3.518 ;
      RECT 23.495 3.244 23.51 3.54 ;
      RECT 23.485 3.252 23.495 3.556 ;
      RECT 23.47 3.261 23.485 3.571 ;
      RECT 23.46 3.271 23.47 3.585 ;
      RECT 23.441 3.284 23.46 3.602 ;
      RECT 23.355 3.329 23.441 3.667 ;
      RECT 23.34 3.374 23.355 3.725 ;
      RECT 23.335 3.383 23.34 3.738 ;
      RECT 23.325 3.39 23.335 3.743 ;
      RECT 23.32 3.395 23.325 3.747 ;
      RECT 23.3 3.405 23.32 3.754 ;
      RECT 23.275 3.425 23.3 3.768 ;
      RECT 23.24 3.45 23.275 3.788 ;
      RECT 23.225 3.473 23.24 3.803 ;
      RECT 23.215 3.483 23.225 3.808 ;
      RECT 23.205 3.491 23.215 3.815 ;
      RECT 23.195 3.5 23.205 3.821 ;
      RECT 23.175 3.512 23.195 3.823 ;
      RECT 23.165 3.525 23.175 3.825 ;
      RECT 23.14 3.54 23.165 3.828 ;
      RECT 23.12 3.557 23.14 3.832 ;
      RECT 23.08 3.585 23.12 3.838 ;
      RECT 23.015 3.632 23.08 3.847 ;
      RECT 23 3.665 23.015 3.855 ;
      RECT 22.995 3.672 23 3.857 ;
      RECT 22.945 3.697 22.995 3.862 ;
      RECT 22.93 3.721 22.945 3.869 ;
      RECT 22.88 3.726 22.93 3.87 ;
      RECT 22.794 3.73 22.88 3.87 ;
      RECT 22.708 3.73 22.794 3.87 ;
      RECT 22.622 3.73 22.708 3.871 ;
      RECT 22.536 3.73 22.622 3.871 ;
      RECT 22.45 3.73 22.536 3.871 ;
      RECT 22.384 3.73 22.45 3.871 ;
      RECT 22.298 3.73 22.384 3.872 ;
      RECT 22.212 3.73 22.298 3.872 ;
      RECT 22.126 3.731 22.212 3.873 ;
      RECT 22.04 3.731 22.126 3.873 ;
      RECT 21.954 3.731 22.04 3.873 ;
      RECT 21.868 3.731 21.954 3.874 ;
      RECT 21.782 3.731 21.868 3.874 ;
      RECT 21.696 3.732 21.782 3.875 ;
      RECT 21.61 3.732 21.696 3.875 ;
      RECT 21.59 3.732 21.61 3.875 ;
      RECT 21.504 3.732 21.59 3.875 ;
      RECT 21.418 3.732 21.504 3.875 ;
      RECT 21.332 3.733 21.418 3.875 ;
      RECT 21.246 3.733 21.332 3.875 ;
      RECT 21.16 3.733 21.246 3.875 ;
      RECT 21.074 3.734 21.16 3.875 ;
      RECT 20.988 3.734 21.074 3.875 ;
      RECT 20.902 3.734 20.988 3.875 ;
      RECT 20.816 3.734 20.902 3.875 ;
      RECT 20.73 3.735 20.816 3.875 ;
      RECT 20.68 3.732 20.73 3.875 ;
      RECT 20.67 3.73 20.68 3.874 ;
      RECT 20.666 3.73 20.67 3.873 ;
      RECT 20.58 3.725 20.666 3.868 ;
      RECT 20.558 3.718 20.58 3.862 ;
      RECT 20.472 3.709 20.558 3.856 ;
      RECT 20.386 3.696 20.472 3.847 ;
      RECT 20.3 3.682 20.386 3.837 ;
      RECT 20.255 3.672 20.3 3.83 ;
      RECT 20.235 2.96 20.255 3.238 ;
      RECT 20.235 3.665 20.255 3.826 ;
      RECT 20.205 2.96 20.235 3.26 ;
      RECT 20.195 3.632 20.235 3.823 ;
      RECT 20.19 2.96 20.205 3.28 ;
      RECT 20.19 3.597 20.195 3.821 ;
      RECT 20.185 2.96 20.19 3.405 ;
      RECT 20.185 3.557 20.19 3.821 ;
      RECT 20.175 2.96 20.185 3.821 ;
      RECT 20.1 2.96 20.175 3.815 ;
      RECT 20.07 2.96 20.1 3.805 ;
      RECT 20.065 2.96 20.07 3.797 ;
      RECT 20.06 3.002 20.065 3.79 ;
      RECT 20.05 3.071 20.06 3.781 ;
      RECT 20.045 3.141 20.05 3.733 ;
      RECT 20.04 3.205 20.045 3.63 ;
      RECT 20.035 3.24 20.04 3.585 ;
      RECT 20.033 3.277 20.035 3.477 ;
      RECT 20.03 3.285 20.033 3.47 ;
      RECT 20.025 3.35 20.03 3.413 ;
      RECT 24.1 2.44 24.38 2.72 ;
      RECT 24.09 2.44 24.38 2.583 ;
      RECT 24.045 2.305 24.305 2.565 ;
      RECT 24.045 2.42 24.36 2.565 ;
      RECT 24.045 2.39 24.355 2.565 ;
      RECT 24.045 2.377 24.345 2.565 ;
      RECT 24.045 2.367 24.34 2.565 ;
      RECT 20.02 2.35 20.28 2.61 ;
      RECT 23.79 1.9 24.05 2.16 ;
      RECT 23.78 1.925 24.05 2.12 ;
      RECT 23.775 1.925 23.78 2.119 ;
      RECT 23.705 1.92 23.775 2.111 ;
      RECT 23.62 1.907 23.705 2.094 ;
      RECT 23.616 1.899 23.62 2.084 ;
      RECT 23.53 1.892 23.616 2.074 ;
      RECT 23.521 1.884 23.53 2.064 ;
      RECT 23.435 1.877 23.521 2.052 ;
      RECT 23.415 1.868 23.435 2.038 ;
      RECT 23.36 1.863 23.415 2.03 ;
      RECT 23.35 1.857 23.36 2.024 ;
      RECT 23.33 1.855 23.35 2.02 ;
      RECT 23.322 1.854 23.33 2.016 ;
      RECT 23.236 1.846 23.322 2.005 ;
      RECT 23.15 1.832 23.236 1.985 ;
      RECT 23.09 1.82 23.15 1.97 ;
      RECT 23.08 1.815 23.09 1.965 ;
      RECT 23.03 1.815 23.08 1.967 ;
      RECT 22.983 1.817 23.03 1.971 ;
      RECT 22.897 1.824 22.983 1.976 ;
      RECT 22.811 1.832 22.897 1.982 ;
      RECT 22.725 1.841 22.811 1.988 ;
      RECT 22.666 1.847 22.725 1.993 ;
      RECT 22.58 1.852 22.666 1.999 ;
      RECT 22.505 1.857 22.58 2.005 ;
      RECT 22.466 1.859 22.505 2.01 ;
      RECT 22.38 1.856 22.466 2.015 ;
      RECT 22.295 1.854 22.38 2.022 ;
      RECT 22.263 1.853 22.295 2.025 ;
      RECT 22.177 1.852 22.263 2.026 ;
      RECT 22.091 1.851 22.177 2.027 ;
      RECT 22.005 1.85 22.091 2.027 ;
      RECT 21.919 1.849 22.005 2.028 ;
      RECT 21.833 1.848 21.919 2.029 ;
      RECT 21.747 1.847 21.833 2.03 ;
      RECT 21.661 1.846 21.747 2.03 ;
      RECT 21.575 1.845 21.661 2.031 ;
      RECT 21.525 1.845 21.575 2.032 ;
      RECT 21.511 1.846 21.525 2.032 ;
      RECT 21.425 1.853 21.511 2.033 ;
      RECT 21.351 1.864 21.425 2.034 ;
      RECT 21.265 1.873 21.351 2.035 ;
      RECT 21.23 1.88 21.265 2.05 ;
      RECT 21.205 1.883 21.23 2.08 ;
      RECT 21.18 1.892 21.205 2.109 ;
      RECT 21.17 1.903 21.18 2.129 ;
      RECT 21.16 1.911 21.17 2.143 ;
      RECT 21.155 1.917 21.16 2.153 ;
      RECT 21.13 1.934 21.155 2.17 ;
      RECT 21.115 1.956 21.13 2.198 ;
      RECT 21.085 1.982 21.115 2.228 ;
      RECT 21.065 2.011 21.085 2.258 ;
      RECT 21.06 2.026 21.065 2.275 ;
      RECT 21.04 2.041 21.06 2.29 ;
      RECT 21.03 2.059 21.04 2.308 ;
      RECT 21.02 2.07 21.03 2.323 ;
      RECT 20.97 2.102 21.02 2.349 ;
      RECT 20.965 2.132 20.97 2.369 ;
      RECT 20.955 2.145 20.965 2.375 ;
      RECT 20.946 2.155 20.955 2.383 ;
      RECT 20.935 2.166 20.946 2.391 ;
      RECT 20.93 2.176 20.935 2.397 ;
      RECT 20.915 2.197 20.93 2.404 ;
      RECT 20.9 2.227 20.915 2.412 ;
      RECT 20.865 2.257 20.9 2.418 ;
      RECT 20.84 2.275 20.865 2.425 ;
      RECT 20.79 2.283 20.84 2.434 ;
      RECT 20.765 2.288 20.79 2.443 ;
      RECT 20.71 2.294 20.765 2.453 ;
      RECT 20.705 2.299 20.71 2.461 ;
      RECT 20.691 2.302 20.705 2.463 ;
      RECT 20.605 2.314 20.691 2.475 ;
      RECT 20.595 2.326 20.605 2.488 ;
      RECT 20.51 2.339 20.595 2.5 ;
      RECT 20.466 2.356 20.51 2.514 ;
      RECT 20.38 2.373 20.466 2.53 ;
      RECT 20.35 2.387 20.38 2.544 ;
      RECT 20.34 2.392 20.35 2.549 ;
      RECT 20.28 2.395 20.34 2.558 ;
      RECT 23.17 2.665 23.43 2.925 ;
      RECT 23.17 2.665 23.45 2.778 ;
      RECT 23.17 2.665 23.475 2.745 ;
      RECT 23.17 2.665 23.48 2.725 ;
      RECT 23.22 2.44 23.5 2.72 ;
      RECT 22.775 3.175 23.035 3.435 ;
      RECT 22.765 3.032 22.96 3.373 ;
      RECT 22.76 3.14 22.975 3.365 ;
      RECT 22.755 3.19 23.035 3.355 ;
      RECT 22.745 3.267 23.035 3.34 ;
      RECT 22.765 3.115 22.975 3.373 ;
      RECT 22.775 2.99 22.96 3.435 ;
      RECT 22.775 2.885 22.94 3.435 ;
      RECT 22.785 2.872 22.94 3.435 ;
      RECT 22.785 2.83 22.93 3.435 ;
      RECT 22.79 2.755 22.93 3.435 ;
      RECT 22.82 2.405 22.93 3.435 ;
      RECT 22.825 2.135 22.95 2.758 ;
      RECT 22.795 2.71 22.95 2.758 ;
      RECT 22.81 2.512 22.93 3.435 ;
      RECT 22.8 2.622 22.95 2.758 ;
      RECT 22.825 2.135 22.965 2.615 ;
      RECT 22.825 2.135 22.985 2.49 ;
      RECT 22.79 2.135 23.05 2.395 ;
      RECT 22.26 2.44 22.54 2.72 ;
      RECT 22.245 2.44 22.54 2.7 ;
      RECT 20.3 3.305 20.56 3.565 ;
      RECT 22.085 3.16 22.345 3.42 ;
      RECT 22.065 3.18 22.345 3.395 ;
      RECT 22.022 3.18 22.065 3.394 ;
      RECT 21.936 3.181 22.022 3.391 ;
      RECT 21.85 3.182 21.936 3.387 ;
      RECT 21.775 3.184 21.85 3.384 ;
      RECT 21.752 3.185 21.775 3.382 ;
      RECT 21.666 3.186 21.752 3.38 ;
      RECT 21.58 3.187 21.666 3.377 ;
      RECT 21.556 3.188 21.58 3.375 ;
      RECT 21.47 3.19 21.556 3.372 ;
      RECT 21.385 3.192 21.47 3.373 ;
      RECT 21.328 3.193 21.385 3.379 ;
      RECT 21.242 3.195 21.328 3.389 ;
      RECT 21.156 3.198 21.242 3.402 ;
      RECT 21.07 3.2 21.156 3.414 ;
      RECT 21.056 3.201 21.07 3.421 ;
      RECT 20.97 3.202 21.056 3.429 ;
      RECT 20.93 3.204 20.97 3.438 ;
      RECT 20.921 3.205 20.93 3.441 ;
      RECT 20.835 3.213 20.921 3.447 ;
      RECT 20.815 3.222 20.835 3.455 ;
      RECT 20.73 3.237 20.815 3.463 ;
      RECT 20.67 3.26 20.73 3.474 ;
      RECT 20.66 3.272 20.67 3.479 ;
      RECT 20.62 3.282 20.66 3.483 ;
      RECT 20.565 3.299 20.62 3.491 ;
      RECT 20.56 3.309 20.565 3.495 ;
      RECT 21.626 2.44 21.685 2.837 ;
      RECT 21.54 2.44 21.745 2.828 ;
      RECT 21.535 2.47 21.745 2.823 ;
      RECT 21.501 2.47 21.745 2.821 ;
      RECT 21.415 2.47 21.745 2.815 ;
      RECT 21.37 2.47 21.765 2.793 ;
      RECT 21.37 2.47 21.785 2.748 ;
      RECT 21.33 2.47 21.785 2.738 ;
      RECT 21.54 2.44 21.82 2.72 ;
      RECT 21.275 2.44 21.535 2.7 ;
      RECT 20.46 1.92 20.72 2.18 ;
      RECT 20.54 1.88 20.82 2.16 ;
      RECT 14.91 6.22 15.23 6.545 ;
      RECT 14.94 5.695 15.11 6.545 ;
      RECT 14.94 5.695 15.115 6.045 ;
      RECT 14.94 5.695 15.915 5.87 ;
      RECT 15.74 1.965 15.915 5.87 ;
      RECT 15.685 1.965 16.035 2.315 ;
      RECT 15.71 6.655 16.035 6.98 ;
      RECT 14.595 6.745 16.035 6.915 ;
      RECT 14.595 2.395 14.755 6.915 ;
      RECT 14.91 2.365 15.23 2.685 ;
      RECT 14.595 2.395 15.23 2.565 ;
      RECT 3.32 3 3.6 3.28 ;
      RECT 3.29 3 3.6 3.265 ;
      RECT 3.285 3 3.6 3.263 ;
      RECT 3.28 1.33 3.45 3.257 ;
      RECT 3.275 2.967 3.545 3.25 ;
      RECT 3.27 3 3.6 3.243 ;
      RECT 3.24 2.97 3.545 3.23 ;
      RECT 3.24 2.997 3.565 3.23 ;
      RECT 3.24 2.987 3.56 3.23 ;
      RECT 3.24 2.972 3.555 3.23 ;
      RECT 3.28 2.962 3.545 3.257 ;
      RECT 3.28 2.957 3.535 3.257 ;
      RECT 3.28 2.956 3.52 3.257 ;
      RECT 13.25 1.34 13.6 1.69 ;
      RECT 13.245 1.34 13.6 1.595 ;
      RECT 3.28 1.33 13.49 1.5 ;
      RECT 12.925 2.85 13.295 3.22 ;
      RECT 13.01 2.235 13.18 3.22 ;
      RECT 9.03 2.455 9.265 2.715 ;
      RECT 12.175 2.235 12.34 2.495 ;
      RECT 12.08 2.225 12.095 2.495 ;
      RECT 12.175 2.235 13.18 2.415 ;
      RECT 10.68 1.795 10.72 1.935 ;
      RECT 12.095 2.23 12.175 2.495 ;
      RECT 12.04 2.225 12.08 2.461 ;
      RECT 12.026 2.225 12.04 2.461 ;
      RECT 11.94 2.23 12.026 2.463 ;
      RECT 11.895 2.237 11.94 2.465 ;
      RECT 11.865 2.237 11.895 2.467 ;
      RECT 11.84 2.232 11.865 2.469 ;
      RECT 11.81 2.228 11.84 2.478 ;
      RECT 11.8 2.225 11.81 2.49 ;
      RECT 11.795 2.225 11.8 2.498 ;
      RECT 11.79 2.225 11.795 2.503 ;
      RECT 11.78 2.224 11.79 2.513 ;
      RECT 11.775 2.223 11.78 2.523 ;
      RECT 11.76 2.222 11.775 2.528 ;
      RECT 11.732 2.219 11.76 2.555 ;
      RECT 11.646 2.211 11.732 2.555 ;
      RECT 11.56 2.2 11.646 2.555 ;
      RECT 11.52 2.185 11.56 2.555 ;
      RECT 11.48 2.159 11.52 2.555 ;
      RECT 11.475 2.141 11.48 2.367 ;
      RECT 11.465 2.137 11.475 2.357 ;
      RECT 11.45 2.127 11.465 2.344 ;
      RECT 11.43 2.111 11.45 2.329 ;
      RECT 11.415 2.096 11.43 2.314 ;
      RECT 11.405 2.085 11.415 2.304 ;
      RECT 11.38 2.069 11.405 2.293 ;
      RECT 11.375 2.056 11.38 2.283 ;
      RECT 11.37 2.052 11.375 2.278 ;
      RECT 11.315 2.038 11.37 2.256 ;
      RECT 11.276 2.019 11.315 2.22 ;
      RECT 11.19 1.993 11.276 2.173 ;
      RECT 11.186 1.975 11.19 2.139 ;
      RECT 11.1 1.956 11.186 2.117 ;
      RECT 11.095 1.938 11.1 2.095 ;
      RECT 11.09 1.936 11.095 2.093 ;
      RECT 11.08 1.935 11.09 2.088 ;
      RECT 11.02 1.922 11.08 2.074 ;
      RECT 10.975 1.9 11.02 2.053 ;
      RECT 10.915 1.877 10.975 2.032 ;
      RECT 10.851 1.852 10.915 2.007 ;
      RECT 10.765 1.822 10.851 1.976 ;
      RECT 10.75 1.802 10.765 1.955 ;
      RECT 10.72 1.797 10.75 1.946 ;
      RECT 10.667 1.795 10.68 1.935 ;
      RECT 10.581 1.795 10.667 1.937 ;
      RECT 10.495 1.795 10.581 1.939 ;
      RECT 10.475 1.795 10.495 1.943 ;
      RECT 10.43 1.797 10.475 1.954 ;
      RECT 10.39 1.807 10.43 1.97 ;
      RECT 10.386 1.816 10.39 1.978 ;
      RECT 10.3 1.836 10.386 1.994 ;
      RECT 10.29 1.855 10.3 2.012 ;
      RECT 10.285 1.857 10.29 2.015 ;
      RECT 10.275 1.861 10.285 2.018 ;
      RECT 10.255 1.866 10.275 2.028 ;
      RECT 10.225 1.876 10.255 2.048 ;
      RECT 10.22 1.883 10.225 2.062 ;
      RECT 10.21 1.887 10.22 2.069 ;
      RECT 10.195 1.895 10.21 2.08 ;
      RECT 10.185 1.905 10.195 2.091 ;
      RECT 10.175 1.912 10.185 2.099 ;
      RECT 10.15 1.925 10.175 2.114 ;
      RECT 10.086 1.961 10.15 2.153 ;
      RECT 10 2.024 10.086 2.217 ;
      RECT 9.965 2.075 10 2.27 ;
      RECT 9.96 2.092 9.965 2.287 ;
      RECT 9.945 2.101 9.96 2.294 ;
      RECT 9.925 2.116 9.945 2.308 ;
      RECT 9.92 2.127 9.925 2.318 ;
      RECT 9.9 2.14 9.92 2.328 ;
      RECT 9.895 2.15 9.9 2.338 ;
      RECT 9.88 2.155 9.895 2.347 ;
      RECT 9.87 2.165 9.88 2.358 ;
      RECT 9.84 2.182 9.87 2.375 ;
      RECT 9.83 2.2 9.84 2.393 ;
      RECT 9.815 2.211 9.83 2.404 ;
      RECT 9.775 2.235 9.815 2.42 ;
      RECT 9.74 2.269 9.775 2.437 ;
      RECT 9.71 2.292 9.74 2.449 ;
      RECT 9.695 2.302 9.71 2.458 ;
      RECT 9.655 2.312 9.695 2.469 ;
      RECT 9.635 2.323 9.655 2.481 ;
      RECT 9.63 2.327 9.635 2.488 ;
      RECT 9.615 2.331 9.63 2.493 ;
      RECT 9.605 2.336 9.615 2.498 ;
      RECT 9.6 2.339 9.605 2.501 ;
      RECT 9.57 2.345 9.6 2.508 ;
      RECT 9.535 2.355 9.57 2.522 ;
      RECT 9.475 2.37 9.535 2.542 ;
      RECT 9.42 2.39 9.475 2.566 ;
      RECT 9.391 2.405 9.42 2.584 ;
      RECT 9.305 2.425 9.391 2.609 ;
      RECT 9.3 2.44 9.305 2.629 ;
      RECT 9.29 2.443 9.3 2.63 ;
      RECT 9.265 2.45 9.29 2.715 ;
      RECT 11.96 2.943 12.24 3.28 ;
      RECT 11.96 2.953 12.245 3.238 ;
      RECT 11.96 2.962 12.25 3.135 ;
      RECT 11.96 2.977 12.255 3.003 ;
      RECT 11.96 2.805 12.22 3.28 ;
      RECT 1.54 6.995 1.83 7.345 ;
      RECT 1.54 7.055 2.955 7.225 ;
      RECT 2.785 6.685 2.955 7.225 ;
      RECT 11.105 6.605 11.455 6.955 ;
      RECT 2.785 6.685 11.455 6.855 ;
      RECT 9.68 3.685 9.69 3.875 ;
      RECT 7.94 3.56 8.22 3.84 ;
      RECT 10.985 2.5 10.99 2.985 ;
      RECT 10.88 2.5 10.94 2.76 ;
      RECT 11.205 3.47 11.21 3.545 ;
      RECT 11.195 3.337 11.205 3.58 ;
      RECT 11.185 3.172 11.195 3.601 ;
      RECT 11.18 3.042 11.185 3.617 ;
      RECT 11.17 2.932 11.18 3.633 ;
      RECT 11.165 2.831 11.17 3.65 ;
      RECT 11.16 2.813 11.165 3.66 ;
      RECT 11.155 2.795 11.16 3.67 ;
      RECT 11.145 2.77 11.155 3.685 ;
      RECT 11.14 2.75 11.145 3.7 ;
      RECT 11.12 2.5 11.14 3.725 ;
      RECT 11.105 2.5 11.12 3.758 ;
      RECT 11.075 2.5 11.105 3.78 ;
      RECT 11.055 2.5 11.075 3.794 ;
      RECT 11.035 2.5 11.055 3.31 ;
      RECT 11.05 3.377 11.055 3.799 ;
      RECT 11.045 3.407 11.05 3.801 ;
      RECT 11.04 3.42 11.045 3.804 ;
      RECT 11.035 3.43 11.04 3.808 ;
      RECT 11.03 2.5 11.035 3.228 ;
      RECT 11.03 3.44 11.035 3.81 ;
      RECT 11.025 2.5 11.03 3.205 ;
      RECT 11.015 3.462 11.03 3.81 ;
      RECT 11.01 2.5 11.025 3.15 ;
      RECT 11.005 3.487 11.015 3.81 ;
      RECT 11.005 2.5 11.01 3.095 ;
      RECT 10.995 2.5 11.005 3.043 ;
      RECT 11 3.5 11.005 3.811 ;
      RECT 10.995 3.512 11 3.812 ;
      RECT 10.99 2.5 10.995 3.003 ;
      RECT 10.99 3.525 10.995 3.813 ;
      RECT 10.975 3.54 10.99 3.814 ;
      RECT 10.98 2.5 10.985 2.965 ;
      RECT 10.975 2.5 10.98 2.93 ;
      RECT 10.97 2.5 10.975 2.905 ;
      RECT 10.965 3.567 10.975 3.816 ;
      RECT 10.96 2.5 10.97 2.863 ;
      RECT 10.96 3.585 10.965 3.817 ;
      RECT 10.955 2.5 10.96 2.823 ;
      RECT 10.955 3.592 10.96 3.818 ;
      RECT 10.95 2.5 10.955 2.795 ;
      RECT 10.945 3.61 10.955 3.819 ;
      RECT 10.94 2.5 10.95 2.775 ;
      RECT 10.935 3.63 10.945 3.821 ;
      RECT 10.925 3.647 10.935 3.822 ;
      RECT 10.89 3.67 10.925 3.825 ;
      RECT 10.835 3.688 10.89 3.831 ;
      RECT 10.749 3.696 10.835 3.84 ;
      RECT 10.663 3.707 10.749 3.851 ;
      RECT 10.577 3.717 10.663 3.862 ;
      RECT 10.491 3.727 10.577 3.874 ;
      RECT 10.405 3.737 10.491 3.885 ;
      RECT 10.385 3.743 10.405 3.891 ;
      RECT 10.305 3.745 10.385 3.895 ;
      RECT 10.3 3.744 10.305 3.9 ;
      RECT 10.292 3.743 10.3 3.9 ;
      RECT 10.206 3.739 10.292 3.898 ;
      RECT 10.12 3.731 10.206 3.895 ;
      RECT 10.034 3.722 10.12 3.891 ;
      RECT 9.948 3.714 10.034 3.888 ;
      RECT 9.862 3.706 9.948 3.884 ;
      RECT 9.776 3.697 9.862 3.881 ;
      RECT 9.69 3.689 9.776 3.877 ;
      RECT 9.635 3.682 9.68 3.875 ;
      RECT 9.55 3.675 9.635 3.873 ;
      RECT 9.476 3.667 9.55 3.869 ;
      RECT 9.39 3.659 9.476 3.866 ;
      RECT 9.387 3.655 9.39 3.864 ;
      RECT 9.301 3.651 9.387 3.863 ;
      RECT 9.215 3.643 9.301 3.86 ;
      RECT 9.13 3.638 9.215 3.857 ;
      RECT 9.044 3.635 9.13 3.854 ;
      RECT 8.958 3.633 9.044 3.851 ;
      RECT 8.872 3.63 8.958 3.848 ;
      RECT 8.786 3.627 8.872 3.845 ;
      RECT 8.7 3.624 8.786 3.842 ;
      RECT 8.624 3.622 8.7 3.839 ;
      RECT 8.538 3.619 8.624 3.836 ;
      RECT 8.452 3.616 8.538 3.834 ;
      RECT 8.366 3.614 8.452 3.831 ;
      RECT 8.28 3.611 8.366 3.828 ;
      RECT 8.22 3.602 8.28 3.826 ;
      RECT 10.73 3.22 10.805 3.48 ;
      RECT 10.71 3.2 10.715 3.48 ;
      RECT 10.03 2.985 10.135 3.28 ;
      RECT 4.475 2.96 4.545 3.22 ;
      RECT 10.37 2.835 10.375 3.206 ;
      RECT 10.36 2.89 10.365 3.206 ;
      RECT 10.665 2.06 10.725 2.32 ;
      RECT 10.72 3.215 10.73 3.48 ;
      RECT 10.715 3.205 10.72 3.48 ;
      RECT 10.635 3.152 10.71 3.48 ;
      RECT 10.66 2.06 10.665 2.34 ;
      RECT 10.65 2.06 10.66 2.36 ;
      RECT 10.635 2.06 10.65 2.39 ;
      RECT 10.62 2.06 10.635 2.433 ;
      RECT 10.615 3.095 10.635 3.48 ;
      RECT 10.605 2.06 10.62 2.47 ;
      RECT 10.6 3.075 10.615 3.48 ;
      RECT 10.6 2.06 10.605 2.493 ;
      RECT 10.59 2.06 10.6 2.518 ;
      RECT 10.56 3.042 10.6 3.48 ;
      RECT 10.565 2.06 10.59 2.568 ;
      RECT 10.56 2.06 10.565 2.623 ;
      RECT 10.555 2.06 10.56 2.665 ;
      RECT 10.545 3.005 10.56 3.48 ;
      RECT 10.55 2.06 10.555 2.708 ;
      RECT 10.545 2.06 10.55 2.773 ;
      RECT 10.54 2.06 10.545 2.795 ;
      RECT 10.54 2.993 10.545 3.345 ;
      RECT 10.535 2.06 10.54 2.863 ;
      RECT 10.535 2.985 10.54 3.328 ;
      RECT 10.53 2.06 10.535 2.908 ;
      RECT 10.525 2.967 10.535 3.305 ;
      RECT 10.525 2.06 10.53 2.945 ;
      RECT 10.515 2.06 10.525 3.285 ;
      RECT 10.51 2.06 10.515 3.268 ;
      RECT 10.505 2.06 10.51 3.253 ;
      RECT 10.5 2.06 10.505 3.238 ;
      RECT 10.48 2.06 10.5 3.228 ;
      RECT 10.475 2.06 10.48 3.218 ;
      RECT 10.465 2.06 10.475 3.214 ;
      RECT 10.46 2.337 10.465 3.213 ;
      RECT 10.455 2.36 10.46 3.212 ;
      RECT 10.45 2.39 10.455 3.211 ;
      RECT 10.445 2.417 10.45 3.21 ;
      RECT 10.44 2.445 10.445 3.21 ;
      RECT 10.435 2.472 10.44 3.21 ;
      RECT 10.43 2.492 10.435 3.21 ;
      RECT 10.425 2.52 10.43 3.21 ;
      RECT 10.415 2.562 10.425 3.21 ;
      RECT 10.405 2.607 10.415 3.209 ;
      RECT 10.4 2.66 10.405 3.208 ;
      RECT 10.395 2.692 10.4 3.207 ;
      RECT 10.39 2.712 10.395 3.206 ;
      RECT 10.385 2.75 10.39 3.206 ;
      RECT 10.38 2.772 10.385 3.206 ;
      RECT 10.375 2.797 10.38 3.206 ;
      RECT 10.365 2.862 10.37 3.206 ;
      RECT 10.35 2.922 10.36 3.206 ;
      RECT 10.335 2.932 10.35 3.206 ;
      RECT 10.315 2.942 10.335 3.206 ;
      RECT 10.285 2.947 10.315 3.203 ;
      RECT 10.225 2.957 10.285 3.2 ;
      RECT 10.205 2.966 10.225 3.205 ;
      RECT 10.18 2.972 10.205 3.218 ;
      RECT 10.16 2.977 10.18 3.233 ;
      RECT 10.135 2.982 10.16 3.28 ;
      RECT 10.006 2.984 10.03 3.28 ;
      RECT 9.92 2.979 10.006 3.28 ;
      RECT 9.88 2.976 9.92 3.28 ;
      RECT 9.83 2.978 9.88 3.26 ;
      RECT 9.8 2.982 9.83 3.26 ;
      RECT 9.721 2.992 9.8 3.26 ;
      RECT 9.635 3.007 9.721 3.261 ;
      RECT 9.585 3.017 9.635 3.262 ;
      RECT 9.577 3.02 9.585 3.262 ;
      RECT 9.491 3.022 9.577 3.263 ;
      RECT 9.405 3.026 9.491 3.263 ;
      RECT 9.319 3.03 9.405 3.264 ;
      RECT 9.233 3.033 9.319 3.265 ;
      RECT 9.147 3.037 9.233 3.265 ;
      RECT 9.061 3.041 9.147 3.266 ;
      RECT 8.975 3.044 9.061 3.267 ;
      RECT 8.889 3.048 8.975 3.267 ;
      RECT 8.803 3.052 8.889 3.268 ;
      RECT 8.717 3.056 8.803 3.269 ;
      RECT 8.631 3.059 8.717 3.269 ;
      RECT 8.545 3.063 8.631 3.27 ;
      RECT 8.515 3.065 8.545 3.27 ;
      RECT 8.429 3.068 8.515 3.271 ;
      RECT 8.343 3.072 8.429 3.272 ;
      RECT 8.257 3.076 8.343 3.273 ;
      RECT 8.171 3.079 8.257 3.273 ;
      RECT 8.085 3.083 8.171 3.274 ;
      RECT 8.05 3.088 8.085 3.275 ;
      RECT 7.995 3.098 8.05 3.282 ;
      RECT 7.97 3.11 7.995 3.292 ;
      RECT 7.935 3.123 7.97 3.3 ;
      RECT 7.895 3.14 7.935 3.323 ;
      RECT 7.875 3.153 7.895 3.35 ;
      RECT 7.845 3.165 7.875 3.378 ;
      RECT 7.84 3.173 7.845 3.398 ;
      RECT 7.835 3.176 7.84 3.408 ;
      RECT 7.785 3.188 7.835 3.442 ;
      RECT 7.775 3.203 7.785 3.475 ;
      RECT 7.765 3.209 7.775 3.488 ;
      RECT 7.755 3.216 7.765 3.5 ;
      RECT 7.73 3.229 7.755 3.518 ;
      RECT 7.715 3.244 7.73 3.54 ;
      RECT 7.705 3.252 7.715 3.556 ;
      RECT 7.69 3.261 7.705 3.571 ;
      RECT 7.68 3.271 7.69 3.585 ;
      RECT 7.661 3.284 7.68 3.602 ;
      RECT 7.575 3.329 7.661 3.667 ;
      RECT 7.56 3.374 7.575 3.725 ;
      RECT 7.555 3.383 7.56 3.738 ;
      RECT 7.545 3.39 7.555 3.743 ;
      RECT 7.54 3.395 7.545 3.747 ;
      RECT 7.52 3.405 7.54 3.754 ;
      RECT 7.495 3.425 7.52 3.768 ;
      RECT 7.46 3.45 7.495 3.788 ;
      RECT 7.445 3.473 7.46 3.803 ;
      RECT 7.435 3.483 7.445 3.808 ;
      RECT 7.425 3.491 7.435 3.815 ;
      RECT 7.415 3.5 7.425 3.821 ;
      RECT 7.395 3.512 7.415 3.823 ;
      RECT 7.385 3.525 7.395 3.825 ;
      RECT 7.36 3.54 7.385 3.828 ;
      RECT 7.34 3.557 7.36 3.832 ;
      RECT 7.3 3.585 7.34 3.838 ;
      RECT 7.235 3.632 7.3 3.847 ;
      RECT 7.22 3.665 7.235 3.855 ;
      RECT 7.215 3.672 7.22 3.857 ;
      RECT 7.165 3.697 7.215 3.862 ;
      RECT 7.15 3.721 7.165 3.869 ;
      RECT 7.1 3.726 7.15 3.87 ;
      RECT 7.014 3.73 7.1 3.87 ;
      RECT 6.928 3.73 7.014 3.87 ;
      RECT 6.842 3.73 6.928 3.871 ;
      RECT 6.756 3.73 6.842 3.871 ;
      RECT 6.67 3.73 6.756 3.871 ;
      RECT 6.604 3.73 6.67 3.871 ;
      RECT 6.518 3.73 6.604 3.872 ;
      RECT 6.432 3.73 6.518 3.872 ;
      RECT 6.346 3.731 6.432 3.873 ;
      RECT 6.26 3.731 6.346 3.873 ;
      RECT 6.174 3.731 6.26 3.873 ;
      RECT 6.088 3.731 6.174 3.874 ;
      RECT 6.002 3.731 6.088 3.874 ;
      RECT 5.916 3.732 6.002 3.875 ;
      RECT 5.83 3.732 5.916 3.875 ;
      RECT 5.81 3.732 5.83 3.875 ;
      RECT 5.724 3.732 5.81 3.875 ;
      RECT 5.638 3.732 5.724 3.875 ;
      RECT 5.552 3.733 5.638 3.875 ;
      RECT 5.466 3.733 5.552 3.875 ;
      RECT 5.38 3.733 5.466 3.875 ;
      RECT 5.294 3.734 5.38 3.875 ;
      RECT 5.208 3.734 5.294 3.875 ;
      RECT 5.122 3.734 5.208 3.875 ;
      RECT 5.036 3.734 5.122 3.875 ;
      RECT 4.95 3.735 5.036 3.875 ;
      RECT 4.9 3.732 4.95 3.875 ;
      RECT 4.89 3.73 4.9 3.874 ;
      RECT 4.886 3.73 4.89 3.873 ;
      RECT 4.8 3.725 4.886 3.868 ;
      RECT 4.778 3.718 4.8 3.862 ;
      RECT 4.692 3.709 4.778 3.856 ;
      RECT 4.606 3.696 4.692 3.847 ;
      RECT 4.52 3.682 4.606 3.837 ;
      RECT 4.475 3.672 4.52 3.83 ;
      RECT 4.455 2.96 4.475 3.238 ;
      RECT 4.455 3.665 4.475 3.826 ;
      RECT 4.425 2.96 4.455 3.26 ;
      RECT 4.415 3.632 4.455 3.823 ;
      RECT 4.41 2.96 4.425 3.28 ;
      RECT 4.41 3.597 4.415 3.821 ;
      RECT 4.405 2.96 4.41 3.405 ;
      RECT 4.405 3.557 4.41 3.821 ;
      RECT 4.395 2.96 4.405 3.821 ;
      RECT 4.32 2.96 4.395 3.815 ;
      RECT 4.29 2.96 4.32 3.805 ;
      RECT 4.285 2.96 4.29 3.797 ;
      RECT 4.28 3.002 4.285 3.79 ;
      RECT 4.27 3.071 4.28 3.781 ;
      RECT 4.265 3.141 4.27 3.733 ;
      RECT 4.26 3.205 4.265 3.63 ;
      RECT 4.255 3.24 4.26 3.585 ;
      RECT 4.253 3.277 4.255 3.477 ;
      RECT 4.25 3.285 4.253 3.47 ;
      RECT 4.245 3.35 4.25 3.413 ;
      RECT 8.32 2.44 8.6 2.72 ;
      RECT 8.31 2.44 8.6 2.583 ;
      RECT 8.265 2.305 8.525 2.565 ;
      RECT 8.265 2.42 8.58 2.565 ;
      RECT 8.265 2.39 8.575 2.565 ;
      RECT 8.265 2.377 8.565 2.565 ;
      RECT 8.265 2.367 8.56 2.565 ;
      RECT 4.24 2.35 4.5 2.61 ;
      RECT 8.01 1.9 8.27 2.16 ;
      RECT 8 1.925 8.27 2.12 ;
      RECT 7.995 1.925 8 2.119 ;
      RECT 7.925 1.92 7.995 2.111 ;
      RECT 7.84 1.907 7.925 2.094 ;
      RECT 7.836 1.899 7.84 2.084 ;
      RECT 7.75 1.892 7.836 2.074 ;
      RECT 7.741 1.884 7.75 2.064 ;
      RECT 7.655 1.877 7.741 2.052 ;
      RECT 7.635 1.868 7.655 2.038 ;
      RECT 7.58 1.863 7.635 2.03 ;
      RECT 7.57 1.857 7.58 2.024 ;
      RECT 7.55 1.855 7.57 2.02 ;
      RECT 7.542 1.854 7.55 2.016 ;
      RECT 7.456 1.846 7.542 2.005 ;
      RECT 7.37 1.832 7.456 1.985 ;
      RECT 7.31 1.82 7.37 1.97 ;
      RECT 7.3 1.815 7.31 1.965 ;
      RECT 7.25 1.815 7.3 1.967 ;
      RECT 7.203 1.817 7.25 1.971 ;
      RECT 7.117 1.824 7.203 1.976 ;
      RECT 7.031 1.832 7.117 1.982 ;
      RECT 6.945 1.841 7.031 1.988 ;
      RECT 6.886 1.847 6.945 1.993 ;
      RECT 6.8 1.852 6.886 1.999 ;
      RECT 6.725 1.857 6.8 2.005 ;
      RECT 6.686 1.859 6.725 2.01 ;
      RECT 6.6 1.856 6.686 2.015 ;
      RECT 6.515 1.854 6.6 2.022 ;
      RECT 6.483 1.853 6.515 2.025 ;
      RECT 6.397 1.852 6.483 2.026 ;
      RECT 6.311 1.851 6.397 2.027 ;
      RECT 6.225 1.85 6.311 2.027 ;
      RECT 6.139 1.849 6.225 2.028 ;
      RECT 6.053 1.848 6.139 2.029 ;
      RECT 5.967 1.847 6.053 2.03 ;
      RECT 5.881 1.846 5.967 2.03 ;
      RECT 5.795 1.845 5.881 2.031 ;
      RECT 5.745 1.845 5.795 2.032 ;
      RECT 5.731 1.846 5.745 2.032 ;
      RECT 5.645 1.853 5.731 2.033 ;
      RECT 5.571 1.864 5.645 2.034 ;
      RECT 5.485 1.873 5.571 2.035 ;
      RECT 5.45 1.88 5.485 2.05 ;
      RECT 5.425 1.883 5.45 2.08 ;
      RECT 5.4 1.892 5.425 2.109 ;
      RECT 5.39 1.903 5.4 2.129 ;
      RECT 5.38 1.911 5.39 2.143 ;
      RECT 5.375 1.917 5.38 2.153 ;
      RECT 5.35 1.934 5.375 2.17 ;
      RECT 5.335 1.956 5.35 2.198 ;
      RECT 5.305 1.982 5.335 2.228 ;
      RECT 5.285 2.011 5.305 2.258 ;
      RECT 5.28 2.026 5.285 2.275 ;
      RECT 5.26 2.041 5.28 2.29 ;
      RECT 5.25 2.059 5.26 2.308 ;
      RECT 5.24 2.07 5.25 2.323 ;
      RECT 5.19 2.102 5.24 2.349 ;
      RECT 5.185 2.132 5.19 2.369 ;
      RECT 5.175 2.145 5.185 2.375 ;
      RECT 5.166 2.155 5.175 2.383 ;
      RECT 5.155 2.166 5.166 2.391 ;
      RECT 5.15 2.176 5.155 2.397 ;
      RECT 5.135 2.197 5.15 2.404 ;
      RECT 5.12 2.227 5.135 2.412 ;
      RECT 5.085 2.257 5.12 2.418 ;
      RECT 5.06 2.275 5.085 2.425 ;
      RECT 5.01 2.283 5.06 2.434 ;
      RECT 4.985 2.288 5.01 2.443 ;
      RECT 4.93 2.294 4.985 2.453 ;
      RECT 4.925 2.299 4.93 2.461 ;
      RECT 4.911 2.302 4.925 2.463 ;
      RECT 4.825 2.314 4.911 2.475 ;
      RECT 4.815 2.326 4.825 2.488 ;
      RECT 4.73 2.339 4.815 2.5 ;
      RECT 4.686 2.356 4.73 2.514 ;
      RECT 4.6 2.373 4.686 2.53 ;
      RECT 4.57 2.387 4.6 2.544 ;
      RECT 4.56 2.392 4.57 2.549 ;
      RECT 4.5 2.395 4.56 2.558 ;
      RECT 7.39 2.665 7.65 2.925 ;
      RECT 7.39 2.665 7.67 2.778 ;
      RECT 7.39 2.665 7.695 2.745 ;
      RECT 7.39 2.665 7.7 2.725 ;
      RECT 7.44 2.44 7.72 2.72 ;
      RECT 6.995 3.175 7.255 3.435 ;
      RECT 6.985 3.032 7.18 3.373 ;
      RECT 6.98 3.14 7.195 3.365 ;
      RECT 6.975 3.19 7.255 3.355 ;
      RECT 6.965 3.267 7.255 3.34 ;
      RECT 6.985 3.115 7.195 3.373 ;
      RECT 6.995 2.99 7.18 3.435 ;
      RECT 6.995 2.885 7.16 3.435 ;
      RECT 7.005 2.872 7.16 3.435 ;
      RECT 7.005 2.83 7.15 3.435 ;
      RECT 7.01 2.755 7.15 3.435 ;
      RECT 7.04 2.405 7.15 3.435 ;
      RECT 7.045 2.135 7.17 2.758 ;
      RECT 7.015 2.71 7.17 2.758 ;
      RECT 7.03 2.512 7.15 3.435 ;
      RECT 7.02 2.622 7.17 2.758 ;
      RECT 7.045 2.135 7.185 2.615 ;
      RECT 7.045 2.135 7.205 2.49 ;
      RECT 7.01 2.135 7.27 2.395 ;
      RECT 6.48 2.44 6.76 2.72 ;
      RECT 6.465 2.44 6.76 2.7 ;
      RECT 4.52 3.305 4.78 3.565 ;
      RECT 6.305 3.16 6.565 3.42 ;
      RECT 6.285 3.18 6.565 3.395 ;
      RECT 6.242 3.18 6.285 3.394 ;
      RECT 6.156 3.181 6.242 3.391 ;
      RECT 6.07 3.182 6.156 3.387 ;
      RECT 5.995 3.184 6.07 3.384 ;
      RECT 5.972 3.185 5.995 3.382 ;
      RECT 5.886 3.186 5.972 3.38 ;
      RECT 5.8 3.187 5.886 3.377 ;
      RECT 5.776 3.188 5.8 3.375 ;
      RECT 5.69 3.19 5.776 3.372 ;
      RECT 5.605 3.192 5.69 3.373 ;
      RECT 5.548 3.193 5.605 3.379 ;
      RECT 5.462 3.195 5.548 3.389 ;
      RECT 5.376 3.198 5.462 3.402 ;
      RECT 5.29 3.2 5.376 3.414 ;
      RECT 5.276 3.201 5.29 3.421 ;
      RECT 5.19 3.202 5.276 3.429 ;
      RECT 5.15 3.204 5.19 3.438 ;
      RECT 5.141 3.205 5.15 3.441 ;
      RECT 5.055 3.213 5.141 3.447 ;
      RECT 5.035 3.222 5.055 3.455 ;
      RECT 4.95 3.237 5.035 3.463 ;
      RECT 4.89 3.26 4.95 3.474 ;
      RECT 4.88 3.272 4.89 3.479 ;
      RECT 4.84 3.282 4.88 3.483 ;
      RECT 4.785 3.299 4.84 3.491 ;
      RECT 4.78 3.309 4.785 3.495 ;
      RECT 5.846 2.44 5.905 2.837 ;
      RECT 5.76 2.44 5.965 2.828 ;
      RECT 5.755 2.47 5.965 2.823 ;
      RECT 5.721 2.47 5.965 2.821 ;
      RECT 5.635 2.47 5.965 2.815 ;
      RECT 5.59 2.47 5.985 2.793 ;
      RECT 5.59 2.47 6.005 2.748 ;
      RECT 5.55 2.47 6.005 2.738 ;
      RECT 5.76 2.44 6.04 2.72 ;
      RECT 5.495 2.44 5.755 2.7 ;
      RECT 4.68 1.92 4.94 2.18 ;
      RECT 4.76 1.88 5.04 2.16 ;
      RECT 0.19 8.5 0.57 8.88 ;
      RECT 0.235 0 0.375 8.88 ;
      RECT 0.19 0 0.57 0.38 ;
      RECT 75.27 0.815 75.64 1.185 ;
      RECT 73.56 7.04 73.93 7.41 ;
      RECT 59.485 0.815 59.855 1.185 ;
      RECT 57.775 7.04 58.145 7.41 ;
      RECT 43.7 0.815 44.07 1.185 ;
      RECT 41.99 7.04 42.36 7.41 ;
      RECT 27.925 0.815 28.295 1.185 ;
      RECT 26.215 7.04 26.585 7.41 ;
      RECT 12.145 0.815 12.515 1.185 ;
      RECT 10.435 7.04 10.805 7.41 ;
    LAYER via1 ;
      RECT 81.295 7.375 81.445 7.525 ;
      RECT 78.925 6.74 79.075 6.89 ;
      RECT 78.91 2.065 79.06 2.215 ;
      RECT 78.12 2.45 78.27 2.6 ;
      RECT 78.12 6.325 78.27 6.475 ;
      RECT 76.475 1.44 76.625 1.59 ;
      RECT 76.16 2.96 76.31 3.11 ;
      RECT 75.38 0.925 75.53 1.075 ;
      RECT 75.26 2.29 75.41 2.44 ;
      RECT 75.14 2.86 75.29 3.01 ;
      RECT 74.31 6.71 74.46 6.86 ;
      RECT 74.06 2.555 74.21 2.705 ;
      RECT 73.725 3.275 73.875 3.425 ;
      RECT 73.67 7.15 73.82 7.3 ;
      RECT 73.645 2.115 73.795 2.265 ;
      RECT 72.21 2.51 72.36 2.66 ;
      RECT 71.445 2.36 71.595 2.51 ;
      RECT 71.19 1.955 71.34 2.105 ;
      RECT 70.57 2.72 70.72 2.87 ;
      RECT 70.19 2.19 70.34 2.34 ;
      RECT 70.175 3.23 70.325 3.38 ;
      RECT 69.645 2.495 69.795 2.645 ;
      RECT 69.485 3.215 69.635 3.365 ;
      RECT 68.675 2.495 68.825 2.645 ;
      RECT 67.86 1.975 68.01 2.125 ;
      RECT 67.7 3.36 67.85 3.51 ;
      RECT 67.465 3.015 67.615 3.165 ;
      RECT 67.42 2.405 67.57 2.555 ;
      RECT 66.42 3.025 66.57 3.175 ;
      RECT 65.485 6.755 65.635 6.905 ;
      RECT 63.14 6.74 63.29 6.89 ;
      RECT 63.125 2.065 63.275 2.215 ;
      RECT 62.335 2.45 62.485 2.6 ;
      RECT 62.335 6.325 62.485 6.475 ;
      RECT 60.69 1.44 60.84 1.59 ;
      RECT 60.375 2.96 60.525 3.11 ;
      RECT 59.595 0.925 59.745 1.075 ;
      RECT 59.475 2.29 59.625 2.44 ;
      RECT 59.355 2.86 59.505 3.01 ;
      RECT 58.525 6.71 58.675 6.86 ;
      RECT 58.275 2.555 58.425 2.705 ;
      RECT 57.94 3.275 58.09 3.425 ;
      RECT 57.885 7.15 58.035 7.3 ;
      RECT 57.86 2.115 58.01 2.265 ;
      RECT 56.425 2.51 56.575 2.66 ;
      RECT 55.66 2.36 55.81 2.51 ;
      RECT 55.405 1.955 55.555 2.105 ;
      RECT 54.785 2.72 54.935 2.87 ;
      RECT 54.405 2.19 54.555 2.34 ;
      RECT 54.39 3.23 54.54 3.38 ;
      RECT 53.86 2.495 54.01 2.645 ;
      RECT 53.7 3.215 53.85 3.365 ;
      RECT 52.89 2.495 53.04 2.645 ;
      RECT 52.075 1.975 52.225 2.125 ;
      RECT 51.915 3.36 52.065 3.51 ;
      RECT 51.68 3.015 51.83 3.165 ;
      RECT 51.635 2.405 51.785 2.555 ;
      RECT 50.635 3.025 50.785 3.175 ;
      RECT 49.7 6.755 49.85 6.905 ;
      RECT 47.355 6.74 47.505 6.89 ;
      RECT 47.34 2.065 47.49 2.215 ;
      RECT 46.55 2.45 46.7 2.6 ;
      RECT 46.55 6.325 46.7 6.475 ;
      RECT 44.905 1.44 45.055 1.59 ;
      RECT 44.59 2.96 44.74 3.11 ;
      RECT 43.81 0.925 43.96 1.075 ;
      RECT 43.69 2.29 43.84 2.44 ;
      RECT 43.57 2.86 43.72 3.01 ;
      RECT 42.795 6.715 42.945 6.865 ;
      RECT 42.49 2.555 42.64 2.705 ;
      RECT 42.155 3.275 42.305 3.425 ;
      RECT 42.1 7.15 42.25 7.3 ;
      RECT 42.075 2.115 42.225 2.265 ;
      RECT 40.64 2.51 40.79 2.66 ;
      RECT 39.875 2.36 40.025 2.51 ;
      RECT 39.62 1.955 39.77 2.105 ;
      RECT 39 2.72 39.15 2.87 ;
      RECT 38.62 2.19 38.77 2.34 ;
      RECT 38.605 3.23 38.755 3.38 ;
      RECT 38.075 2.495 38.225 2.645 ;
      RECT 37.915 3.215 38.065 3.365 ;
      RECT 37.105 2.495 37.255 2.645 ;
      RECT 36.29 1.975 36.44 2.125 ;
      RECT 36.13 3.36 36.28 3.51 ;
      RECT 35.895 3.015 36.045 3.165 ;
      RECT 35.85 2.405 36 2.555 ;
      RECT 34.85 3.025 35 3.175 ;
      RECT 33.97 6.76 34.12 6.91 ;
      RECT 31.58 6.74 31.73 6.89 ;
      RECT 31.565 2.065 31.715 2.215 ;
      RECT 30.775 2.45 30.925 2.6 ;
      RECT 30.775 6.325 30.925 6.475 ;
      RECT 29.13 1.44 29.28 1.59 ;
      RECT 28.815 2.96 28.965 3.11 ;
      RECT 28.035 0.925 28.185 1.075 ;
      RECT 27.915 2.29 28.065 2.44 ;
      RECT 27.795 2.86 27.945 3.01 ;
      RECT 27.015 6.71 27.165 6.86 ;
      RECT 26.715 2.555 26.865 2.705 ;
      RECT 26.38 3.275 26.53 3.425 ;
      RECT 26.325 7.15 26.475 7.3 ;
      RECT 26.3 2.115 26.45 2.265 ;
      RECT 24.865 2.51 25.015 2.66 ;
      RECT 24.1 2.36 24.25 2.51 ;
      RECT 23.845 1.955 23.995 2.105 ;
      RECT 23.225 2.72 23.375 2.87 ;
      RECT 22.845 2.19 22.995 2.34 ;
      RECT 22.83 3.23 22.98 3.38 ;
      RECT 22.3 2.495 22.45 2.645 ;
      RECT 22.14 3.215 22.29 3.365 ;
      RECT 21.33 2.495 21.48 2.645 ;
      RECT 20.515 1.975 20.665 2.125 ;
      RECT 20.355 3.36 20.505 3.51 ;
      RECT 20.12 3.015 20.27 3.165 ;
      RECT 20.075 2.405 20.225 2.555 ;
      RECT 19.075 3.025 19.225 3.175 ;
      RECT 18.19 6.755 18.34 6.905 ;
      RECT 15.8 6.74 15.95 6.89 ;
      RECT 15.785 2.065 15.935 2.215 ;
      RECT 14.995 2.45 15.145 2.6 ;
      RECT 14.995 6.325 15.145 6.475 ;
      RECT 13.35 1.44 13.5 1.59 ;
      RECT 13.035 2.96 13.185 3.11 ;
      RECT 12.255 0.925 12.405 1.075 ;
      RECT 12.135 2.29 12.285 2.44 ;
      RECT 12.015 2.86 12.165 3.01 ;
      RECT 11.205 6.705 11.355 6.855 ;
      RECT 10.935 2.555 11.085 2.705 ;
      RECT 10.6 3.275 10.75 3.425 ;
      RECT 10.545 7.15 10.695 7.3 ;
      RECT 10.52 2.115 10.67 2.265 ;
      RECT 9.085 2.51 9.235 2.66 ;
      RECT 8.32 2.36 8.47 2.51 ;
      RECT 8.065 1.955 8.215 2.105 ;
      RECT 7.445 2.72 7.595 2.87 ;
      RECT 7.065 2.19 7.215 2.34 ;
      RECT 7.05 3.23 7.2 3.38 ;
      RECT 6.52 2.495 6.67 2.645 ;
      RECT 6.36 3.215 6.51 3.365 ;
      RECT 5.55 2.495 5.7 2.645 ;
      RECT 4.735 1.975 4.885 2.125 ;
      RECT 4.575 3.36 4.725 3.51 ;
      RECT 4.34 3.015 4.49 3.165 ;
      RECT 4.295 2.405 4.445 2.555 ;
      RECT 3.295 3.025 3.445 3.175 ;
      RECT 1.61 7.095 1.76 7.245 ;
      RECT 1.235 6.355 1.385 6.505 ;
      RECT 0.305 0.115 0.455 0.265 ;
      RECT 0.305 8.615 0.455 8.765 ;
    LAYER met1 ;
      RECT 66.17 1.26 75.83 1.74 ;
      RECT 50.385 1.26 60.045 1.74 ;
      RECT 34.6 1.26 44.26 1.74 ;
      RECT 18.825 1.26 28.485 1.74 ;
      RECT 3.045 1.26 12.705 1.74 ;
      RECT 66.17 1.26 75.885 1.59 ;
      RECT 50.385 1.26 60.1 1.59 ;
      RECT 34.6 1.26 44.315 1.59 ;
      RECT 18.825 1.26 28.54 1.59 ;
      RECT 3.045 1.26 12.76 1.59 ;
      RECT 66.285 0 76 1.585 ;
      RECT 50.5 0 60.215 1.585 ;
      RECT 34.715 0 44.43 1.585 ;
      RECT 18.94 0 28.655 1.585 ;
      RECT 3.16 0 12.875 1.585 ;
      RECT 0.205 0 0.555 0.335 ;
      RECT 0 0 0.805 0.315 ;
      RECT 81.585 0 81.765 0.305 ;
      RECT 65.8 0 79.635 0.305 ;
      RECT 50.015 0 63.85 0.305 ;
      RECT 34.24 0 48.065 0.305 ;
      RECT 18.46 0 32.29 0.305 ;
      RECT 0 0 16.51 0.305 ;
      RECT 0 0 81.765 0.3 ;
      RECT 0 8.58 81.765 8.88 ;
      RECT 81.585 8.575 81.765 8.88 ;
      RECT 65.8 8.575 79.635 8.88 ;
      RECT 50.015 8.575 63.85 8.88 ;
      RECT 34.24 8.575 48.065 8.88 ;
      RECT 18.46 8.575 32.29 8.88 ;
      RECT 0 8.575 16.51 8.88 ;
      RECT 72.855 6.315 73.025 8.88 ;
      RECT 57.07 6.315 57.24 8.88 ;
      RECT 41.285 6.315 41.455 8.88 ;
      RECT 25.51 6.315 25.68 8.88 ;
      RECT 9.73 6.315 9.9 8.88 ;
      RECT 0 8.565 0.805 8.88 ;
      RECT 0.205 8.545 0.555 8.88 ;
      RECT 73.225 6.285 73.515 6.515 ;
      RECT 57.44 6.285 57.73 6.515 ;
      RECT 41.655 6.285 41.945 6.515 ;
      RECT 25.88 6.285 26.17 6.515 ;
      RECT 10.1 6.285 10.39 6.515 ;
      RECT 72.855 6.315 73.515 6.485 ;
      RECT 57.07 6.315 57.73 6.485 ;
      RECT 41.285 6.315 41.945 6.485 ;
      RECT 25.51 6.315 26.17 6.485 ;
      RECT 9.73 6.315 10.39 6.485 ;
      RECT 81.16 7.77 81.45 8 ;
      RECT 81.22 6.29 81.39 8 ;
      RECT 81.195 7.275 81.545 7.625 ;
      RECT 81.16 6.29 81.45 6.52 ;
      RECT 80.755 2.395 80.86 2.965 ;
      RECT 80.755 2.73 81.08 2.96 ;
      RECT 80.755 2.76 81.25 2.93 ;
      RECT 80.755 2.395 80.945 2.96 ;
      RECT 80.17 2.36 80.46 2.59 ;
      RECT 80.17 2.395 80.945 2.565 ;
      RECT 80.23 0.88 80.4 2.59 ;
      RECT 80.17 0.88 80.46 1.11 ;
      RECT 80.17 7.77 80.46 8 ;
      RECT 80.23 6.29 80.4 8 ;
      RECT 80.17 6.29 80.46 6.52 ;
      RECT 80.17 6.325 81.025 6.485 ;
      RECT 80.855 5.92 81.025 6.485 ;
      RECT 80.17 6.32 80.565 6.485 ;
      RECT 80.79 5.92 81.08 6.15 ;
      RECT 80.79 5.95 81.25 6.12 ;
      RECT 79.8 2.73 80.09 2.96 ;
      RECT 79.8 2.76 80.26 2.93 ;
      RECT 79.865 1.655 80.03 2.96 ;
      RECT 78.38 1.625 78.67 1.855 ;
      RECT 78.38 1.655 80.03 1.825 ;
      RECT 78.44 0.885 78.61 1.855 ;
      RECT 78.38 0.885 78.67 1.115 ;
      RECT 78.38 7.765 78.67 7.995 ;
      RECT 78.44 7.025 78.61 7.995 ;
      RECT 78.44 7.12 80.03 7.29 ;
      RECT 79.86 5.92 80.03 7.29 ;
      RECT 78.38 7.025 78.67 7.255 ;
      RECT 79.8 5.92 80.09 6.15 ;
      RECT 79.8 5.95 80.26 6.12 ;
      RECT 78.81 1.965 79.16 2.315 ;
      RECT 76.475 2.025 79.16 2.195 ;
      RECT 76.475 1.34 76.645 2.195 ;
      RECT 76.375 1.34 76.725 1.69 ;
      RECT 78.835 6.655 79.16 6.98 ;
      RECT 74.21 6.61 74.56 6.96 ;
      RECT 78.81 6.655 79.16 6.885 ;
      RECT 74.03 6.655 74.56 6.885 ;
      RECT 73.86 6.685 79.16 6.855 ;
      RECT 78.035 2.365 78.355 2.685 ;
      RECT 78.005 2.365 78.355 2.595 ;
      RECT 77.835 2.395 78.355 2.565 ;
      RECT 78.035 6.255 78.355 6.545 ;
      RECT 78.005 6.285 78.355 6.515 ;
      RECT 77.835 6.315 78.355 6.485 ;
      RECT 74.67 2.465 74.855 2.675 ;
      RECT 74.66 2.47 74.87 2.668 ;
      RECT 74.66 2.47 74.956 2.645 ;
      RECT 74.66 2.47 75.015 2.62 ;
      RECT 74.66 2.47 75.07 2.6 ;
      RECT 74.66 2.47 75.08 2.588 ;
      RECT 74.66 2.47 75.275 2.527 ;
      RECT 74.66 2.47 75.305 2.51 ;
      RECT 74.66 2.47 75.325 2.5 ;
      RECT 75.205 2.235 75.465 2.495 ;
      RECT 75.19 2.325 75.205 2.542 ;
      RECT 74.725 2.457 75.465 2.495 ;
      RECT 75.176 2.336 75.19 2.548 ;
      RECT 74.765 2.45 75.465 2.495 ;
      RECT 75.09 2.376 75.176 2.567 ;
      RECT 75.015 2.437 75.465 2.495 ;
      RECT 75.085 2.412 75.09 2.584 ;
      RECT 75.07 2.422 75.465 2.495 ;
      RECT 75.08 2.417 75.085 2.586 ;
      RECT 75.375 2.922 75.38 3.014 ;
      RECT 75.37 2.9 75.375 3.031 ;
      RECT 75.365 2.89 75.37 3.043 ;
      RECT 75.355 2.881 75.365 3.053 ;
      RECT 75.35 2.876 75.355 3.061 ;
      RECT 75.345 2.735 75.35 3.064 ;
      RECT 75.311 2.735 75.345 3.075 ;
      RECT 75.225 2.735 75.311 3.11 ;
      RECT 75.145 2.735 75.225 3.158 ;
      RECT 75.116 2.735 75.145 3.182 ;
      RECT 75.03 2.735 75.116 3.188 ;
      RECT 75.025 2.919 75.03 3.193 ;
      RECT 74.99 2.93 75.025 3.196 ;
      RECT 74.965 2.945 74.99 3.2 ;
      RECT 74.951 2.954 74.965 3.202 ;
      RECT 74.865 2.981 74.951 3.208 ;
      RECT 74.8 3.022 74.865 3.217 ;
      RECT 74.785 3.042 74.8 3.222 ;
      RECT 74.755 3.052 74.785 3.225 ;
      RECT 74.75 3.062 74.755 3.228 ;
      RECT 74.72 3.067 74.75 3.23 ;
      RECT 74.7 3.072 74.72 3.234 ;
      RECT 74.615 3.075 74.7 3.241 ;
      RECT 74.6 3.072 74.615 3.247 ;
      RECT 74.59 3.069 74.6 3.249 ;
      RECT 74.57 3.066 74.59 3.251 ;
      RECT 74.55 3.062 74.57 3.252 ;
      RECT 74.535 3.058 74.55 3.254 ;
      RECT 74.525 3.055 74.535 3.255 ;
      RECT 74.485 3.049 74.525 3.253 ;
      RECT 74.475 3.044 74.485 3.251 ;
      RECT 74.46 3.041 74.475 3.247 ;
      RECT 74.435 3.036 74.46 3.24 ;
      RECT 74.385 3.027 74.435 3.228 ;
      RECT 74.315 3.013 74.385 3.21 ;
      RECT 74.257 2.998 74.315 3.192 ;
      RECT 74.171 2.981 74.257 3.172 ;
      RECT 74.085 2.96 74.171 3.147 ;
      RECT 74.035 2.945 74.085 3.128 ;
      RECT 74.031 2.939 74.035 3.12 ;
      RECT 73.945 2.929 74.031 3.107 ;
      RECT 73.91 2.914 73.945 3.09 ;
      RECT 73.895 2.907 73.91 3.083 ;
      RECT 73.835 2.895 73.895 3.071 ;
      RECT 73.815 2.882 73.835 3.059 ;
      RECT 73.775 2.873 73.815 3.051 ;
      RECT 73.77 2.865 73.775 3.044 ;
      RECT 73.69 2.855 73.77 3.03 ;
      RECT 73.675 2.842 73.69 3.015 ;
      RECT 73.67 2.84 73.675 3.013 ;
      RECT 73.591 2.828 73.67 3 ;
      RECT 73.505 2.803 73.591 2.975 ;
      RECT 73.49 2.772 73.505 2.96 ;
      RECT 73.475 2.747 73.49 2.956 ;
      RECT 73.46 2.74 73.475 2.952 ;
      RECT 73.285 2.745 73.29 2.948 ;
      RECT 73.28 2.75 73.285 2.943 ;
      RECT 73.29 2.74 73.46 2.95 ;
      RECT 74.005 2.5 74.11 2.76 ;
      RECT 74.82 2.025 74.825 2.25 ;
      RECT 74.95 2.025 75.005 2.235 ;
      RECT 75.005 2.03 75.015 2.228 ;
      RECT 74.911 2.025 74.95 2.238 ;
      RECT 74.825 2.025 74.911 2.245 ;
      RECT 74.805 2.03 74.82 2.251 ;
      RECT 74.795 2.07 74.805 2.253 ;
      RECT 74.765 2.08 74.795 2.255 ;
      RECT 74.76 2.085 74.765 2.257 ;
      RECT 74.735 2.09 74.76 2.259 ;
      RECT 74.72 2.095 74.735 2.261 ;
      RECT 74.705 2.097 74.72 2.263 ;
      RECT 74.7 2.102 74.705 2.265 ;
      RECT 74.65 2.11 74.7 2.268 ;
      RECT 74.625 2.119 74.65 2.273 ;
      RECT 74.615 2.126 74.625 2.278 ;
      RECT 74.61 2.129 74.615 2.282 ;
      RECT 74.59 2.132 74.61 2.291 ;
      RECT 74.56 2.14 74.59 2.311 ;
      RECT 74.531 2.153 74.56 2.333 ;
      RECT 74.445 2.187 74.531 2.377 ;
      RECT 74.44 2.213 74.445 2.415 ;
      RECT 74.435 2.217 74.44 2.424 ;
      RECT 74.4 2.23 74.435 2.457 ;
      RECT 74.39 2.244 74.4 2.495 ;
      RECT 74.385 2.248 74.39 2.508 ;
      RECT 74.38 2.252 74.385 2.513 ;
      RECT 74.37 2.26 74.38 2.525 ;
      RECT 74.365 2.267 74.37 2.54 ;
      RECT 74.34 2.28 74.365 2.565 ;
      RECT 74.3 2.309 74.34 2.62 ;
      RECT 74.285 2.334 74.3 2.675 ;
      RECT 74.275 2.345 74.285 2.698 ;
      RECT 74.27 2.352 74.275 2.71 ;
      RECT 74.265 2.356 74.27 2.718 ;
      RECT 74.21 2.384 74.265 2.76 ;
      RECT 74.19 2.42 74.21 2.76 ;
      RECT 74.175 2.435 74.19 2.76 ;
      RECT 74.12 2.467 74.175 2.76 ;
      RECT 74.11 2.497 74.12 2.76 ;
      RECT 73.72 2.112 73.905 2.35 ;
      RECT 73.705 2.114 73.915 2.345 ;
      RECT 73.59 2.06 73.85 2.32 ;
      RECT 73.585 2.097 73.85 2.274 ;
      RECT 73.58 2.107 73.85 2.271 ;
      RECT 73.575 2.147 73.915 2.265 ;
      RECT 73.57 2.18 73.915 2.255 ;
      RECT 73.58 2.122 73.93 2.193 ;
      RECT 73.877 3.22 73.89 3.75 ;
      RECT 73.791 3.22 73.89 3.749 ;
      RECT 73.791 3.22 73.895 3.748 ;
      RECT 73.705 3.22 73.895 3.746 ;
      RECT 73.7 3.22 73.895 3.743 ;
      RECT 73.7 3.22 73.905 3.741 ;
      RECT 73.695 3.512 73.905 3.738 ;
      RECT 73.695 3.522 73.91 3.735 ;
      RECT 73.695 3.59 73.915 3.731 ;
      RECT 73.685 3.595 73.915 3.73 ;
      RECT 73.685 3.687 73.92 3.727 ;
      RECT 73.67 3.22 73.93 3.48 ;
      RECT 73.6 7.765 73.89 7.995 ;
      RECT 73.66 7.025 73.83 7.995 ;
      RECT 73.575 7.055 73.915 7.4 ;
      RECT 73.6 7.025 73.89 7.4 ;
      RECT 72.9 2.21 72.945 3.745 ;
      RECT 73.1 2.21 73.13 2.425 ;
      RECT 71.475 1.95 71.595 2.16 ;
      RECT 71.135 1.9 71.395 2.16 ;
      RECT 71.135 1.945 71.43 2.15 ;
      RECT 73.14 2.226 73.145 2.28 ;
      RECT 73.135 2.219 73.14 2.413 ;
      RECT 73.13 2.213 73.135 2.42 ;
      RECT 73.085 2.21 73.1 2.433 ;
      RECT 73.08 2.21 73.085 2.455 ;
      RECT 73.075 2.21 73.08 2.503 ;
      RECT 73.07 2.21 73.075 2.523 ;
      RECT 73.06 2.21 73.07 2.63 ;
      RECT 73.055 2.21 73.06 2.693 ;
      RECT 73.05 2.21 73.055 2.75 ;
      RECT 73.045 2.21 73.05 2.758 ;
      RECT 73.03 2.21 73.045 2.865 ;
      RECT 73.02 2.21 73.03 3 ;
      RECT 73.01 2.21 73.02 3.11 ;
      RECT 73 2.21 73.01 3.167 ;
      RECT 72.995 2.21 73 3.207 ;
      RECT 72.99 2.21 72.995 3.243 ;
      RECT 72.98 2.21 72.99 3.283 ;
      RECT 72.975 2.21 72.98 3.325 ;
      RECT 72.955 2.21 72.975 3.39 ;
      RECT 72.96 3.535 72.965 3.715 ;
      RECT 72.955 3.517 72.96 3.723 ;
      RECT 72.95 2.21 72.955 3.453 ;
      RECT 72.95 3.497 72.955 3.73 ;
      RECT 72.945 2.21 72.95 3.74 ;
      RECT 72.89 2.21 72.9 2.51 ;
      RECT 72.895 2.757 72.9 3.745 ;
      RECT 72.89 2.822 72.895 3.745 ;
      RECT 72.885 2.211 72.89 2.5 ;
      RECT 72.88 2.887 72.89 3.745 ;
      RECT 72.875 2.212 72.885 2.49 ;
      RECT 72.865 3 72.88 3.745 ;
      RECT 72.87 2.213 72.875 2.48 ;
      RECT 72.85 2.214 72.87 2.458 ;
      RECT 72.855 3.097 72.865 3.745 ;
      RECT 72.85 3.172 72.855 3.745 ;
      RECT 72.84 2.213 72.85 2.435 ;
      RECT 72.845 3.215 72.85 3.745 ;
      RECT 72.84 3.242 72.845 3.745 ;
      RECT 72.83 2.211 72.84 2.423 ;
      RECT 72.835 3.285 72.84 3.745 ;
      RECT 72.83 3.312 72.835 3.745 ;
      RECT 72.82 2.21 72.83 2.41 ;
      RECT 72.825 3.327 72.83 3.745 ;
      RECT 72.785 3.385 72.825 3.745 ;
      RECT 72.815 2.209 72.82 2.395 ;
      RECT 72.81 2.207 72.815 2.388 ;
      RECT 72.8 2.204 72.81 2.378 ;
      RECT 72.795 2.201 72.8 2.363 ;
      RECT 72.78 2.197 72.795 2.356 ;
      RECT 72.775 3.44 72.785 3.745 ;
      RECT 72.775 2.194 72.78 2.351 ;
      RECT 72.76 2.19 72.775 2.345 ;
      RECT 72.77 3.457 72.775 3.745 ;
      RECT 72.76 3.52 72.77 3.745 ;
      RECT 72.68 2.175 72.76 2.325 ;
      RECT 72.755 3.527 72.76 3.74 ;
      RECT 72.75 3.535 72.755 3.73 ;
      RECT 72.67 2.161 72.68 2.309 ;
      RECT 72.655 2.157 72.67 2.307 ;
      RECT 72.645 2.152 72.655 2.303 ;
      RECT 72.62 2.145 72.645 2.295 ;
      RECT 72.615 2.14 72.62 2.29 ;
      RECT 72.605 2.14 72.615 2.288 ;
      RECT 72.595 2.138 72.605 2.286 ;
      RECT 72.565 2.13 72.595 2.28 ;
      RECT 72.55 2.122 72.565 2.273 ;
      RECT 72.53 2.117 72.55 2.266 ;
      RECT 72.525 2.113 72.53 2.261 ;
      RECT 72.495 2.106 72.525 2.255 ;
      RECT 72.47 2.097 72.495 2.245 ;
      RECT 72.44 2.09 72.47 2.237 ;
      RECT 72.415 2.08 72.44 2.228 ;
      RECT 72.4 2.072 72.415 2.222 ;
      RECT 72.375 2.067 72.4 2.217 ;
      RECT 72.365 2.063 72.375 2.212 ;
      RECT 72.345 2.058 72.365 2.207 ;
      RECT 72.31 2.053 72.345 2.2 ;
      RECT 72.25 2.048 72.31 2.193 ;
      RECT 72.237 2.044 72.25 2.191 ;
      RECT 72.151 2.039 72.237 2.188 ;
      RECT 72.065 2.029 72.151 2.184 ;
      RECT 72.024 2.022 72.065 2.181 ;
      RECT 71.938 2.015 72.024 2.178 ;
      RECT 71.852 2.005 71.938 2.174 ;
      RECT 71.766 1.995 71.852 2.169 ;
      RECT 71.68 1.985 71.766 2.165 ;
      RECT 71.67 1.97 71.68 2.163 ;
      RECT 71.66 1.955 71.67 2.163 ;
      RECT 71.595 1.95 71.66 2.162 ;
      RECT 71.43 1.947 71.475 2.155 ;
      RECT 72.675 2.852 72.68 3.043 ;
      RECT 72.67 2.847 72.675 3.05 ;
      RECT 72.656 2.845 72.67 3.056 ;
      RECT 72.57 2.845 72.656 3.058 ;
      RECT 72.566 2.845 72.57 3.061 ;
      RECT 72.48 2.845 72.566 3.079 ;
      RECT 72.47 2.85 72.48 3.098 ;
      RECT 72.46 2.905 72.47 3.102 ;
      RECT 72.435 2.92 72.46 3.109 ;
      RECT 72.395 2.94 72.435 3.122 ;
      RECT 72.39 2.952 72.395 3.132 ;
      RECT 72.375 2.958 72.39 3.137 ;
      RECT 72.37 2.963 72.375 3.141 ;
      RECT 72.35 2.97 72.37 3.146 ;
      RECT 72.28 2.995 72.35 3.163 ;
      RECT 72.24 3.023 72.28 3.183 ;
      RECT 72.235 3.033 72.24 3.191 ;
      RECT 72.215 3.04 72.235 3.193 ;
      RECT 72.21 3.047 72.215 3.196 ;
      RECT 72.18 3.055 72.21 3.199 ;
      RECT 72.175 3.06 72.18 3.203 ;
      RECT 72.101 3.064 72.175 3.211 ;
      RECT 72.015 3.073 72.101 3.227 ;
      RECT 72.011 3.078 72.015 3.236 ;
      RECT 71.925 3.083 72.011 3.246 ;
      RECT 71.885 3.091 71.925 3.258 ;
      RECT 71.835 3.097 71.885 3.265 ;
      RECT 71.75 3.106 71.835 3.28 ;
      RECT 71.675 3.117 71.75 3.298 ;
      RECT 71.64 3.124 71.675 3.308 ;
      RECT 71.565 3.132 71.64 3.313 ;
      RECT 71.51 3.141 71.565 3.313 ;
      RECT 71.485 3.146 71.51 3.311 ;
      RECT 71.475 3.149 71.485 3.309 ;
      RECT 71.44 3.151 71.475 3.307 ;
      RECT 71.41 3.153 71.44 3.303 ;
      RECT 71.365 3.152 71.41 3.299 ;
      RECT 71.345 3.147 71.365 3.296 ;
      RECT 71.295 3.132 71.345 3.293 ;
      RECT 71.285 3.117 71.295 3.288 ;
      RECT 71.235 3.102 71.285 3.278 ;
      RECT 71.185 3.077 71.235 3.258 ;
      RECT 71.175 3.062 71.185 3.24 ;
      RECT 71.17 3.06 71.175 3.234 ;
      RECT 71.15 3.055 71.17 3.229 ;
      RECT 71.145 3.047 71.15 3.223 ;
      RECT 71.13 3.041 71.145 3.216 ;
      RECT 71.125 3.036 71.13 3.208 ;
      RECT 71.105 3.031 71.125 3.2 ;
      RECT 71.09 3.024 71.105 3.193 ;
      RECT 71.075 3.018 71.09 3.184 ;
      RECT 71.07 3.012 71.075 3.177 ;
      RECT 71.025 2.987 71.07 3.163 ;
      RECT 71.01 2.957 71.025 3.145 ;
      RECT 70.995 2.94 71.01 3.136 ;
      RECT 70.97 2.92 70.995 3.124 ;
      RECT 70.93 2.89 70.97 3.104 ;
      RECT 70.92 2.86 70.93 3.089 ;
      RECT 70.905 2.85 70.92 3.082 ;
      RECT 70.85 2.815 70.905 3.061 ;
      RECT 70.835 2.778 70.85 3.04 ;
      RECT 70.825 2.765 70.835 3.032 ;
      RECT 70.775 2.735 70.825 3.014 ;
      RECT 70.76 2.665 70.775 2.995 ;
      RECT 70.715 2.665 70.76 2.978 ;
      RECT 70.69 2.665 70.715 2.96 ;
      RECT 70.68 2.665 70.69 2.953 ;
      RECT 70.601 2.665 70.68 2.946 ;
      RECT 70.515 2.665 70.601 2.938 ;
      RECT 70.5 2.697 70.515 2.933 ;
      RECT 70.425 2.707 70.5 2.929 ;
      RECT 70.405 2.717 70.425 2.924 ;
      RECT 70.38 2.717 70.405 2.921 ;
      RECT 70.37 2.707 70.38 2.92 ;
      RECT 70.36 2.68 70.37 2.919 ;
      RECT 70.32 2.675 70.36 2.917 ;
      RECT 70.275 2.675 70.32 2.913 ;
      RECT 70.25 2.675 70.275 2.908 ;
      RECT 70.2 2.675 70.25 2.895 ;
      RECT 70.16 2.68 70.17 2.88 ;
      RECT 70.17 2.675 70.2 2.885 ;
      RECT 72.155 2.455 72.415 2.715 ;
      RECT 72.15 2.477 72.415 2.673 ;
      RECT 71.39 2.305 71.61 2.67 ;
      RECT 71.372 2.392 71.61 2.669 ;
      RECT 71.355 2.397 71.61 2.666 ;
      RECT 71.355 2.397 71.63 2.665 ;
      RECT 71.325 2.407 71.63 2.663 ;
      RECT 71.32 2.422 71.63 2.659 ;
      RECT 71.32 2.422 71.635 2.658 ;
      RECT 71.315 2.48 71.635 2.656 ;
      RECT 71.315 2.48 71.645 2.653 ;
      RECT 71.31 2.545 71.645 2.648 ;
      RECT 71.39 2.305 71.65 2.565 ;
      RECT 70.135 2.135 70.395 2.395 ;
      RECT 70.135 2.178 70.481 2.369 ;
      RECT 70.135 2.178 70.525 2.368 ;
      RECT 70.135 2.178 70.545 2.366 ;
      RECT 70.135 2.178 70.645 2.365 ;
      RECT 70.135 2.178 70.665 2.363 ;
      RECT 70.135 2.178 70.675 2.358 ;
      RECT 70.545 2.145 70.735 2.355 ;
      RECT 70.545 2.147 70.74 2.353 ;
      RECT 70.535 2.152 70.745 2.345 ;
      RECT 70.481 2.176 70.745 2.345 ;
      RECT 70.525 2.17 70.535 2.367 ;
      RECT 70.535 2.15 70.74 2.353 ;
      RECT 69.49 3.21 69.695 3.44 ;
      RECT 69.43 3.16 69.485 3.42 ;
      RECT 69.49 3.16 69.69 3.44 ;
      RECT 70.46 3.475 70.465 3.502 ;
      RECT 70.45 3.385 70.46 3.507 ;
      RECT 70.445 3.307 70.45 3.513 ;
      RECT 70.435 3.297 70.445 3.52 ;
      RECT 70.43 3.287 70.435 3.526 ;
      RECT 70.42 3.282 70.43 3.528 ;
      RECT 70.405 3.274 70.42 3.536 ;
      RECT 70.39 3.265 70.405 3.548 ;
      RECT 70.38 3.257 70.39 3.558 ;
      RECT 70.345 3.175 70.38 3.576 ;
      RECT 70.31 3.175 70.345 3.595 ;
      RECT 70.295 3.175 70.31 3.603 ;
      RECT 70.24 3.175 70.295 3.603 ;
      RECT 70.206 3.175 70.24 3.594 ;
      RECT 70.12 3.175 70.206 3.57 ;
      RECT 70.11 3.235 70.12 3.552 ;
      RECT 70.07 3.237 70.11 3.543 ;
      RECT 70.065 3.239 70.07 3.533 ;
      RECT 70.045 3.241 70.065 3.528 ;
      RECT 70.035 3.244 70.045 3.523 ;
      RECT 70.025 3.245 70.035 3.518 ;
      RECT 70.001 3.246 70.025 3.51 ;
      RECT 69.915 3.251 70.001 3.488 ;
      RECT 69.86 3.25 69.915 3.461 ;
      RECT 69.845 3.243 69.86 3.448 ;
      RECT 69.81 3.238 69.845 3.444 ;
      RECT 69.755 3.23 69.81 3.443 ;
      RECT 69.695 3.217 69.755 3.441 ;
      RECT 69.485 3.16 69.49 3.428 ;
      RECT 69.56 2.53 69.745 2.74 ;
      RECT 69.55 2.535 69.76 2.733 ;
      RECT 69.59 2.44 69.85 2.7 ;
      RECT 69.545 2.597 69.85 2.623 ;
      RECT 68.89 2.39 68.895 3.19 ;
      RECT 68.835 2.44 68.865 3.19 ;
      RECT 68.825 2.44 68.83 2.75 ;
      RECT 68.81 2.44 68.815 2.745 ;
      RECT 68.355 2.485 68.37 2.7 ;
      RECT 68.285 2.485 68.37 2.695 ;
      RECT 69.55 2.065 69.62 2.275 ;
      RECT 69.62 2.072 69.63 2.27 ;
      RECT 69.516 2.065 69.55 2.282 ;
      RECT 69.43 2.065 69.516 2.306 ;
      RECT 69.42 2.07 69.43 2.325 ;
      RECT 69.415 2.082 69.42 2.328 ;
      RECT 69.4 2.097 69.415 2.332 ;
      RECT 69.395 2.115 69.4 2.336 ;
      RECT 69.355 2.125 69.395 2.345 ;
      RECT 69.34 2.132 69.355 2.357 ;
      RECT 69.325 2.137 69.34 2.362 ;
      RECT 69.31 2.14 69.325 2.367 ;
      RECT 69.3 2.142 69.31 2.371 ;
      RECT 69.265 2.149 69.3 2.379 ;
      RECT 69.23 2.157 69.265 2.393 ;
      RECT 69.22 2.163 69.23 2.402 ;
      RECT 69.215 2.165 69.22 2.404 ;
      RECT 69.195 2.168 69.215 2.41 ;
      RECT 69.165 2.175 69.195 2.421 ;
      RECT 69.155 2.181 69.165 2.428 ;
      RECT 69.13 2.184 69.155 2.435 ;
      RECT 69.12 2.188 69.13 2.443 ;
      RECT 69.115 2.189 69.12 2.465 ;
      RECT 69.11 2.19 69.115 2.48 ;
      RECT 69.105 2.191 69.11 2.495 ;
      RECT 69.1 2.192 69.105 2.51 ;
      RECT 69.095 2.193 69.1 2.54 ;
      RECT 69.085 2.195 69.095 2.573 ;
      RECT 69.07 2.199 69.085 2.62 ;
      RECT 69.06 2.202 69.07 2.665 ;
      RECT 69.055 2.205 69.06 2.693 ;
      RECT 69.045 2.207 69.055 2.72 ;
      RECT 69.04 2.21 69.045 2.755 ;
      RECT 69.01 2.215 69.04 2.813 ;
      RECT 69.005 2.22 69.01 2.898 ;
      RECT 69 2.222 69.005 2.933 ;
      RECT 68.995 2.224 69 3.015 ;
      RECT 68.99 2.226 68.995 3.103 ;
      RECT 68.98 2.228 68.99 3.185 ;
      RECT 68.965 2.242 68.98 3.19 ;
      RECT 68.93 2.287 68.965 3.19 ;
      RECT 68.92 2.327 68.93 3.19 ;
      RECT 68.905 2.355 68.92 3.19 ;
      RECT 68.9 2.372 68.905 3.19 ;
      RECT 68.895 2.38 68.9 3.19 ;
      RECT 68.885 2.395 68.89 3.19 ;
      RECT 68.88 2.402 68.885 3.19 ;
      RECT 68.87 2.422 68.88 3.19 ;
      RECT 68.865 2.435 68.87 3.19 ;
      RECT 68.83 2.44 68.835 2.775 ;
      RECT 68.815 2.83 68.835 3.19 ;
      RECT 68.815 2.44 68.825 2.748 ;
      RECT 68.81 2.87 68.815 3.19 ;
      RECT 68.76 2.44 68.81 2.743 ;
      RECT 68.805 2.907 68.81 3.19 ;
      RECT 68.795 2.93 68.805 3.19 ;
      RECT 68.79 2.975 68.795 3.19 ;
      RECT 68.78 2.985 68.79 3.183 ;
      RECT 68.706 2.44 68.76 2.737 ;
      RECT 68.62 2.44 68.706 2.73 ;
      RECT 68.571 2.487 68.62 2.723 ;
      RECT 68.485 2.495 68.571 2.716 ;
      RECT 68.47 2.492 68.485 2.711 ;
      RECT 68.456 2.485 68.47 2.71 ;
      RECT 68.37 2.485 68.456 2.705 ;
      RECT 68.275 2.49 68.285 2.69 ;
      RECT 67.865 1.92 67.88 2.32 ;
      RECT 68.06 1.92 68.065 2.18 ;
      RECT 67.805 1.92 67.85 2.18 ;
      RECT 68.26 3.225 68.265 3.43 ;
      RECT 68.255 3.215 68.26 3.435 ;
      RECT 68.25 3.202 68.255 3.44 ;
      RECT 68.245 3.182 68.25 3.44 ;
      RECT 68.22 3.135 68.245 3.44 ;
      RECT 68.185 3.05 68.22 3.44 ;
      RECT 68.18 2.987 68.185 3.44 ;
      RECT 68.175 2.972 68.18 3.44 ;
      RECT 68.16 2.932 68.175 3.44 ;
      RECT 68.155 2.907 68.16 3.44 ;
      RECT 68.145 2.89 68.155 3.44 ;
      RECT 68.11 2.812 68.145 3.44 ;
      RECT 68.105 2.755 68.11 3.44 ;
      RECT 68.1 2.742 68.105 3.44 ;
      RECT 68.09 2.72 68.1 3.44 ;
      RECT 68.08 2.685 68.09 3.44 ;
      RECT 68.07 2.655 68.08 3.44 ;
      RECT 68.06 2.57 68.07 3.083 ;
      RECT 68.067 3.215 68.07 3.44 ;
      RECT 68.065 3.225 68.067 3.44 ;
      RECT 68.055 3.235 68.065 3.435 ;
      RECT 68.05 1.92 68.06 2.315 ;
      RECT 68.055 2.447 68.06 3.058 ;
      RECT 68.05 2.345 68.055 3.041 ;
      RECT 68.04 1.92 68.05 3.017 ;
      RECT 68.035 1.92 68.04 2.988 ;
      RECT 68.03 1.92 68.035 2.978 ;
      RECT 68.01 1.92 68.03 2.94 ;
      RECT 68.005 1.92 68.01 2.898 ;
      RECT 68 1.92 68.005 2.878 ;
      RECT 67.97 1.92 68 2.828 ;
      RECT 67.96 1.92 67.97 2.775 ;
      RECT 67.955 1.92 67.96 2.748 ;
      RECT 67.95 1.92 67.955 2.733 ;
      RECT 67.94 1.92 67.95 2.71 ;
      RECT 67.93 1.92 67.94 2.685 ;
      RECT 67.925 1.92 67.93 2.625 ;
      RECT 67.915 1.92 67.925 2.563 ;
      RECT 67.91 1.92 67.915 2.483 ;
      RECT 67.905 1.92 67.91 2.448 ;
      RECT 67.9 1.92 67.905 2.423 ;
      RECT 67.895 1.92 67.9 2.408 ;
      RECT 67.89 1.92 67.895 2.378 ;
      RECT 67.885 1.92 67.89 2.355 ;
      RECT 67.88 1.92 67.885 2.328 ;
      RECT 67.85 1.92 67.865 2.315 ;
      RECT 67.005 3.455 67.19 3.665 ;
      RECT 66.995 3.46 67.205 3.658 ;
      RECT 66.995 3.46 67.225 3.63 ;
      RECT 66.995 3.46 67.24 3.609 ;
      RECT 66.995 3.46 67.255 3.607 ;
      RECT 66.995 3.46 67.265 3.606 ;
      RECT 66.995 3.46 67.295 3.603 ;
      RECT 67.645 3.305 67.905 3.565 ;
      RECT 67.605 3.352 67.905 3.548 ;
      RECT 67.596 3.36 67.605 3.551 ;
      RECT 67.19 3.453 67.905 3.548 ;
      RECT 67.51 3.378 67.596 3.558 ;
      RECT 67.205 3.45 67.905 3.548 ;
      RECT 67.451 3.4 67.51 3.57 ;
      RECT 67.225 3.446 67.905 3.548 ;
      RECT 67.365 3.412 67.451 3.581 ;
      RECT 67.24 3.442 67.905 3.548 ;
      RECT 67.31 3.425 67.365 3.593 ;
      RECT 67.255 3.44 67.905 3.548 ;
      RECT 67.295 3.431 67.31 3.599 ;
      RECT 67.265 3.436 67.905 3.548 ;
      RECT 67.41 2.96 67.67 3.22 ;
      RECT 67.41 2.98 67.78 3.19 ;
      RECT 67.41 2.985 67.79 3.185 ;
      RECT 67.601 2.399 67.68 2.63 ;
      RECT 67.515 2.402 67.73 2.625 ;
      RECT 67.51 2.402 67.73 2.62 ;
      RECT 67.51 2.407 67.74 2.618 ;
      RECT 67.485 2.407 67.74 2.615 ;
      RECT 67.485 2.415 67.75 2.613 ;
      RECT 67.365 2.35 67.625 2.61 ;
      RECT 67.365 2.397 67.675 2.61 ;
      RECT 66.62 2.97 66.625 3.23 ;
      RECT 66.45 2.74 66.455 3.23 ;
      RECT 66.335 2.98 66.34 3.205 ;
      RECT 67.045 2.075 67.05 2.285 ;
      RECT 67.05 2.08 67.065 2.28 ;
      RECT 66.985 2.075 67.045 2.293 ;
      RECT 66.97 2.075 66.985 2.303 ;
      RECT 66.92 2.075 66.97 2.32 ;
      RECT 66.9 2.075 66.92 2.343 ;
      RECT 66.885 2.075 66.9 2.355 ;
      RECT 66.865 2.075 66.885 2.365 ;
      RECT 66.855 2.08 66.865 2.374 ;
      RECT 66.85 2.09 66.855 2.379 ;
      RECT 66.845 2.102 66.85 2.383 ;
      RECT 66.835 2.125 66.845 2.388 ;
      RECT 66.83 2.14 66.835 2.392 ;
      RECT 66.825 2.157 66.83 2.395 ;
      RECT 66.82 2.165 66.825 2.398 ;
      RECT 66.81 2.17 66.82 2.402 ;
      RECT 66.805 2.177 66.81 2.407 ;
      RECT 66.795 2.182 66.805 2.411 ;
      RECT 66.77 2.194 66.795 2.422 ;
      RECT 66.75 2.211 66.77 2.438 ;
      RECT 66.725 2.228 66.75 2.46 ;
      RECT 66.69 2.251 66.725 2.518 ;
      RECT 66.67 2.273 66.69 2.58 ;
      RECT 66.665 2.283 66.67 2.615 ;
      RECT 66.655 2.29 66.665 2.653 ;
      RECT 66.65 2.297 66.655 2.673 ;
      RECT 66.645 2.308 66.65 2.71 ;
      RECT 66.64 2.316 66.645 2.775 ;
      RECT 66.63 2.327 66.64 2.828 ;
      RECT 66.625 2.345 66.63 2.898 ;
      RECT 66.62 2.355 66.625 2.935 ;
      RECT 66.615 2.365 66.62 3.23 ;
      RECT 66.61 2.377 66.615 3.23 ;
      RECT 66.605 2.387 66.61 3.23 ;
      RECT 66.595 2.397 66.605 3.23 ;
      RECT 66.585 2.42 66.595 3.23 ;
      RECT 66.57 2.455 66.585 3.23 ;
      RECT 66.53 2.517 66.57 3.23 ;
      RECT 66.525 2.57 66.53 3.23 ;
      RECT 66.5 2.605 66.525 3.23 ;
      RECT 66.485 2.65 66.5 3.23 ;
      RECT 66.48 2.672 66.485 3.23 ;
      RECT 66.47 2.685 66.48 3.23 ;
      RECT 66.46 2.71 66.47 3.23 ;
      RECT 66.455 2.732 66.46 3.23 ;
      RECT 66.43 2.77 66.45 3.23 ;
      RECT 66.39 2.827 66.43 3.23 ;
      RECT 66.385 2.877 66.39 3.23 ;
      RECT 66.38 2.895 66.385 3.23 ;
      RECT 66.375 2.907 66.38 3.23 ;
      RECT 66.365 2.925 66.375 3.23 ;
      RECT 66.355 2.945 66.365 3.205 ;
      RECT 66.35 2.962 66.355 3.205 ;
      RECT 66.34 2.975 66.35 3.205 ;
      RECT 66.31 2.985 66.335 3.205 ;
      RECT 66.3 2.992 66.31 3.205 ;
      RECT 66.285 3.002 66.3 3.2 ;
      RECT 65.375 7.77 65.665 8 ;
      RECT 65.435 6.29 65.605 8 ;
      RECT 65.385 6.655 65.735 7.005 ;
      RECT 65.375 6.29 65.665 6.52 ;
      RECT 64.97 2.395 65.075 2.965 ;
      RECT 64.97 2.73 65.295 2.96 ;
      RECT 64.97 2.76 65.465 2.93 ;
      RECT 64.97 2.395 65.16 2.96 ;
      RECT 64.385 2.36 64.675 2.59 ;
      RECT 64.385 2.395 65.16 2.565 ;
      RECT 64.445 0.88 64.615 2.59 ;
      RECT 64.385 0.88 64.675 1.11 ;
      RECT 64.385 7.77 64.675 8 ;
      RECT 64.445 6.29 64.615 8 ;
      RECT 64.385 6.29 64.675 6.52 ;
      RECT 64.385 6.325 65.24 6.485 ;
      RECT 65.07 5.92 65.24 6.485 ;
      RECT 64.385 6.32 64.78 6.485 ;
      RECT 65.005 5.92 65.295 6.15 ;
      RECT 65.005 5.95 65.465 6.12 ;
      RECT 64.015 2.73 64.305 2.96 ;
      RECT 64.015 2.76 64.475 2.93 ;
      RECT 64.08 1.655 64.245 2.96 ;
      RECT 62.595 1.625 62.885 1.855 ;
      RECT 62.595 1.655 64.245 1.825 ;
      RECT 62.655 0.885 62.825 1.855 ;
      RECT 62.595 0.885 62.885 1.115 ;
      RECT 62.595 7.765 62.885 7.995 ;
      RECT 62.655 7.025 62.825 7.995 ;
      RECT 62.655 7.12 64.245 7.29 ;
      RECT 64.075 5.92 64.245 7.29 ;
      RECT 62.595 7.025 62.885 7.255 ;
      RECT 64.015 5.92 64.305 6.15 ;
      RECT 64.015 5.95 64.475 6.12 ;
      RECT 63.025 1.965 63.375 2.315 ;
      RECT 60.69 2.025 63.375 2.195 ;
      RECT 60.69 1.34 60.86 2.195 ;
      RECT 60.59 1.34 60.94 1.69 ;
      RECT 63.05 6.655 63.375 6.98 ;
      RECT 58.425 6.61 58.775 6.96 ;
      RECT 63.025 6.655 63.375 6.885 ;
      RECT 58.245 6.655 58.775 6.885 ;
      RECT 58.075 6.685 63.375 6.855 ;
      RECT 62.25 2.365 62.57 2.685 ;
      RECT 62.22 2.365 62.57 2.595 ;
      RECT 62.05 2.395 62.57 2.565 ;
      RECT 62.25 6.255 62.57 6.545 ;
      RECT 62.22 6.285 62.57 6.515 ;
      RECT 62.05 6.315 62.57 6.485 ;
      RECT 58.885 2.465 59.07 2.675 ;
      RECT 58.875 2.47 59.085 2.668 ;
      RECT 58.875 2.47 59.171 2.645 ;
      RECT 58.875 2.47 59.23 2.62 ;
      RECT 58.875 2.47 59.285 2.6 ;
      RECT 58.875 2.47 59.295 2.588 ;
      RECT 58.875 2.47 59.49 2.527 ;
      RECT 58.875 2.47 59.52 2.51 ;
      RECT 58.875 2.47 59.54 2.5 ;
      RECT 59.42 2.235 59.68 2.495 ;
      RECT 59.405 2.325 59.42 2.542 ;
      RECT 58.94 2.457 59.68 2.495 ;
      RECT 59.391 2.336 59.405 2.548 ;
      RECT 58.98 2.45 59.68 2.495 ;
      RECT 59.305 2.376 59.391 2.567 ;
      RECT 59.23 2.437 59.68 2.495 ;
      RECT 59.3 2.412 59.305 2.584 ;
      RECT 59.285 2.422 59.68 2.495 ;
      RECT 59.295 2.417 59.3 2.586 ;
      RECT 59.59 2.922 59.595 3.014 ;
      RECT 59.585 2.9 59.59 3.031 ;
      RECT 59.58 2.89 59.585 3.043 ;
      RECT 59.57 2.881 59.58 3.053 ;
      RECT 59.565 2.876 59.57 3.061 ;
      RECT 59.56 2.735 59.565 3.064 ;
      RECT 59.526 2.735 59.56 3.075 ;
      RECT 59.44 2.735 59.526 3.11 ;
      RECT 59.36 2.735 59.44 3.158 ;
      RECT 59.331 2.735 59.36 3.182 ;
      RECT 59.245 2.735 59.331 3.188 ;
      RECT 59.24 2.919 59.245 3.193 ;
      RECT 59.205 2.93 59.24 3.196 ;
      RECT 59.18 2.945 59.205 3.2 ;
      RECT 59.166 2.954 59.18 3.202 ;
      RECT 59.08 2.981 59.166 3.208 ;
      RECT 59.015 3.022 59.08 3.217 ;
      RECT 59 3.042 59.015 3.222 ;
      RECT 58.97 3.052 59 3.225 ;
      RECT 58.965 3.062 58.97 3.228 ;
      RECT 58.935 3.067 58.965 3.23 ;
      RECT 58.915 3.072 58.935 3.234 ;
      RECT 58.83 3.075 58.915 3.241 ;
      RECT 58.815 3.072 58.83 3.247 ;
      RECT 58.805 3.069 58.815 3.249 ;
      RECT 58.785 3.066 58.805 3.251 ;
      RECT 58.765 3.062 58.785 3.252 ;
      RECT 58.75 3.058 58.765 3.254 ;
      RECT 58.74 3.055 58.75 3.255 ;
      RECT 58.7 3.049 58.74 3.253 ;
      RECT 58.69 3.044 58.7 3.251 ;
      RECT 58.675 3.041 58.69 3.247 ;
      RECT 58.65 3.036 58.675 3.24 ;
      RECT 58.6 3.027 58.65 3.228 ;
      RECT 58.53 3.013 58.6 3.21 ;
      RECT 58.472 2.998 58.53 3.192 ;
      RECT 58.386 2.981 58.472 3.172 ;
      RECT 58.3 2.96 58.386 3.147 ;
      RECT 58.25 2.945 58.3 3.128 ;
      RECT 58.246 2.939 58.25 3.12 ;
      RECT 58.16 2.929 58.246 3.107 ;
      RECT 58.125 2.914 58.16 3.09 ;
      RECT 58.11 2.907 58.125 3.083 ;
      RECT 58.05 2.895 58.11 3.071 ;
      RECT 58.03 2.882 58.05 3.059 ;
      RECT 57.99 2.873 58.03 3.051 ;
      RECT 57.985 2.865 57.99 3.044 ;
      RECT 57.905 2.855 57.985 3.03 ;
      RECT 57.89 2.842 57.905 3.015 ;
      RECT 57.885 2.84 57.89 3.013 ;
      RECT 57.806 2.828 57.885 3 ;
      RECT 57.72 2.803 57.806 2.975 ;
      RECT 57.705 2.772 57.72 2.96 ;
      RECT 57.69 2.747 57.705 2.956 ;
      RECT 57.675 2.74 57.69 2.952 ;
      RECT 57.5 2.745 57.505 2.948 ;
      RECT 57.495 2.75 57.5 2.943 ;
      RECT 57.505 2.74 57.675 2.95 ;
      RECT 58.22 2.5 58.325 2.76 ;
      RECT 59.035 2.025 59.04 2.25 ;
      RECT 59.165 2.025 59.22 2.235 ;
      RECT 59.22 2.03 59.23 2.228 ;
      RECT 59.126 2.025 59.165 2.238 ;
      RECT 59.04 2.025 59.126 2.245 ;
      RECT 59.02 2.03 59.035 2.251 ;
      RECT 59.01 2.07 59.02 2.253 ;
      RECT 58.98 2.08 59.01 2.255 ;
      RECT 58.975 2.085 58.98 2.257 ;
      RECT 58.95 2.09 58.975 2.259 ;
      RECT 58.935 2.095 58.95 2.261 ;
      RECT 58.92 2.097 58.935 2.263 ;
      RECT 58.915 2.102 58.92 2.265 ;
      RECT 58.865 2.11 58.915 2.268 ;
      RECT 58.84 2.119 58.865 2.273 ;
      RECT 58.83 2.126 58.84 2.278 ;
      RECT 58.825 2.129 58.83 2.282 ;
      RECT 58.805 2.132 58.825 2.291 ;
      RECT 58.775 2.14 58.805 2.311 ;
      RECT 58.746 2.153 58.775 2.333 ;
      RECT 58.66 2.187 58.746 2.377 ;
      RECT 58.655 2.213 58.66 2.415 ;
      RECT 58.65 2.217 58.655 2.424 ;
      RECT 58.615 2.23 58.65 2.457 ;
      RECT 58.605 2.244 58.615 2.495 ;
      RECT 58.6 2.248 58.605 2.508 ;
      RECT 58.595 2.252 58.6 2.513 ;
      RECT 58.585 2.26 58.595 2.525 ;
      RECT 58.58 2.267 58.585 2.54 ;
      RECT 58.555 2.28 58.58 2.565 ;
      RECT 58.515 2.309 58.555 2.62 ;
      RECT 58.5 2.334 58.515 2.675 ;
      RECT 58.49 2.345 58.5 2.698 ;
      RECT 58.485 2.352 58.49 2.71 ;
      RECT 58.48 2.356 58.485 2.718 ;
      RECT 58.425 2.384 58.48 2.76 ;
      RECT 58.405 2.42 58.425 2.76 ;
      RECT 58.39 2.435 58.405 2.76 ;
      RECT 58.335 2.467 58.39 2.76 ;
      RECT 58.325 2.497 58.335 2.76 ;
      RECT 57.935 2.112 58.12 2.35 ;
      RECT 57.92 2.114 58.13 2.345 ;
      RECT 57.805 2.06 58.065 2.32 ;
      RECT 57.8 2.097 58.065 2.274 ;
      RECT 57.795 2.107 58.065 2.271 ;
      RECT 57.79 2.147 58.13 2.265 ;
      RECT 57.785 2.18 58.13 2.255 ;
      RECT 57.795 2.122 58.145 2.193 ;
      RECT 58.092 3.22 58.105 3.75 ;
      RECT 58.006 3.22 58.105 3.749 ;
      RECT 58.006 3.22 58.11 3.748 ;
      RECT 57.92 3.22 58.11 3.746 ;
      RECT 57.915 3.22 58.11 3.743 ;
      RECT 57.915 3.22 58.12 3.741 ;
      RECT 57.91 3.512 58.12 3.738 ;
      RECT 57.91 3.522 58.125 3.735 ;
      RECT 57.91 3.59 58.13 3.731 ;
      RECT 57.9 3.595 58.13 3.73 ;
      RECT 57.9 3.687 58.135 3.727 ;
      RECT 57.885 3.22 58.145 3.48 ;
      RECT 57.815 7.765 58.105 7.995 ;
      RECT 57.875 7.025 58.045 7.995 ;
      RECT 57.79 7.055 58.13 7.4 ;
      RECT 57.815 7.025 58.105 7.4 ;
      RECT 57.115 2.21 57.16 3.745 ;
      RECT 57.315 2.21 57.345 2.425 ;
      RECT 55.69 1.95 55.81 2.16 ;
      RECT 55.35 1.9 55.61 2.16 ;
      RECT 55.35 1.945 55.645 2.15 ;
      RECT 57.355 2.226 57.36 2.28 ;
      RECT 57.35 2.219 57.355 2.413 ;
      RECT 57.345 2.213 57.35 2.42 ;
      RECT 57.3 2.21 57.315 2.433 ;
      RECT 57.295 2.21 57.3 2.455 ;
      RECT 57.29 2.21 57.295 2.503 ;
      RECT 57.285 2.21 57.29 2.523 ;
      RECT 57.275 2.21 57.285 2.63 ;
      RECT 57.27 2.21 57.275 2.693 ;
      RECT 57.265 2.21 57.27 2.75 ;
      RECT 57.26 2.21 57.265 2.758 ;
      RECT 57.245 2.21 57.26 2.865 ;
      RECT 57.235 2.21 57.245 3 ;
      RECT 57.225 2.21 57.235 3.11 ;
      RECT 57.215 2.21 57.225 3.167 ;
      RECT 57.21 2.21 57.215 3.207 ;
      RECT 57.205 2.21 57.21 3.243 ;
      RECT 57.195 2.21 57.205 3.283 ;
      RECT 57.19 2.21 57.195 3.325 ;
      RECT 57.17 2.21 57.19 3.39 ;
      RECT 57.175 3.535 57.18 3.715 ;
      RECT 57.17 3.517 57.175 3.723 ;
      RECT 57.165 2.21 57.17 3.453 ;
      RECT 57.165 3.497 57.17 3.73 ;
      RECT 57.16 2.21 57.165 3.74 ;
      RECT 57.105 2.21 57.115 2.51 ;
      RECT 57.11 2.757 57.115 3.745 ;
      RECT 57.105 2.822 57.11 3.745 ;
      RECT 57.1 2.211 57.105 2.5 ;
      RECT 57.095 2.887 57.105 3.745 ;
      RECT 57.09 2.212 57.1 2.49 ;
      RECT 57.08 3 57.095 3.745 ;
      RECT 57.085 2.213 57.09 2.48 ;
      RECT 57.065 2.214 57.085 2.458 ;
      RECT 57.07 3.097 57.08 3.745 ;
      RECT 57.065 3.172 57.07 3.745 ;
      RECT 57.055 2.213 57.065 2.435 ;
      RECT 57.06 3.215 57.065 3.745 ;
      RECT 57.055 3.242 57.06 3.745 ;
      RECT 57.045 2.211 57.055 2.423 ;
      RECT 57.05 3.285 57.055 3.745 ;
      RECT 57.045 3.312 57.05 3.745 ;
      RECT 57.035 2.21 57.045 2.41 ;
      RECT 57.04 3.327 57.045 3.745 ;
      RECT 57 3.385 57.04 3.745 ;
      RECT 57.03 2.209 57.035 2.395 ;
      RECT 57.025 2.207 57.03 2.388 ;
      RECT 57.015 2.204 57.025 2.378 ;
      RECT 57.01 2.201 57.015 2.363 ;
      RECT 56.995 2.197 57.01 2.356 ;
      RECT 56.99 3.44 57 3.745 ;
      RECT 56.99 2.194 56.995 2.351 ;
      RECT 56.975 2.19 56.99 2.345 ;
      RECT 56.985 3.457 56.99 3.745 ;
      RECT 56.975 3.52 56.985 3.745 ;
      RECT 56.895 2.175 56.975 2.325 ;
      RECT 56.97 3.527 56.975 3.74 ;
      RECT 56.965 3.535 56.97 3.73 ;
      RECT 56.885 2.161 56.895 2.309 ;
      RECT 56.87 2.157 56.885 2.307 ;
      RECT 56.86 2.152 56.87 2.303 ;
      RECT 56.835 2.145 56.86 2.295 ;
      RECT 56.83 2.14 56.835 2.29 ;
      RECT 56.82 2.14 56.83 2.288 ;
      RECT 56.81 2.138 56.82 2.286 ;
      RECT 56.78 2.13 56.81 2.28 ;
      RECT 56.765 2.122 56.78 2.273 ;
      RECT 56.745 2.117 56.765 2.266 ;
      RECT 56.74 2.113 56.745 2.261 ;
      RECT 56.71 2.106 56.74 2.255 ;
      RECT 56.685 2.097 56.71 2.245 ;
      RECT 56.655 2.09 56.685 2.237 ;
      RECT 56.63 2.08 56.655 2.228 ;
      RECT 56.615 2.072 56.63 2.222 ;
      RECT 56.59 2.067 56.615 2.217 ;
      RECT 56.58 2.063 56.59 2.212 ;
      RECT 56.56 2.058 56.58 2.207 ;
      RECT 56.525 2.053 56.56 2.2 ;
      RECT 56.465 2.048 56.525 2.193 ;
      RECT 56.452 2.044 56.465 2.191 ;
      RECT 56.366 2.039 56.452 2.188 ;
      RECT 56.28 2.029 56.366 2.184 ;
      RECT 56.239 2.022 56.28 2.181 ;
      RECT 56.153 2.015 56.239 2.178 ;
      RECT 56.067 2.005 56.153 2.174 ;
      RECT 55.981 1.995 56.067 2.169 ;
      RECT 55.895 1.985 55.981 2.165 ;
      RECT 55.885 1.97 55.895 2.163 ;
      RECT 55.875 1.955 55.885 2.163 ;
      RECT 55.81 1.95 55.875 2.162 ;
      RECT 55.645 1.947 55.69 2.155 ;
      RECT 56.89 2.852 56.895 3.043 ;
      RECT 56.885 2.847 56.89 3.05 ;
      RECT 56.871 2.845 56.885 3.056 ;
      RECT 56.785 2.845 56.871 3.058 ;
      RECT 56.781 2.845 56.785 3.061 ;
      RECT 56.695 2.845 56.781 3.079 ;
      RECT 56.685 2.85 56.695 3.098 ;
      RECT 56.675 2.905 56.685 3.102 ;
      RECT 56.65 2.92 56.675 3.109 ;
      RECT 56.61 2.94 56.65 3.122 ;
      RECT 56.605 2.952 56.61 3.132 ;
      RECT 56.59 2.958 56.605 3.137 ;
      RECT 56.585 2.963 56.59 3.141 ;
      RECT 56.565 2.97 56.585 3.146 ;
      RECT 56.495 2.995 56.565 3.163 ;
      RECT 56.455 3.023 56.495 3.183 ;
      RECT 56.45 3.033 56.455 3.191 ;
      RECT 56.43 3.04 56.45 3.193 ;
      RECT 56.425 3.047 56.43 3.196 ;
      RECT 56.395 3.055 56.425 3.199 ;
      RECT 56.39 3.06 56.395 3.203 ;
      RECT 56.316 3.064 56.39 3.211 ;
      RECT 56.23 3.073 56.316 3.227 ;
      RECT 56.226 3.078 56.23 3.236 ;
      RECT 56.14 3.083 56.226 3.246 ;
      RECT 56.1 3.091 56.14 3.258 ;
      RECT 56.05 3.097 56.1 3.265 ;
      RECT 55.965 3.106 56.05 3.28 ;
      RECT 55.89 3.117 55.965 3.298 ;
      RECT 55.855 3.124 55.89 3.308 ;
      RECT 55.78 3.132 55.855 3.313 ;
      RECT 55.725 3.141 55.78 3.313 ;
      RECT 55.7 3.146 55.725 3.311 ;
      RECT 55.69 3.149 55.7 3.309 ;
      RECT 55.655 3.151 55.69 3.307 ;
      RECT 55.625 3.153 55.655 3.303 ;
      RECT 55.58 3.152 55.625 3.299 ;
      RECT 55.56 3.147 55.58 3.296 ;
      RECT 55.51 3.132 55.56 3.293 ;
      RECT 55.5 3.117 55.51 3.288 ;
      RECT 55.45 3.102 55.5 3.278 ;
      RECT 55.4 3.077 55.45 3.258 ;
      RECT 55.39 3.062 55.4 3.24 ;
      RECT 55.385 3.06 55.39 3.234 ;
      RECT 55.365 3.055 55.385 3.229 ;
      RECT 55.36 3.047 55.365 3.223 ;
      RECT 55.345 3.041 55.36 3.216 ;
      RECT 55.34 3.036 55.345 3.208 ;
      RECT 55.32 3.031 55.34 3.2 ;
      RECT 55.305 3.024 55.32 3.193 ;
      RECT 55.29 3.018 55.305 3.184 ;
      RECT 55.285 3.012 55.29 3.177 ;
      RECT 55.24 2.987 55.285 3.163 ;
      RECT 55.225 2.957 55.24 3.145 ;
      RECT 55.21 2.94 55.225 3.136 ;
      RECT 55.185 2.92 55.21 3.124 ;
      RECT 55.145 2.89 55.185 3.104 ;
      RECT 55.135 2.86 55.145 3.089 ;
      RECT 55.12 2.85 55.135 3.082 ;
      RECT 55.065 2.815 55.12 3.061 ;
      RECT 55.05 2.778 55.065 3.04 ;
      RECT 55.04 2.765 55.05 3.032 ;
      RECT 54.99 2.735 55.04 3.014 ;
      RECT 54.975 2.665 54.99 2.995 ;
      RECT 54.93 2.665 54.975 2.978 ;
      RECT 54.905 2.665 54.93 2.96 ;
      RECT 54.895 2.665 54.905 2.953 ;
      RECT 54.816 2.665 54.895 2.946 ;
      RECT 54.73 2.665 54.816 2.938 ;
      RECT 54.715 2.697 54.73 2.933 ;
      RECT 54.64 2.707 54.715 2.929 ;
      RECT 54.62 2.717 54.64 2.924 ;
      RECT 54.595 2.717 54.62 2.921 ;
      RECT 54.585 2.707 54.595 2.92 ;
      RECT 54.575 2.68 54.585 2.919 ;
      RECT 54.535 2.675 54.575 2.917 ;
      RECT 54.49 2.675 54.535 2.913 ;
      RECT 54.465 2.675 54.49 2.908 ;
      RECT 54.415 2.675 54.465 2.895 ;
      RECT 54.375 2.68 54.385 2.88 ;
      RECT 54.385 2.675 54.415 2.885 ;
      RECT 56.37 2.455 56.63 2.715 ;
      RECT 56.365 2.477 56.63 2.673 ;
      RECT 55.605 2.305 55.825 2.67 ;
      RECT 55.587 2.392 55.825 2.669 ;
      RECT 55.57 2.397 55.825 2.666 ;
      RECT 55.57 2.397 55.845 2.665 ;
      RECT 55.54 2.407 55.845 2.663 ;
      RECT 55.535 2.422 55.845 2.659 ;
      RECT 55.535 2.422 55.85 2.658 ;
      RECT 55.53 2.48 55.85 2.656 ;
      RECT 55.53 2.48 55.86 2.653 ;
      RECT 55.525 2.545 55.86 2.648 ;
      RECT 55.605 2.305 55.865 2.565 ;
      RECT 54.35 2.135 54.61 2.395 ;
      RECT 54.35 2.178 54.696 2.369 ;
      RECT 54.35 2.178 54.74 2.368 ;
      RECT 54.35 2.178 54.76 2.366 ;
      RECT 54.35 2.178 54.86 2.365 ;
      RECT 54.35 2.178 54.88 2.363 ;
      RECT 54.35 2.178 54.89 2.358 ;
      RECT 54.76 2.145 54.95 2.355 ;
      RECT 54.76 2.147 54.955 2.353 ;
      RECT 54.75 2.152 54.96 2.345 ;
      RECT 54.696 2.176 54.96 2.345 ;
      RECT 54.74 2.17 54.75 2.367 ;
      RECT 54.75 2.15 54.955 2.353 ;
      RECT 53.705 3.21 53.91 3.44 ;
      RECT 53.645 3.16 53.7 3.42 ;
      RECT 53.705 3.16 53.905 3.44 ;
      RECT 54.675 3.475 54.68 3.502 ;
      RECT 54.665 3.385 54.675 3.507 ;
      RECT 54.66 3.307 54.665 3.513 ;
      RECT 54.65 3.297 54.66 3.52 ;
      RECT 54.645 3.287 54.65 3.526 ;
      RECT 54.635 3.282 54.645 3.528 ;
      RECT 54.62 3.274 54.635 3.536 ;
      RECT 54.605 3.265 54.62 3.548 ;
      RECT 54.595 3.257 54.605 3.558 ;
      RECT 54.56 3.175 54.595 3.576 ;
      RECT 54.525 3.175 54.56 3.595 ;
      RECT 54.51 3.175 54.525 3.603 ;
      RECT 54.455 3.175 54.51 3.603 ;
      RECT 54.421 3.175 54.455 3.594 ;
      RECT 54.335 3.175 54.421 3.57 ;
      RECT 54.325 3.235 54.335 3.552 ;
      RECT 54.285 3.237 54.325 3.543 ;
      RECT 54.28 3.239 54.285 3.533 ;
      RECT 54.26 3.241 54.28 3.528 ;
      RECT 54.25 3.244 54.26 3.523 ;
      RECT 54.24 3.245 54.25 3.518 ;
      RECT 54.216 3.246 54.24 3.51 ;
      RECT 54.13 3.251 54.216 3.488 ;
      RECT 54.075 3.25 54.13 3.461 ;
      RECT 54.06 3.243 54.075 3.448 ;
      RECT 54.025 3.238 54.06 3.444 ;
      RECT 53.97 3.23 54.025 3.443 ;
      RECT 53.91 3.217 53.97 3.441 ;
      RECT 53.7 3.16 53.705 3.428 ;
      RECT 53.775 2.53 53.96 2.74 ;
      RECT 53.765 2.535 53.975 2.733 ;
      RECT 53.805 2.44 54.065 2.7 ;
      RECT 53.76 2.597 54.065 2.623 ;
      RECT 53.105 2.39 53.11 3.19 ;
      RECT 53.05 2.44 53.08 3.19 ;
      RECT 53.04 2.44 53.045 2.75 ;
      RECT 53.025 2.44 53.03 2.745 ;
      RECT 52.57 2.485 52.585 2.7 ;
      RECT 52.5 2.485 52.585 2.695 ;
      RECT 53.765 2.065 53.835 2.275 ;
      RECT 53.835 2.072 53.845 2.27 ;
      RECT 53.731 2.065 53.765 2.282 ;
      RECT 53.645 2.065 53.731 2.306 ;
      RECT 53.635 2.07 53.645 2.325 ;
      RECT 53.63 2.082 53.635 2.328 ;
      RECT 53.615 2.097 53.63 2.332 ;
      RECT 53.61 2.115 53.615 2.336 ;
      RECT 53.57 2.125 53.61 2.345 ;
      RECT 53.555 2.132 53.57 2.357 ;
      RECT 53.54 2.137 53.555 2.362 ;
      RECT 53.525 2.14 53.54 2.367 ;
      RECT 53.515 2.142 53.525 2.371 ;
      RECT 53.48 2.149 53.515 2.379 ;
      RECT 53.445 2.157 53.48 2.393 ;
      RECT 53.435 2.163 53.445 2.402 ;
      RECT 53.43 2.165 53.435 2.404 ;
      RECT 53.41 2.168 53.43 2.41 ;
      RECT 53.38 2.175 53.41 2.421 ;
      RECT 53.37 2.181 53.38 2.428 ;
      RECT 53.345 2.184 53.37 2.435 ;
      RECT 53.335 2.188 53.345 2.443 ;
      RECT 53.33 2.189 53.335 2.465 ;
      RECT 53.325 2.19 53.33 2.48 ;
      RECT 53.32 2.191 53.325 2.495 ;
      RECT 53.315 2.192 53.32 2.51 ;
      RECT 53.31 2.193 53.315 2.54 ;
      RECT 53.3 2.195 53.31 2.573 ;
      RECT 53.285 2.199 53.3 2.62 ;
      RECT 53.275 2.202 53.285 2.665 ;
      RECT 53.27 2.205 53.275 2.693 ;
      RECT 53.26 2.207 53.27 2.72 ;
      RECT 53.255 2.21 53.26 2.755 ;
      RECT 53.225 2.215 53.255 2.813 ;
      RECT 53.22 2.22 53.225 2.898 ;
      RECT 53.215 2.222 53.22 2.933 ;
      RECT 53.21 2.224 53.215 3.015 ;
      RECT 53.205 2.226 53.21 3.103 ;
      RECT 53.195 2.228 53.205 3.185 ;
      RECT 53.18 2.242 53.195 3.19 ;
      RECT 53.145 2.287 53.18 3.19 ;
      RECT 53.135 2.327 53.145 3.19 ;
      RECT 53.12 2.355 53.135 3.19 ;
      RECT 53.115 2.372 53.12 3.19 ;
      RECT 53.11 2.38 53.115 3.19 ;
      RECT 53.1 2.395 53.105 3.19 ;
      RECT 53.095 2.402 53.1 3.19 ;
      RECT 53.085 2.422 53.095 3.19 ;
      RECT 53.08 2.435 53.085 3.19 ;
      RECT 53.045 2.44 53.05 2.775 ;
      RECT 53.03 2.83 53.05 3.19 ;
      RECT 53.03 2.44 53.04 2.748 ;
      RECT 53.025 2.87 53.03 3.19 ;
      RECT 52.975 2.44 53.025 2.743 ;
      RECT 53.02 2.907 53.025 3.19 ;
      RECT 53.01 2.93 53.02 3.19 ;
      RECT 53.005 2.975 53.01 3.19 ;
      RECT 52.995 2.985 53.005 3.183 ;
      RECT 52.921 2.44 52.975 2.737 ;
      RECT 52.835 2.44 52.921 2.73 ;
      RECT 52.786 2.487 52.835 2.723 ;
      RECT 52.7 2.495 52.786 2.716 ;
      RECT 52.685 2.492 52.7 2.711 ;
      RECT 52.671 2.485 52.685 2.71 ;
      RECT 52.585 2.485 52.671 2.705 ;
      RECT 52.49 2.49 52.5 2.69 ;
      RECT 52.08 1.92 52.095 2.32 ;
      RECT 52.275 1.92 52.28 2.18 ;
      RECT 52.02 1.92 52.065 2.18 ;
      RECT 52.475 3.225 52.48 3.43 ;
      RECT 52.47 3.215 52.475 3.435 ;
      RECT 52.465 3.202 52.47 3.44 ;
      RECT 52.46 3.182 52.465 3.44 ;
      RECT 52.435 3.135 52.46 3.44 ;
      RECT 52.4 3.05 52.435 3.44 ;
      RECT 52.395 2.987 52.4 3.44 ;
      RECT 52.39 2.972 52.395 3.44 ;
      RECT 52.375 2.932 52.39 3.44 ;
      RECT 52.37 2.907 52.375 3.44 ;
      RECT 52.36 2.89 52.37 3.44 ;
      RECT 52.325 2.812 52.36 3.44 ;
      RECT 52.32 2.755 52.325 3.44 ;
      RECT 52.315 2.742 52.32 3.44 ;
      RECT 52.305 2.72 52.315 3.44 ;
      RECT 52.295 2.685 52.305 3.44 ;
      RECT 52.285 2.655 52.295 3.44 ;
      RECT 52.275 2.57 52.285 3.083 ;
      RECT 52.282 3.215 52.285 3.44 ;
      RECT 52.28 3.225 52.282 3.44 ;
      RECT 52.27 3.235 52.28 3.435 ;
      RECT 52.265 1.92 52.275 2.315 ;
      RECT 52.27 2.447 52.275 3.058 ;
      RECT 52.265 2.345 52.27 3.041 ;
      RECT 52.255 1.92 52.265 3.017 ;
      RECT 52.25 1.92 52.255 2.988 ;
      RECT 52.245 1.92 52.25 2.978 ;
      RECT 52.225 1.92 52.245 2.94 ;
      RECT 52.22 1.92 52.225 2.898 ;
      RECT 52.215 1.92 52.22 2.878 ;
      RECT 52.185 1.92 52.215 2.828 ;
      RECT 52.175 1.92 52.185 2.775 ;
      RECT 52.17 1.92 52.175 2.748 ;
      RECT 52.165 1.92 52.17 2.733 ;
      RECT 52.155 1.92 52.165 2.71 ;
      RECT 52.145 1.92 52.155 2.685 ;
      RECT 52.14 1.92 52.145 2.625 ;
      RECT 52.13 1.92 52.14 2.563 ;
      RECT 52.125 1.92 52.13 2.483 ;
      RECT 52.12 1.92 52.125 2.448 ;
      RECT 52.115 1.92 52.12 2.423 ;
      RECT 52.11 1.92 52.115 2.408 ;
      RECT 52.105 1.92 52.11 2.378 ;
      RECT 52.1 1.92 52.105 2.355 ;
      RECT 52.095 1.92 52.1 2.328 ;
      RECT 52.065 1.92 52.08 2.315 ;
      RECT 51.22 3.455 51.405 3.665 ;
      RECT 51.21 3.46 51.42 3.658 ;
      RECT 51.21 3.46 51.44 3.63 ;
      RECT 51.21 3.46 51.455 3.609 ;
      RECT 51.21 3.46 51.47 3.607 ;
      RECT 51.21 3.46 51.48 3.606 ;
      RECT 51.21 3.46 51.51 3.603 ;
      RECT 51.86 3.305 52.12 3.565 ;
      RECT 51.82 3.352 52.12 3.548 ;
      RECT 51.811 3.36 51.82 3.551 ;
      RECT 51.405 3.453 52.12 3.548 ;
      RECT 51.725 3.378 51.811 3.558 ;
      RECT 51.42 3.45 52.12 3.548 ;
      RECT 51.666 3.4 51.725 3.57 ;
      RECT 51.44 3.446 52.12 3.548 ;
      RECT 51.58 3.412 51.666 3.581 ;
      RECT 51.455 3.442 52.12 3.548 ;
      RECT 51.525 3.425 51.58 3.593 ;
      RECT 51.47 3.44 52.12 3.548 ;
      RECT 51.51 3.431 51.525 3.599 ;
      RECT 51.48 3.436 52.12 3.548 ;
      RECT 51.625 2.96 51.885 3.22 ;
      RECT 51.625 2.98 51.995 3.19 ;
      RECT 51.625 2.985 52.005 3.185 ;
      RECT 51.816 2.399 51.895 2.63 ;
      RECT 51.73 2.402 51.945 2.625 ;
      RECT 51.725 2.402 51.945 2.62 ;
      RECT 51.725 2.407 51.955 2.618 ;
      RECT 51.7 2.407 51.955 2.615 ;
      RECT 51.7 2.415 51.965 2.613 ;
      RECT 51.58 2.35 51.84 2.61 ;
      RECT 51.58 2.397 51.89 2.61 ;
      RECT 50.835 2.97 50.84 3.23 ;
      RECT 50.665 2.74 50.67 3.23 ;
      RECT 50.55 2.98 50.555 3.205 ;
      RECT 51.26 2.075 51.265 2.285 ;
      RECT 51.265 2.08 51.28 2.28 ;
      RECT 51.2 2.075 51.26 2.293 ;
      RECT 51.185 2.075 51.2 2.303 ;
      RECT 51.135 2.075 51.185 2.32 ;
      RECT 51.115 2.075 51.135 2.343 ;
      RECT 51.1 2.075 51.115 2.355 ;
      RECT 51.08 2.075 51.1 2.365 ;
      RECT 51.07 2.08 51.08 2.374 ;
      RECT 51.065 2.09 51.07 2.379 ;
      RECT 51.06 2.102 51.065 2.383 ;
      RECT 51.05 2.125 51.06 2.388 ;
      RECT 51.045 2.14 51.05 2.392 ;
      RECT 51.04 2.157 51.045 2.395 ;
      RECT 51.035 2.165 51.04 2.398 ;
      RECT 51.025 2.17 51.035 2.402 ;
      RECT 51.02 2.177 51.025 2.407 ;
      RECT 51.01 2.182 51.02 2.411 ;
      RECT 50.985 2.194 51.01 2.422 ;
      RECT 50.965 2.211 50.985 2.438 ;
      RECT 50.94 2.228 50.965 2.46 ;
      RECT 50.905 2.251 50.94 2.518 ;
      RECT 50.885 2.273 50.905 2.58 ;
      RECT 50.88 2.283 50.885 2.615 ;
      RECT 50.87 2.29 50.88 2.653 ;
      RECT 50.865 2.297 50.87 2.673 ;
      RECT 50.86 2.308 50.865 2.71 ;
      RECT 50.855 2.316 50.86 2.775 ;
      RECT 50.845 2.327 50.855 2.828 ;
      RECT 50.84 2.345 50.845 2.898 ;
      RECT 50.835 2.355 50.84 2.935 ;
      RECT 50.83 2.365 50.835 3.23 ;
      RECT 50.825 2.377 50.83 3.23 ;
      RECT 50.82 2.387 50.825 3.23 ;
      RECT 50.81 2.397 50.82 3.23 ;
      RECT 50.8 2.42 50.81 3.23 ;
      RECT 50.785 2.455 50.8 3.23 ;
      RECT 50.745 2.517 50.785 3.23 ;
      RECT 50.74 2.57 50.745 3.23 ;
      RECT 50.715 2.605 50.74 3.23 ;
      RECT 50.7 2.65 50.715 3.23 ;
      RECT 50.695 2.672 50.7 3.23 ;
      RECT 50.685 2.685 50.695 3.23 ;
      RECT 50.675 2.71 50.685 3.23 ;
      RECT 50.67 2.732 50.675 3.23 ;
      RECT 50.645 2.77 50.665 3.23 ;
      RECT 50.605 2.827 50.645 3.23 ;
      RECT 50.6 2.877 50.605 3.23 ;
      RECT 50.595 2.895 50.6 3.23 ;
      RECT 50.59 2.907 50.595 3.23 ;
      RECT 50.58 2.925 50.59 3.23 ;
      RECT 50.57 2.945 50.58 3.205 ;
      RECT 50.565 2.962 50.57 3.205 ;
      RECT 50.555 2.975 50.565 3.205 ;
      RECT 50.525 2.985 50.55 3.205 ;
      RECT 50.515 2.992 50.525 3.205 ;
      RECT 50.5 3.002 50.515 3.2 ;
      RECT 49.59 7.77 49.88 8 ;
      RECT 49.65 6.29 49.82 8 ;
      RECT 49.6 6.655 49.95 7.005 ;
      RECT 49.59 6.29 49.88 6.52 ;
      RECT 49.185 2.395 49.29 2.965 ;
      RECT 49.185 2.73 49.51 2.96 ;
      RECT 49.185 2.76 49.68 2.93 ;
      RECT 49.185 2.395 49.375 2.96 ;
      RECT 48.6 2.36 48.89 2.59 ;
      RECT 48.6 2.395 49.375 2.565 ;
      RECT 48.66 0.88 48.83 2.59 ;
      RECT 48.6 0.88 48.89 1.11 ;
      RECT 48.6 7.77 48.89 8 ;
      RECT 48.66 6.29 48.83 8 ;
      RECT 48.6 6.29 48.89 6.52 ;
      RECT 48.6 6.325 49.455 6.485 ;
      RECT 49.285 5.92 49.455 6.485 ;
      RECT 48.6 6.32 48.995 6.485 ;
      RECT 49.22 5.92 49.51 6.15 ;
      RECT 49.22 5.95 49.68 6.12 ;
      RECT 48.23 2.73 48.52 2.96 ;
      RECT 48.23 2.76 48.69 2.93 ;
      RECT 48.295 1.655 48.46 2.96 ;
      RECT 46.81 1.625 47.1 1.855 ;
      RECT 46.81 1.655 48.46 1.825 ;
      RECT 46.87 0.885 47.04 1.855 ;
      RECT 46.81 0.885 47.1 1.115 ;
      RECT 46.81 7.765 47.1 7.995 ;
      RECT 46.87 7.025 47.04 7.995 ;
      RECT 46.87 7.12 48.46 7.29 ;
      RECT 48.29 5.92 48.46 7.29 ;
      RECT 46.81 7.025 47.1 7.255 ;
      RECT 48.23 5.92 48.52 6.15 ;
      RECT 48.23 5.95 48.69 6.12 ;
      RECT 47.24 1.965 47.59 2.315 ;
      RECT 44.905 2.025 47.59 2.195 ;
      RECT 44.905 1.34 45.075 2.195 ;
      RECT 44.805 1.34 45.155 1.69 ;
      RECT 47.265 6.655 47.59 6.98 ;
      RECT 42.695 6.615 43.045 6.965 ;
      RECT 47.24 6.655 47.59 6.885 ;
      RECT 42.46 6.655 43.045 6.885 ;
      RECT 42.29 6.685 47.59 6.855 ;
      RECT 46.465 2.365 46.785 2.685 ;
      RECT 46.435 2.365 46.785 2.595 ;
      RECT 46.265 2.395 46.785 2.565 ;
      RECT 46.465 6.255 46.785 6.545 ;
      RECT 46.435 6.285 46.785 6.515 ;
      RECT 46.265 6.315 46.785 6.485 ;
      RECT 43.1 2.465 43.285 2.675 ;
      RECT 43.09 2.47 43.3 2.668 ;
      RECT 43.09 2.47 43.386 2.645 ;
      RECT 43.09 2.47 43.445 2.62 ;
      RECT 43.09 2.47 43.5 2.6 ;
      RECT 43.09 2.47 43.51 2.588 ;
      RECT 43.09 2.47 43.705 2.527 ;
      RECT 43.09 2.47 43.735 2.51 ;
      RECT 43.09 2.47 43.755 2.5 ;
      RECT 43.635 2.235 43.895 2.495 ;
      RECT 43.62 2.325 43.635 2.542 ;
      RECT 43.155 2.457 43.895 2.495 ;
      RECT 43.606 2.336 43.62 2.548 ;
      RECT 43.195 2.45 43.895 2.495 ;
      RECT 43.52 2.376 43.606 2.567 ;
      RECT 43.445 2.437 43.895 2.495 ;
      RECT 43.515 2.412 43.52 2.584 ;
      RECT 43.5 2.422 43.895 2.495 ;
      RECT 43.51 2.417 43.515 2.586 ;
      RECT 43.805 2.922 43.81 3.014 ;
      RECT 43.8 2.9 43.805 3.031 ;
      RECT 43.795 2.89 43.8 3.043 ;
      RECT 43.785 2.881 43.795 3.053 ;
      RECT 43.78 2.876 43.785 3.061 ;
      RECT 43.775 2.735 43.78 3.064 ;
      RECT 43.741 2.735 43.775 3.075 ;
      RECT 43.655 2.735 43.741 3.11 ;
      RECT 43.575 2.735 43.655 3.158 ;
      RECT 43.546 2.735 43.575 3.182 ;
      RECT 43.46 2.735 43.546 3.188 ;
      RECT 43.455 2.919 43.46 3.193 ;
      RECT 43.42 2.93 43.455 3.196 ;
      RECT 43.395 2.945 43.42 3.2 ;
      RECT 43.381 2.954 43.395 3.202 ;
      RECT 43.295 2.981 43.381 3.208 ;
      RECT 43.23 3.022 43.295 3.217 ;
      RECT 43.215 3.042 43.23 3.222 ;
      RECT 43.185 3.052 43.215 3.225 ;
      RECT 43.18 3.062 43.185 3.228 ;
      RECT 43.15 3.067 43.18 3.23 ;
      RECT 43.13 3.072 43.15 3.234 ;
      RECT 43.045 3.075 43.13 3.241 ;
      RECT 43.03 3.072 43.045 3.247 ;
      RECT 43.02 3.069 43.03 3.249 ;
      RECT 43 3.066 43.02 3.251 ;
      RECT 42.98 3.062 43 3.252 ;
      RECT 42.965 3.058 42.98 3.254 ;
      RECT 42.955 3.055 42.965 3.255 ;
      RECT 42.915 3.049 42.955 3.253 ;
      RECT 42.905 3.044 42.915 3.251 ;
      RECT 42.89 3.041 42.905 3.247 ;
      RECT 42.865 3.036 42.89 3.24 ;
      RECT 42.815 3.027 42.865 3.228 ;
      RECT 42.745 3.013 42.815 3.21 ;
      RECT 42.687 2.998 42.745 3.192 ;
      RECT 42.601 2.981 42.687 3.172 ;
      RECT 42.515 2.96 42.601 3.147 ;
      RECT 42.465 2.945 42.515 3.128 ;
      RECT 42.461 2.939 42.465 3.12 ;
      RECT 42.375 2.929 42.461 3.107 ;
      RECT 42.34 2.914 42.375 3.09 ;
      RECT 42.325 2.907 42.34 3.083 ;
      RECT 42.265 2.895 42.325 3.071 ;
      RECT 42.245 2.882 42.265 3.059 ;
      RECT 42.205 2.873 42.245 3.051 ;
      RECT 42.2 2.865 42.205 3.044 ;
      RECT 42.12 2.855 42.2 3.03 ;
      RECT 42.105 2.842 42.12 3.015 ;
      RECT 42.1 2.84 42.105 3.013 ;
      RECT 42.021 2.828 42.1 3 ;
      RECT 41.935 2.803 42.021 2.975 ;
      RECT 41.92 2.772 41.935 2.96 ;
      RECT 41.905 2.747 41.92 2.956 ;
      RECT 41.89 2.74 41.905 2.952 ;
      RECT 41.715 2.745 41.72 2.948 ;
      RECT 41.71 2.75 41.715 2.943 ;
      RECT 41.72 2.74 41.89 2.95 ;
      RECT 42.435 2.5 42.54 2.76 ;
      RECT 43.25 2.025 43.255 2.25 ;
      RECT 43.38 2.025 43.435 2.235 ;
      RECT 43.435 2.03 43.445 2.228 ;
      RECT 43.341 2.025 43.38 2.238 ;
      RECT 43.255 2.025 43.341 2.245 ;
      RECT 43.235 2.03 43.25 2.251 ;
      RECT 43.225 2.07 43.235 2.253 ;
      RECT 43.195 2.08 43.225 2.255 ;
      RECT 43.19 2.085 43.195 2.257 ;
      RECT 43.165 2.09 43.19 2.259 ;
      RECT 43.15 2.095 43.165 2.261 ;
      RECT 43.135 2.097 43.15 2.263 ;
      RECT 43.13 2.102 43.135 2.265 ;
      RECT 43.08 2.11 43.13 2.268 ;
      RECT 43.055 2.119 43.08 2.273 ;
      RECT 43.045 2.126 43.055 2.278 ;
      RECT 43.04 2.129 43.045 2.282 ;
      RECT 43.02 2.132 43.04 2.291 ;
      RECT 42.99 2.14 43.02 2.311 ;
      RECT 42.961 2.153 42.99 2.333 ;
      RECT 42.875 2.187 42.961 2.377 ;
      RECT 42.87 2.213 42.875 2.415 ;
      RECT 42.865 2.217 42.87 2.424 ;
      RECT 42.83 2.23 42.865 2.457 ;
      RECT 42.82 2.244 42.83 2.495 ;
      RECT 42.815 2.248 42.82 2.508 ;
      RECT 42.81 2.252 42.815 2.513 ;
      RECT 42.8 2.26 42.81 2.525 ;
      RECT 42.795 2.267 42.8 2.54 ;
      RECT 42.77 2.28 42.795 2.565 ;
      RECT 42.73 2.309 42.77 2.62 ;
      RECT 42.715 2.334 42.73 2.675 ;
      RECT 42.705 2.345 42.715 2.698 ;
      RECT 42.7 2.352 42.705 2.71 ;
      RECT 42.695 2.356 42.7 2.718 ;
      RECT 42.64 2.384 42.695 2.76 ;
      RECT 42.62 2.42 42.64 2.76 ;
      RECT 42.605 2.435 42.62 2.76 ;
      RECT 42.55 2.467 42.605 2.76 ;
      RECT 42.54 2.497 42.55 2.76 ;
      RECT 42.15 2.112 42.335 2.35 ;
      RECT 42.135 2.114 42.345 2.345 ;
      RECT 42.02 2.06 42.28 2.32 ;
      RECT 42.015 2.097 42.28 2.274 ;
      RECT 42.01 2.107 42.28 2.271 ;
      RECT 42.005 2.147 42.345 2.265 ;
      RECT 42 2.18 42.345 2.255 ;
      RECT 42.01 2.122 42.36 2.193 ;
      RECT 42.307 3.22 42.32 3.75 ;
      RECT 42.221 3.22 42.32 3.749 ;
      RECT 42.221 3.22 42.325 3.748 ;
      RECT 42.135 3.22 42.325 3.746 ;
      RECT 42.13 3.22 42.325 3.743 ;
      RECT 42.13 3.22 42.335 3.741 ;
      RECT 42.125 3.512 42.335 3.738 ;
      RECT 42.125 3.522 42.34 3.735 ;
      RECT 42.125 3.59 42.345 3.731 ;
      RECT 42.115 3.595 42.345 3.73 ;
      RECT 42.115 3.687 42.35 3.727 ;
      RECT 42.1 3.22 42.36 3.48 ;
      RECT 42.03 7.765 42.32 7.995 ;
      RECT 42.09 7.025 42.26 7.995 ;
      RECT 42.005 7.055 42.345 7.4 ;
      RECT 42.03 7.025 42.32 7.4 ;
      RECT 41.33 2.21 41.375 3.745 ;
      RECT 41.53 2.21 41.56 2.425 ;
      RECT 39.905 1.95 40.025 2.16 ;
      RECT 39.565 1.9 39.825 2.16 ;
      RECT 39.565 1.945 39.86 2.15 ;
      RECT 41.57 2.226 41.575 2.28 ;
      RECT 41.565 2.219 41.57 2.413 ;
      RECT 41.56 2.213 41.565 2.42 ;
      RECT 41.515 2.21 41.53 2.433 ;
      RECT 41.51 2.21 41.515 2.455 ;
      RECT 41.505 2.21 41.51 2.503 ;
      RECT 41.5 2.21 41.505 2.523 ;
      RECT 41.49 2.21 41.5 2.63 ;
      RECT 41.485 2.21 41.49 2.693 ;
      RECT 41.48 2.21 41.485 2.75 ;
      RECT 41.475 2.21 41.48 2.758 ;
      RECT 41.46 2.21 41.475 2.865 ;
      RECT 41.45 2.21 41.46 3 ;
      RECT 41.44 2.21 41.45 3.11 ;
      RECT 41.43 2.21 41.44 3.167 ;
      RECT 41.425 2.21 41.43 3.207 ;
      RECT 41.42 2.21 41.425 3.243 ;
      RECT 41.41 2.21 41.42 3.283 ;
      RECT 41.405 2.21 41.41 3.325 ;
      RECT 41.385 2.21 41.405 3.39 ;
      RECT 41.39 3.535 41.395 3.715 ;
      RECT 41.385 3.517 41.39 3.723 ;
      RECT 41.38 2.21 41.385 3.453 ;
      RECT 41.38 3.497 41.385 3.73 ;
      RECT 41.375 2.21 41.38 3.74 ;
      RECT 41.32 2.21 41.33 2.51 ;
      RECT 41.325 2.757 41.33 3.745 ;
      RECT 41.32 2.822 41.325 3.745 ;
      RECT 41.315 2.211 41.32 2.5 ;
      RECT 41.31 2.887 41.32 3.745 ;
      RECT 41.305 2.212 41.315 2.49 ;
      RECT 41.295 3 41.31 3.745 ;
      RECT 41.3 2.213 41.305 2.48 ;
      RECT 41.28 2.214 41.3 2.458 ;
      RECT 41.285 3.097 41.295 3.745 ;
      RECT 41.28 3.172 41.285 3.745 ;
      RECT 41.27 2.213 41.28 2.435 ;
      RECT 41.275 3.215 41.28 3.745 ;
      RECT 41.27 3.242 41.275 3.745 ;
      RECT 41.26 2.211 41.27 2.423 ;
      RECT 41.265 3.285 41.27 3.745 ;
      RECT 41.26 3.312 41.265 3.745 ;
      RECT 41.25 2.21 41.26 2.41 ;
      RECT 41.255 3.327 41.26 3.745 ;
      RECT 41.215 3.385 41.255 3.745 ;
      RECT 41.245 2.209 41.25 2.395 ;
      RECT 41.24 2.207 41.245 2.388 ;
      RECT 41.23 2.204 41.24 2.378 ;
      RECT 41.225 2.201 41.23 2.363 ;
      RECT 41.21 2.197 41.225 2.356 ;
      RECT 41.205 3.44 41.215 3.745 ;
      RECT 41.205 2.194 41.21 2.351 ;
      RECT 41.19 2.19 41.205 2.345 ;
      RECT 41.2 3.457 41.205 3.745 ;
      RECT 41.19 3.52 41.2 3.745 ;
      RECT 41.11 2.175 41.19 2.325 ;
      RECT 41.185 3.527 41.19 3.74 ;
      RECT 41.18 3.535 41.185 3.73 ;
      RECT 41.1 2.161 41.11 2.309 ;
      RECT 41.085 2.157 41.1 2.307 ;
      RECT 41.075 2.152 41.085 2.303 ;
      RECT 41.05 2.145 41.075 2.295 ;
      RECT 41.045 2.14 41.05 2.29 ;
      RECT 41.035 2.14 41.045 2.288 ;
      RECT 41.025 2.138 41.035 2.286 ;
      RECT 40.995 2.13 41.025 2.28 ;
      RECT 40.98 2.122 40.995 2.273 ;
      RECT 40.96 2.117 40.98 2.266 ;
      RECT 40.955 2.113 40.96 2.261 ;
      RECT 40.925 2.106 40.955 2.255 ;
      RECT 40.9 2.097 40.925 2.245 ;
      RECT 40.87 2.09 40.9 2.237 ;
      RECT 40.845 2.08 40.87 2.228 ;
      RECT 40.83 2.072 40.845 2.222 ;
      RECT 40.805 2.067 40.83 2.217 ;
      RECT 40.795 2.063 40.805 2.212 ;
      RECT 40.775 2.058 40.795 2.207 ;
      RECT 40.74 2.053 40.775 2.2 ;
      RECT 40.68 2.048 40.74 2.193 ;
      RECT 40.667 2.044 40.68 2.191 ;
      RECT 40.581 2.039 40.667 2.188 ;
      RECT 40.495 2.029 40.581 2.184 ;
      RECT 40.454 2.022 40.495 2.181 ;
      RECT 40.368 2.015 40.454 2.178 ;
      RECT 40.282 2.005 40.368 2.174 ;
      RECT 40.196 1.995 40.282 2.169 ;
      RECT 40.11 1.985 40.196 2.165 ;
      RECT 40.1 1.97 40.11 2.163 ;
      RECT 40.09 1.955 40.1 2.163 ;
      RECT 40.025 1.95 40.09 2.162 ;
      RECT 39.86 1.947 39.905 2.155 ;
      RECT 41.105 2.852 41.11 3.043 ;
      RECT 41.1 2.847 41.105 3.05 ;
      RECT 41.086 2.845 41.1 3.056 ;
      RECT 41 2.845 41.086 3.058 ;
      RECT 40.996 2.845 41 3.061 ;
      RECT 40.91 2.845 40.996 3.079 ;
      RECT 40.9 2.85 40.91 3.098 ;
      RECT 40.89 2.905 40.9 3.102 ;
      RECT 40.865 2.92 40.89 3.109 ;
      RECT 40.825 2.94 40.865 3.122 ;
      RECT 40.82 2.952 40.825 3.132 ;
      RECT 40.805 2.958 40.82 3.137 ;
      RECT 40.8 2.963 40.805 3.141 ;
      RECT 40.78 2.97 40.8 3.146 ;
      RECT 40.71 2.995 40.78 3.163 ;
      RECT 40.67 3.023 40.71 3.183 ;
      RECT 40.665 3.033 40.67 3.191 ;
      RECT 40.645 3.04 40.665 3.193 ;
      RECT 40.64 3.047 40.645 3.196 ;
      RECT 40.61 3.055 40.64 3.199 ;
      RECT 40.605 3.06 40.61 3.203 ;
      RECT 40.531 3.064 40.605 3.211 ;
      RECT 40.445 3.073 40.531 3.227 ;
      RECT 40.441 3.078 40.445 3.236 ;
      RECT 40.355 3.083 40.441 3.246 ;
      RECT 40.315 3.091 40.355 3.258 ;
      RECT 40.265 3.097 40.315 3.265 ;
      RECT 40.18 3.106 40.265 3.28 ;
      RECT 40.105 3.117 40.18 3.298 ;
      RECT 40.07 3.124 40.105 3.308 ;
      RECT 39.995 3.132 40.07 3.313 ;
      RECT 39.94 3.141 39.995 3.313 ;
      RECT 39.915 3.146 39.94 3.311 ;
      RECT 39.905 3.149 39.915 3.309 ;
      RECT 39.87 3.151 39.905 3.307 ;
      RECT 39.84 3.153 39.87 3.303 ;
      RECT 39.795 3.152 39.84 3.299 ;
      RECT 39.775 3.147 39.795 3.296 ;
      RECT 39.725 3.132 39.775 3.293 ;
      RECT 39.715 3.117 39.725 3.288 ;
      RECT 39.665 3.102 39.715 3.278 ;
      RECT 39.615 3.077 39.665 3.258 ;
      RECT 39.605 3.062 39.615 3.24 ;
      RECT 39.6 3.06 39.605 3.234 ;
      RECT 39.58 3.055 39.6 3.229 ;
      RECT 39.575 3.047 39.58 3.223 ;
      RECT 39.56 3.041 39.575 3.216 ;
      RECT 39.555 3.036 39.56 3.208 ;
      RECT 39.535 3.031 39.555 3.2 ;
      RECT 39.52 3.024 39.535 3.193 ;
      RECT 39.505 3.018 39.52 3.184 ;
      RECT 39.5 3.012 39.505 3.177 ;
      RECT 39.455 2.987 39.5 3.163 ;
      RECT 39.44 2.957 39.455 3.145 ;
      RECT 39.425 2.94 39.44 3.136 ;
      RECT 39.4 2.92 39.425 3.124 ;
      RECT 39.36 2.89 39.4 3.104 ;
      RECT 39.35 2.86 39.36 3.089 ;
      RECT 39.335 2.85 39.35 3.082 ;
      RECT 39.28 2.815 39.335 3.061 ;
      RECT 39.265 2.778 39.28 3.04 ;
      RECT 39.255 2.765 39.265 3.032 ;
      RECT 39.205 2.735 39.255 3.014 ;
      RECT 39.19 2.665 39.205 2.995 ;
      RECT 39.145 2.665 39.19 2.978 ;
      RECT 39.12 2.665 39.145 2.96 ;
      RECT 39.11 2.665 39.12 2.953 ;
      RECT 39.031 2.665 39.11 2.946 ;
      RECT 38.945 2.665 39.031 2.938 ;
      RECT 38.93 2.697 38.945 2.933 ;
      RECT 38.855 2.707 38.93 2.929 ;
      RECT 38.835 2.717 38.855 2.924 ;
      RECT 38.81 2.717 38.835 2.921 ;
      RECT 38.8 2.707 38.81 2.92 ;
      RECT 38.79 2.68 38.8 2.919 ;
      RECT 38.75 2.675 38.79 2.917 ;
      RECT 38.705 2.675 38.75 2.913 ;
      RECT 38.68 2.675 38.705 2.908 ;
      RECT 38.63 2.675 38.68 2.895 ;
      RECT 38.59 2.68 38.6 2.88 ;
      RECT 38.6 2.675 38.63 2.885 ;
      RECT 40.585 2.455 40.845 2.715 ;
      RECT 40.58 2.477 40.845 2.673 ;
      RECT 39.82 2.305 40.04 2.67 ;
      RECT 39.802 2.392 40.04 2.669 ;
      RECT 39.785 2.397 40.04 2.666 ;
      RECT 39.785 2.397 40.06 2.665 ;
      RECT 39.755 2.407 40.06 2.663 ;
      RECT 39.75 2.422 40.06 2.659 ;
      RECT 39.75 2.422 40.065 2.658 ;
      RECT 39.745 2.48 40.065 2.656 ;
      RECT 39.745 2.48 40.075 2.653 ;
      RECT 39.74 2.545 40.075 2.648 ;
      RECT 39.82 2.305 40.08 2.565 ;
      RECT 38.565 2.135 38.825 2.395 ;
      RECT 38.565 2.178 38.911 2.369 ;
      RECT 38.565 2.178 38.955 2.368 ;
      RECT 38.565 2.178 38.975 2.366 ;
      RECT 38.565 2.178 39.075 2.365 ;
      RECT 38.565 2.178 39.095 2.363 ;
      RECT 38.565 2.178 39.105 2.358 ;
      RECT 38.975 2.145 39.165 2.355 ;
      RECT 38.975 2.147 39.17 2.353 ;
      RECT 38.965 2.152 39.175 2.345 ;
      RECT 38.911 2.176 39.175 2.345 ;
      RECT 38.955 2.17 38.965 2.367 ;
      RECT 38.965 2.15 39.17 2.353 ;
      RECT 37.92 3.21 38.125 3.44 ;
      RECT 37.86 3.16 37.915 3.42 ;
      RECT 37.92 3.16 38.12 3.44 ;
      RECT 38.89 3.475 38.895 3.502 ;
      RECT 38.88 3.385 38.89 3.507 ;
      RECT 38.875 3.307 38.88 3.513 ;
      RECT 38.865 3.297 38.875 3.52 ;
      RECT 38.86 3.287 38.865 3.526 ;
      RECT 38.85 3.282 38.86 3.528 ;
      RECT 38.835 3.274 38.85 3.536 ;
      RECT 38.82 3.265 38.835 3.548 ;
      RECT 38.81 3.257 38.82 3.558 ;
      RECT 38.775 3.175 38.81 3.576 ;
      RECT 38.74 3.175 38.775 3.595 ;
      RECT 38.725 3.175 38.74 3.603 ;
      RECT 38.67 3.175 38.725 3.603 ;
      RECT 38.636 3.175 38.67 3.594 ;
      RECT 38.55 3.175 38.636 3.57 ;
      RECT 38.54 3.235 38.55 3.552 ;
      RECT 38.5 3.237 38.54 3.543 ;
      RECT 38.495 3.239 38.5 3.533 ;
      RECT 38.475 3.241 38.495 3.528 ;
      RECT 38.465 3.244 38.475 3.523 ;
      RECT 38.455 3.245 38.465 3.518 ;
      RECT 38.431 3.246 38.455 3.51 ;
      RECT 38.345 3.251 38.431 3.488 ;
      RECT 38.29 3.25 38.345 3.461 ;
      RECT 38.275 3.243 38.29 3.448 ;
      RECT 38.24 3.238 38.275 3.444 ;
      RECT 38.185 3.23 38.24 3.443 ;
      RECT 38.125 3.217 38.185 3.441 ;
      RECT 37.915 3.16 37.92 3.428 ;
      RECT 37.99 2.53 38.175 2.74 ;
      RECT 37.98 2.535 38.19 2.733 ;
      RECT 38.02 2.44 38.28 2.7 ;
      RECT 37.975 2.597 38.28 2.623 ;
      RECT 37.32 2.39 37.325 3.19 ;
      RECT 37.265 2.44 37.295 3.19 ;
      RECT 37.255 2.44 37.26 2.75 ;
      RECT 37.24 2.44 37.245 2.745 ;
      RECT 36.785 2.485 36.8 2.7 ;
      RECT 36.715 2.485 36.8 2.695 ;
      RECT 37.98 2.065 38.05 2.275 ;
      RECT 38.05 2.072 38.06 2.27 ;
      RECT 37.946 2.065 37.98 2.282 ;
      RECT 37.86 2.065 37.946 2.306 ;
      RECT 37.85 2.07 37.86 2.325 ;
      RECT 37.845 2.082 37.85 2.328 ;
      RECT 37.83 2.097 37.845 2.332 ;
      RECT 37.825 2.115 37.83 2.336 ;
      RECT 37.785 2.125 37.825 2.345 ;
      RECT 37.77 2.132 37.785 2.357 ;
      RECT 37.755 2.137 37.77 2.362 ;
      RECT 37.74 2.14 37.755 2.367 ;
      RECT 37.73 2.142 37.74 2.371 ;
      RECT 37.695 2.149 37.73 2.379 ;
      RECT 37.66 2.157 37.695 2.393 ;
      RECT 37.65 2.163 37.66 2.402 ;
      RECT 37.645 2.165 37.65 2.404 ;
      RECT 37.625 2.168 37.645 2.41 ;
      RECT 37.595 2.175 37.625 2.421 ;
      RECT 37.585 2.181 37.595 2.428 ;
      RECT 37.56 2.184 37.585 2.435 ;
      RECT 37.55 2.188 37.56 2.443 ;
      RECT 37.545 2.189 37.55 2.465 ;
      RECT 37.54 2.19 37.545 2.48 ;
      RECT 37.535 2.191 37.54 2.495 ;
      RECT 37.53 2.192 37.535 2.51 ;
      RECT 37.525 2.193 37.53 2.54 ;
      RECT 37.515 2.195 37.525 2.573 ;
      RECT 37.5 2.199 37.515 2.62 ;
      RECT 37.49 2.202 37.5 2.665 ;
      RECT 37.485 2.205 37.49 2.693 ;
      RECT 37.475 2.207 37.485 2.72 ;
      RECT 37.47 2.21 37.475 2.755 ;
      RECT 37.44 2.215 37.47 2.813 ;
      RECT 37.435 2.22 37.44 2.898 ;
      RECT 37.43 2.222 37.435 2.933 ;
      RECT 37.425 2.224 37.43 3.015 ;
      RECT 37.42 2.226 37.425 3.103 ;
      RECT 37.41 2.228 37.42 3.185 ;
      RECT 37.395 2.242 37.41 3.19 ;
      RECT 37.36 2.287 37.395 3.19 ;
      RECT 37.35 2.327 37.36 3.19 ;
      RECT 37.335 2.355 37.35 3.19 ;
      RECT 37.33 2.372 37.335 3.19 ;
      RECT 37.325 2.38 37.33 3.19 ;
      RECT 37.315 2.395 37.32 3.19 ;
      RECT 37.31 2.402 37.315 3.19 ;
      RECT 37.3 2.422 37.31 3.19 ;
      RECT 37.295 2.435 37.3 3.19 ;
      RECT 37.26 2.44 37.265 2.775 ;
      RECT 37.245 2.83 37.265 3.19 ;
      RECT 37.245 2.44 37.255 2.748 ;
      RECT 37.24 2.87 37.245 3.19 ;
      RECT 37.19 2.44 37.24 2.743 ;
      RECT 37.235 2.907 37.24 3.19 ;
      RECT 37.225 2.93 37.235 3.19 ;
      RECT 37.22 2.975 37.225 3.19 ;
      RECT 37.21 2.985 37.22 3.183 ;
      RECT 37.136 2.44 37.19 2.737 ;
      RECT 37.05 2.44 37.136 2.73 ;
      RECT 37.001 2.487 37.05 2.723 ;
      RECT 36.915 2.495 37.001 2.716 ;
      RECT 36.9 2.492 36.915 2.711 ;
      RECT 36.886 2.485 36.9 2.71 ;
      RECT 36.8 2.485 36.886 2.705 ;
      RECT 36.705 2.49 36.715 2.69 ;
      RECT 36.295 1.92 36.31 2.32 ;
      RECT 36.49 1.92 36.495 2.18 ;
      RECT 36.235 1.92 36.28 2.18 ;
      RECT 36.69 3.225 36.695 3.43 ;
      RECT 36.685 3.215 36.69 3.435 ;
      RECT 36.68 3.202 36.685 3.44 ;
      RECT 36.675 3.182 36.68 3.44 ;
      RECT 36.65 3.135 36.675 3.44 ;
      RECT 36.615 3.05 36.65 3.44 ;
      RECT 36.61 2.987 36.615 3.44 ;
      RECT 36.605 2.972 36.61 3.44 ;
      RECT 36.59 2.932 36.605 3.44 ;
      RECT 36.585 2.907 36.59 3.44 ;
      RECT 36.575 2.89 36.585 3.44 ;
      RECT 36.54 2.812 36.575 3.44 ;
      RECT 36.535 2.755 36.54 3.44 ;
      RECT 36.53 2.742 36.535 3.44 ;
      RECT 36.52 2.72 36.53 3.44 ;
      RECT 36.51 2.685 36.52 3.44 ;
      RECT 36.5 2.655 36.51 3.44 ;
      RECT 36.49 2.57 36.5 3.083 ;
      RECT 36.497 3.215 36.5 3.44 ;
      RECT 36.495 3.225 36.497 3.44 ;
      RECT 36.485 3.235 36.495 3.435 ;
      RECT 36.48 1.92 36.49 2.315 ;
      RECT 36.485 2.447 36.49 3.058 ;
      RECT 36.48 2.345 36.485 3.041 ;
      RECT 36.47 1.92 36.48 3.017 ;
      RECT 36.465 1.92 36.47 2.988 ;
      RECT 36.46 1.92 36.465 2.978 ;
      RECT 36.44 1.92 36.46 2.94 ;
      RECT 36.435 1.92 36.44 2.898 ;
      RECT 36.43 1.92 36.435 2.878 ;
      RECT 36.4 1.92 36.43 2.828 ;
      RECT 36.39 1.92 36.4 2.775 ;
      RECT 36.385 1.92 36.39 2.748 ;
      RECT 36.38 1.92 36.385 2.733 ;
      RECT 36.37 1.92 36.38 2.71 ;
      RECT 36.36 1.92 36.37 2.685 ;
      RECT 36.355 1.92 36.36 2.625 ;
      RECT 36.345 1.92 36.355 2.563 ;
      RECT 36.34 1.92 36.345 2.483 ;
      RECT 36.335 1.92 36.34 2.448 ;
      RECT 36.33 1.92 36.335 2.423 ;
      RECT 36.325 1.92 36.33 2.408 ;
      RECT 36.32 1.92 36.325 2.378 ;
      RECT 36.315 1.92 36.32 2.355 ;
      RECT 36.31 1.92 36.315 2.328 ;
      RECT 36.28 1.92 36.295 2.315 ;
      RECT 35.435 3.455 35.62 3.665 ;
      RECT 35.425 3.46 35.635 3.658 ;
      RECT 35.425 3.46 35.655 3.63 ;
      RECT 35.425 3.46 35.67 3.609 ;
      RECT 35.425 3.46 35.685 3.607 ;
      RECT 35.425 3.46 35.695 3.606 ;
      RECT 35.425 3.46 35.725 3.603 ;
      RECT 36.075 3.305 36.335 3.565 ;
      RECT 36.035 3.352 36.335 3.548 ;
      RECT 36.026 3.36 36.035 3.551 ;
      RECT 35.62 3.453 36.335 3.548 ;
      RECT 35.94 3.378 36.026 3.558 ;
      RECT 35.635 3.45 36.335 3.548 ;
      RECT 35.881 3.4 35.94 3.57 ;
      RECT 35.655 3.446 36.335 3.548 ;
      RECT 35.795 3.412 35.881 3.581 ;
      RECT 35.67 3.442 36.335 3.548 ;
      RECT 35.74 3.425 35.795 3.593 ;
      RECT 35.685 3.44 36.335 3.548 ;
      RECT 35.725 3.431 35.74 3.599 ;
      RECT 35.695 3.436 36.335 3.548 ;
      RECT 35.84 2.96 36.1 3.22 ;
      RECT 35.84 2.98 36.21 3.19 ;
      RECT 35.84 2.985 36.22 3.185 ;
      RECT 36.031 2.399 36.11 2.63 ;
      RECT 35.945 2.402 36.16 2.625 ;
      RECT 35.94 2.402 36.16 2.62 ;
      RECT 35.94 2.407 36.17 2.618 ;
      RECT 35.915 2.407 36.17 2.615 ;
      RECT 35.915 2.415 36.18 2.613 ;
      RECT 35.795 2.35 36.055 2.61 ;
      RECT 35.795 2.397 36.105 2.61 ;
      RECT 35.05 2.97 35.055 3.23 ;
      RECT 34.88 2.74 34.885 3.23 ;
      RECT 34.765 2.98 34.77 3.205 ;
      RECT 35.475 2.075 35.48 2.285 ;
      RECT 35.48 2.08 35.495 2.28 ;
      RECT 35.415 2.075 35.475 2.293 ;
      RECT 35.4 2.075 35.415 2.303 ;
      RECT 35.35 2.075 35.4 2.32 ;
      RECT 35.33 2.075 35.35 2.343 ;
      RECT 35.315 2.075 35.33 2.355 ;
      RECT 35.295 2.075 35.315 2.365 ;
      RECT 35.285 2.08 35.295 2.374 ;
      RECT 35.28 2.09 35.285 2.379 ;
      RECT 35.275 2.102 35.28 2.383 ;
      RECT 35.265 2.125 35.275 2.388 ;
      RECT 35.26 2.14 35.265 2.392 ;
      RECT 35.255 2.157 35.26 2.395 ;
      RECT 35.25 2.165 35.255 2.398 ;
      RECT 35.24 2.17 35.25 2.402 ;
      RECT 35.235 2.177 35.24 2.407 ;
      RECT 35.225 2.182 35.235 2.411 ;
      RECT 35.2 2.194 35.225 2.422 ;
      RECT 35.18 2.211 35.2 2.438 ;
      RECT 35.155 2.228 35.18 2.46 ;
      RECT 35.12 2.251 35.155 2.518 ;
      RECT 35.1 2.273 35.12 2.58 ;
      RECT 35.095 2.283 35.1 2.615 ;
      RECT 35.085 2.29 35.095 2.653 ;
      RECT 35.08 2.297 35.085 2.673 ;
      RECT 35.075 2.308 35.08 2.71 ;
      RECT 35.07 2.316 35.075 2.775 ;
      RECT 35.06 2.327 35.07 2.828 ;
      RECT 35.055 2.345 35.06 2.898 ;
      RECT 35.05 2.355 35.055 2.935 ;
      RECT 35.045 2.365 35.05 3.23 ;
      RECT 35.04 2.377 35.045 3.23 ;
      RECT 35.035 2.387 35.04 3.23 ;
      RECT 35.025 2.397 35.035 3.23 ;
      RECT 35.015 2.42 35.025 3.23 ;
      RECT 35 2.455 35.015 3.23 ;
      RECT 34.96 2.517 35 3.23 ;
      RECT 34.955 2.57 34.96 3.23 ;
      RECT 34.93 2.605 34.955 3.23 ;
      RECT 34.915 2.65 34.93 3.23 ;
      RECT 34.91 2.672 34.915 3.23 ;
      RECT 34.9 2.685 34.91 3.23 ;
      RECT 34.89 2.71 34.9 3.23 ;
      RECT 34.885 2.732 34.89 3.23 ;
      RECT 34.86 2.77 34.88 3.23 ;
      RECT 34.82 2.827 34.86 3.23 ;
      RECT 34.815 2.877 34.82 3.23 ;
      RECT 34.81 2.895 34.815 3.23 ;
      RECT 34.805 2.907 34.81 3.23 ;
      RECT 34.795 2.925 34.805 3.23 ;
      RECT 34.785 2.945 34.795 3.205 ;
      RECT 34.78 2.962 34.785 3.205 ;
      RECT 34.77 2.975 34.78 3.205 ;
      RECT 34.74 2.985 34.765 3.205 ;
      RECT 34.73 2.992 34.74 3.205 ;
      RECT 34.715 3.002 34.73 3.2 ;
      RECT 33.815 7.77 34.105 8 ;
      RECT 33.875 6.29 34.045 8 ;
      RECT 33.865 6.66 34.22 7.015 ;
      RECT 33.815 6.29 34.105 6.52 ;
      RECT 33.41 2.395 33.515 2.965 ;
      RECT 33.41 2.73 33.735 2.96 ;
      RECT 33.41 2.76 33.905 2.93 ;
      RECT 33.41 2.395 33.6 2.96 ;
      RECT 32.825 2.36 33.115 2.59 ;
      RECT 32.825 2.395 33.6 2.565 ;
      RECT 32.885 0.88 33.055 2.59 ;
      RECT 32.825 0.88 33.115 1.11 ;
      RECT 32.825 7.77 33.115 8 ;
      RECT 32.885 6.29 33.055 8 ;
      RECT 32.825 6.29 33.115 6.52 ;
      RECT 32.825 6.325 33.68 6.485 ;
      RECT 33.51 5.92 33.68 6.485 ;
      RECT 32.825 6.32 33.22 6.485 ;
      RECT 33.445 5.92 33.735 6.15 ;
      RECT 33.445 5.95 33.905 6.12 ;
      RECT 32.455 2.73 32.745 2.96 ;
      RECT 32.455 2.76 32.915 2.93 ;
      RECT 32.52 1.655 32.685 2.96 ;
      RECT 31.035 1.625 31.325 1.855 ;
      RECT 31.035 1.655 32.685 1.825 ;
      RECT 31.095 0.885 31.265 1.855 ;
      RECT 31.035 0.885 31.325 1.115 ;
      RECT 31.035 7.765 31.325 7.995 ;
      RECT 31.095 7.025 31.265 7.995 ;
      RECT 31.095 7.12 32.685 7.29 ;
      RECT 32.515 5.92 32.685 7.29 ;
      RECT 31.035 7.025 31.325 7.255 ;
      RECT 32.455 5.92 32.745 6.15 ;
      RECT 32.455 5.95 32.915 6.12 ;
      RECT 31.465 1.965 31.815 2.315 ;
      RECT 29.13 2.025 31.815 2.195 ;
      RECT 29.13 1.34 29.3 2.195 ;
      RECT 29.03 1.34 29.38 1.69 ;
      RECT 31.49 6.655 31.815 6.98 ;
      RECT 26.915 6.61 27.265 6.96 ;
      RECT 31.465 6.655 31.815 6.885 ;
      RECT 26.685 6.655 27.265 6.885 ;
      RECT 26.515 6.685 31.815 6.855 ;
      RECT 30.69 2.365 31.01 2.685 ;
      RECT 30.66 2.365 31.01 2.595 ;
      RECT 30.49 2.395 31.01 2.565 ;
      RECT 30.69 6.255 31.01 6.545 ;
      RECT 30.66 6.285 31.01 6.515 ;
      RECT 30.49 6.315 31.01 6.485 ;
      RECT 27.325 2.465 27.51 2.675 ;
      RECT 27.315 2.47 27.525 2.668 ;
      RECT 27.315 2.47 27.611 2.645 ;
      RECT 27.315 2.47 27.67 2.62 ;
      RECT 27.315 2.47 27.725 2.6 ;
      RECT 27.315 2.47 27.735 2.588 ;
      RECT 27.315 2.47 27.93 2.527 ;
      RECT 27.315 2.47 27.96 2.51 ;
      RECT 27.315 2.47 27.98 2.5 ;
      RECT 27.86 2.235 28.12 2.495 ;
      RECT 27.845 2.325 27.86 2.542 ;
      RECT 27.38 2.457 28.12 2.495 ;
      RECT 27.831 2.336 27.845 2.548 ;
      RECT 27.42 2.45 28.12 2.495 ;
      RECT 27.745 2.376 27.831 2.567 ;
      RECT 27.67 2.437 28.12 2.495 ;
      RECT 27.74 2.412 27.745 2.584 ;
      RECT 27.725 2.422 28.12 2.495 ;
      RECT 27.735 2.417 27.74 2.586 ;
      RECT 28.03 2.922 28.035 3.014 ;
      RECT 28.025 2.9 28.03 3.031 ;
      RECT 28.02 2.89 28.025 3.043 ;
      RECT 28.01 2.881 28.02 3.053 ;
      RECT 28.005 2.876 28.01 3.061 ;
      RECT 28 2.735 28.005 3.064 ;
      RECT 27.966 2.735 28 3.075 ;
      RECT 27.88 2.735 27.966 3.11 ;
      RECT 27.8 2.735 27.88 3.158 ;
      RECT 27.771 2.735 27.8 3.182 ;
      RECT 27.685 2.735 27.771 3.188 ;
      RECT 27.68 2.919 27.685 3.193 ;
      RECT 27.645 2.93 27.68 3.196 ;
      RECT 27.62 2.945 27.645 3.2 ;
      RECT 27.606 2.954 27.62 3.202 ;
      RECT 27.52 2.981 27.606 3.208 ;
      RECT 27.455 3.022 27.52 3.217 ;
      RECT 27.44 3.042 27.455 3.222 ;
      RECT 27.41 3.052 27.44 3.225 ;
      RECT 27.405 3.062 27.41 3.228 ;
      RECT 27.375 3.067 27.405 3.23 ;
      RECT 27.355 3.072 27.375 3.234 ;
      RECT 27.27 3.075 27.355 3.241 ;
      RECT 27.255 3.072 27.27 3.247 ;
      RECT 27.245 3.069 27.255 3.249 ;
      RECT 27.225 3.066 27.245 3.251 ;
      RECT 27.205 3.062 27.225 3.252 ;
      RECT 27.19 3.058 27.205 3.254 ;
      RECT 27.18 3.055 27.19 3.255 ;
      RECT 27.14 3.049 27.18 3.253 ;
      RECT 27.13 3.044 27.14 3.251 ;
      RECT 27.115 3.041 27.13 3.247 ;
      RECT 27.09 3.036 27.115 3.24 ;
      RECT 27.04 3.027 27.09 3.228 ;
      RECT 26.97 3.013 27.04 3.21 ;
      RECT 26.912 2.998 26.97 3.192 ;
      RECT 26.826 2.981 26.912 3.172 ;
      RECT 26.74 2.96 26.826 3.147 ;
      RECT 26.69 2.945 26.74 3.128 ;
      RECT 26.686 2.939 26.69 3.12 ;
      RECT 26.6 2.929 26.686 3.107 ;
      RECT 26.565 2.914 26.6 3.09 ;
      RECT 26.55 2.907 26.565 3.083 ;
      RECT 26.49 2.895 26.55 3.071 ;
      RECT 26.47 2.882 26.49 3.059 ;
      RECT 26.43 2.873 26.47 3.051 ;
      RECT 26.425 2.865 26.43 3.044 ;
      RECT 26.345 2.855 26.425 3.03 ;
      RECT 26.33 2.842 26.345 3.015 ;
      RECT 26.325 2.84 26.33 3.013 ;
      RECT 26.246 2.828 26.325 3 ;
      RECT 26.16 2.803 26.246 2.975 ;
      RECT 26.145 2.772 26.16 2.96 ;
      RECT 26.13 2.747 26.145 2.956 ;
      RECT 26.115 2.74 26.13 2.952 ;
      RECT 25.94 2.745 25.945 2.948 ;
      RECT 25.935 2.75 25.94 2.943 ;
      RECT 25.945 2.74 26.115 2.95 ;
      RECT 26.66 2.5 26.765 2.76 ;
      RECT 27.475 2.025 27.48 2.25 ;
      RECT 27.605 2.025 27.66 2.235 ;
      RECT 27.66 2.03 27.67 2.228 ;
      RECT 27.566 2.025 27.605 2.238 ;
      RECT 27.48 2.025 27.566 2.245 ;
      RECT 27.46 2.03 27.475 2.251 ;
      RECT 27.45 2.07 27.46 2.253 ;
      RECT 27.42 2.08 27.45 2.255 ;
      RECT 27.415 2.085 27.42 2.257 ;
      RECT 27.39 2.09 27.415 2.259 ;
      RECT 27.375 2.095 27.39 2.261 ;
      RECT 27.36 2.097 27.375 2.263 ;
      RECT 27.355 2.102 27.36 2.265 ;
      RECT 27.305 2.11 27.355 2.268 ;
      RECT 27.28 2.119 27.305 2.273 ;
      RECT 27.27 2.126 27.28 2.278 ;
      RECT 27.265 2.129 27.27 2.282 ;
      RECT 27.245 2.132 27.265 2.291 ;
      RECT 27.215 2.14 27.245 2.311 ;
      RECT 27.186 2.153 27.215 2.333 ;
      RECT 27.1 2.187 27.186 2.377 ;
      RECT 27.095 2.213 27.1 2.415 ;
      RECT 27.09 2.217 27.095 2.424 ;
      RECT 27.055 2.23 27.09 2.457 ;
      RECT 27.045 2.244 27.055 2.495 ;
      RECT 27.04 2.248 27.045 2.508 ;
      RECT 27.035 2.252 27.04 2.513 ;
      RECT 27.025 2.26 27.035 2.525 ;
      RECT 27.02 2.267 27.025 2.54 ;
      RECT 26.995 2.28 27.02 2.565 ;
      RECT 26.955 2.309 26.995 2.62 ;
      RECT 26.94 2.334 26.955 2.675 ;
      RECT 26.93 2.345 26.94 2.698 ;
      RECT 26.925 2.352 26.93 2.71 ;
      RECT 26.92 2.356 26.925 2.718 ;
      RECT 26.865 2.384 26.92 2.76 ;
      RECT 26.845 2.42 26.865 2.76 ;
      RECT 26.83 2.435 26.845 2.76 ;
      RECT 26.775 2.467 26.83 2.76 ;
      RECT 26.765 2.497 26.775 2.76 ;
      RECT 26.375 2.112 26.56 2.35 ;
      RECT 26.36 2.114 26.57 2.345 ;
      RECT 26.245 2.06 26.505 2.32 ;
      RECT 26.24 2.097 26.505 2.274 ;
      RECT 26.235 2.107 26.505 2.271 ;
      RECT 26.23 2.147 26.57 2.265 ;
      RECT 26.225 2.18 26.57 2.255 ;
      RECT 26.235 2.122 26.585 2.193 ;
      RECT 26.532 3.22 26.545 3.75 ;
      RECT 26.446 3.22 26.545 3.749 ;
      RECT 26.446 3.22 26.55 3.748 ;
      RECT 26.36 3.22 26.55 3.746 ;
      RECT 26.355 3.22 26.55 3.743 ;
      RECT 26.355 3.22 26.56 3.741 ;
      RECT 26.35 3.512 26.56 3.738 ;
      RECT 26.35 3.522 26.565 3.735 ;
      RECT 26.35 3.59 26.57 3.731 ;
      RECT 26.34 3.595 26.57 3.73 ;
      RECT 26.34 3.687 26.575 3.727 ;
      RECT 26.325 3.22 26.585 3.48 ;
      RECT 26.255 7.765 26.545 7.995 ;
      RECT 26.315 7.025 26.485 7.995 ;
      RECT 26.23 7.055 26.57 7.4 ;
      RECT 26.255 7.025 26.545 7.4 ;
      RECT 25.555 2.21 25.6 3.745 ;
      RECT 25.755 2.21 25.785 2.425 ;
      RECT 24.13 1.95 24.25 2.16 ;
      RECT 23.79 1.9 24.05 2.16 ;
      RECT 23.79 1.945 24.085 2.15 ;
      RECT 25.795 2.226 25.8 2.28 ;
      RECT 25.79 2.219 25.795 2.413 ;
      RECT 25.785 2.213 25.79 2.42 ;
      RECT 25.74 2.21 25.755 2.433 ;
      RECT 25.735 2.21 25.74 2.455 ;
      RECT 25.73 2.21 25.735 2.503 ;
      RECT 25.725 2.21 25.73 2.523 ;
      RECT 25.715 2.21 25.725 2.63 ;
      RECT 25.71 2.21 25.715 2.693 ;
      RECT 25.705 2.21 25.71 2.75 ;
      RECT 25.7 2.21 25.705 2.758 ;
      RECT 25.685 2.21 25.7 2.865 ;
      RECT 25.675 2.21 25.685 3 ;
      RECT 25.665 2.21 25.675 3.11 ;
      RECT 25.655 2.21 25.665 3.167 ;
      RECT 25.65 2.21 25.655 3.207 ;
      RECT 25.645 2.21 25.65 3.243 ;
      RECT 25.635 2.21 25.645 3.283 ;
      RECT 25.63 2.21 25.635 3.325 ;
      RECT 25.61 2.21 25.63 3.39 ;
      RECT 25.615 3.535 25.62 3.715 ;
      RECT 25.61 3.517 25.615 3.723 ;
      RECT 25.605 2.21 25.61 3.453 ;
      RECT 25.605 3.497 25.61 3.73 ;
      RECT 25.6 2.21 25.605 3.74 ;
      RECT 25.545 2.21 25.555 2.51 ;
      RECT 25.55 2.757 25.555 3.745 ;
      RECT 25.545 2.822 25.55 3.745 ;
      RECT 25.54 2.211 25.545 2.5 ;
      RECT 25.535 2.887 25.545 3.745 ;
      RECT 25.53 2.212 25.54 2.49 ;
      RECT 25.52 3 25.535 3.745 ;
      RECT 25.525 2.213 25.53 2.48 ;
      RECT 25.505 2.214 25.525 2.458 ;
      RECT 25.51 3.097 25.52 3.745 ;
      RECT 25.505 3.172 25.51 3.745 ;
      RECT 25.495 2.213 25.505 2.435 ;
      RECT 25.5 3.215 25.505 3.745 ;
      RECT 25.495 3.242 25.5 3.745 ;
      RECT 25.485 2.211 25.495 2.423 ;
      RECT 25.49 3.285 25.495 3.745 ;
      RECT 25.485 3.312 25.49 3.745 ;
      RECT 25.475 2.21 25.485 2.41 ;
      RECT 25.48 3.327 25.485 3.745 ;
      RECT 25.44 3.385 25.48 3.745 ;
      RECT 25.47 2.209 25.475 2.395 ;
      RECT 25.465 2.207 25.47 2.388 ;
      RECT 25.455 2.204 25.465 2.378 ;
      RECT 25.45 2.201 25.455 2.363 ;
      RECT 25.435 2.197 25.45 2.356 ;
      RECT 25.43 3.44 25.44 3.745 ;
      RECT 25.43 2.194 25.435 2.351 ;
      RECT 25.415 2.19 25.43 2.345 ;
      RECT 25.425 3.457 25.43 3.745 ;
      RECT 25.415 3.52 25.425 3.745 ;
      RECT 25.335 2.175 25.415 2.325 ;
      RECT 25.41 3.527 25.415 3.74 ;
      RECT 25.405 3.535 25.41 3.73 ;
      RECT 25.325 2.161 25.335 2.309 ;
      RECT 25.31 2.157 25.325 2.307 ;
      RECT 25.3 2.152 25.31 2.303 ;
      RECT 25.275 2.145 25.3 2.295 ;
      RECT 25.27 2.14 25.275 2.29 ;
      RECT 25.26 2.14 25.27 2.288 ;
      RECT 25.25 2.138 25.26 2.286 ;
      RECT 25.22 2.13 25.25 2.28 ;
      RECT 25.205 2.122 25.22 2.273 ;
      RECT 25.185 2.117 25.205 2.266 ;
      RECT 25.18 2.113 25.185 2.261 ;
      RECT 25.15 2.106 25.18 2.255 ;
      RECT 25.125 2.097 25.15 2.245 ;
      RECT 25.095 2.09 25.125 2.237 ;
      RECT 25.07 2.08 25.095 2.228 ;
      RECT 25.055 2.072 25.07 2.222 ;
      RECT 25.03 2.067 25.055 2.217 ;
      RECT 25.02 2.063 25.03 2.212 ;
      RECT 25 2.058 25.02 2.207 ;
      RECT 24.965 2.053 25 2.2 ;
      RECT 24.905 2.048 24.965 2.193 ;
      RECT 24.892 2.044 24.905 2.191 ;
      RECT 24.806 2.039 24.892 2.188 ;
      RECT 24.72 2.029 24.806 2.184 ;
      RECT 24.679 2.022 24.72 2.181 ;
      RECT 24.593 2.015 24.679 2.178 ;
      RECT 24.507 2.005 24.593 2.174 ;
      RECT 24.421 1.995 24.507 2.169 ;
      RECT 24.335 1.985 24.421 2.165 ;
      RECT 24.325 1.97 24.335 2.163 ;
      RECT 24.315 1.955 24.325 2.163 ;
      RECT 24.25 1.95 24.315 2.162 ;
      RECT 24.085 1.947 24.13 2.155 ;
      RECT 25.33 2.852 25.335 3.043 ;
      RECT 25.325 2.847 25.33 3.05 ;
      RECT 25.311 2.845 25.325 3.056 ;
      RECT 25.225 2.845 25.311 3.058 ;
      RECT 25.221 2.845 25.225 3.061 ;
      RECT 25.135 2.845 25.221 3.079 ;
      RECT 25.125 2.85 25.135 3.098 ;
      RECT 25.115 2.905 25.125 3.102 ;
      RECT 25.09 2.92 25.115 3.109 ;
      RECT 25.05 2.94 25.09 3.122 ;
      RECT 25.045 2.952 25.05 3.132 ;
      RECT 25.03 2.958 25.045 3.137 ;
      RECT 25.025 2.963 25.03 3.141 ;
      RECT 25.005 2.97 25.025 3.146 ;
      RECT 24.935 2.995 25.005 3.163 ;
      RECT 24.895 3.023 24.935 3.183 ;
      RECT 24.89 3.033 24.895 3.191 ;
      RECT 24.87 3.04 24.89 3.193 ;
      RECT 24.865 3.047 24.87 3.196 ;
      RECT 24.835 3.055 24.865 3.199 ;
      RECT 24.83 3.06 24.835 3.203 ;
      RECT 24.756 3.064 24.83 3.211 ;
      RECT 24.67 3.073 24.756 3.227 ;
      RECT 24.666 3.078 24.67 3.236 ;
      RECT 24.58 3.083 24.666 3.246 ;
      RECT 24.54 3.091 24.58 3.258 ;
      RECT 24.49 3.097 24.54 3.265 ;
      RECT 24.405 3.106 24.49 3.28 ;
      RECT 24.33 3.117 24.405 3.298 ;
      RECT 24.295 3.124 24.33 3.308 ;
      RECT 24.22 3.132 24.295 3.313 ;
      RECT 24.165 3.141 24.22 3.313 ;
      RECT 24.14 3.146 24.165 3.311 ;
      RECT 24.13 3.149 24.14 3.309 ;
      RECT 24.095 3.151 24.13 3.307 ;
      RECT 24.065 3.153 24.095 3.303 ;
      RECT 24.02 3.152 24.065 3.299 ;
      RECT 24 3.147 24.02 3.296 ;
      RECT 23.95 3.132 24 3.293 ;
      RECT 23.94 3.117 23.95 3.288 ;
      RECT 23.89 3.102 23.94 3.278 ;
      RECT 23.84 3.077 23.89 3.258 ;
      RECT 23.83 3.062 23.84 3.24 ;
      RECT 23.825 3.06 23.83 3.234 ;
      RECT 23.805 3.055 23.825 3.229 ;
      RECT 23.8 3.047 23.805 3.223 ;
      RECT 23.785 3.041 23.8 3.216 ;
      RECT 23.78 3.036 23.785 3.208 ;
      RECT 23.76 3.031 23.78 3.2 ;
      RECT 23.745 3.024 23.76 3.193 ;
      RECT 23.73 3.018 23.745 3.184 ;
      RECT 23.725 3.012 23.73 3.177 ;
      RECT 23.68 2.987 23.725 3.163 ;
      RECT 23.665 2.957 23.68 3.145 ;
      RECT 23.65 2.94 23.665 3.136 ;
      RECT 23.625 2.92 23.65 3.124 ;
      RECT 23.585 2.89 23.625 3.104 ;
      RECT 23.575 2.86 23.585 3.089 ;
      RECT 23.56 2.85 23.575 3.082 ;
      RECT 23.505 2.815 23.56 3.061 ;
      RECT 23.49 2.778 23.505 3.04 ;
      RECT 23.48 2.765 23.49 3.032 ;
      RECT 23.43 2.735 23.48 3.014 ;
      RECT 23.415 2.665 23.43 2.995 ;
      RECT 23.37 2.665 23.415 2.978 ;
      RECT 23.345 2.665 23.37 2.96 ;
      RECT 23.335 2.665 23.345 2.953 ;
      RECT 23.256 2.665 23.335 2.946 ;
      RECT 23.17 2.665 23.256 2.938 ;
      RECT 23.155 2.697 23.17 2.933 ;
      RECT 23.08 2.707 23.155 2.929 ;
      RECT 23.06 2.717 23.08 2.924 ;
      RECT 23.035 2.717 23.06 2.921 ;
      RECT 23.025 2.707 23.035 2.92 ;
      RECT 23.015 2.68 23.025 2.919 ;
      RECT 22.975 2.675 23.015 2.917 ;
      RECT 22.93 2.675 22.975 2.913 ;
      RECT 22.905 2.675 22.93 2.908 ;
      RECT 22.855 2.675 22.905 2.895 ;
      RECT 22.815 2.68 22.825 2.88 ;
      RECT 22.825 2.675 22.855 2.885 ;
      RECT 24.81 2.455 25.07 2.715 ;
      RECT 24.805 2.477 25.07 2.673 ;
      RECT 24.045 2.305 24.265 2.67 ;
      RECT 24.027 2.392 24.265 2.669 ;
      RECT 24.01 2.397 24.265 2.666 ;
      RECT 24.01 2.397 24.285 2.665 ;
      RECT 23.98 2.407 24.285 2.663 ;
      RECT 23.975 2.422 24.285 2.659 ;
      RECT 23.975 2.422 24.29 2.658 ;
      RECT 23.97 2.48 24.29 2.656 ;
      RECT 23.97 2.48 24.3 2.653 ;
      RECT 23.965 2.545 24.3 2.648 ;
      RECT 24.045 2.305 24.305 2.565 ;
      RECT 22.79 2.135 23.05 2.395 ;
      RECT 22.79 2.178 23.136 2.369 ;
      RECT 22.79 2.178 23.18 2.368 ;
      RECT 22.79 2.178 23.2 2.366 ;
      RECT 22.79 2.178 23.3 2.365 ;
      RECT 22.79 2.178 23.32 2.363 ;
      RECT 22.79 2.178 23.33 2.358 ;
      RECT 23.2 2.145 23.39 2.355 ;
      RECT 23.2 2.147 23.395 2.353 ;
      RECT 23.19 2.152 23.4 2.345 ;
      RECT 23.136 2.176 23.4 2.345 ;
      RECT 23.18 2.17 23.19 2.367 ;
      RECT 23.19 2.15 23.395 2.353 ;
      RECT 22.145 3.21 22.35 3.44 ;
      RECT 22.085 3.16 22.14 3.42 ;
      RECT 22.145 3.16 22.345 3.44 ;
      RECT 23.115 3.475 23.12 3.502 ;
      RECT 23.105 3.385 23.115 3.507 ;
      RECT 23.1 3.307 23.105 3.513 ;
      RECT 23.09 3.297 23.1 3.52 ;
      RECT 23.085 3.287 23.09 3.526 ;
      RECT 23.075 3.282 23.085 3.528 ;
      RECT 23.06 3.274 23.075 3.536 ;
      RECT 23.045 3.265 23.06 3.548 ;
      RECT 23.035 3.257 23.045 3.558 ;
      RECT 23 3.175 23.035 3.576 ;
      RECT 22.965 3.175 23 3.595 ;
      RECT 22.95 3.175 22.965 3.603 ;
      RECT 22.895 3.175 22.95 3.603 ;
      RECT 22.861 3.175 22.895 3.594 ;
      RECT 22.775 3.175 22.861 3.57 ;
      RECT 22.765 3.235 22.775 3.552 ;
      RECT 22.725 3.237 22.765 3.543 ;
      RECT 22.72 3.239 22.725 3.533 ;
      RECT 22.7 3.241 22.72 3.528 ;
      RECT 22.69 3.244 22.7 3.523 ;
      RECT 22.68 3.245 22.69 3.518 ;
      RECT 22.656 3.246 22.68 3.51 ;
      RECT 22.57 3.251 22.656 3.488 ;
      RECT 22.515 3.25 22.57 3.461 ;
      RECT 22.5 3.243 22.515 3.448 ;
      RECT 22.465 3.238 22.5 3.444 ;
      RECT 22.41 3.23 22.465 3.443 ;
      RECT 22.35 3.217 22.41 3.441 ;
      RECT 22.14 3.16 22.145 3.428 ;
      RECT 22.215 2.53 22.4 2.74 ;
      RECT 22.205 2.535 22.415 2.733 ;
      RECT 22.245 2.44 22.505 2.7 ;
      RECT 22.2 2.597 22.505 2.623 ;
      RECT 21.545 2.39 21.55 3.19 ;
      RECT 21.49 2.44 21.52 3.19 ;
      RECT 21.48 2.44 21.485 2.75 ;
      RECT 21.465 2.44 21.47 2.745 ;
      RECT 21.01 2.485 21.025 2.7 ;
      RECT 20.94 2.485 21.025 2.695 ;
      RECT 22.205 2.065 22.275 2.275 ;
      RECT 22.275 2.072 22.285 2.27 ;
      RECT 22.171 2.065 22.205 2.282 ;
      RECT 22.085 2.065 22.171 2.306 ;
      RECT 22.075 2.07 22.085 2.325 ;
      RECT 22.07 2.082 22.075 2.328 ;
      RECT 22.055 2.097 22.07 2.332 ;
      RECT 22.05 2.115 22.055 2.336 ;
      RECT 22.01 2.125 22.05 2.345 ;
      RECT 21.995 2.132 22.01 2.357 ;
      RECT 21.98 2.137 21.995 2.362 ;
      RECT 21.965 2.14 21.98 2.367 ;
      RECT 21.955 2.142 21.965 2.371 ;
      RECT 21.92 2.149 21.955 2.379 ;
      RECT 21.885 2.157 21.92 2.393 ;
      RECT 21.875 2.163 21.885 2.402 ;
      RECT 21.87 2.165 21.875 2.404 ;
      RECT 21.85 2.168 21.87 2.41 ;
      RECT 21.82 2.175 21.85 2.421 ;
      RECT 21.81 2.181 21.82 2.428 ;
      RECT 21.785 2.184 21.81 2.435 ;
      RECT 21.775 2.188 21.785 2.443 ;
      RECT 21.77 2.189 21.775 2.465 ;
      RECT 21.765 2.19 21.77 2.48 ;
      RECT 21.76 2.191 21.765 2.495 ;
      RECT 21.755 2.192 21.76 2.51 ;
      RECT 21.75 2.193 21.755 2.54 ;
      RECT 21.74 2.195 21.75 2.573 ;
      RECT 21.725 2.199 21.74 2.62 ;
      RECT 21.715 2.202 21.725 2.665 ;
      RECT 21.71 2.205 21.715 2.693 ;
      RECT 21.7 2.207 21.71 2.72 ;
      RECT 21.695 2.21 21.7 2.755 ;
      RECT 21.665 2.215 21.695 2.813 ;
      RECT 21.66 2.22 21.665 2.898 ;
      RECT 21.655 2.222 21.66 2.933 ;
      RECT 21.65 2.224 21.655 3.015 ;
      RECT 21.645 2.226 21.65 3.103 ;
      RECT 21.635 2.228 21.645 3.185 ;
      RECT 21.62 2.242 21.635 3.19 ;
      RECT 21.585 2.287 21.62 3.19 ;
      RECT 21.575 2.327 21.585 3.19 ;
      RECT 21.56 2.355 21.575 3.19 ;
      RECT 21.555 2.372 21.56 3.19 ;
      RECT 21.55 2.38 21.555 3.19 ;
      RECT 21.54 2.395 21.545 3.19 ;
      RECT 21.535 2.402 21.54 3.19 ;
      RECT 21.525 2.422 21.535 3.19 ;
      RECT 21.52 2.435 21.525 3.19 ;
      RECT 21.485 2.44 21.49 2.775 ;
      RECT 21.47 2.83 21.49 3.19 ;
      RECT 21.47 2.44 21.48 2.748 ;
      RECT 21.465 2.87 21.47 3.19 ;
      RECT 21.415 2.44 21.465 2.743 ;
      RECT 21.46 2.907 21.465 3.19 ;
      RECT 21.45 2.93 21.46 3.19 ;
      RECT 21.445 2.975 21.45 3.19 ;
      RECT 21.435 2.985 21.445 3.183 ;
      RECT 21.361 2.44 21.415 2.737 ;
      RECT 21.275 2.44 21.361 2.73 ;
      RECT 21.226 2.487 21.275 2.723 ;
      RECT 21.14 2.495 21.226 2.716 ;
      RECT 21.125 2.492 21.14 2.711 ;
      RECT 21.111 2.485 21.125 2.71 ;
      RECT 21.025 2.485 21.111 2.705 ;
      RECT 20.93 2.49 20.94 2.69 ;
      RECT 20.52 1.92 20.535 2.32 ;
      RECT 20.715 1.92 20.72 2.18 ;
      RECT 20.46 1.92 20.505 2.18 ;
      RECT 20.915 3.225 20.92 3.43 ;
      RECT 20.91 3.215 20.915 3.435 ;
      RECT 20.905 3.202 20.91 3.44 ;
      RECT 20.9 3.182 20.905 3.44 ;
      RECT 20.875 3.135 20.9 3.44 ;
      RECT 20.84 3.05 20.875 3.44 ;
      RECT 20.835 2.987 20.84 3.44 ;
      RECT 20.83 2.972 20.835 3.44 ;
      RECT 20.815 2.932 20.83 3.44 ;
      RECT 20.81 2.907 20.815 3.44 ;
      RECT 20.8 2.89 20.81 3.44 ;
      RECT 20.765 2.812 20.8 3.44 ;
      RECT 20.76 2.755 20.765 3.44 ;
      RECT 20.755 2.742 20.76 3.44 ;
      RECT 20.745 2.72 20.755 3.44 ;
      RECT 20.735 2.685 20.745 3.44 ;
      RECT 20.725 2.655 20.735 3.44 ;
      RECT 20.715 2.57 20.725 3.083 ;
      RECT 20.722 3.215 20.725 3.44 ;
      RECT 20.72 3.225 20.722 3.44 ;
      RECT 20.71 3.235 20.72 3.435 ;
      RECT 20.705 1.92 20.715 2.315 ;
      RECT 20.71 2.447 20.715 3.058 ;
      RECT 20.705 2.345 20.71 3.041 ;
      RECT 20.695 1.92 20.705 3.017 ;
      RECT 20.69 1.92 20.695 2.988 ;
      RECT 20.685 1.92 20.69 2.978 ;
      RECT 20.665 1.92 20.685 2.94 ;
      RECT 20.66 1.92 20.665 2.898 ;
      RECT 20.655 1.92 20.66 2.878 ;
      RECT 20.625 1.92 20.655 2.828 ;
      RECT 20.615 1.92 20.625 2.775 ;
      RECT 20.61 1.92 20.615 2.748 ;
      RECT 20.605 1.92 20.61 2.733 ;
      RECT 20.595 1.92 20.605 2.71 ;
      RECT 20.585 1.92 20.595 2.685 ;
      RECT 20.58 1.92 20.585 2.625 ;
      RECT 20.57 1.92 20.58 2.563 ;
      RECT 20.565 1.92 20.57 2.483 ;
      RECT 20.56 1.92 20.565 2.448 ;
      RECT 20.555 1.92 20.56 2.423 ;
      RECT 20.55 1.92 20.555 2.408 ;
      RECT 20.545 1.92 20.55 2.378 ;
      RECT 20.54 1.92 20.545 2.355 ;
      RECT 20.535 1.92 20.54 2.328 ;
      RECT 20.505 1.92 20.52 2.315 ;
      RECT 19.66 3.455 19.845 3.665 ;
      RECT 19.65 3.46 19.86 3.658 ;
      RECT 19.65 3.46 19.88 3.63 ;
      RECT 19.65 3.46 19.895 3.609 ;
      RECT 19.65 3.46 19.91 3.607 ;
      RECT 19.65 3.46 19.92 3.606 ;
      RECT 19.65 3.46 19.95 3.603 ;
      RECT 20.3 3.305 20.56 3.565 ;
      RECT 20.26 3.352 20.56 3.548 ;
      RECT 20.251 3.36 20.26 3.551 ;
      RECT 19.845 3.453 20.56 3.548 ;
      RECT 20.165 3.378 20.251 3.558 ;
      RECT 19.86 3.45 20.56 3.548 ;
      RECT 20.106 3.4 20.165 3.57 ;
      RECT 19.88 3.446 20.56 3.548 ;
      RECT 20.02 3.412 20.106 3.581 ;
      RECT 19.895 3.442 20.56 3.548 ;
      RECT 19.965 3.425 20.02 3.593 ;
      RECT 19.91 3.44 20.56 3.548 ;
      RECT 19.95 3.431 19.965 3.599 ;
      RECT 19.92 3.436 20.56 3.548 ;
      RECT 20.065 2.96 20.325 3.22 ;
      RECT 20.065 2.98 20.435 3.19 ;
      RECT 20.065 2.985 20.445 3.185 ;
      RECT 20.256 2.399 20.335 2.63 ;
      RECT 20.17 2.402 20.385 2.625 ;
      RECT 20.165 2.402 20.385 2.62 ;
      RECT 20.165 2.407 20.395 2.618 ;
      RECT 20.14 2.407 20.395 2.615 ;
      RECT 20.14 2.415 20.405 2.613 ;
      RECT 20.02 2.35 20.28 2.61 ;
      RECT 20.02 2.397 20.33 2.61 ;
      RECT 19.275 2.97 19.28 3.23 ;
      RECT 19.105 2.74 19.11 3.23 ;
      RECT 18.99 2.98 18.995 3.205 ;
      RECT 19.7 2.075 19.705 2.285 ;
      RECT 19.705 2.08 19.72 2.28 ;
      RECT 19.64 2.075 19.7 2.293 ;
      RECT 19.625 2.075 19.64 2.303 ;
      RECT 19.575 2.075 19.625 2.32 ;
      RECT 19.555 2.075 19.575 2.343 ;
      RECT 19.54 2.075 19.555 2.355 ;
      RECT 19.52 2.075 19.54 2.365 ;
      RECT 19.51 2.08 19.52 2.374 ;
      RECT 19.505 2.09 19.51 2.379 ;
      RECT 19.5 2.102 19.505 2.383 ;
      RECT 19.49 2.125 19.5 2.388 ;
      RECT 19.485 2.14 19.49 2.392 ;
      RECT 19.48 2.157 19.485 2.395 ;
      RECT 19.475 2.165 19.48 2.398 ;
      RECT 19.465 2.17 19.475 2.402 ;
      RECT 19.46 2.177 19.465 2.407 ;
      RECT 19.45 2.182 19.46 2.411 ;
      RECT 19.425 2.194 19.45 2.422 ;
      RECT 19.405 2.211 19.425 2.438 ;
      RECT 19.38 2.228 19.405 2.46 ;
      RECT 19.345 2.251 19.38 2.518 ;
      RECT 19.325 2.273 19.345 2.58 ;
      RECT 19.32 2.283 19.325 2.615 ;
      RECT 19.31 2.29 19.32 2.653 ;
      RECT 19.305 2.297 19.31 2.673 ;
      RECT 19.3 2.308 19.305 2.71 ;
      RECT 19.295 2.316 19.3 2.775 ;
      RECT 19.285 2.327 19.295 2.828 ;
      RECT 19.28 2.345 19.285 2.898 ;
      RECT 19.275 2.355 19.28 2.935 ;
      RECT 19.27 2.365 19.275 3.23 ;
      RECT 19.265 2.377 19.27 3.23 ;
      RECT 19.26 2.387 19.265 3.23 ;
      RECT 19.25 2.397 19.26 3.23 ;
      RECT 19.24 2.42 19.25 3.23 ;
      RECT 19.225 2.455 19.24 3.23 ;
      RECT 19.185 2.517 19.225 3.23 ;
      RECT 19.18 2.57 19.185 3.23 ;
      RECT 19.155 2.605 19.18 3.23 ;
      RECT 19.14 2.65 19.155 3.23 ;
      RECT 19.135 2.672 19.14 3.23 ;
      RECT 19.125 2.685 19.135 3.23 ;
      RECT 19.115 2.71 19.125 3.23 ;
      RECT 19.11 2.732 19.115 3.23 ;
      RECT 19.085 2.77 19.105 3.23 ;
      RECT 19.045 2.827 19.085 3.23 ;
      RECT 19.04 2.877 19.045 3.23 ;
      RECT 19.035 2.895 19.04 3.23 ;
      RECT 19.03 2.907 19.035 3.23 ;
      RECT 19.02 2.925 19.03 3.23 ;
      RECT 19.01 2.945 19.02 3.205 ;
      RECT 19.005 2.962 19.01 3.205 ;
      RECT 18.995 2.975 19.005 3.205 ;
      RECT 18.965 2.985 18.99 3.205 ;
      RECT 18.955 2.992 18.965 3.205 ;
      RECT 18.94 3.002 18.955 3.2 ;
      RECT 18.035 7.77 18.325 8 ;
      RECT 18.095 6.29 18.265 8 ;
      RECT 18.09 6.655 18.44 7.005 ;
      RECT 18.035 6.29 18.325 6.52 ;
      RECT 17.63 2.395 17.735 2.965 ;
      RECT 17.63 2.73 17.955 2.96 ;
      RECT 17.63 2.76 18.125 2.93 ;
      RECT 17.63 2.395 17.82 2.96 ;
      RECT 17.045 2.36 17.335 2.59 ;
      RECT 17.045 2.395 17.82 2.565 ;
      RECT 17.105 0.88 17.275 2.59 ;
      RECT 17.045 0.88 17.335 1.11 ;
      RECT 17.045 7.77 17.335 8 ;
      RECT 17.105 6.29 17.275 8 ;
      RECT 17.045 6.29 17.335 6.52 ;
      RECT 17.045 6.325 17.9 6.485 ;
      RECT 17.73 5.92 17.9 6.485 ;
      RECT 17.045 6.32 17.44 6.485 ;
      RECT 17.665 5.92 17.955 6.15 ;
      RECT 17.665 5.95 18.125 6.12 ;
      RECT 16.675 2.73 16.965 2.96 ;
      RECT 16.675 2.76 17.135 2.93 ;
      RECT 16.74 1.655 16.905 2.96 ;
      RECT 15.255 1.625 15.545 1.855 ;
      RECT 15.255 1.655 16.905 1.825 ;
      RECT 15.315 0.885 15.485 1.855 ;
      RECT 15.255 0.885 15.545 1.115 ;
      RECT 15.255 7.765 15.545 7.995 ;
      RECT 15.315 7.025 15.485 7.995 ;
      RECT 15.315 7.12 16.905 7.29 ;
      RECT 16.735 5.92 16.905 7.29 ;
      RECT 15.255 7.025 15.545 7.255 ;
      RECT 16.675 5.92 16.965 6.15 ;
      RECT 16.675 5.95 17.135 6.12 ;
      RECT 15.685 1.965 16.035 2.315 ;
      RECT 13.35 2.025 16.035 2.195 ;
      RECT 13.35 1.34 13.52 2.195 ;
      RECT 13.25 1.34 13.6 1.69 ;
      RECT 15.71 6.655 16.035 6.98 ;
      RECT 11.105 6.605 11.455 6.955 ;
      RECT 15.685 6.655 16.035 6.885 ;
      RECT 10.905 6.655 11.455 6.885 ;
      RECT 10.735 6.685 16.035 6.855 ;
      RECT 14.91 2.365 15.23 2.685 ;
      RECT 14.88 2.365 15.23 2.595 ;
      RECT 14.71 2.395 15.23 2.565 ;
      RECT 14.91 6.255 15.23 6.545 ;
      RECT 14.88 6.285 15.23 6.515 ;
      RECT 14.71 6.315 15.23 6.485 ;
      RECT 11.545 2.465 11.73 2.675 ;
      RECT 11.535 2.47 11.745 2.668 ;
      RECT 11.535 2.47 11.831 2.645 ;
      RECT 11.535 2.47 11.89 2.62 ;
      RECT 11.535 2.47 11.945 2.6 ;
      RECT 11.535 2.47 11.955 2.588 ;
      RECT 11.535 2.47 12.15 2.527 ;
      RECT 11.535 2.47 12.18 2.51 ;
      RECT 11.535 2.47 12.2 2.5 ;
      RECT 12.08 2.235 12.34 2.495 ;
      RECT 12.065 2.325 12.08 2.542 ;
      RECT 11.6 2.457 12.34 2.495 ;
      RECT 12.051 2.336 12.065 2.548 ;
      RECT 11.64 2.45 12.34 2.495 ;
      RECT 11.965 2.376 12.051 2.567 ;
      RECT 11.89 2.437 12.34 2.495 ;
      RECT 11.96 2.412 11.965 2.584 ;
      RECT 11.945 2.422 12.34 2.495 ;
      RECT 11.955 2.417 11.96 2.586 ;
      RECT 12.25 2.922 12.255 3.014 ;
      RECT 12.245 2.9 12.25 3.031 ;
      RECT 12.24 2.89 12.245 3.043 ;
      RECT 12.23 2.881 12.24 3.053 ;
      RECT 12.225 2.876 12.23 3.061 ;
      RECT 12.22 2.735 12.225 3.064 ;
      RECT 12.186 2.735 12.22 3.075 ;
      RECT 12.1 2.735 12.186 3.11 ;
      RECT 12.02 2.735 12.1 3.158 ;
      RECT 11.991 2.735 12.02 3.182 ;
      RECT 11.905 2.735 11.991 3.188 ;
      RECT 11.9 2.919 11.905 3.193 ;
      RECT 11.865 2.93 11.9 3.196 ;
      RECT 11.84 2.945 11.865 3.2 ;
      RECT 11.826 2.954 11.84 3.202 ;
      RECT 11.74 2.981 11.826 3.208 ;
      RECT 11.675 3.022 11.74 3.217 ;
      RECT 11.66 3.042 11.675 3.222 ;
      RECT 11.63 3.052 11.66 3.225 ;
      RECT 11.625 3.062 11.63 3.228 ;
      RECT 11.595 3.067 11.625 3.23 ;
      RECT 11.575 3.072 11.595 3.234 ;
      RECT 11.49 3.075 11.575 3.241 ;
      RECT 11.475 3.072 11.49 3.247 ;
      RECT 11.465 3.069 11.475 3.249 ;
      RECT 11.445 3.066 11.465 3.251 ;
      RECT 11.425 3.062 11.445 3.252 ;
      RECT 11.41 3.058 11.425 3.254 ;
      RECT 11.4 3.055 11.41 3.255 ;
      RECT 11.36 3.049 11.4 3.253 ;
      RECT 11.35 3.044 11.36 3.251 ;
      RECT 11.335 3.041 11.35 3.247 ;
      RECT 11.31 3.036 11.335 3.24 ;
      RECT 11.26 3.027 11.31 3.228 ;
      RECT 11.19 3.013 11.26 3.21 ;
      RECT 11.132 2.998 11.19 3.192 ;
      RECT 11.046 2.981 11.132 3.172 ;
      RECT 10.96 2.96 11.046 3.147 ;
      RECT 10.91 2.945 10.96 3.128 ;
      RECT 10.906 2.939 10.91 3.12 ;
      RECT 10.82 2.929 10.906 3.107 ;
      RECT 10.785 2.914 10.82 3.09 ;
      RECT 10.77 2.907 10.785 3.083 ;
      RECT 10.71 2.895 10.77 3.071 ;
      RECT 10.69 2.882 10.71 3.059 ;
      RECT 10.65 2.873 10.69 3.051 ;
      RECT 10.645 2.865 10.65 3.044 ;
      RECT 10.565 2.855 10.645 3.03 ;
      RECT 10.55 2.842 10.565 3.015 ;
      RECT 10.545 2.84 10.55 3.013 ;
      RECT 10.466 2.828 10.545 3 ;
      RECT 10.38 2.803 10.466 2.975 ;
      RECT 10.365 2.772 10.38 2.96 ;
      RECT 10.35 2.747 10.365 2.956 ;
      RECT 10.335 2.74 10.35 2.952 ;
      RECT 10.16 2.745 10.165 2.948 ;
      RECT 10.155 2.75 10.16 2.943 ;
      RECT 10.165 2.74 10.335 2.95 ;
      RECT 10.88 2.5 10.985 2.76 ;
      RECT 11.695 2.025 11.7 2.25 ;
      RECT 11.825 2.025 11.88 2.235 ;
      RECT 11.88 2.03 11.89 2.228 ;
      RECT 11.786 2.025 11.825 2.238 ;
      RECT 11.7 2.025 11.786 2.245 ;
      RECT 11.68 2.03 11.695 2.251 ;
      RECT 11.67 2.07 11.68 2.253 ;
      RECT 11.64 2.08 11.67 2.255 ;
      RECT 11.635 2.085 11.64 2.257 ;
      RECT 11.61 2.09 11.635 2.259 ;
      RECT 11.595 2.095 11.61 2.261 ;
      RECT 11.58 2.097 11.595 2.263 ;
      RECT 11.575 2.102 11.58 2.265 ;
      RECT 11.525 2.11 11.575 2.268 ;
      RECT 11.5 2.119 11.525 2.273 ;
      RECT 11.49 2.126 11.5 2.278 ;
      RECT 11.485 2.129 11.49 2.282 ;
      RECT 11.465 2.132 11.485 2.291 ;
      RECT 11.435 2.14 11.465 2.311 ;
      RECT 11.406 2.153 11.435 2.333 ;
      RECT 11.32 2.187 11.406 2.377 ;
      RECT 11.315 2.213 11.32 2.415 ;
      RECT 11.31 2.217 11.315 2.424 ;
      RECT 11.275 2.23 11.31 2.457 ;
      RECT 11.265 2.244 11.275 2.495 ;
      RECT 11.26 2.248 11.265 2.508 ;
      RECT 11.255 2.252 11.26 2.513 ;
      RECT 11.245 2.26 11.255 2.525 ;
      RECT 11.24 2.267 11.245 2.54 ;
      RECT 11.215 2.28 11.24 2.565 ;
      RECT 11.175 2.309 11.215 2.62 ;
      RECT 11.16 2.334 11.175 2.675 ;
      RECT 11.15 2.345 11.16 2.698 ;
      RECT 11.145 2.352 11.15 2.71 ;
      RECT 11.14 2.356 11.145 2.718 ;
      RECT 11.085 2.384 11.14 2.76 ;
      RECT 11.065 2.42 11.085 2.76 ;
      RECT 11.05 2.435 11.065 2.76 ;
      RECT 10.995 2.467 11.05 2.76 ;
      RECT 10.985 2.497 10.995 2.76 ;
      RECT 10.595 2.112 10.78 2.35 ;
      RECT 10.58 2.114 10.79 2.345 ;
      RECT 10.465 2.06 10.725 2.32 ;
      RECT 10.46 2.097 10.725 2.274 ;
      RECT 10.455 2.107 10.725 2.271 ;
      RECT 10.45 2.147 10.79 2.265 ;
      RECT 10.445 2.18 10.79 2.255 ;
      RECT 10.455 2.122 10.805 2.193 ;
      RECT 10.752 3.22 10.765 3.75 ;
      RECT 10.666 3.22 10.765 3.749 ;
      RECT 10.666 3.22 10.77 3.748 ;
      RECT 10.58 3.22 10.77 3.746 ;
      RECT 10.575 3.22 10.77 3.743 ;
      RECT 10.575 3.22 10.78 3.741 ;
      RECT 10.57 3.512 10.78 3.738 ;
      RECT 10.57 3.522 10.785 3.735 ;
      RECT 10.57 3.59 10.79 3.731 ;
      RECT 10.56 3.595 10.79 3.73 ;
      RECT 10.56 3.687 10.795 3.727 ;
      RECT 10.545 3.22 10.805 3.48 ;
      RECT 10.475 7.765 10.765 7.995 ;
      RECT 10.535 7.025 10.705 7.995 ;
      RECT 10.45 7.055 10.79 7.4 ;
      RECT 10.475 7.025 10.765 7.4 ;
      RECT 9.775 2.21 9.82 3.745 ;
      RECT 9.975 2.21 10.005 2.425 ;
      RECT 8.35 1.95 8.47 2.16 ;
      RECT 8.01 1.9 8.27 2.16 ;
      RECT 8.01 1.945 8.305 2.15 ;
      RECT 10.015 2.226 10.02 2.28 ;
      RECT 10.01 2.219 10.015 2.413 ;
      RECT 10.005 2.213 10.01 2.42 ;
      RECT 9.96 2.21 9.975 2.433 ;
      RECT 9.955 2.21 9.96 2.455 ;
      RECT 9.95 2.21 9.955 2.503 ;
      RECT 9.945 2.21 9.95 2.523 ;
      RECT 9.935 2.21 9.945 2.63 ;
      RECT 9.93 2.21 9.935 2.693 ;
      RECT 9.925 2.21 9.93 2.75 ;
      RECT 9.92 2.21 9.925 2.758 ;
      RECT 9.905 2.21 9.92 2.865 ;
      RECT 9.895 2.21 9.905 3 ;
      RECT 9.885 2.21 9.895 3.11 ;
      RECT 9.875 2.21 9.885 3.167 ;
      RECT 9.87 2.21 9.875 3.207 ;
      RECT 9.865 2.21 9.87 3.243 ;
      RECT 9.855 2.21 9.865 3.283 ;
      RECT 9.85 2.21 9.855 3.325 ;
      RECT 9.83 2.21 9.85 3.39 ;
      RECT 9.835 3.535 9.84 3.715 ;
      RECT 9.83 3.517 9.835 3.723 ;
      RECT 9.825 2.21 9.83 3.453 ;
      RECT 9.825 3.497 9.83 3.73 ;
      RECT 9.82 2.21 9.825 3.74 ;
      RECT 9.765 2.21 9.775 2.51 ;
      RECT 9.77 2.757 9.775 3.745 ;
      RECT 9.765 2.822 9.77 3.745 ;
      RECT 9.76 2.211 9.765 2.5 ;
      RECT 9.755 2.887 9.765 3.745 ;
      RECT 9.75 2.212 9.76 2.49 ;
      RECT 9.74 3 9.755 3.745 ;
      RECT 9.745 2.213 9.75 2.48 ;
      RECT 9.725 2.214 9.745 2.458 ;
      RECT 9.73 3.097 9.74 3.745 ;
      RECT 9.725 3.172 9.73 3.745 ;
      RECT 9.715 2.213 9.725 2.435 ;
      RECT 9.72 3.215 9.725 3.745 ;
      RECT 9.715 3.242 9.72 3.745 ;
      RECT 9.705 2.211 9.715 2.423 ;
      RECT 9.71 3.285 9.715 3.745 ;
      RECT 9.705 3.312 9.71 3.745 ;
      RECT 9.695 2.21 9.705 2.41 ;
      RECT 9.7 3.327 9.705 3.745 ;
      RECT 9.66 3.385 9.7 3.745 ;
      RECT 9.69 2.209 9.695 2.395 ;
      RECT 9.685 2.207 9.69 2.388 ;
      RECT 9.675 2.204 9.685 2.378 ;
      RECT 9.67 2.201 9.675 2.363 ;
      RECT 9.655 2.197 9.67 2.356 ;
      RECT 9.65 3.44 9.66 3.745 ;
      RECT 9.65 2.194 9.655 2.351 ;
      RECT 9.635 2.19 9.65 2.345 ;
      RECT 9.645 3.457 9.65 3.745 ;
      RECT 9.635 3.52 9.645 3.745 ;
      RECT 9.555 2.175 9.635 2.325 ;
      RECT 9.63 3.527 9.635 3.74 ;
      RECT 9.625 3.535 9.63 3.73 ;
      RECT 9.545 2.161 9.555 2.309 ;
      RECT 9.53 2.157 9.545 2.307 ;
      RECT 9.52 2.152 9.53 2.303 ;
      RECT 9.495 2.145 9.52 2.295 ;
      RECT 9.49 2.14 9.495 2.29 ;
      RECT 9.48 2.14 9.49 2.288 ;
      RECT 9.47 2.138 9.48 2.286 ;
      RECT 9.44 2.13 9.47 2.28 ;
      RECT 9.425 2.122 9.44 2.273 ;
      RECT 9.405 2.117 9.425 2.266 ;
      RECT 9.4 2.113 9.405 2.261 ;
      RECT 9.37 2.106 9.4 2.255 ;
      RECT 9.345 2.097 9.37 2.245 ;
      RECT 9.315 2.09 9.345 2.237 ;
      RECT 9.29 2.08 9.315 2.228 ;
      RECT 9.275 2.072 9.29 2.222 ;
      RECT 9.25 2.067 9.275 2.217 ;
      RECT 9.24 2.063 9.25 2.212 ;
      RECT 9.22 2.058 9.24 2.207 ;
      RECT 9.185 2.053 9.22 2.2 ;
      RECT 9.125 2.048 9.185 2.193 ;
      RECT 9.112 2.044 9.125 2.191 ;
      RECT 9.026 2.039 9.112 2.188 ;
      RECT 8.94 2.029 9.026 2.184 ;
      RECT 8.899 2.022 8.94 2.181 ;
      RECT 8.813 2.015 8.899 2.178 ;
      RECT 8.727 2.005 8.813 2.174 ;
      RECT 8.641 1.995 8.727 2.169 ;
      RECT 8.555 1.985 8.641 2.165 ;
      RECT 8.545 1.97 8.555 2.163 ;
      RECT 8.535 1.955 8.545 2.163 ;
      RECT 8.47 1.95 8.535 2.162 ;
      RECT 8.305 1.947 8.35 2.155 ;
      RECT 9.55 2.852 9.555 3.043 ;
      RECT 9.545 2.847 9.55 3.05 ;
      RECT 9.531 2.845 9.545 3.056 ;
      RECT 9.445 2.845 9.531 3.058 ;
      RECT 9.441 2.845 9.445 3.061 ;
      RECT 9.355 2.845 9.441 3.079 ;
      RECT 9.345 2.85 9.355 3.098 ;
      RECT 9.335 2.905 9.345 3.102 ;
      RECT 9.31 2.92 9.335 3.109 ;
      RECT 9.27 2.94 9.31 3.122 ;
      RECT 9.265 2.952 9.27 3.132 ;
      RECT 9.25 2.958 9.265 3.137 ;
      RECT 9.245 2.963 9.25 3.141 ;
      RECT 9.225 2.97 9.245 3.146 ;
      RECT 9.155 2.995 9.225 3.163 ;
      RECT 9.115 3.023 9.155 3.183 ;
      RECT 9.11 3.033 9.115 3.191 ;
      RECT 9.09 3.04 9.11 3.193 ;
      RECT 9.085 3.047 9.09 3.196 ;
      RECT 9.055 3.055 9.085 3.199 ;
      RECT 9.05 3.06 9.055 3.203 ;
      RECT 8.976 3.064 9.05 3.211 ;
      RECT 8.89 3.073 8.976 3.227 ;
      RECT 8.886 3.078 8.89 3.236 ;
      RECT 8.8 3.083 8.886 3.246 ;
      RECT 8.76 3.091 8.8 3.258 ;
      RECT 8.71 3.097 8.76 3.265 ;
      RECT 8.625 3.106 8.71 3.28 ;
      RECT 8.55 3.117 8.625 3.298 ;
      RECT 8.515 3.124 8.55 3.308 ;
      RECT 8.44 3.132 8.515 3.313 ;
      RECT 8.385 3.141 8.44 3.313 ;
      RECT 8.36 3.146 8.385 3.311 ;
      RECT 8.35 3.149 8.36 3.309 ;
      RECT 8.315 3.151 8.35 3.307 ;
      RECT 8.285 3.153 8.315 3.303 ;
      RECT 8.24 3.152 8.285 3.299 ;
      RECT 8.22 3.147 8.24 3.296 ;
      RECT 8.17 3.132 8.22 3.293 ;
      RECT 8.16 3.117 8.17 3.288 ;
      RECT 8.11 3.102 8.16 3.278 ;
      RECT 8.06 3.077 8.11 3.258 ;
      RECT 8.05 3.062 8.06 3.24 ;
      RECT 8.045 3.06 8.05 3.234 ;
      RECT 8.025 3.055 8.045 3.229 ;
      RECT 8.02 3.047 8.025 3.223 ;
      RECT 8.005 3.041 8.02 3.216 ;
      RECT 8 3.036 8.005 3.208 ;
      RECT 7.98 3.031 8 3.2 ;
      RECT 7.965 3.024 7.98 3.193 ;
      RECT 7.95 3.018 7.965 3.184 ;
      RECT 7.945 3.012 7.95 3.177 ;
      RECT 7.9 2.987 7.945 3.163 ;
      RECT 7.885 2.957 7.9 3.145 ;
      RECT 7.87 2.94 7.885 3.136 ;
      RECT 7.845 2.92 7.87 3.124 ;
      RECT 7.805 2.89 7.845 3.104 ;
      RECT 7.795 2.86 7.805 3.089 ;
      RECT 7.78 2.85 7.795 3.082 ;
      RECT 7.725 2.815 7.78 3.061 ;
      RECT 7.71 2.778 7.725 3.04 ;
      RECT 7.7 2.765 7.71 3.032 ;
      RECT 7.65 2.735 7.7 3.014 ;
      RECT 7.635 2.665 7.65 2.995 ;
      RECT 7.59 2.665 7.635 2.978 ;
      RECT 7.565 2.665 7.59 2.96 ;
      RECT 7.555 2.665 7.565 2.953 ;
      RECT 7.476 2.665 7.555 2.946 ;
      RECT 7.39 2.665 7.476 2.938 ;
      RECT 7.375 2.697 7.39 2.933 ;
      RECT 7.3 2.707 7.375 2.929 ;
      RECT 7.28 2.717 7.3 2.924 ;
      RECT 7.255 2.717 7.28 2.921 ;
      RECT 7.245 2.707 7.255 2.92 ;
      RECT 7.235 2.68 7.245 2.919 ;
      RECT 7.195 2.675 7.235 2.917 ;
      RECT 7.15 2.675 7.195 2.913 ;
      RECT 7.125 2.675 7.15 2.908 ;
      RECT 7.075 2.675 7.125 2.895 ;
      RECT 7.035 2.68 7.045 2.88 ;
      RECT 7.045 2.675 7.075 2.885 ;
      RECT 9.03 2.455 9.29 2.715 ;
      RECT 9.025 2.477 9.29 2.673 ;
      RECT 8.265 2.305 8.485 2.67 ;
      RECT 8.247 2.392 8.485 2.669 ;
      RECT 8.23 2.397 8.485 2.666 ;
      RECT 8.23 2.397 8.505 2.665 ;
      RECT 8.2 2.407 8.505 2.663 ;
      RECT 8.195 2.422 8.505 2.659 ;
      RECT 8.195 2.422 8.51 2.658 ;
      RECT 8.19 2.48 8.51 2.656 ;
      RECT 8.19 2.48 8.52 2.653 ;
      RECT 8.185 2.545 8.52 2.648 ;
      RECT 8.265 2.305 8.525 2.565 ;
      RECT 7.01 2.135 7.27 2.395 ;
      RECT 7.01 2.178 7.356 2.369 ;
      RECT 7.01 2.178 7.4 2.368 ;
      RECT 7.01 2.178 7.42 2.366 ;
      RECT 7.01 2.178 7.52 2.365 ;
      RECT 7.01 2.178 7.54 2.363 ;
      RECT 7.01 2.178 7.55 2.358 ;
      RECT 7.42 2.145 7.61 2.355 ;
      RECT 7.42 2.147 7.615 2.353 ;
      RECT 7.41 2.152 7.62 2.345 ;
      RECT 7.356 2.176 7.62 2.345 ;
      RECT 7.4 2.17 7.41 2.367 ;
      RECT 7.41 2.15 7.615 2.353 ;
      RECT 6.365 3.21 6.57 3.44 ;
      RECT 6.305 3.16 6.36 3.42 ;
      RECT 6.365 3.16 6.565 3.44 ;
      RECT 7.335 3.475 7.34 3.502 ;
      RECT 7.325 3.385 7.335 3.507 ;
      RECT 7.32 3.307 7.325 3.513 ;
      RECT 7.31 3.297 7.32 3.52 ;
      RECT 7.305 3.287 7.31 3.526 ;
      RECT 7.295 3.282 7.305 3.528 ;
      RECT 7.28 3.274 7.295 3.536 ;
      RECT 7.265 3.265 7.28 3.548 ;
      RECT 7.255 3.257 7.265 3.558 ;
      RECT 7.22 3.175 7.255 3.576 ;
      RECT 7.185 3.175 7.22 3.595 ;
      RECT 7.17 3.175 7.185 3.603 ;
      RECT 7.115 3.175 7.17 3.603 ;
      RECT 7.081 3.175 7.115 3.594 ;
      RECT 6.995 3.175 7.081 3.57 ;
      RECT 6.985 3.235 6.995 3.552 ;
      RECT 6.945 3.237 6.985 3.543 ;
      RECT 6.94 3.239 6.945 3.533 ;
      RECT 6.92 3.241 6.94 3.528 ;
      RECT 6.91 3.244 6.92 3.523 ;
      RECT 6.9 3.245 6.91 3.518 ;
      RECT 6.876 3.246 6.9 3.51 ;
      RECT 6.79 3.251 6.876 3.488 ;
      RECT 6.735 3.25 6.79 3.461 ;
      RECT 6.72 3.243 6.735 3.448 ;
      RECT 6.685 3.238 6.72 3.444 ;
      RECT 6.63 3.23 6.685 3.443 ;
      RECT 6.57 3.217 6.63 3.441 ;
      RECT 6.36 3.16 6.365 3.428 ;
      RECT 6.435 2.53 6.62 2.74 ;
      RECT 6.425 2.535 6.635 2.733 ;
      RECT 6.465 2.44 6.725 2.7 ;
      RECT 6.42 2.597 6.725 2.623 ;
      RECT 5.765 2.39 5.77 3.19 ;
      RECT 5.71 2.44 5.74 3.19 ;
      RECT 5.7 2.44 5.705 2.75 ;
      RECT 5.685 2.44 5.69 2.745 ;
      RECT 5.23 2.485 5.245 2.7 ;
      RECT 5.16 2.485 5.245 2.695 ;
      RECT 6.425 2.065 6.495 2.275 ;
      RECT 6.495 2.072 6.505 2.27 ;
      RECT 6.391 2.065 6.425 2.282 ;
      RECT 6.305 2.065 6.391 2.306 ;
      RECT 6.295 2.07 6.305 2.325 ;
      RECT 6.29 2.082 6.295 2.328 ;
      RECT 6.275 2.097 6.29 2.332 ;
      RECT 6.27 2.115 6.275 2.336 ;
      RECT 6.23 2.125 6.27 2.345 ;
      RECT 6.215 2.132 6.23 2.357 ;
      RECT 6.2 2.137 6.215 2.362 ;
      RECT 6.185 2.14 6.2 2.367 ;
      RECT 6.175 2.142 6.185 2.371 ;
      RECT 6.14 2.149 6.175 2.379 ;
      RECT 6.105 2.157 6.14 2.393 ;
      RECT 6.095 2.163 6.105 2.402 ;
      RECT 6.09 2.165 6.095 2.404 ;
      RECT 6.07 2.168 6.09 2.41 ;
      RECT 6.04 2.175 6.07 2.421 ;
      RECT 6.03 2.181 6.04 2.428 ;
      RECT 6.005 2.184 6.03 2.435 ;
      RECT 5.995 2.188 6.005 2.443 ;
      RECT 5.99 2.189 5.995 2.465 ;
      RECT 5.985 2.19 5.99 2.48 ;
      RECT 5.98 2.191 5.985 2.495 ;
      RECT 5.975 2.192 5.98 2.51 ;
      RECT 5.97 2.193 5.975 2.54 ;
      RECT 5.96 2.195 5.97 2.573 ;
      RECT 5.945 2.199 5.96 2.62 ;
      RECT 5.935 2.202 5.945 2.665 ;
      RECT 5.93 2.205 5.935 2.693 ;
      RECT 5.92 2.207 5.93 2.72 ;
      RECT 5.915 2.21 5.92 2.755 ;
      RECT 5.885 2.215 5.915 2.813 ;
      RECT 5.88 2.22 5.885 2.898 ;
      RECT 5.875 2.222 5.88 2.933 ;
      RECT 5.87 2.224 5.875 3.015 ;
      RECT 5.865 2.226 5.87 3.103 ;
      RECT 5.855 2.228 5.865 3.185 ;
      RECT 5.84 2.242 5.855 3.19 ;
      RECT 5.805 2.287 5.84 3.19 ;
      RECT 5.795 2.327 5.805 3.19 ;
      RECT 5.78 2.355 5.795 3.19 ;
      RECT 5.775 2.372 5.78 3.19 ;
      RECT 5.77 2.38 5.775 3.19 ;
      RECT 5.76 2.395 5.765 3.19 ;
      RECT 5.755 2.402 5.76 3.19 ;
      RECT 5.745 2.422 5.755 3.19 ;
      RECT 5.74 2.435 5.745 3.19 ;
      RECT 5.705 2.44 5.71 2.775 ;
      RECT 5.69 2.83 5.71 3.19 ;
      RECT 5.69 2.44 5.7 2.748 ;
      RECT 5.685 2.87 5.69 3.19 ;
      RECT 5.635 2.44 5.685 2.743 ;
      RECT 5.68 2.907 5.685 3.19 ;
      RECT 5.67 2.93 5.68 3.19 ;
      RECT 5.665 2.975 5.67 3.19 ;
      RECT 5.655 2.985 5.665 3.183 ;
      RECT 5.581 2.44 5.635 2.737 ;
      RECT 5.495 2.44 5.581 2.73 ;
      RECT 5.446 2.487 5.495 2.723 ;
      RECT 5.36 2.495 5.446 2.716 ;
      RECT 5.345 2.492 5.36 2.711 ;
      RECT 5.331 2.485 5.345 2.71 ;
      RECT 5.245 2.485 5.331 2.705 ;
      RECT 5.15 2.49 5.16 2.69 ;
      RECT 4.74 1.92 4.755 2.32 ;
      RECT 4.935 1.92 4.94 2.18 ;
      RECT 4.68 1.92 4.725 2.18 ;
      RECT 5.135 3.225 5.14 3.43 ;
      RECT 5.13 3.215 5.135 3.435 ;
      RECT 5.125 3.202 5.13 3.44 ;
      RECT 5.12 3.182 5.125 3.44 ;
      RECT 5.095 3.135 5.12 3.44 ;
      RECT 5.06 3.05 5.095 3.44 ;
      RECT 5.055 2.987 5.06 3.44 ;
      RECT 5.05 2.972 5.055 3.44 ;
      RECT 5.035 2.932 5.05 3.44 ;
      RECT 5.03 2.907 5.035 3.44 ;
      RECT 5.02 2.89 5.03 3.44 ;
      RECT 4.985 2.812 5.02 3.44 ;
      RECT 4.98 2.755 4.985 3.44 ;
      RECT 4.975 2.742 4.98 3.44 ;
      RECT 4.965 2.72 4.975 3.44 ;
      RECT 4.955 2.685 4.965 3.44 ;
      RECT 4.945 2.655 4.955 3.44 ;
      RECT 4.935 2.57 4.945 3.083 ;
      RECT 4.942 3.215 4.945 3.44 ;
      RECT 4.94 3.225 4.942 3.44 ;
      RECT 4.93 3.235 4.94 3.435 ;
      RECT 4.925 1.92 4.935 2.315 ;
      RECT 4.93 2.447 4.935 3.058 ;
      RECT 4.925 2.345 4.93 3.041 ;
      RECT 4.915 1.92 4.925 3.017 ;
      RECT 4.91 1.92 4.915 2.988 ;
      RECT 4.905 1.92 4.91 2.978 ;
      RECT 4.885 1.92 4.905 2.94 ;
      RECT 4.88 1.92 4.885 2.898 ;
      RECT 4.875 1.92 4.88 2.878 ;
      RECT 4.845 1.92 4.875 2.828 ;
      RECT 4.835 1.92 4.845 2.775 ;
      RECT 4.83 1.92 4.835 2.748 ;
      RECT 4.825 1.92 4.83 2.733 ;
      RECT 4.815 1.92 4.825 2.71 ;
      RECT 4.805 1.92 4.815 2.685 ;
      RECT 4.8 1.92 4.805 2.625 ;
      RECT 4.79 1.92 4.8 2.563 ;
      RECT 4.785 1.92 4.79 2.483 ;
      RECT 4.78 1.92 4.785 2.448 ;
      RECT 4.775 1.92 4.78 2.423 ;
      RECT 4.77 1.92 4.775 2.408 ;
      RECT 4.765 1.92 4.77 2.378 ;
      RECT 4.76 1.92 4.765 2.355 ;
      RECT 4.755 1.92 4.76 2.328 ;
      RECT 4.725 1.92 4.74 2.315 ;
      RECT 3.88 3.455 4.065 3.665 ;
      RECT 3.87 3.46 4.08 3.658 ;
      RECT 3.87 3.46 4.1 3.63 ;
      RECT 3.87 3.46 4.115 3.609 ;
      RECT 3.87 3.46 4.13 3.607 ;
      RECT 3.87 3.46 4.14 3.606 ;
      RECT 3.87 3.46 4.17 3.603 ;
      RECT 4.52 3.305 4.78 3.565 ;
      RECT 4.48 3.352 4.78 3.548 ;
      RECT 4.471 3.36 4.48 3.551 ;
      RECT 4.065 3.453 4.78 3.548 ;
      RECT 4.385 3.378 4.471 3.558 ;
      RECT 4.08 3.45 4.78 3.548 ;
      RECT 4.326 3.4 4.385 3.57 ;
      RECT 4.1 3.446 4.78 3.548 ;
      RECT 4.24 3.412 4.326 3.581 ;
      RECT 4.115 3.442 4.78 3.548 ;
      RECT 4.185 3.425 4.24 3.593 ;
      RECT 4.13 3.44 4.78 3.548 ;
      RECT 4.17 3.431 4.185 3.599 ;
      RECT 4.14 3.436 4.78 3.548 ;
      RECT 4.285 2.96 4.545 3.22 ;
      RECT 4.285 2.98 4.655 3.19 ;
      RECT 4.285 2.985 4.665 3.185 ;
      RECT 4.476 2.399 4.555 2.63 ;
      RECT 4.39 2.402 4.605 2.625 ;
      RECT 4.385 2.402 4.605 2.62 ;
      RECT 4.385 2.407 4.615 2.618 ;
      RECT 4.36 2.407 4.615 2.615 ;
      RECT 4.36 2.415 4.625 2.613 ;
      RECT 4.24 2.35 4.5 2.61 ;
      RECT 4.24 2.397 4.55 2.61 ;
      RECT 3.495 2.97 3.5 3.23 ;
      RECT 3.325 2.74 3.33 3.23 ;
      RECT 3.21 2.98 3.215 3.205 ;
      RECT 3.92 2.075 3.925 2.285 ;
      RECT 3.925 2.08 3.94 2.28 ;
      RECT 3.86 2.075 3.92 2.293 ;
      RECT 3.845 2.075 3.86 2.303 ;
      RECT 3.795 2.075 3.845 2.32 ;
      RECT 3.775 2.075 3.795 2.343 ;
      RECT 3.76 2.075 3.775 2.355 ;
      RECT 3.74 2.075 3.76 2.365 ;
      RECT 3.73 2.08 3.74 2.374 ;
      RECT 3.725 2.09 3.73 2.379 ;
      RECT 3.72 2.102 3.725 2.383 ;
      RECT 3.71 2.125 3.72 2.388 ;
      RECT 3.705 2.14 3.71 2.392 ;
      RECT 3.7 2.157 3.705 2.395 ;
      RECT 3.695 2.165 3.7 2.398 ;
      RECT 3.685 2.17 3.695 2.402 ;
      RECT 3.68 2.177 3.685 2.407 ;
      RECT 3.67 2.182 3.68 2.411 ;
      RECT 3.645 2.194 3.67 2.422 ;
      RECT 3.625 2.211 3.645 2.438 ;
      RECT 3.6 2.228 3.625 2.46 ;
      RECT 3.565 2.251 3.6 2.518 ;
      RECT 3.545 2.273 3.565 2.58 ;
      RECT 3.54 2.283 3.545 2.615 ;
      RECT 3.53 2.29 3.54 2.653 ;
      RECT 3.525 2.297 3.53 2.673 ;
      RECT 3.52 2.308 3.525 2.71 ;
      RECT 3.515 2.316 3.52 2.775 ;
      RECT 3.505 2.327 3.515 2.828 ;
      RECT 3.5 2.345 3.505 2.898 ;
      RECT 3.495 2.355 3.5 2.935 ;
      RECT 3.49 2.365 3.495 3.23 ;
      RECT 3.485 2.377 3.49 3.23 ;
      RECT 3.48 2.387 3.485 3.23 ;
      RECT 3.47 2.397 3.48 3.23 ;
      RECT 3.46 2.42 3.47 3.23 ;
      RECT 3.445 2.455 3.46 3.23 ;
      RECT 3.405 2.517 3.445 3.23 ;
      RECT 3.4 2.57 3.405 3.23 ;
      RECT 3.375 2.605 3.4 3.23 ;
      RECT 3.36 2.65 3.375 3.23 ;
      RECT 3.355 2.672 3.36 3.23 ;
      RECT 3.345 2.685 3.355 3.23 ;
      RECT 3.335 2.71 3.345 3.23 ;
      RECT 3.33 2.732 3.335 3.23 ;
      RECT 3.305 2.77 3.325 3.23 ;
      RECT 3.265 2.827 3.305 3.23 ;
      RECT 3.26 2.877 3.265 3.23 ;
      RECT 3.255 2.895 3.26 3.23 ;
      RECT 3.25 2.907 3.255 3.23 ;
      RECT 3.24 2.925 3.25 3.23 ;
      RECT 3.23 2.945 3.24 3.205 ;
      RECT 3.225 2.962 3.23 3.205 ;
      RECT 3.215 2.975 3.225 3.205 ;
      RECT 3.185 2.985 3.21 3.205 ;
      RECT 3.175 2.992 3.185 3.205 ;
      RECT 3.16 3.002 3.175 3.2 ;
      RECT 1.54 7.765 1.83 7.995 ;
      RECT 1.6 7.025 1.77 7.995 ;
      RECT 1.51 7.025 1.86 7.315 ;
      RECT 1.135 6.285 1.485 6.575 ;
      RECT 0.995 6.315 1.485 6.485 ;
      RECT 76.05 2.85 76.42 3.22 ;
      RECT 60.265 2.85 60.635 3.22 ;
      RECT 44.48 2.85 44.85 3.22 ;
      RECT 28.705 2.85 29.075 3.22 ;
      RECT 12.925 2.85 13.295 3.22 ;
    LAYER mcon ;
      RECT 81.22 6.32 81.39 6.49 ;
      RECT 81.225 6.315 81.395 6.485 ;
      RECT 65.435 6.32 65.605 6.49 ;
      RECT 65.44 6.315 65.61 6.485 ;
      RECT 49.65 6.32 49.82 6.49 ;
      RECT 49.655 6.315 49.825 6.485 ;
      RECT 33.875 6.32 34.045 6.49 ;
      RECT 33.88 6.315 34.05 6.485 ;
      RECT 18.095 6.32 18.265 6.49 ;
      RECT 18.1 6.315 18.27 6.485 ;
      RECT 81.22 7.8 81.39 7.97 ;
      RECT 80.87 0.1 81.04 0.27 ;
      RECT 80.87 8.61 81.04 8.78 ;
      RECT 80.85 2.76 81.02 2.93 ;
      RECT 80.85 5.95 81.02 6.12 ;
      RECT 80.23 0.91 80.4 1.08 ;
      RECT 80.23 2.39 80.4 2.56 ;
      RECT 80.23 6.32 80.4 6.49 ;
      RECT 80.23 7.8 80.4 7.97 ;
      RECT 79.88 0.1 80.05 0.27 ;
      RECT 79.88 8.61 80.05 8.78 ;
      RECT 79.86 2.76 80.03 2.93 ;
      RECT 79.86 5.95 80.03 6.12 ;
      RECT 79.18 0.105 79.35 0.275 ;
      RECT 79.18 8.605 79.35 8.775 ;
      RECT 78.87 2.025 79.04 2.195 ;
      RECT 78.87 6.685 79.04 6.855 ;
      RECT 78.5 0.105 78.67 0.275 ;
      RECT 78.5 8.605 78.67 8.775 ;
      RECT 78.44 0.915 78.61 1.085 ;
      RECT 78.44 1.655 78.61 1.825 ;
      RECT 78.44 7.055 78.61 7.225 ;
      RECT 78.44 7.795 78.61 7.965 ;
      RECT 78.065 2.395 78.235 2.565 ;
      RECT 78.065 6.315 78.235 6.485 ;
      RECT 77.82 0.105 77.99 0.275 ;
      RECT 77.82 8.605 77.99 8.775 ;
      RECT 77.14 0.105 77.31 0.275 ;
      RECT 77.14 8.605 77.31 8.775 ;
      RECT 75.515 1.415 75.685 1.585 ;
      RECT 75.145 2.875 75.315 3.045 ;
      RECT 75.055 1.415 75.225 1.585 ;
      RECT 74.825 2.045 74.995 2.215 ;
      RECT 74.68 2.485 74.85 2.655 ;
      RECT 74.595 1.415 74.765 1.585 ;
      RECT 74.4 8.605 74.57 8.775 ;
      RECT 74.135 1.415 74.305 1.585 ;
      RECT 74.09 6.685 74.26 6.855 ;
      RECT 74.07 2.525 74.24 2.695 ;
      RECT 73.725 2.16 73.895 2.33 ;
      RECT 73.72 8.605 73.89 8.775 ;
      RECT 73.715 3.52 73.885 3.69 ;
      RECT 73.675 1.415 73.845 1.585 ;
      RECT 73.66 7.055 73.83 7.225 ;
      RECT 73.66 7.795 73.83 7.965 ;
      RECT 73.3 2.76 73.47 2.93 ;
      RECT 73.285 6.315 73.455 6.485 ;
      RECT 73.215 1.415 73.385 1.585 ;
      RECT 73.04 8.605 73.21 8.775 ;
      RECT 72.95 2.235 73.12 2.405 ;
      RECT 72.77 3.55 72.94 3.72 ;
      RECT 72.755 1.415 72.925 1.585 ;
      RECT 72.49 2.865 72.66 3.035 ;
      RECT 72.36 8.605 72.53 8.775 ;
      RECT 72.295 1.415 72.465 1.585 ;
      RECT 72.17 2.49 72.34 2.66 ;
      RECT 71.835 1.415 72.005 1.585 ;
      RECT 71.48 1.97 71.65 2.14 ;
      RECT 71.405 2.44 71.575 2.61 ;
      RECT 71.375 1.415 71.545 1.585 ;
      RECT 70.915 1.415 71.085 1.585 ;
      RECT 70.555 2.165 70.725 2.335 ;
      RECT 70.455 1.415 70.625 1.585 ;
      RECT 70.215 3.36 70.385 3.53 ;
      RECT 70.18 2.695 70.35 2.865 ;
      RECT 69.995 1.415 70.165 1.585 ;
      RECT 69.57 2.55 69.74 2.72 ;
      RECT 69.535 1.415 69.705 1.585 ;
      RECT 69.5 3.25 69.67 3.42 ;
      RECT 69.44 2.085 69.61 2.255 ;
      RECT 69.075 1.415 69.245 1.585 ;
      RECT 68.8 3 68.97 3.17 ;
      RECT 68.615 1.415 68.785 1.585 ;
      RECT 68.295 2.505 68.465 2.675 ;
      RECT 68.155 1.415 68.325 1.585 ;
      RECT 68.075 3.25 68.245 3.42 ;
      RECT 67.87 2.13 68.04 2.3 ;
      RECT 67.695 1.415 67.865 1.585 ;
      RECT 67.6 3 67.77 3.17 ;
      RECT 67.56 2.43 67.73 2.6 ;
      RECT 67.235 1.415 67.405 1.585 ;
      RECT 67.015 3.475 67.185 3.645 ;
      RECT 66.875 2.095 67.045 2.265 ;
      RECT 66.775 1.415 66.945 1.585 ;
      RECT 66.315 1.415 66.485 1.585 ;
      RECT 66.305 3.015 66.475 3.185 ;
      RECT 65.435 7.8 65.605 7.97 ;
      RECT 65.085 0.1 65.255 0.27 ;
      RECT 65.085 8.61 65.255 8.78 ;
      RECT 65.065 2.76 65.235 2.93 ;
      RECT 65.065 5.95 65.235 6.12 ;
      RECT 64.445 0.91 64.615 1.08 ;
      RECT 64.445 2.39 64.615 2.56 ;
      RECT 64.445 6.32 64.615 6.49 ;
      RECT 64.445 7.8 64.615 7.97 ;
      RECT 64.095 0.1 64.265 0.27 ;
      RECT 64.095 8.61 64.265 8.78 ;
      RECT 64.075 2.76 64.245 2.93 ;
      RECT 64.075 5.95 64.245 6.12 ;
      RECT 63.395 0.105 63.565 0.275 ;
      RECT 63.395 8.605 63.565 8.775 ;
      RECT 63.085 2.025 63.255 2.195 ;
      RECT 63.085 6.685 63.255 6.855 ;
      RECT 62.715 0.105 62.885 0.275 ;
      RECT 62.715 8.605 62.885 8.775 ;
      RECT 62.655 0.915 62.825 1.085 ;
      RECT 62.655 1.655 62.825 1.825 ;
      RECT 62.655 7.055 62.825 7.225 ;
      RECT 62.655 7.795 62.825 7.965 ;
      RECT 62.28 2.395 62.45 2.565 ;
      RECT 62.28 6.315 62.45 6.485 ;
      RECT 62.035 0.105 62.205 0.275 ;
      RECT 62.035 8.605 62.205 8.775 ;
      RECT 61.355 0.105 61.525 0.275 ;
      RECT 61.355 8.605 61.525 8.775 ;
      RECT 59.73 1.415 59.9 1.585 ;
      RECT 59.36 2.875 59.53 3.045 ;
      RECT 59.27 1.415 59.44 1.585 ;
      RECT 59.04 2.045 59.21 2.215 ;
      RECT 58.895 2.485 59.065 2.655 ;
      RECT 58.81 1.415 58.98 1.585 ;
      RECT 58.615 8.605 58.785 8.775 ;
      RECT 58.35 1.415 58.52 1.585 ;
      RECT 58.305 6.685 58.475 6.855 ;
      RECT 58.285 2.525 58.455 2.695 ;
      RECT 57.94 2.16 58.11 2.33 ;
      RECT 57.935 8.605 58.105 8.775 ;
      RECT 57.93 3.52 58.1 3.69 ;
      RECT 57.89 1.415 58.06 1.585 ;
      RECT 57.875 7.055 58.045 7.225 ;
      RECT 57.875 7.795 58.045 7.965 ;
      RECT 57.515 2.76 57.685 2.93 ;
      RECT 57.5 6.315 57.67 6.485 ;
      RECT 57.43 1.415 57.6 1.585 ;
      RECT 57.255 8.605 57.425 8.775 ;
      RECT 57.165 2.235 57.335 2.405 ;
      RECT 56.985 3.55 57.155 3.72 ;
      RECT 56.97 1.415 57.14 1.585 ;
      RECT 56.705 2.865 56.875 3.035 ;
      RECT 56.575 8.605 56.745 8.775 ;
      RECT 56.51 1.415 56.68 1.585 ;
      RECT 56.385 2.49 56.555 2.66 ;
      RECT 56.05 1.415 56.22 1.585 ;
      RECT 55.695 1.97 55.865 2.14 ;
      RECT 55.62 2.44 55.79 2.61 ;
      RECT 55.59 1.415 55.76 1.585 ;
      RECT 55.13 1.415 55.3 1.585 ;
      RECT 54.77 2.165 54.94 2.335 ;
      RECT 54.67 1.415 54.84 1.585 ;
      RECT 54.43 3.36 54.6 3.53 ;
      RECT 54.395 2.695 54.565 2.865 ;
      RECT 54.21 1.415 54.38 1.585 ;
      RECT 53.785 2.55 53.955 2.72 ;
      RECT 53.75 1.415 53.92 1.585 ;
      RECT 53.715 3.25 53.885 3.42 ;
      RECT 53.655 2.085 53.825 2.255 ;
      RECT 53.29 1.415 53.46 1.585 ;
      RECT 53.015 3 53.185 3.17 ;
      RECT 52.83 1.415 53 1.585 ;
      RECT 52.51 2.505 52.68 2.675 ;
      RECT 52.37 1.415 52.54 1.585 ;
      RECT 52.29 3.25 52.46 3.42 ;
      RECT 52.085 2.13 52.255 2.3 ;
      RECT 51.91 1.415 52.08 1.585 ;
      RECT 51.815 3 51.985 3.17 ;
      RECT 51.775 2.43 51.945 2.6 ;
      RECT 51.45 1.415 51.62 1.585 ;
      RECT 51.23 3.475 51.4 3.645 ;
      RECT 51.09 2.095 51.26 2.265 ;
      RECT 50.99 1.415 51.16 1.585 ;
      RECT 50.53 1.415 50.7 1.585 ;
      RECT 50.52 3.015 50.69 3.185 ;
      RECT 49.65 7.8 49.82 7.97 ;
      RECT 49.3 0.1 49.47 0.27 ;
      RECT 49.3 8.61 49.47 8.78 ;
      RECT 49.28 2.76 49.45 2.93 ;
      RECT 49.28 5.95 49.45 6.12 ;
      RECT 48.66 0.91 48.83 1.08 ;
      RECT 48.66 2.39 48.83 2.56 ;
      RECT 48.66 6.32 48.83 6.49 ;
      RECT 48.66 7.8 48.83 7.97 ;
      RECT 48.31 0.1 48.48 0.27 ;
      RECT 48.31 8.61 48.48 8.78 ;
      RECT 48.29 2.76 48.46 2.93 ;
      RECT 48.29 5.95 48.46 6.12 ;
      RECT 47.61 0.105 47.78 0.275 ;
      RECT 47.61 8.605 47.78 8.775 ;
      RECT 47.3 2.025 47.47 2.195 ;
      RECT 47.3 6.685 47.47 6.855 ;
      RECT 46.93 0.105 47.1 0.275 ;
      RECT 46.93 8.605 47.1 8.775 ;
      RECT 46.87 0.915 47.04 1.085 ;
      RECT 46.87 1.655 47.04 1.825 ;
      RECT 46.87 7.055 47.04 7.225 ;
      RECT 46.87 7.795 47.04 7.965 ;
      RECT 46.495 2.395 46.665 2.565 ;
      RECT 46.495 6.315 46.665 6.485 ;
      RECT 46.25 0.105 46.42 0.275 ;
      RECT 46.25 8.605 46.42 8.775 ;
      RECT 45.57 0.105 45.74 0.275 ;
      RECT 45.57 8.605 45.74 8.775 ;
      RECT 43.945 1.415 44.115 1.585 ;
      RECT 43.575 2.875 43.745 3.045 ;
      RECT 43.485 1.415 43.655 1.585 ;
      RECT 43.255 2.045 43.425 2.215 ;
      RECT 43.11 2.485 43.28 2.655 ;
      RECT 43.025 1.415 43.195 1.585 ;
      RECT 42.83 8.605 43 8.775 ;
      RECT 42.565 1.415 42.735 1.585 ;
      RECT 42.52 6.685 42.69 6.855 ;
      RECT 42.5 2.525 42.67 2.695 ;
      RECT 42.155 2.16 42.325 2.33 ;
      RECT 42.15 8.605 42.32 8.775 ;
      RECT 42.145 3.52 42.315 3.69 ;
      RECT 42.105 1.415 42.275 1.585 ;
      RECT 42.09 7.055 42.26 7.225 ;
      RECT 42.09 7.795 42.26 7.965 ;
      RECT 41.73 2.76 41.9 2.93 ;
      RECT 41.715 6.315 41.885 6.485 ;
      RECT 41.645 1.415 41.815 1.585 ;
      RECT 41.47 8.605 41.64 8.775 ;
      RECT 41.38 2.235 41.55 2.405 ;
      RECT 41.2 3.55 41.37 3.72 ;
      RECT 41.185 1.415 41.355 1.585 ;
      RECT 40.92 2.865 41.09 3.035 ;
      RECT 40.79 8.605 40.96 8.775 ;
      RECT 40.725 1.415 40.895 1.585 ;
      RECT 40.6 2.49 40.77 2.66 ;
      RECT 40.265 1.415 40.435 1.585 ;
      RECT 39.91 1.97 40.08 2.14 ;
      RECT 39.835 2.44 40.005 2.61 ;
      RECT 39.805 1.415 39.975 1.585 ;
      RECT 39.345 1.415 39.515 1.585 ;
      RECT 38.985 2.165 39.155 2.335 ;
      RECT 38.885 1.415 39.055 1.585 ;
      RECT 38.645 3.36 38.815 3.53 ;
      RECT 38.61 2.695 38.78 2.865 ;
      RECT 38.425 1.415 38.595 1.585 ;
      RECT 38 2.55 38.17 2.72 ;
      RECT 37.965 1.415 38.135 1.585 ;
      RECT 37.93 3.25 38.1 3.42 ;
      RECT 37.87 2.085 38.04 2.255 ;
      RECT 37.505 1.415 37.675 1.585 ;
      RECT 37.23 3 37.4 3.17 ;
      RECT 37.045 1.415 37.215 1.585 ;
      RECT 36.725 2.505 36.895 2.675 ;
      RECT 36.585 1.415 36.755 1.585 ;
      RECT 36.505 3.25 36.675 3.42 ;
      RECT 36.3 2.13 36.47 2.3 ;
      RECT 36.125 1.415 36.295 1.585 ;
      RECT 36.03 3 36.2 3.17 ;
      RECT 35.99 2.43 36.16 2.6 ;
      RECT 35.665 1.415 35.835 1.585 ;
      RECT 35.445 3.475 35.615 3.645 ;
      RECT 35.305 2.095 35.475 2.265 ;
      RECT 35.205 1.415 35.375 1.585 ;
      RECT 34.745 1.415 34.915 1.585 ;
      RECT 34.735 3.015 34.905 3.185 ;
      RECT 33.875 7.8 34.045 7.97 ;
      RECT 33.525 0.1 33.695 0.27 ;
      RECT 33.525 8.61 33.695 8.78 ;
      RECT 33.505 2.76 33.675 2.93 ;
      RECT 33.505 5.95 33.675 6.12 ;
      RECT 32.885 0.91 33.055 1.08 ;
      RECT 32.885 2.39 33.055 2.56 ;
      RECT 32.885 6.32 33.055 6.49 ;
      RECT 32.885 7.8 33.055 7.97 ;
      RECT 32.535 0.1 32.705 0.27 ;
      RECT 32.535 8.61 32.705 8.78 ;
      RECT 32.515 2.76 32.685 2.93 ;
      RECT 32.515 5.95 32.685 6.12 ;
      RECT 31.835 0.105 32.005 0.275 ;
      RECT 31.835 8.605 32.005 8.775 ;
      RECT 31.525 2.025 31.695 2.195 ;
      RECT 31.525 6.685 31.695 6.855 ;
      RECT 31.155 0.105 31.325 0.275 ;
      RECT 31.155 8.605 31.325 8.775 ;
      RECT 31.095 0.915 31.265 1.085 ;
      RECT 31.095 1.655 31.265 1.825 ;
      RECT 31.095 7.055 31.265 7.225 ;
      RECT 31.095 7.795 31.265 7.965 ;
      RECT 30.72 2.395 30.89 2.565 ;
      RECT 30.72 6.315 30.89 6.485 ;
      RECT 30.475 0.105 30.645 0.275 ;
      RECT 30.475 8.605 30.645 8.775 ;
      RECT 29.795 0.105 29.965 0.275 ;
      RECT 29.795 8.605 29.965 8.775 ;
      RECT 28.17 1.415 28.34 1.585 ;
      RECT 27.8 2.875 27.97 3.045 ;
      RECT 27.71 1.415 27.88 1.585 ;
      RECT 27.48 2.045 27.65 2.215 ;
      RECT 27.335 2.485 27.505 2.655 ;
      RECT 27.25 1.415 27.42 1.585 ;
      RECT 27.055 8.605 27.225 8.775 ;
      RECT 26.79 1.415 26.96 1.585 ;
      RECT 26.745 6.685 26.915 6.855 ;
      RECT 26.725 2.525 26.895 2.695 ;
      RECT 26.38 2.16 26.55 2.33 ;
      RECT 26.375 8.605 26.545 8.775 ;
      RECT 26.37 3.52 26.54 3.69 ;
      RECT 26.33 1.415 26.5 1.585 ;
      RECT 26.315 7.055 26.485 7.225 ;
      RECT 26.315 7.795 26.485 7.965 ;
      RECT 25.955 2.76 26.125 2.93 ;
      RECT 25.94 6.315 26.11 6.485 ;
      RECT 25.87 1.415 26.04 1.585 ;
      RECT 25.695 8.605 25.865 8.775 ;
      RECT 25.605 2.235 25.775 2.405 ;
      RECT 25.425 3.55 25.595 3.72 ;
      RECT 25.41 1.415 25.58 1.585 ;
      RECT 25.145 2.865 25.315 3.035 ;
      RECT 25.015 8.605 25.185 8.775 ;
      RECT 24.95 1.415 25.12 1.585 ;
      RECT 24.825 2.49 24.995 2.66 ;
      RECT 24.49 1.415 24.66 1.585 ;
      RECT 24.135 1.97 24.305 2.14 ;
      RECT 24.06 2.44 24.23 2.61 ;
      RECT 24.03 1.415 24.2 1.585 ;
      RECT 23.57 1.415 23.74 1.585 ;
      RECT 23.21 2.165 23.38 2.335 ;
      RECT 23.11 1.415 23.28 1.585 ;
      RECT 22.87 3.36 23.04 3.53 ;
      RECT 22.835 2.695 23.005 2.865 ;
      RECT 22.65 1.415 22.82 1.585 ;
      RECT 22.225 2.55 22.395 2.72 ;
      RECT 22.19 1.415 22.36 1.585 ;
      RECT 22.155 3.25 22.325 3.42 ;
      RECT 22.095 2.085 22.265 2.255 ;
      RECT 21.73 1.415 21.9 1.585 ;
      RECT 21.455 3 21.625 3.17 ;
      RECT 21.27 1.415 21.44 1.585 ;
      RECT 20.95 2.505 21.12 2.675 ;
      RECT 20.81 1.415 20.98 1.585 ;
      RECT 20.73 3.25 20.9 3.42 ;
      RECT 20.525 2.13 20.695 2.3 ;
      RECT 20.35 1.415 20.52 1.585 ;
      RECT 20.255 3 20.425 3.17 ;
      RECT 20.215 2.43 20.385 2.6 ;
      RECT 19.89 1.415 20.06 1.585 ;
      RECT 19.67 3.475 19.84 3.645 ;
      RECT 19.53 2.095 19.7 2.265 ;
      RECT 19.43 1.415 19.6 1.585 ;
      RECT 18.97 1.415 19.14 1.585 ;
      RECT 18.96 3.015 19.13 3.185 ;
      RECT 18.095 7.8 18.265 7.97 ;
      RECT 17.745 0.1 17.915 0.27 ;
      RECT 17.745 8.61 17.915 8.78 ;
      RECT 17.725 2.76 17.895 2.93 ;
      RECT 17.725 5.95 17.895 6.12 ;
      RECT 17.105 0.91 17.275 1.08 ;
      RECT 17.105 2.39 17.275 2.56 ;
      RECT 17.105 6.32 17.275 6.49 ;
      RECT 17.105 7.8 17.275 7.97 ;
      RECT 16.755 0.1 16.925 0.27 ;
      RECT 16.755 8.61 16.925 8.78 ;
      RECT 16.735 2.76 16.905 2.93 ;
      RECT 16.735 5.95 16.905 6.12 ;
      RECT 16.055 0.105 16.225 0.275 ;
      RECT 16.055 8.605 16.225 8.775 ;
      RECT 15.745 2.025 15.915 2.195 ;
      RECT 15.745 6.685 15.915 6.855 ;
      RECT 15.375 0.105 15.545 0.275 ;
      RECT 15.375 8.605 15.545 8.775 ;
      RECT 15.315 0.915 15.485 1.085 ;
      RECT 15.315 1.655 15.485 1.825 ;
      RECT 15.315 7.055 15.485 7.225 ;
      RECT 15.315 7.795 15.485 7.965 ;
      RECT 14.94 2.395 15.11 2.565 ;
      RECT 14.94 6.315 15.11 6.485 ;
      RECT 14.695 0.105 14.865 0.275 ;
      RECT 14.695 8.605 14.865 8.775 ;
      RECT 14.015 0.105 14.185 0.275 ;
      RECT 14.015 8.605 14.185 8.775 ;
      RECT 12.39 1.415 12.56 1.585 ;
      RECT 12.02 2.875 12.19 3.045 ;
      RECT 11.93 1.415 12.1 1.585 ;
      RECT 11.7 2.045 11.87 2.215 ;
      RECT 11.555 2.485 11.725 2.655 ;
      RECT 11.47 1.415 11.64 1.585 ;
      RECT 11.275 8.605 11.445 8.775 ;
      RECT 11.01 1.415 11.18 1.585 ;
      RECT 10.965 6.685 11.135 6.855 ;
      RECT 10.945 2.525 11.115 2.695 ;
      RECT 10.6 2.16 10.77 2.33 ;
      RECT 10.595 8.605 10.765 8.775 ;
      RECT 10.59 3.52 10.76 3.69 ;
      RECT 10.55 1.415 10.72 1.585 ;
      RECT 10.535 7.055 10.705 7.225 ;
      RECT 10.535 7.795 10.705 7.965 ;
      RECT 10.175 2.76 10.345 2.93 ;
      RECT 10.16 6.315 10.33 6.485 ;
      RECT 10.09 1.415 10.26 1.585 ;
      RECT 9.915 8.605 10.085 8.775 ;
      RECT 9.825 2.235 9.995 2.405 ;
      RECT 9.645 3.55 9.815 3.72 ;
      RECT 9.63 1.415 9.8 1.585 ;
      RECT 9.365 2.865 9.535 3.035 ;
      RECT 9.235 8.605 9.405 8.775 ;
      RECT 9.17 1.415 9.34 1.585 ;
      RECT 9.045 2.49 9.215 2.66 ;
      RECT 8.71 1.415 8.88 1.585 ;
      RECT 8.355 1.97 8.525 2.14 ;
      RECT 8.28 2.44 8.45 2.61 ;
      RECT 8.25 1.415 8.42 1.585 ;
      RECT 7.79 1.415 7.96 1.585 ;
      RECT 7.43 2.165 7.6 2.335 ;
      RECT 7.33 1.415 7.5 1.585 ;
      RECT 7.09 3.36 7.26 3.53 ;
      RECT 7.055 2.695 7.225 2.865 ;
      RECT 6.87 1.415 7.04 1.585 ;
      RECT 6.445 2.55 6.615 2.72 ;
      RECT 6.41 1.415 6.58 1.585 ;
      RECT 6.375 3.25 6.545 3.42 ;
      RECT 6.315 2.085 6.485 2.255 ;
      RECT 5.95 1.415 6.12 1.585 ;
      RECT 5.675 3 5.845 3.17 ;
      RECT 5.49 1.415 5.66 1.585 ;
      RECT 5.17 2.505 5.34 2.675 ;
      RECT 5.03 1.415 5.2 1.585 ;
      RECT 4.95 3.25 5.12 3.42 ;
      RECT 4.745 2.13 4.915 2.3 ;
      RECT 4.57 1.415 4.74 1.585 ;
      RECT 4.475 3 4.645 3.17 ;
      RECT 4.435 2.43 4.605 2.6 ;
      RECT 4.11 1.415 4.28 1.585 ;
      RECT 3.89 3.475 4.06 3.645 ;
      RECT 3.75 2.095 3.92 2.265 ;
      RECT 3.65 1.415 3.82 1.585 ;
      RECT 3.19 1.415 3.36 1.585 ;
      RECT 3.18 3.015 3.35 3.185 ;
      RECT 2.34 8.605 2.51 8.775 ;
      RECT 1.66 8.605 1.83 8.775 ;
      RECT 1.6 7.055 1.77 7.225 ;
      RECT 1.6 7.795 1.77 7.965 ;
      RECT 1.225 6.315 1.395 6.485 ;
      RECT 0.98 8.605 1.15 8.775 ;
      RECT 0.3 8.605 0.47 8.775 ;
    LAYER li1 ;
      RECT 74.3 0 74.47 2.085 ;
      RECT 72.34 0 72.51 2.085 ;
      RECT 69.9 0 70.07 2.085 ;
      RECT 68.94 0 69.11 2.085 ;
      RECT 68.42 0 68.59 2.085 ;
      RECT 67.46 0 67.63 2.085 ;
      RECT 66.5 0 66.67 2.085 ;
      RECT 58.515 0 58.685 2.085 ;
      RECT 56.555 0 56.725 2.085 ;
      RECT 54.115 0 54.285 2.085 ;
      RECT 53.155 0 53.325 2.085 ;
      RECT 52.635 0 52.805 2.085 ;
      RECT 51.675 0 51.845 2.085 ;
      RECT 50.715 0 50.885 2.085 ;
      RECT 42.73 0 42.9 2.085 ;
      RECT 40.77 0 40.94 2.085 ;
      RECT 38.33 0 38.5 2.085 ;
      RECT 37.37 0 37.54 2.085 ;
      RECT 36.85 0 37.02 2.085 ;
      RECT 35.89 0 36.06 2.085 ;
      RECT 34.93 0 35.1 2.085 ;
      RECT 26.955 0 27.125 2.085 ;
      RECT 24.995 0 25.165 2.085 ;
      RECT 22.555 0 22.725 2.085 ;
      RECT 21.595 0 21.765 2.085 ;
      RECT 21.075 0 21.245 2.085 ;
      RECT 20.115 0 20.285 2.085 ;
      RECT 19.155 0 19.325 2.085 ;
      RECT 11.175 0 11.345 2.085 ;
      RECT 9.215 0 9.385 2.085 ;
      RECT 6.775 0 6.945 2.085 ;
      RECT 5.815 0 5.985 2.085 ;
      RECT 5.295 0 5.465 2.085 ;
      RECT 4.335 0 4.505 2.085 ;
      RECT 3.375 0 3.545 2.085 ;
      RECT 66.285 0 75.885 1.59 ;
      RECT 50.5 0 60.1 1.59 ;
      RECT 34.715 0 44.315 1.59 ;
      RECT 18.94 0 28.54 1.59 ;
      RECT 3.16 0 12.76 1.59 ;
      RECT 66.17 1.415 76 1.585 ;
      RECT 66.285 0 76 1.585 ;
      RECT 50.385 1.415 60.215 1.585 ;
      RECT 50.5 0 60.215 1.585 ;
      RECT 34.6 1.415 44.43 1.585 ;
      RECT 34.715 0 44.43 1.585 ;
      RECT 18.825 1.415 28.655 1.585 ;
      RECT 18.94 0 28.655 1.585 ;
      RECT 3.045 1.415 12.875 1.585 ;
      RECT 3.16 0 12.875 1.585 ;
      RECT 77.06 0 77.23 0.935 ;
      RECT 61.275 0 61.445 0.935 ;
      RECT 45.49 0 45.66 0.935 ;
      RECT 29.715 0 29.885 0.935 ;
      RECT 13.935 0 14.105 0.935 ;
      RECT 80.79 0 80.96 0.93 ;
      RECT 79.8 0 79.97 0.93 ;
      RECT 65.005 0 65.175 0.93 ;
      RECT 64.015 0 64.185 0.93 ;
      RECT 49.22 0 49.39 0.93 ;
      RECT 48.23 0 48.4 0.93 ;
      RECT 33.445 0 33.615 0.93 ;
      RECT 32.455 0 32.625 0.93 ;
      RECT 17.665 0 17.835 0.93 ;
      RECT 16.675 0 16.845 0.93 ;
      RECT 0.295 0.245 0.465 0.335 ;
      RECT 0 0.245 0.805 0.315 ;
      RECT 81.585 0 81.765 0.305 ;
      RECT 65.8 0 79.635 0.305 ;
      RECT 50.015 0 63.85 0.305 ;
      RECT 34.24 0 48.065 0.305 ;
      RECT 18.46 0 32.29 0.305 ;
      RECT 0 0.245 16.51 0.305 ;
      RECT 0.465 0 81.765 0.3 ;
      RECT 0 0 0.295 0.315 ;
      RECT 0 0 81.765 0.075 ;
      RECT 0 8.58 81.765 8.88 ;
      RECT 81.585 8.575 81.765 8.88 ;
      RECT 80.79 7.95 80.96 8.88 ;
      RECT 79.8 7.95 79.97 8.88 ;
      RECT 65.8 8.575 79.635 8.88 ;
      RECT 65.005 7.95 65.175 8.88 ;
      RECT 64.015 7.95 64.185 8.88 ;
      RECT 50.015 8.575 63.85 8.88 ;
      RECT 49.22 7.95 49.39 8.88 ;
      RECT 48.23 7.95 48.4 8.88 ;
      RECT 34.24 8.575 48.065 8.88 ;
      RECT 33.445 7.95 33.615 8.88 ;
      RECT 32.455 7.95 32.625 8.88 ;
      RECT 18.46 8.575 32.29 8.88 ;
      RECT 17.665 7.95 17.835 8.88 ;
      RECT 16.675 7.95 16.845 8.88 ;
      RECT 0 8.575 16.51 8.88 ;
      RECT 77.06 7.945 77.23 8.88 ;
      RECT 72.28 7.945 72.45 8.88 ;
      RECT 61.275 7.945 61.445 8.88 ;
      RECT 56.495 7.945 56.665 8.88 ;
      RECT 45.49 7.945 45.66 8.88 ;
      RECT 40.71 7.945 40.88 8.88 ;
      RECT 29.715 7.945 29.885 8.88 ;
      RECT 24.935 7.945 25.105 8.88 ;
      RECT 13.935 7.945 14.105 8.88 ;
      RECT 9.155 7.945 9.325 8.88 ;
      RECT 0 8.565 0.805 8.88 ;
      RECT 0.22 8.545 0.465 8.88 ;
      RECT 0.22 7.945 0.39 8.88 ;
      RECT 81.22 5.02 81.39 6.49 ;
      RECT 81.22 6.315 81.395 6.485 ;
      RECT 80.85 1.74 81.02 2.93 ;
      RECT 80.85 1.74 81.32 1.91 ;
      RECT 80.85 6.97 81.32 7.14 ;
      RECT 80.85 5.95 81.02 7.14 ;
      RECT 79.86 1.74 80.03 2.93 ;
      RECT 79.86 1.74 80.33 1.91 ;
      RECT 79.86 6.97 80.33 7.14 ;
      RECT 79.86 5.95 80.03 7.14 ;
      RECT 78.01 2.635 78.18 3.865 ;
      RECT 78.065 0.855 78.235 2.805 ;
      RECT 78.01 0.575 78.18 1.025 ;
      RECT 78.01 7.855 78.18 8.305 ;
      RECT 78.065 6.075 78.235 8.025 ;
      RECT 78.01 5.015 78.18 6.245 ;
      RECT 77.49 0.575 77.66 3.865 ;
      RECT 77.49 2.075 77.895 2.405 ;
      RECT 77.49 1.235 77.895 1.565 ;
      RECT 77.49 5.015 77.66 8.305 ;
      RECT 77.49 7.315 77.895 7.645 ;
      RECT 77.49 6.475 77.895 6.805 ;
      RECT 74.825 1.975 75.555 2.215 ;
      RECT 75.367 1.77 75.555 2.215 ;
      RECT 75.195 1.782 75.57 2.209 ;
      RECT 75.11 1.797 75.59 2.194 ;
      RECT 75.11 1.812 75.595 2.184 ;
      RECT 75.065 1.832 75.61 2.176 ;
      RECT 75.042 1.867 75.625 2.13 ;
      RECT 74.956 1.89 75.63 2.09 ;
      RECT 74.956 1.908 75.64 2.06 ;
      RECT 74.825 1.977 75.645 2.023 ;
      RECT 74.87 1.92 75.64 2.06 ;
      RECT 74.956 1.872 75.625 2.13 ;
      RECT 75.042 1.841 75.61 2.176 ;
      RECT 75.065 1.822 75.595 2.184 ;
      RECT 75.11 1.795 75.57 2.209 ;
      RECT 75.195 1.777 75.555 2.215 ;
      RECT 75.281 1.771 75.555 2.215 ;
      RECT 75.367 1.766 75.5 2.215 ;
      RECT 75.453 1.761 75.5 2.215 ;
      RECT 75.145 2.659 75.315 3.045 ;
      RECT 75.14 2.659 75.315 3.04 ;
      RECT 75.115 2.659 75.315 3.005 ;
      RECT 75.115 2.687 75.325 2.995 ;
      RECT 75.095 2.687 75.325 2.955 ;
      RECT 75.09 2.687 75.325 2.928 ;
      RECT 75.09 2.705 75.33 2.92 ;
      RECT 75.035 2.705 75.33 2.855 ;
      RECT 75.035 2.722 75.34 2.838 ;
      RECT 75.025 2.722 75.34 2.778 ;
      RECT 75.025 2.739 75.345 2.775 ;
      RECT 75.02 2.575 75.19 2.753 ;
      RECT 75.02 2.609 75.276 2.753 ;
      RECT 75.015 3.375 75.02 3.388 ;
      RECT 75.01 3.27 75.015 3.393 ;
      RECT 74.985 3.13 75.01 3.408 ;
      RECT 74.95 3.081 74.985 3.44 ;
      RECT 74.945 3.049 74.95 3.46 ;
      RECT 74.94 3.04 74.945 3.46 ;
      RECT 74.86 3.005 74.94 3.46 ;
      RECT 74.797 2.975 74.86 3.46 ;
      RECT 74.711 2.963 74.797 3.46 ;
      RECT 74.625 2.949 74.711 3.46 ;
      RECT 74.545 2.936 74.625 3.446 ;
      RECT 74.51 2.928 74.545 3.426 ;
      RECT 74.5 2.925 74.51 3.417 ;
      RECT 74.47 2.92 74.5 3.404 ;
      RECT 74.42 2.895 74.47 3.38 ;
      RECT 74.406 2.869 74.42 3.362 ;
      RECT 74.32 2.829 74.406 3.338 ;
      RECT 74.275 2.777 74.32 3.307 ;
      RECT 74.265 2.752 74.275 3.294 ;
      RECT 74.26 2.533 74.265 2.555 ;
      RECT 74.255 2.735 74.265 3.29 ;
      RECT 74.255 2.531 74.26 2.645 ;
      RECT 74.245 2.527 74.255 3.286 ;
      RECT 74.201 2.525 74.245 3.274 ;
      RECT 74.115 2.525 74.201 3.245 ;
      RECT 74.085 2.525 74.115 3.218 ;
      RECT 74.07 2.525 74.085 3.206 ;
      RECT 74.03 2.537 74.07 3.191 ;
      RECT 74.01 2.556 74.03 3.17 ;
      RECT 74 2.566 74.01 3.154 ;
      RECT 73.99 2.572 74 3.143 ;
      RECT 73.97 2.582 73.99 3.126 ;
      RECT 73.965 2.591 73.97 3.113 ;
      RECT 73.96 2.595 73.965 3.063 ;
      RECT 73.95 2.601 73.96 2.98 ;
      RECT 73.945 2.605 73.95 2.894 ;
      RECT 73.94 2.625 73.945 2.831 ;
      RECT 73.935 2.648 73.94 2.778 ;
      RECT 73.93 2.666 73.935 2.723 ;
      RECT 74.54 2.485 74.71 2.745 ;
      RECT 74.71 2.45 74.755 2.731 ;
      RECT 74.671 2.452 74.76 2.714 ;
      RECT 74.56 2.469 74.846 2.685 ;
      RECT 74.56 2.484 74.85 2.657 ;
      RECT 74.56 2.465 74.76 2.714 ;
      RECT 74.585 2.453 74.71 2.745 ;
      RECT 74.671 2.451 74.755 2.731 ;
      RECT 73.725 1.84 73.895 2.33 ;
      RECT 73.725 1.84 73.93 2.31 ;
      RECT 73.86 1.76 73.97 2.27 ;
      RECT 73.841 1.764 73.99 2.24 ;
      RECT 73.755 1.772 74.01 2.223 ;
      RECT 73.755 1.778 74.015 2.213 ;
      RECT 73.755 1.787 74.035 2.201 ;
      RECT 73.73 1.812 74.065 2.179 ;
      RECT 73.73 1.832 74.07 2.159 ;
      RECT 73.725 1.845 74.08 2.139 ;
      RECT 73.725 1.912 74.085 2.12 ;
      RECT 73.725 2.045 74.09 2.107 ;
      RECT 73.72 1.85 74.08 1.94 ;
      RECT 73.73 1.807 74.035 2.201 ;
      RECT 73.841 1.762 73.97 2.27 ;
      RECT 73.715 3.515 74.015 3.77 ;
      RECT 73.8 3.481 74.015 3.77 ;
      RECT 73.8 3.484 74.02 3.63 ;
      RECT 73.735 3.505 74.02 3.63 ;
      RECT 73.77 3.495 74.015 3.77 ;
      RECT 73.765 3.5 74.02 3.63 ;
      RECT 73.8 3.479 74.001 3.77 ;
      RECT 73.886 3.47 74.001 3.77 ;
      RECT 73.886 3.464 73.915 3.77 ;
      RECT 73.375 3.105 73.385 3.595 ;
      RECT 73.035 3.04 73.045 3.34 ;
      RECT 73.55 3.212 73.555 3.431 ;
      RECT 73.54 3.192 73.55 3.448 ;
      RECT 73.53 3.172 73.54 3.478 ;
      RECT 73.525 3.162 73.53 3.493 ;
      RECT 73.52 3.158 73.525 3.498 ;
      RECT 73.505 3.15 73.52 3.505 ;
      RECT 73.465 3.13 73.505 3.53 ;
      RECT 73.44 3.112 73.465 3.563 ;
      RECT 73.435 3.11 73.44 3.576 ;
      RECT 73.415 3.107 73.435 3.58 ;
      RECT 73.385 3.105 73.415 3.59 ;
      RECT 73.315 3.107 73.375 3.591 ;
      RECT 73.295 3.107 73.315 3.585 ;
      RECT 73.27 3.105 73.295 3.582 ;
      RECT 73.235 3.1 73.27 3.578 ;
      RECT 73.215 3.094 73.235 3.565 ;
      RECT 73.205 3.091 73.215 3.553 ;
      RECT 73.185 3.088 73.205 3.538 ;
      RECT 73.165 3.084 73.185 3.52 ;
      RECT 73.16 3.081 73.165 3.51 ;
      RECT 73.155 3.08 73.16 3.508 ;
      RECT 73.145 3.077 73.155 3.5 ;
      RECT 73.135 3.071 73.145 3.483 ;
      RECT 73.125 3.065 73.135 3.465 ;
      RECT 73.115 3.059 73.125 3.453 ;
      RECT 73.105 3.053 73.115 3.433 ;
      RECT 73.1 3.049 73.105 3.418 ;
      RECT 73.095 3.047 73.1 3.41 ;
      RECT 73.09 3.045 73.095 3.403 ;
      RECT 73.085 3.043 73.09 3.393 ;
      RECT 73.08 3.041 73.085 3.387 ;
      RECT 73.07 3.04 73.08 3.377 ;
      RECT 73.06 3.04 73.07 3.368 ;
      RECT 73.045 3.04 73.06 3.353 ;
      RECT 73.005 3.04 73.035 3.337 ;
      RECT 72.985 3.042 73.005 3.332 ;
      RECT 72.98 3.047 72.985 3.33 ;
      RECT 72.95 3.055 72.98 3.328 ;
      RECT 72.92 3.07 72.95 3.327 ;
      RECT 72.875 3.092 72.92 3.332 ;
      RECT 72.87 3.107 72.875 3.336 ;
      RECT 72.855 3.112 72.87 3.338 ;
      RECT 72.85 3.116 72.855 3.34 ;
      RECT 72.79 3.139 72.85 3.349 ;
      RECT 72.77 3.165 72.79 3.362 ;
      RECT 72.76 3.172 72.77 3.366 ;
      RECT 72.745 3.179 72.76 3.369 ;
      RECT 72.725 3.189 72.745 3.372 ;
      RECT 72.72 3.197 72.725 3.375 ;
      RECT 72.675 3.202 72.72 3.382 ;
      RECT 72.665 3.205 72.675 3.389 ;
      RECT 72.655 3.205 72.665 3.393 ;
      RECT 72.62 3.207 72.655 3.405 ;
      RECT 72.6 3.21 72.62 3.418 ;
      RECT 72.56 3.213 72.6 3.429 ;
      RECT 72.545 3.215 72.56 3.442 ;
      RECT 72.535 3.215 72.545 3.447 ;
      RECT 72.51 3.216 72.535 3.455 ;
      RECT 72.5 3.218 72.51 3.46 ;
      RECT 72.495 3.219 72.5 3.463 ;
      RECT 72.47 3.217 72.495 3.466 ;
      RECT 72.455 3.215 72.47 3.467 ;
      RECT 72.435 3.212 72.455 3.469 ;
      RECT 72.415 3.207 72.435 3.469 ;
      RECT 72.355 3.202 72.415 3.466 ;
      RECT 72.32 3.177 72.355 3.462 ;
      RECT 72.31 3.154 72.32 3.46 ;
      RECT 72.28 3.131 72.31 3.46 ;
      RECT 72.27 3.11 72.28 3.46 ;
      RECT 72.245 3.092 72.27 3.458 ;
      RECT 72.23 3.07 72.245 3.455 ;
      RECT 72.215 3.052 72.23 3.453 ;
      RECT 72.195 3.042 72.215 3.451 ;
      RECT 72.18 3.037 72.195 3.45 ;
      RECT 72.165 3.035 72.18 3.449 ;
      RECT 72.135 3.036 72.165 3.447 ;
      RECT 72.115 3.039 72.135 3.445 ;
      RECT 72.058 3.043 72.115 3.445 ;
      RECT 71.972 3.052 72.058 3.445 ;
      RECT 71.886 3.063 71.972 3.445 ;
      RECT 71.8 3.074 71.886 3.445 ;
      RECT 71.78 3.081 71.8 3.453 ;
      RECT 71.77 3.084 71.78 3.46 ;
      RECT 71.705 3.089 71.77 3.478 ;
      RECT 71.675 3.096 71.705 3.503 ;
      RECT 71.665 3.099 71.675 3.51 ;
      RECT 71.62 3.103 71.665 3.515 ;
      RECT 71.59 3.108 71.62 3.52 ;
      RECT 71.589 3.11 71.59 3.52 ;
      RECT 71.503 3.116 71.589 3.52 ;
      RECT 71.417 3.127 71.503 3.52 ;
      RECT 71.331 3.139 71.417 3.52 ;
      RECT 71.245 3.15 71.331 3.52 ;
      RECT 71.23 3.157 71.245 3.515 ;
      RECT 71.225 3.159 71.23 3.509 ;
      RECT 71.205 3.17 71.225 3.504 ;
      RECT 71.195 3.188 71.205 3.498 ;
      RECT 71.19 3.2 71.195 3.298 ;
      RECT 73.485 1.953 73.505 2.04 ;
      RECT 73.48 1.888 73.485 2.072 ;
      RECT 73.47 1.855 73.48 2.077 ;
      RECT 73.465 1.835 73.47 2.083 ;
      RECT 73.435 1.835 73.465 2.1 ;
      RECT 73.386 1.835 73.435 2.136 ;
      RECT 73.3 1.835 73.386 2.194 ;
      RECT 73.271 1.845 73.3 2.243 ;
      RECT 73.185 1.887 73.271 2.296 ;
      RECT 73.165 1.925 73.185 2.343 ;
      RECT 73.14 1.942 73.165 2.363 ;
      RECT 73.13 1.956 73.14 2.383 ;
      RECT 73.125 1.962 73.13 2.393 ;
      RECT 73.12 1.966 73.125 2.4 ;
      RECT 73.07 1.986 73.12 2.405 ;
      RECT 73.005 2.03 73.07 2.405 ;
      RECT 72.98 2.08 73.005 2.405 ;
      RECT 72.97 2.11 72.98 2.405 ;
      RECT 72.965 2.137 72.97 2.405 ;
      RECT 72.96 2.155 72.965 2.405 ;
      RECT 72.95 2.197 72.96 2.405 ;
      RECT 73.3 2.755 73.47 2.93 ;
      RECT 73.24 2.583 73.3 2.918 ;
      RECT 73.23 2.576 73.24 2.901 ;
      RECT 73.185 2.755 73.47 2.881 ;
      RECT 73.166 2.755 73.47 2.859 ;
      RECT 73.08 2.755 73.47 2.824 ;
      RECT 73.06 2.575 73.23 2.78 ;
      RECT 73.06 2.722 73.465 2.78 ;
      RECT 73.06 2.67 73.44 2.78 ;
      RECT 73.06 2.625 73.405 2.78 ;
      RECT 73.06 2.607 73.37 2.78 ;
      RECT 73.06 2.597 73.365 2.78 ;
      RECT 73.23 7.855 73.4 8.305 ;
      RECT 73.285 6.075 73.455 8.025 ;
      RECT 73.23 5.015 73.4 6.245 ;
      RECT 72.71 5.015 72.88 8.305 ;
      RECT 72.71 7.315 73.115 7.645 ;
      RECT 72.71 6.475 73.115 6.805 ;
      RECT 72.78 3.555 72.97 3.78 ;
      RECT 72.77 3.556 72.975 3.775 ;
      RECT 72.77 3.558 72.985 3.755 ;
      RECT 72.77 3.562 72.99 3.74 ;
      RECT 72.77 3.549 72.94 3.775 ;
      RECT 72.77 3.552 72.965 3.775 ;
      RECT 72.78 3.548 72.94 3.78 ;
      RECT 72.866 3.546 72.94 3.78 ;
      RECT 72.49 2.797 72.66 3.035 ;
      RECT 72.49 2.797 72.746 2.949 ;
      RECT 72.49 2.797 72.75 2.859 ;
      RECT 72.54 2.57 72.76 2.838 ;
      RECT 72.535 2.587 72.765 2.811 ;
      RECT 72.5 2.745 72.765 2.811 ;
      RECT 72.52 2.595 72.66 3.035 ;
      RECT 72.51 2.677 72.77 2.794 ;
      RECT 72.505 2.725 72.77 2.794 ;
      RECT 72.51 2.635 72.765 2.811 ;
      RECT 72.535 2.572 72.76 2.838 ;
      RECT 72.1 2.547 72.27 2.745 ;
      RECT 72.1 2.547 72.315 2.72 ;
      RECT 72.17 2.49 72.34 2.678 ;
      RECT 72.145 2.505 72.34 2.678 ;
      RECT 71.76 2.551 71.79 2.745 ;
      RECT 71.755 2.523 71.76 2.745 ;
      RECT 71.725 2.497 71.755 2.747 ;
      RECT 71.7 2.455 71.725 2.75 ;
      RECT 71.69 2.427 71.7 2.752 ;
      RECT 71.655 2.407 71.69 2.754 ;
      RECT 71.59 2.392 71.655 2.76 ;
      RECT 71.54 2.39 71.59 2.766 ;
      RECT 71.517 2.392 71.54 2.771 ;
      RECT 71.431 2.403 71.517 2.777 ;
      RECT 71.345 2.421 71.431 2.787 ;
      RECT 71.33 2.432 71.345 2.793 ;
      RECT 71.26 2.455 71.33 2.799 ;
      RECT 71.205 2.487 71.26 2.807 ;
      RECT 71.165 2.51 71.205 2.813 ;
      RECT 71.151 2.523 71.165 2.816 ;
      RECT 71.065 2.545 71.151 2.822 ;
      RECT 71.05 2.57 71.065 2.828 ;
      RECT 71.01 2.585 71.05 2.832 ;
      RECT 70.96 2.6 71.01 2.837 ;
      RECT 70.935 2.607 70.96 2.841 ;
      RECT 70.875 2.602 70.935 2.845 ;
      RECT 70.86 2.593 70.875 2.849 ;
      RECT 70.79 2.583 70.86 2.845 ;
      RECT 70.765 2.575 70.785 2.835 ;
      RECT 70.706 2.575 70.765 2.813 ;
      RECT 70.62 2.575 70.706 2.77 ;
      RECT 70.785 2.575 70.79 2.84 ;
      RECT 71.48 1.806 71.65 2.14 ;
      RECT 71.45 1.806 71.65 2.135 ;
      RECT 71.39 1.773 71.45 2.123 ;
      RECT 71.39 1.829 71.66 2.118 ;
      RECT 71.365 1.829 71.66 2.112 ;
      RECT 71.36 1.77 71.39 2.109 ;
      RECT 71.345 1.776 71.48 2.107 ;
      RECT 71.34 1.784 71.565 2.095 ;
      RECT 71.34 1.836 71.675 2.048 ;
      RECT 71.325 1.792 71.565 2.043 ;
      RECT 71.325 1.862 71.685 1.984 ;
      RECT 71.295 1.812 71.65 1.945 ;
      RECT 71.295 1.902 71.695 1.941 ;
      RECT 71.345 1.781 71.565 2.107 ;
      RECT 70.685 2.111 70.74 2.375 ;
      RECT 70.685 2.111 70.805 2.374 ;
      RECT 70.685 2.111 70.83 2.373 ;
      RECT 70.685 2.111 70.895 2.372 ;
      RECT 70.83 2.077 70.91 2.371 ;
      RECT 70.645 2.121 71.055 2.37 ;
      RECT 70.685 2.118 71.055 2.37 ;
      RECT 70.645 2.126 71.06 2.363 ;
      RECT 70.63 2.128 71.06 2.362 ;
      RECT 70.63 2.135 71.065 2.358 ;
      RECT 70.61 2.134 71.06 2.354 ;
      RECT 70.61 2.142 71.07 2.353 ;
      RECT 70.605 2.139 71.065 2.349 ;
      RECT 70.605 2.152 71.08 2.348 ;
      RECT 70.59 2.142 71.07 2.347 ;
      RECT 70.555 2.155 71.08 2.34 ;
      RECT 70.74 2.11 71.05 2.37 ;
      RECT 70.74 2.095 71 2.37 ;
      RECT 70.805 2.082 70.935 2.37 ;
      RECT 70.35 3.171 70.365 3.564 ;
      RECT 70.315 3.176 70.365 3.563 ;
      RECT 70.35 3.175 70.41 3.562 ;
      RECT 70.295 3.186 70.41 3.561 ;
      RECT 70.31 3.182 70.41 3.561 ;
      RECT 70.275 3.192 70.485 3.558 ;
      RECT 70.275 3.211 70.53 3.556 ;
      RECT 70.275 3.218 70.535 3.553 ;
      RECT 70.26 3.195 70.485 3.55 ;
      RECT 70.24 3.2 70.485 3.543 ;
      RECT 70.235 3.204 70.485 3.539 ;
      RECT 70.235 3.221 70.545 3.538 ;
      RECT 70.215 3.215 70.53 3.534 ;
      RECT 70.215 3.224 70.55 3.528 ;
      RECT 70.21 3.23 70.55 3.3 ;
      RECT 70.275 3.19 70.41 3.558 ;
      RECT 70.15 2.553 70.35 2.865 ;
      RECT 70.225 2.531 70.35 2.865 ;
      RECT 70.165 2.55 70.355 2.85 ;
      RECT 70.135 2.561 70.355 2.848 ;
      RECT 70.15 2.556 70.36 2.814 ;
      RECT 70.135 2.66 70.365 2.781 ;
      RECT 70.165 2.532 70.35 2.865 ;
      RECT 70.225 2.51 70.325 2.865 ;
      RECT 70.25 2.507 70.325 2.865 ;
      RECT 70.25 2.502 70.27 2.865 ;
      RECT 69.655 2.57 69.83 2.745 ;
      RECT 69.65 2.57 69.83 2.743 ;
      RECT 69.625 2.57 69.83 2.738 ;
      RECT 69.57 2.55 69.74 2.728 ;
      RECT 69.57 2.557 69.805 2.728 ;
      RECT 69.655 3.237 69.67 3.42 ;
      RECT 69.645 3.215 69.655 3.42 ;
      RECT 69.63 3.195 69.645 3.42 ;
      RECT 69.62 3.17 69.63 3.42 ;
      RECT 69.59 3.135 69.62 3.42 ;
      RECT 69.555 3.075 69.59 3.42 ;
      RECT 69.55 3.037 69.555 3.42 ;
      RECT 69.5 2.988 69.55 3.42 ;
      RECT 69.49 2.938 69.5 3.408 ;
      RECT 69.475 2.917 69.49 3.368 ;
      RECT 69.455 2.885 69.475 3.318 ;
      RECT 69.43 2.841 69.455 3.258 ;
      RECT 69.425 2.813 69.43 3.213 ;
      RECT 69.42 2.804 69.425 3.199 ;
      RECT 69.415 2.797 69.42 3.186 ;
      RECT 69.41 2.792 69.415 3.175 ;
      RECT 69.405 2.777 69.41 3.165 ;
      RECT 69.4 2.755 69.405 3.152 ;
      RECT 69.39 2.715 69.4 3.127 ;
      RECT 69.365 2.645 69.39 3.083 ;
      RECT 69.36 2.585 69.365 3.048 ;
      RECT 69.345 2.565 69.36 3.015 ;
      RECT 69.34 2.565 69.345 2.99 ;
      RECT 69.31 2.565 69.34 2.945 ;
      RECT 69.265 2.565 69.31 2.885 ;
      RECT 69.19 2.565 69.265 2.833 ;
      RECT 69.185 2.565 69.19 2.798 ;
      RECT 69.18 2.565 69.185 2.788 ;
      RECT 69.175 2.565 69.18 2.768 ;
      RECT 69.44 1.785 69.61 2.255 ;
      RECT 69.385 1.778 69.58 2.239 ;
      RECT 69.385 1.792 69.615 2.238 ;
      RECT 69.37 1.793 69.615 2.219 ;
      RECT 69.365 1.811 69.615 2.205 ;
      RECT 69.37 1.794 69.62 2.203 ;
      RECT 69.355 1.825 69.62 2.188 ;
      RECT 69.37 1.8 69.625 2.173 ;
      RECT 69.35 1.84 69.625 2.17 ;
      RECT 69.365 1.812 69.63 2.155 ;
      RECT 69.365 1.824 69.635 2.135 ;
      RECT 69.35 1.84 69.64 2.118 ;
      RECT 69.35 1.85 69.645 1.973 ;
      RECT 69.345 1.85 69.645 1.93 ;
      RECT 69.345 1.865 69.65 1.908 ;
      RECT 69.44 1.775 69.58 2.255 ;
      RECT 69.44 1.773 69.55 2.255 ;
      RECT 69.526 1.77 69.55 2.255 ;
      RECT 69.185 3.437 69.19 3.483 ;
      RECT 69.175 3.285 69.185 3.507 ;
      RECT 69.17 3.13 69.175 3.532 ;
      RECT 69.155 3.092 69.17 3.543 ;
      RECT 69.15 3.075 69.155 3.55 ;
      RECT 69.14 3.063 69.15 3.557 ;
      RECT 69.135 3.054 69.14 3.559 ;
      RECT 69.13 3.052 69.135 3.563 ;
      RECT 69.085 3.043 69.13 3.578 ;
      RECT 69.08 3.035 69.085 3.592 ;
      RECT 69.075 3.032 69.08 3.596 ;
      RECT 69.06 3.027 69.075 3.604 ;
      RECT 69.005 3.017 69.06 3.615 ;
      RECT 68.97 3.005 69.005 3.616 ;
      RECT 68.961 3 68.97 3.61 ;
      RECT 68.875 3 68.961 3.6 ;
      RECT 68.845 3 68.875 3.578 ;
      RECT 68.835 3 68.84 3.558 ;
      RECT 68.83 3 68.835 3.52 ;
      RECT 68.825 3 68.83 3.478 ;
      RECT 68.82 3 68.825 3.438 ;
      RECT 68.815 3 68.82 3.368 ;
      RECT 68.805 3 68.815 3.29 ;
      RECT 68.8 3 68.805 3.19 ;
      RECT 68.84 3 68.845 3.56 ;
      RECT 68.335 3.082 68.425 3.56 ;
      RECT 68.32 3.085 68.44 3.558 ;
      RECT 68.335 3.084 68.44 3.558 ;
      RECT 68.3 3.091 68.465 3.548 ;
      RECT 68.32 3.085 68.465 3.548 ;
      RECT 68.285 3.097 68.465 3.536 ;
      RECT 68.32 3.088 68.515 3.529 ;
      RECT 68.271 3.105 68.515 3.527 ;
      RECT 68.3 3.095 68.525 3.515 ;
      RECT 68.271 3.116 68.555 3.506 ;
      RECT 68.185 3.14 68.555 3.5 ;
      RECT 68.185 3.153 68.595 3.483 ;
      RECT 68.18 3.175 68.595 3.476 ;
      RECT 68.15 3.19 68.595 3.466 ;
      RECT 68.145 3.201 68.595 3.456 ;
      RECT 68.115 3.214 68.595 3.447 ;
      RECT 68.1 3.232 68.595 3.436 ;
      RECT 68.075 3.245 68.595 3.426 ;
      RECT 68.335 3.081 68.345 3.56 ;
      RECT 68.381 2.505 68.42 2.75 ;
      RECT 68.295 2.505 68.43 2.748 ;
      RECT 68.18 2.53 68.43 2.745 ;
      RECT 68.18 2.53 68.435 2.743 ;
      RECT 68.18 2.53 68.45 2.738 ;
      RECT 68.286 2.505 68.465 2.718 ;
      RECT 68.2 2.513 68.465 2.718 ;
      RECT 67.87 1.865 68.04 2.3 ;
      RECT 67.86 1.899 68.04 2.283 ;
      RECT 67.94 1.835 68.11 2.27 ;
      RECT 67.845 1.91 68.11 2.248 ;
      RECT 67.94 1.845 68.115 2.238 ;
      RECT 67.87 1.897 68.145 2.223 ;
      RECT 67.83 1.923 68.145 2.208 ;
      RECT 67.83 1.965 68.155 2.188 ;
      RECT 67.825 1.99 68.16 2.17 ;
      RECT 67.825 2 68.165 2.155 ;
      RECT 67.82 1.937 68.145 2.153 ;
      RECT 67.82 2.01 68.17 2.138 ;
      RECT 67.815 1.947 68.145 2.135 ;
      RECT 67.81 2.031 68.175 2.118 ;
      RECT 67.81 2.063 68.18 2.098 ;
      RECT 67.805 1.977 68.155 2.09 ;
      RECT 67.81 1.962 68.145 2.118 ;
      RECT 67.825 1.932 68.145 2.17 ;
      RECT 67.67 2.519 67.895 2.775 ;
      RECT 67.67 2.552 67.915 2.765 ;
      RECT 67.635 2.552 67.915 2.763 ;
      RECT 67.635 2.565 67.92 2.753 ;
      RECT 67.635 2.585 67.93 2.745 ;
      RECT 67.635 2.682 67.935 2.738 ;
      RECT 67.615 2.43 67.745 2.728 ;
      RECT 67.57 2.585 67.93 2.67 ;
      RECT 67.56 2.43 67.745 2.615 ;
      RECT 67.56 2.462 67.831 2.615 ;
      RECT 67.525 2.992 67.545 3.17 ;
      RECT 67.49 2.945 67.525 3.17 ;
      RECT 67.475 2.885 67.49 3.17 ;
      RECT 67.45 2.832 67.475 3.17 ;
      RECT 67.435 2.785 67.45 3.17 ;
      RECT 67.415 2.762 67.435 3.17 ;
      RECT 67.39 2.727 67.415 3.17 ;
      RECT 67.38 2.573 67.39 3.17 ;
      RECT 67.35 2.568 67.38 3.161 ;
      RECT 67.345 2.565 67.35 3.151 ;
      RECT 67.33 2.565 67.345 3.125 ;
      RECT 67.325 2.565 67.33 3.088 ;
      RECT 67.3 2.565 67.325 3.04 ;
      RECT 67.28 2.565 67.3 2.965 ;
      RECT 67.27 2.565 67.28 2.925 ;
      RECT 67.265 2.565 67.27 2.9 ;
      RECT 67.26 2.565 67.265 2.883 ;
      RECT 67.255 2.565 67.26 2.865 ;
      RECT 67.25 2.566 67.255 2.855 ;
      RECT 67.24 2.568 67.25 2.823 ;
      RECT 67.23 2.57 67.24 2.79 ;
      RECT 67.22 2.573 67.23 2.763 ;
      RECT 67.545 3 67.77 3.17 ;
      RECT 66.875 1.812 67.045 2.265 ;
      RECT 66.875 1.812 67.135 2.231 ;
      RECT 66.875 1.812 67.165 2.215 ;
      RECT 66.875 1.812 67.195 2.188 ;
      RECT 67.131 1.79 67.21 2.17 ;
      RECT 66.91 1.797 67.215 2.155 ;
      RECT 66.91 1.805 67.225 2.118 ;
      RECT 66.87 1.832 67.225 2.09 ;
      RECT 66.855 1.845 67.225 2.055 ;
      RECT 66.875 1.82 67.245 2.045 ;
      RECT 66.85 1.885 67.245 2.015 ;
      RECT 66.85 1.915 67.25 1.998 ;
      RECT 66.845 1.945 67.25 1.985 ;
      RECT 66.91 1.794 67.21 2.17 ;
      RECT 67.045 1.791 67.131 2.249 ;
      RECT 66.996 1.792 67.21 2.17 ;
      RECT 67.14 3.452 67.185 3.645 ;
      RECT 67.13 3.422 67.14 3.645 ;
      RECT 67.125 3.407 67.13 3.645 ;
      RECT 67.085 3.317 67.125 3.645 ;
      RECT 67.08 3.23 67.085 3.645 ;
      RECT 67.07 3.2 67.08 3.645 ;
      RECT 67.065 3.16 67.07 3.645 ;
      RECT 67.055 3.122 67.065 3.645 ;
      RECT 67.05 3.087 67.055 3.645 ;
      RECT 67.03 3.04 67.05 3.645 ;
      RECT 67.015 2.965 67.03 3.645 ;
      RECT 67.01 2.92 67.015 3.64 ;
      RECT 67.005 2.9 67.01 3.613 ;
      RECT 67 2.88 67.005 3.598 ;
      RECT 66.995 2.855 67 3.578 ;
      RECT 66.99 2.833 66.995 3.563 ;
      RECT 66.985 2.811 66.99 3.545 ;
      RECT 66.98 2.79 66.985 3.535 ;
      RECT 66.97 2.762 66.98 3.505 ;
      RECT 66.96 2.725 66.97 3.473 ;
      RECT 66.95 2.685 66.96 3.44 ;
      RECT 66.94 2.663 66.95 3.41 ;
      RECT 66.91 2.615 66.94 3.342 ;
      RECT 66.895 2.575 66.91 3.269 ;
      RECT 66.885 2.575 66.895 3.235 ;
      RECT 66.88 2.575 66.885 3.21 ;
      RECT 66.875 2.575 66.88 3.195 ;
      RECT 66.87 2.575 66.875 3.173 ;
      RECT 66.865 2.575 66.87 3.16 ;
      RECT 66.85 2.575 66.865 3.125 ;
      RECT 66.83 2.575 66.85 3.065 ;
      RECT 66.82 2.575 66.83 3.015 ;
      RECT 66.8 2.575 66.82 2.963 ;
      RECT 66.78 2.575 66.8 2.92 ;
      RECT 66.77 2.575 66.78 2.908 ;
      RECT 66.74 2.575 66.77 2.895 ;
      RECT 66.71 2.596 66.74 2.875 ;
      RECT 66.7 2.624 66.71 2.855 ;
      RECT 66.685 2.641 66.7 2.823 ;
      RECT 66.68 2.655 66.685 2.79 ;
      RECT 66.675 2.663 66.68 2.763 ;
      RECT 66.67 2.671 66.675 2.725 ;
      RECT 66.675 3.195 66.68 3.53 ;
      RECT 66.64 3.182 66.675 3.529 ;
      RECT 66.57 3.122 66.64 3.528 ;
      RECT 66.49 3.065 66.57 3.527 ;
      RECT 66.355 3.025 66.49 3.526 ;
      RECT 66.355 3.212 66.69 3.515 ;
      RECT 66.315 3.212 66.69 3.505 ;
      RECT 66.315 3.23 66.695 3.5 ;
      RECT 66.315 3.32 66.7 3.49 ;
      RECT 66.31 3.015 66.475 3.47 ;
      RECT 66.305 3.015 66.475 3.213 ;
      RECT 66.305 3.172 66.67 3.213 ;
      RECT 66.305 3.16 66.665 3.213 ;
      RECT 65.435 5.02 65.605 6.49 ;
      RECT 65.435 6.315 65.61 6.485 ;
      RECT 65.065 1.74 65.235 2.93 ;
      RECT 65.065 1.74 65.535 1.91 ;
      RECT 65.065 6.97 65.535 7.14 ;
      RECT 65.065 5.95 65.235 7.14 ;
      RECT 64.075 1.74 64.245 2.93 ;
      RECT 64.075 1.74 64.545 1.91 ;
      RECT 64.075 6.97 64.545 7.14 ;
      RECT 64.075 5.95 64.245 7.14 ;
      RECT 62.225 2.635 62.395 3.865 ;
      RECT 62.28 0.855 62.45 2.805 ;
      RECT 62.225 0.575 62.395 1.025 ;
      RECT 62.225 7.855 62.395 8.305 ;
      RECT 62.28 6.075 62.45 8.025 ;
      RECT 62.225 5.015 62.395 6.245 ;
      RECT 61.705 0.575 61.875 3.865 ;
      RECT 61.705 2.075 62.11 2.405 ;
      RECT 61.705 1.235 62.11 1.565 ;
      RECT 61.705 5.015 61.875 8.305 ;
      RECT 61.705 7.315 62.11 7.645 ;
      RECT 61.705 6.475 62.11 6.805 ;
      RECT 59.04 1.975 59.77 2.215 ;
      RECT 59.582 1.77 59.77 2.215 ;
      RECT 59.41 1.782 59.785 2.209 ;
      RECT 59.325 1.797 59.805 2.194 ;
      RECT 59.325 1.812 59.81 2.184 ;
      RECT 59.28 1.832 59.825 2.176 ;
      RECT 59.257 1.867 59.84 2.13 ;
      RECT 59.171 1.89 59.845 2.09 ;
      RECT 59.171 1.908 59.855 2.06 ;
      RECT 59.04 1.977 59.86 2.023 ;
      RECT 59.085 1.92 59.855 2.06 ;
      RECT 59.171 1.872 59.84 2.13 ;
      RECT 59.257 1.841 59.825 2.176 ;
      RECT 59.28 1.822 59.81 2.184 ;
      RECT 59.325 1.795 59.785 2.209 ;
      RECT 59.41 1.777 59.77 2.215 ;
      RECT 59.496 1.771 59.77 2.215 ;
      RECT 59.582 1.766 59.715 2.215 ;
      RECT 59.668 1.761 59.715 2.215 ;
      RECT 59.36 2.659 59.53 3.045 ;
      RECT 59.355 2.659 59.53 3.04 ;
      RECT 59.33 2.659 59.53 3.005 ;
      RECT 59.33 2.687 59.54 2.995 ;
      RECT 59.31 2.687 59.54 2.955 ;
      RECT 59.305 2.687 59.54 2.928 ;
      RECT 59.305 2.705 59.545 2.92 ;
      RECT 59.25 2.705 59.545 2.855 ;
      RECT 59.25 2.722 59.555 2.838 ;
      RECT 59.24 2.722 59.555 2.778 ;
      RECT 59.24 2.739 59.56 2.775 ;
      RECT 59.235 2.575 59.405 2.753 ;
      RECT 59.235 2.609 59.491 2.753 ;
      RECT 59.23 3.375 59.235 3.388 ;
      RECT 59.225 3.27 59.23 3.393 ;
      RECT 59.2 3.13 59.225 3.408 ;
      RECT 59.165 3.081 59.2 3.44 ;
      RECT 59.16 3.049 59.165 3.46 ;
      RECT 59.155 3.04 59.16 3.46 ;
      RECT 59.075 3.005 59.155 3.46 ;
      RECT 59.012 2.975 59.075 3.46 ;
      RECT 58.926 2.963 59.012 3.46 ;
      RECT 58.84 2.949 58.926 3.46 ;
      RECT 58.76 2.936 58.84 3.446 ;
      RECT 58.725 2.928 58.76 3.426 ;
      RECT 58.715 2.925 58.725 3.417 ;
      RECT 58.685 2.92 58.715 3.404 ;
      RECT 58.635 2.895 58.685 3.38 ;
      RECT 58.621 2.869 58.635 3.362 ;
      RECT 58.535 2.829 58.621 3.338 ;
      RECT 58.49 2.777 58.535 3.307 ;
      RECT 58.48 2.752 58.49 3.294 ;
      RECT 58.475 2.533 58.48 2.555 ;
      RECT 58.47 2.735 58.48 3.29 ;
      RECT 58.47 2.531 58.475 2.645 ;
      RECT 58.46 2.527 58.47 3.286 ;
      RECT 58.416 2.525 58.46 3.274 ;
      RECT 58.33 2.525 58.416 3.245 ;
      RECT 58.3 2.525 58.33 3.218 ;
      RECT 58.285 2.525 58.3 3.206 ;
      RECT 58.245 2.537 58.285 3.191 ;
      RECT 58.225 2.556 58.245 3.17 ;
      RECT 58.215 2.566 58.225 3.154 ;
      RECT 58.205 2.572 58.215 3.143 ;
      RECT 58.185 2.582 58.205 3.126 ;
      RECT 58.18 2.591 58.185 3.113 ;
      RECT 58.175 2.595 58.18 3.063 ;
      RECT 58.165 2.601 58.175 2.98 ;
      RECT 58.16 2.605 58.165 2.894 ;
      RECT 58.155 2.625 58.16 2.831 ;
      RECT 58.15 2.648 58.155 2.778 ;
      RECT 58.145 2.666 58.15 2.723 ;
      RECT 58.755 2.485 58.925 2.745 ;
      RECT 58.925 2.45 58.97 2.731 ;
      RECT 58.886 2.452 58.975 2.714 ;
      RECT 58.775 2.469 59.061 2.685 ;
      RECT 58.775 2.484 59.065 2.657 ;
      RECT 58.775 2.465 58.975 2.714 ;
      RECT 58.8 2.453 58.925 2.745 ;
      RECT 58.886 2.451 58.97 2.731 ;
      RECT 57.94 1.84 58.11 2.33 ;
      RECT 57.94 1.84 58.145 2.31 ;
      RECT 58.075 1.76 58.185 2.27 ;
      RECT 58.056 1.764 58.205 2.24 ;
      RECT 57.97 1.772 58.225 2.223 ;
      RECT 57.97 1.778 58.23 2.213 ;
      RECT 57.97 1.787 58.25 2.201 ;
      RECT 57.945 1.812 58.28 2.179 ;
      RECT 57.945 1.832 58.285 2.159 ;
      RECT 57.94 1.845 58.295 2.139 ;
      RECT 57.94 1.912 58.3 2.12 ;
      RECT 57.94 2.045 58.305 2.107 ;
      RECT 57.935 1.85 58.295 1.94 ;
      RECT 57.945 1.807 58.25 2.201 ;
      RECT 58.056 1.762 58.185 2.27 ;
      RECT 57.93 3.515 58.23 3.77 ;
      RECT 58.015 3.481 58.23 3.77 ;
      RECT 58.015 3.484 58.235 3.63 ;
      RECT 57.95 3.505 58.235 3.63 ;
      RECT 57.985 3.495 58.23 3.77 ;
      RECT 57.98 3.5 58.235 3.63 ;
      RECT 58.015 3.479 58.216 3.77 ;
      RECT 58.101 3.47 58.216 3.77 ;
      RECT 58.101 3.464 58.13 3.77 ;
      RECT 57.59 3.105 57.6 3.595 ;
      RECT 57.25 3.04 57.26 3.34 ;
      RECT 57.765 3.212 57.77 3.431 ;
      RECT 57.755 3.192 57.765 3.448 ;
      RECT 57.745 3.172 57.755 3.478 ;
      RECT 57.74 3.162 57.745 3.493 ;
      RECT 57.735 3.158 57.74 3.498 ;
      RECT 57.72 3.15 57.735 3.505 ;
      RECT 57.68 3.13 57.72 3.53 ;
      RECT 57.655 3.112 57.68 3.563 ;
      RECT 57.65 3.11 57.655 3.576 ;
      RECT 57.63 3.107 57.65 3.58 ;
      RECT 57.6 3.105 57.63 3.59 ;
      RECT 57.53 3.107 57.59 3.591 ;
      RECT 57.51 3.107 57.53 3.585 ;
      RECT 57.485 3.105 57.51 3.582 ;
      RECT 57.45 3.1 57.485 3.578 ;
      RECT 57.43 3.094 57.45 3.565 ;
      RECT 57.42 3.091 57.43 3.553 ;
      RECT 57.4 3.088 57.42 3.538 ;
      RECT 57.38 3.084 57.4 3.52 ;
      RECT 57.375 3.081 57.38 3.51 ;
      RECT 57.37 3.08 57.375 3.508 ;
      RECT 57.36 3.077 57.37 3.5 ;
      RECT 57.35 3.071 57.36 3.483 ;
      RECT 57.34 3.065 57.35 3.465 ;
      RECT 57.33 3.059 57.34 3.453 ;
      RECT 57.32 3.053 57.33 3.433 ;
      RECT 57.315 3.049 57.32 3.418 ;
      RECT 57.31 3.047 57.315 3.41 ;
      RECT 57.305 3.045 57.31 3.403 ;
      RECT 57.3 3.043 57.305 3.393 ;
      RECT 57.295 3.041 57.3 3.387 ;
      RECT 57.285 3.04 57.295 3.377 ;
      RECT 57.275 3.04 57.285 3.368 ;
      RECT 57.26 3.04 57.275 3.353 ;
      RECT 57.22 3.04 57.25 3.337 ;
      RECT 57.2 3.042 57.22 3.332 ;
      RECT 57.195 3.047 57.2 3.33 ;
      RECT 57.165 3.055 57.195 3.328 ;
      RECT 57.135 3.07 57.165 3.327 ;
      RECT 57.09 3.092 57.135 3.332 ;
      RECT 57.085 3.107 57.09 3.336 ;
      RECT 57.07 3.112 57.085 3.338 ;
      RECT 57.065 3.116 57.07 3.34 ;
      RECT 57.005 3.139 57.065 3.349 ;
      RECT 56.985 3.165 57.005 3.362 ;
      RECT 56.975 3.172 56.985 3.366 ;
      RECT 56.96 3.179 56.975 3.369 ;
      RECT 56.94 3.189 56.96 3.372 ;
      RECT 56.935 3.197 56.94 3.375 ;
      RECT 56.89 3.202 56.935 3.382 ;
      RECT 56.88 3.205 56.89 3.389 ;
      RECT 56.87 3.205 56.88 3.393 ;
      RECT 56.835 3.207 56.87 3.405 ;
      RECT 56.815 3.21 56.835 3.418 ;
      RECT 56.775 3.213 56.815 3.429 ;
      RECT 56.76 3.215 56.775 3.442 ;
      RECT 56.75 3.215 56.76 3.447 ;
      RECT 56.725 3.216 56.75 3.455 ;
      RECT 56.715 3.218 56.725 3.46 ;
      RECT 56.71 3.219 56.715 3.463 ;
      RECT 56.685 3.217 56.71 3.466 ;
      RECT 56.67 3.215 56.685 3.467 ;
      RECT 56.65 3.212 56.67 3.469 ;
      RECT 56.63 3.207 56.65 3.469 ;
      RECT 56.57 3.202 56.63 3.466 ;
      RECT 56.535 3.177 56.57 3.462 ;
      RECT 56.525 3.154 56.535 3.46 ;
      RECT 56.495 3.131 56.525 3.46 ;
      RECT 56.485 3.11 56.495 3.46 ;
      RECT 56.46 3.092 56.485 3.458 ;
      RECT 56.445 3.07 56.46 3.455 ;
      RECT 56.43 3.052 56.445 3.453 ;
      RECT 56.41 3.042 56.43 3.451 ;
      RECT 56.395 3.037 56.41 3.45 ;
      RECT 56.38 3.035 56.395 3.449 ;
      RECT 56.35 3.036 56.38 3.447 ;
      RECT 56.33 3.039 56.35 3.445 ;
      RECT 56.273 3.043 56.33 3.445 ;
      RECT 56.187 3.052 56.273 3.445 ;
      RECT 56.101 3.063 56.187 3.445 ;
      RECT 56.015 3.074 56.101 3.445 ;
      RECT 55.995 3.081 56.015 3.453 ;
      RECT 55.985 3.084 55.995 3.46 ;
      RECT 55.92 3.089 55.985 3.478 ;
      RECT 55.89 3.096 55.92 3.503 ;
      RECT 55.88 3.099 55.89 3.51 ;
      RECT 55.835 3.103 55.88 3.515 ;
      RECT 55.805 3.108 55.835 3.52 ;
      RECT 55.804 3.11 55.805 3.52 ;
      RECT 55.718 3.116 55.804 3.52 ;
      RECT 55.632 3.127 55.718 3.52 ;
      RECT 55.546 3.139 55.632 3.52 ;
      RECT 55.46 3.15 55.546 3.52 ;
      RECT 55.445 3.157 55.46 3.515 ;
      RECT 55.44 3.159 55.445 3.509 ;
      RECT 55.42 3.17 55.44 3.504 ;
      RECT 55.41 3.188 55.42 3.498 ;
      RECT 55.405 3.2 55.41 3.298 ;
      RECT 57.7 1.953 57.72 2.04 ;
      RECT 57.695 1.888 57.7 2.072 ;
      RECT 57.685 1.855 57.695 2.077 ;
      RECT 57.68 1.835 57.685 2.083 ;
      RECT 57.65 1.835 57.68 2.1 ;
      RECT 57.601 1.835 57.65 2.136 ;
      RECT 57.515 1.835 57.601 2.194 ;
      RECT 57.486 1.845 57.515 2.243 ;
      RECT 57.4 1.887 57.486 2.296 ;
      RECT 57.38 1.925 57.4 2.343 ;
      RECT 57.355 1.942 57.38 2.363 ;
      RECT 57.345 1.956 57.355 2.383 ;
      RECT 57.34 1.962 57.345 2.393 ;
      RECT 57.335 1.966 57.34 2.4 ;
      RECT 57.285 1.986 57.335 2.405 ;
      RECT 57.22 2.03 57.285 2.405 ;
      RECT 57.195 2.08 57.22 2.405 ;
      RECT 57.185 2.11 57.195 2.405 ;
      RECT 57.18 2.137 57.185 2.405 ;
      RECT 57.175 2.155 57.18 2.405 ;
      RECT 57.165 2.197 57.175 2.405 ;
      RECT 57.515 2.755 57.685 2.93 ;
      RECT 57.455 2.583 57.515 2.918 ;
      RECT 57.445 2.576 57.455 2.901 ;
      RECT 57.4 2.755 57.685 2.881 ;
      RECT 57.381 2.755 57.685 2.859 ;
      RECT 57.295 2.755 57.685 2.824 ;
      RECT 57.275 2.575 57.445 2.78 ;
      RECT 57.275 2.722 57.68 2.78 ;
      RECT 57.275 2.67 57.655 2.78 ;
      RECT 57.275 2.625 57.62 2.78 ;
      RECT 57.275 2.607 57.585 2.78 ;
      RECT 57.275 2.597 57.58 2.78 ;
      RECT 57.445 7.855 57.615 8.305 ;
      RECT 57.5 6.075 57.67 8.025 ;
      RECT 57.445 5.015 57.615 6.245 ;
      RECT 56.925 5.015 57.095 8.305 ;
      RECT 56.925 7.315 57.33 7.645 ;
      RECT 56.925 6.475 57.33 6.805 ;
      RECT 56.995 3.555 57.185 3.78 ;
      RECT 56.985 3.556 57.19 3.775 ;
      RECT 56.985 3.558 57.2 3.755 ;
      RECT 56.985 3.562 57.205 3.74 ;
      RECT 56.985 3.549 57.155 3.775 ;
      RECT 56.985 3.552 57.18 3.775 ;
      RECT 56.995 3.548 57.155 3.78 ;
      RECT 57.081 3.546 57.155 3.78 ;
      RECT 56.705 2.797 56.875 3.035 ;
      RECT 56.705 2.797 56.961 2.949 ;
      RECT 56.705 2.797 56.965 2.859 ;
      RECT 56.755 2.57 56.975 2.838 ;
      RECT 56.75 2.587 56.98 2.811 ;
      RECT 56.715 2.745 56.98 2.811 ;
      RECT 56.735 2.595 56.875 3.035 ;
      RECT 56.725 2.677 56.985 2.794 ;
      RECT 56.72 2.725 56.985 2.794 ;
      RECT 56.725 2.635 56.98 2.811 ;
      RECT 56.75 2.572 56.975 2.838 ;
      RECT 56.315 2.547 56.485 2.745 ;
      RECT 56.315 2.547 56.53 2.72 ;
      RECT 56.385 2.49 56.555 2.678 ;
      RECT 56.36 2.505 56.555 2.678 ;
      RECT 55.975 2.551 56.005 2.745 ;
      RECT 55.97 2.523 55.975 2.745 ;
      RECT 55.94 2.497 55.97 2.747 ;
      RECT 55.915 2.455 55.94 2.75 ;
      RECT 55.905 2.427 55.915 2.752 ;
      RECT 55.87 2.407 55.905 2.754 ;
      RECT 55.805 2.392 55.87 2.76 ;
      RECT 55.755 2.39 55.805 2.766 ;
      RECT 55.732 2.392 55.755 2.771 ;
      RECT 55.646 2.403 55.732 2.777 ;
      RECT 55.56 2.421 55.646 2.787 ;
      RECT 55.545 2.432 55.56 2.793 ;
      RECT 55.475 2.455 55.545 2.799 ;
      RECT 55.42 2.487 55.475 2.807 ;
      RECT 55.38 2.51 55.42 2.813 ;
      RECT 55.366 2.523 55.38 2.816 ;
      RECT 55.28 2.545 55.366 2.822 ;
      RECT 55.265 2.57 55.28 2.828 ;
      RECT 55.225 2.585 55.265 2.832 ;
      RECT 55.175 2.6 55.225 2.837 ;
      RECT 55.15 2.607 55.175 2.841 ;
      RECT 55.09 2.602 55.15 2.845 ;
      RECT 55.075 2.593 55.09 2.849 ;
      RECT 55.005 2.583 55.075 2.845 ;
      RECT 54.98 2.575 55 2.835 ;
      RECT 54.921 2.575 54.98 2.813 ;
      RECT 54.835 2.575 54.921 2.77 ;
      RECT 55 2.575 55.005 2.84 ;
      RECT 55.695 1.806 55.865 2.14 ;
      RECT 55.665 1.806 55.865 2.135 ;
      RECT 55.605 1.773 55.665 2.123 ;
      RECT 55.605 1.829 55.875 2.118 ;
      RECT 55.58 1.829 55.875 2.112 ;
      RECT 55.575 1.77 55.605 2.109 ;
      RECT 55.56 1.776 55.695 2.107 ;
      RECT 55.555 1.784 55.78 2.095 ;
      RECT 55.555 1.836 55.89 2.048 ;
      RECT 55.54 1.792 55.78 2.043 ;
      RECT 55.54 1.862 55.9 1.984 ;
      RECT 55.51 1.812 55.865 1.945 ;
      RECT 55.51 1.902 55.91 1.941 ;
      RECT 55.56 1.781 55.78 2.107 ;
      RECT 54.9 2.111 54.955 2.375 ;
      RECT 54.9 2.111 55.02 2.374 ;
      RECT 54.9 2.111 55.045 2.373 ;
      RECT 54.9 2.111 55.11 2.372 ;
      RECT 55.045 2.077 55.125 2.371 ;
      RECT 54.86 2.121 55.27 2.37 ;
      RECT 54.9 2.118 55.27 2.37 ;
      RECT 54.86 2.126 55.275 2.363 ;
      RECT 54.845 2.128 55.275 2.362 ;
      RECT 54.845 2.135 55.28 2.358 ;
      RECT 54.825 2.134 55.275 2.354 ;
      RECT 54.825 2.142 55.285 2.353 ;
      RECT 54.82 2.139 55.28 2.349 ;
      RECT 54.82 2.152 55.295 2.348 ;
      RECT 54.805 2.142 55.285 2.347 ;
      RECT 54.77 2.155 55.295 2.34 ;
      RECT 54.955 2.11 55.265 2.37 ;
      RECT 54.955 2.095 55.215 2.37 ;
      RECT 55.02 2.082 55.15 2.37 ;
      RECT 54.565 3.171 54.58 3.564 ;
      RECT 54.53 3.176 54.58 3.563 ;
      RECT 54.565 3.175 54.625 3.562 ;
      RECT 54.51 3.186 54.625 3.561 ;
      RECT 54.525 3.182 54.625 3.561 ;
      RECT 54.49 3.192 54.7 3.558 ;
      RECT 54.49 3.211 54.745 3.556 ;
      RECT 54.49 3.218 54.75 3.553 ;
      RECT 54.475 3.195 54.7 3.55 ;
      RECT 54.455 3.2 54.7 3.543 ;
      RECT 54.45 3.204 54.7 3.539 ;
      RECT 54.45 3.221 54.76 3.538 ;
      RECT 54.43 3.215 54.745 3.534 ;
      RECT 54.43 3.224 54.765 3.528 ;
      RECT 54.425 3.23 54.765 3.3 ;
      RECT 54.49 3.19 54.625 3.558 ;
      RECT 54.365 2.553 54.565 2.865 ;
      RECT 54.44 2.531 54.565 2.865 ;
      RECT 54.38 2.55 54.57 2.85 ;
      RECT 54.35 2.561 54.57 2.848 ;
      RECT 54.365 2.556 54.575 2.814 ;
      RECT 54.35 2.66 54.58 2.781 ;
      RECT 54.38 2.532 54.565 2.865 ;
      RECT 54.44 2.51 54.54 2.865 ;
      RECT 54.465 2.507 54.54 2.865 ;
      RECT 54.465 2.502 54.485 2.865 ;
      RECT 53.87 2.57 54.045 2.745 ;
      RECT 53.865 2.57 54.045 2.743 ;
      RECT 53.84 2.57 54.045 2.738 ;
      RECT 53.785 2.55 53.955 2.728 ;
      RECT 53.785 2.557 54.02 2.728 ;
      RECT 53.87 3.237 53.885 3.42 ;
      RECT 53.86 3.215 53.87 3.42 ;
      RECT 53.845 3.195 53.86 3.42 ;
      RECT 53.835 3.17 53.845 3.42 ;
      RECT 53.805 3.135 53.835 3.42 ;
      RECT 53.77 3.075 53.805 3.42 ;
      RECT 53.765 3.037 53.77 3.42 ;
      RECT 53.715 2.988 53.765 3.42 ;
      RECT 53.705 2.938 53.715 3.408 ;
      RECT 53.69 2.917 53.705 3.368 ;
      RECT 53.67 2.885 53.69 3.318 ;
      RECT 53.645 2.841 53.67 3.258 ;
      RECT 53.64 2.813 53.645 3.213 ;
      RECT 53.635 2.804 53.64 3.199 ;
      RECT 53.63 2.797 53.635 3.186 ;
      RECT 53.625 2.792 53.63 3.175 ;
      RECT 53.62 2.777 53.625 3.165 ;
      RECT 53.615 2.755 53.62 3.152 ;
      RECT 53.605 2.715 53.615 3.127 ;
      RECT 53.58 2.645 53.605 3.083 ;
      RECT 53.575 2.585 53.58 3.048 ;
      RECT 53.56 2.565 53.575 3.015 ;
      RECT 53.555 2.565 53.56 2.99 ;
      RECT 53.525 2.565 53.555 2.945 ;
      RECT 53.48 2.565 53.525 2.885 ;
      RECT 53.405 2.565 53.48 2.833 ;
      RECT 53.4 2.565 53.405 2.798 ;
      RECT 53.395 2.565 53.4 2.788 ;
      RECT 53.39 2.565 53.395 2.768 ;
      RECT 53.655 1.785 53.825 2.255 ;
      RECT 53.6 1.778 53.795 2.239 ;
      RECT 53.6 1.792 53.83 2.238 ;
      RECT 53.585 1.793 53.83 2.219 ;
      RECT 53.58 1.811 53.83 2.205 ;
      RECT 53.585 1.794 53.835 2.203 ;
      RECT 53.57 1.825 53.835 2.188 ;
      RECT 53.585 1.8 53.84 2.173 ;
      RECT 53.565 1.84 53.84 2.17 ;
      RECT 53.58 1.812 53.845 2.155 ;
      RECT 53.58 1.824 53.85 2.135 ;
      RECT 53.565 1.84 53.855 2.118 ;
      RECT 53.565 1.85 53.86 1.973 ;
      RECT 53.56 1.85 53.86 1.93 ;
      RECT 53.56 1.865 53.865 1.908 ;
      RECT 53.655 1.775 53.795 2.255 ;
      RECT 53.655 1.773 53.765 2.255 ;
      RECT 53.741 1.77 53.765 2.255 ;
      RECT 53.4 3.437 53.405 3.483 ;
      RECT 53.39 3.285 53.4 3.507 ;
      RECT 53.385 3.13 53.39 3.532 ;
      RECT 53.37 3.092 53.385 3.543 ;
      RECT 53.365 3.075 53.37 3.55 ;
      RECT 53.355 3.063 53.365 3.557 ;
      RECT 53.35 3.054 53.355 3.559 ;
      RECT 53.345 3.052 53.35 3.563 ;
      RECT 53.3 3.043 53.345 3.578 ;
      RECT 53.295 3.035 53.3 3.592 ;
      RECT 53.29 3.032 53.295 3.596 ;
      RECT 53.275 3.027 53.29 3.604 ;
      RECT 53.22 3.017 53.275 3.615 ;
      RECT 53.185 3.005 53.22 3.616 ;
      RECT 53.176 3 53.185 3.61 ;
      RECT 53.09 3 53.176 3.6 ;
      RECT 53.06 3 53.09 3.578 ;
      RECT 53.05 3 53.055 3.558 ;
      RECT 53.045 3 53.05 3.52 ;
      RECT 53.04 3 53.045 3.478 ;
      RECT 53.035 3 53.04 3.438 ;
      RECT 53.03 3 53.035 3.368 ;
      RECT 53.02 3 53.03 3.29 ;
      RECT 53.015 3 53.02 3.19 ;
      RECT 53.055 3 53.06 3.56 ;
      RECT 52.55 3.082 52.64 3.56 ;
      RECT 52.535 3.085 52.655 3.558 ;
      RECT 52.55 3.084 52.655 3.558 ;
      RECT 52.515 3.091 52.68 3.548 ;
      RECT 52.535 3.085 52.68 3.548 ;
      RECT 52.5 3.097 52.68 3.536 ;
      RECT 52.535 3.088 52.73 3.529 ;
      RECT 52.486 3.105 52.73 3.527 ;
      RECT 52.515 3.095 52.74 3.515 ;
      RECT 52.486 3.116 52.77 3.506 ;
      RECT 52.4 3.14 52.77 3.5 ;
      RECT 52.4 3.153 52.81 3.483 ;
      RECT 52.395 3.175 52.81 3.476 ;
      RECT 52.365 3.19 52.81 3.466 ;
      RECT 52.36 3.201 52.81 3.456 ;
      RECT 52.33 3.214 52.81 3.447 ;
      RECT 52.315 3.232 52.81 3.436 ;
      RECT 52.29 3.245 52.81 3.426 ;
      RECT 52.55 3.081 52.56 3.56 ;
      RECT 52.596 2.505 52.635 2.75 ;
      RECT 52.51 2.505 52.645 2.748 ;
      RECT 52.395 2.53 52.645 2.745 ;
      RECT 52.395 2.53 52.65 2.743 ;
      RECT 52.395 2.53 52.665 2.738 ;
      RECT 52.501 2.505 52.68 2.718 ;
      RECT 52.415 2.513 52.68 2.718 ;
      RECT 52.085 1.865 52.255 2.3 ;
      RECT 52.075 1.899 52.255 2.283 ;
      RECT 52.155 1.835 52.325 2.27 ;
      RECT 52.06 1.91 52.325 2.248 ;
      RECT 52.155 1.845 52.33 2.238 ;
      RECT 52.085 1.897 52.36 2.223 ;
      RECT 52.045 1.923 52.36 2.208 ;
      RECT 52.045 1.965 52.37 2.188 ;
      RECT 52.04 1.99 52.375 2.17 ;
      RECT 52.04 2 52.38 2.155 ;
      RECT 52.035 1.937 52.36 2.153 ;
      RECT 52.035 2.01 52.385 2.138 ;
      RECT 52.03 1.947 52.36 2.135 ;
      RECT 52.025 2.031 52.39 2.118 ;
      RECT 52.025 2.063 52.395 2.098 ;
      RECT 52.02 1.977 52.37 2.09 ;
      RECT 52.025 1.962 52.36 2.118 ;
      RECT 52.04 1.932 52.36 2.17 ;
      RECT 51.885 2.519 52.11 2.775 ;
      RECT 51.885 2.552 52.13 2.765 ;
      RECT 51.85 2.552 52.13 2.763 ;
      RECT 51.85 2.565 52.135 2.753 ;
      RECT 51.85 2.585 52.145 2.745 ;
      RECT 51.85 2.682 52.15 2.738 ;
      RECT 51.83 2.43 51.96 2.728 ;
      RECT 51.785 2.585 52.145 2.67 ;
      RECT 51.775 2.43 51.96 2.615 ;
      RECT 51.775 2.462 52.046 2.615 ;
      RECT 51.74 2.992 51.76 3.17 ;
      RECT 51.705 2.945 51.74 3.17 ;
      RECT 51.69 2.885 51.705 3.17 ;
      RECT 51.665 2.832 51.69 3.17 ;
      RECT 51.65 2.785 51.665 3.17 ;
      RECT 51.63 2.762 51.65 3.17 ;
      RECT 51.605 2.727 51.63 3.17 ;
      RECT 51.595 2.573 51.605 3.17 ;
      RECT 51.565 2.568 51.595 3.161 ;
      RECT 51.56 2.565 51.565 3.151 ;
      RECT 51.545 2.565 51.56 3.125 ;
      RECT 51.54 2.565 51.545 3.088 ;
      RECT 51.515 2.565 51.54 3.04 ;
      RECT 51.495 2.565 51.515 2.965 ;
      RECT 51.485 2.565 51.495 2.925 ;
      RECT 51.48 2.565 51.485 2.9 ;
      RECT 51.475 2.565 51.48 2.883 ;
      RECT 51.47 2.565 51.475 2.865 ;
      RECT 51.465 2.566 51.47 2.855 ;
      RECT 51.455 2.568 51.465 2.823 ;
      RECT 51.445 2.57 51.455 2.79 ;
      RECT 51.435 2.573 51.445 2.763 ;
      RECT 51.76 3 51.985 3.17 ;
      RECT 51.09 1.812 51.26 2.265 ;
      RECT 51.09 1.812 51.35 2.231 ;
      RECT 51.09 1.812 51.38 2.215 ;
      RECT 51.09 1.812 51.41 2.188 ;
      RECT 51.346 1.79 51.425 2.17 ;
      RECT 51.125 1.797 51.43 2.155 ;
      RECT 51.125 1.805 51.44 2.118 ;
      RECT 51.085 1.832 51.44 2.09 ;
      RECT 51.07 1.845 51.44 2.055 ;
      RECT 51.09 1.82 51.46 2.045 ;
      RECT 51.065 1.885 51.46 2.015 ;
      RECT 51.065 1.915 51.465 1.998 ;
      RECT 51.06 1.945 51.465 1.985 ;
      RECT 51.125 1.794 51.425 2.17 ;
      RECT 51.26 1.791 51.346 2.249 ;
      RECT 51.211 1.792 51.425 2.17 ;
      RECT 51.355 3.452 51.4 3.645 ;
      RECT 51.345 3.422 51.355 3.645 ;
      RECT 51.34 3.407 51.345 3.645 ;
      RECT 51.3 3.317 51.34 3.645 ;
      RECT 51.295 3.23 51.3 3.645 ;
      RECT 51.285 3.2 51.295 3.645 ;
      RECT 51.28 3.16 51.285 3.645 ;
      RECT 51.27 3.122 51.28 3.645 ;
      RECT 51.265 3.087 51.27 3.645 ;
      RECT 51.245 3.04 51.265 3.645 ;
      RECT 51.23 2.965 51.245 3.645 ;
      RECT 51.225 2.92 51.23 3.64 ;
      RECT 51.22 2.9 51.225 3.613 ;
      RECT 51.215 2.88 51.22 3.598 ;
      RECT 51.21 2.855 51.215 3.578 ;
      RECT 51.205 2.833 51.21 3.563 ;
      RECT 51.2 2.811 51.205 3.545 ;
      RECT 51.195 2.79 51.2 3.535 ;
      RECT 51.185 2.762 51.195 3.505 ;
      RECT 51.175 2.725 51.185 3.473 ;
      RECT 51.165 2.685 51.175 3.44 ;
      RECT 51.155 2.663 51.165 3.41 ;
      RECT 51.125 2.615 51.155 3.342 ;
      RECT 51.11 2.575 51.125 3.269 ;
      RECT 51.1 2.575 51.11 3.235 ;
      RECT 51.095 2.575 51.1 3.21 ;
      RECT 51.09 2.575 51.095 3.195 ;
      RECT 51.085 2.575 51.09 3.173 ;
      RECT 51.08 2.575 51.085 3.16 ;
      RECT 51.065 2.575 51.08 3.125 ;
      RECT 51.045 2.575 51.065 3.065 ;
      RECT 51.035 2.575 51.045 3.015 ;
      RECT 51.015 2.575 51.035 2.963 ;
      RECT 50.995 2.575 51.015 2.92 ;
      RECT 50.985 2.575 50.995 2.908 ;
      RECT 50.955 2.575 50.985 2.895 ;
      RECT 50.925 2.596 50.955 2.875 ;
      RECT 50.915 2.624 50.925 2.855 ;
      RECT 50.9 2.641 50.915 2.823 ;
      RECT 50.895 2.655 50.9 2.79 ;
      RECT 50.89 2.663 50.895 2.763 ;
      RECT 50.885 2.671 50.89 2.725 ;
      RECT 50.89 3.195 50.895 3.53 ;
      RECT 50.855 3.182 50.89 3.529 ;
      RECT 50.785 3.122 50.855 3.528 ;
      RECT 50.705 3.065 50.785 3.527 ;
      RECT 50.57 3.025 50.705 3.526 ;
      RECT 50.57 3.212 50.905 3.515 ;
      RECT 50.53 3.212 50.905 3.505 ;
      RECT 50.53 3.23 50.91 3.5 ;
      RECT 50.53 3.32 50.915 3.49 ;
      RECT 50.525 3.015 50.69 3.47 ;
      RECT 50.52 3.015 50.69 3.213 ;
      RECT 50.52 3.172 50.885 3.213 ;
      RECT 50.52 3.16 50.88 3.213 ;
      RECT 49.65 5.02 49.82 6.49 ;
      RECT 49.65 6.315 49.825 6.485 ;
      RECT 49.28 1.74 49.45 2.93 ;
      RECT 49.28 1.74 49.75 1.91 ;
      RECT 49.28 6.97 49.75 7.14 ;
      RECT 49.28 5.95 49.45 7.14 ;
      RECT 48.29 1.74 48.46 2.93 ;
      RECT 48.29 1.74 48.76 1.91 ;
      RECT 48.29 6.97 48.76 7.14 ;
      RECT 48.29 5.95 48.46 7.14 ;
      RECT 46.44 2.635 46.61 3.865 ;
      RECT 46.495 0.855 46.665 2.805 ;
      RECT 46.44 0.575 46.61 1.025 ;
      RECT 46.44 7.855 46.61 8.305 ;
      RECT 46.495 6.075 46.665 8.025 ;
      RECT 46.44 5.015 46.61 6.245 ;
      RECT 45.92 0.575 46.09 3.865 ;
      RECT 45.92 2.075 46.325 2.405 ;
      RECT 45.92 1.235 46.325 1.565 ;
      RECT 45.92 5.015 46.09 8.305 ;
      RECT 45.92 7.315 46.325 7.645 ;
      RECT 45.92 6.475 46.325 6.805 ;
      RECT 43.255 1.975 43.985 2.215 ;
      RECT 43.797 1.77 43.985 2.215 ;
      RECT 43.625 1.782 44 2.209 ;
      RECT 43.54 1.797 44.02 2.194 ;
      RECT 43.54 1.812 44.025 2.184 ;
      RECT 43.495 1.832 44.04 2.176 ;
      RECT 43.472 1.867 44.055 2.13 ;
      RECT 43.386 1.89 44.06 2.09 ;
      RECT 43.386 1.908 44.07 2.06 ;
      RECT 43.255 1.977 44.075 2.023 ;
      RECT 43.3 1.92 44.07 2.06 ;
      RECT 43.386 1.872 44.055 2.13 ;
      RECT 43.472 1.841 44.04 2.176 ;
      RECT 43.495 1.822 44.025 2.184 ;
      RECT 43.54 1.795 44 2.209 ;
      RECT 43.625 1.777 43.985 2.215 ;
      RECT 43.711 1.771 43.985 2.215 ;
      RECT 43.797 1.766 43.93 2.215 ;
      RECT 43.883 1.761 43.93 2.215 ;
      RECT 43.575 2.659 43.745 3.045 ;
      RECT 43.57 2.659 43.745 3.04 ;
      RECT 43.545 2.659 43.745 3.005 ;
      RECT 43.545 2.687 43.755 2.995 ;
      RECT 43.525 2.687 43.755 2.955 ;
      RECT 43.52 2.687 43.755 2.928 ;
      RECT 43.52 2.705 43.76 2.92 ;
      RECT 43.465 2.705 43.76 2.855 ;
      RECT 43.465 2.722 43.77 2.838 ;
      RECT 43.455 2.722 43.77 2.778 ;
      RECT 43.455 2.739 43.775 2.775 ;
      RECT 43.45 2.575 43.62 2.753 ;
      RECT 43.45 2.609 43.706 2.753 ;
      RECT 43.445 3.375 43.45 3.388 ;
      RECT 43.44 3.27 43.445 3.393 ;
      RECT 43.415 3.13 43.44 3.408 ;
      RECT 43.38 3.081 43.415 3.44 ;
      RECT 43.375 3.049 43.38 3.46 ;
      RECT 43.37 3.04 43.375 3.46 ;
      RECT 43.29 3.005 43.37 3.46 ;
      RECT 43.227 2.975 43.29 3.46 ;
      RECT 43.141 2.963 43.227 3.46 ;
      RECT 43.055 2.949 43.141 3.46 ;
      RECT 42.975 2.936 43.055 3.446 ;
      RECT 42.94 2.928 42.975 3.426 ;
      RECT 42.93 2.925 42.94 3.417 ;
      RECT 42.9 2.92 42.93 3.404 ;
      RECT 42.85 2.895 42.9 3.38 ;
      RECT 42.836 2.869 42.85 3.362 ;
      RECT 42.75 2.829 42.836 3.338 ;
      RECT 42.705 2.777 42.75 3.307 ;
      RECT 42.695 2.752 42.705 3.294 ;
      RECT 42.69 2.533 42.695 2.555 ;
      RECT 42.685 2.735 42.695 3.29 ;
      RECT 42.685 2.531 42.69 2.645 ;
      RECT 42.675 2.527 42.685 3.286 ;
      RECT 42.631 2.525 42.675 3.274 ;
      RECT 42.545 2.525 42.631 3.245 ;
      RECT 42.515 2.525 42.545 3.218 ;
      RECT 42.5 2.525 42.515 3.206 ;
      RECT 42.46 2.537 42.5 3.191 ;
      RECT 42.44 2.556 42.46 3.17 ;
      RECT 42.43 2.566 42.44 3.154 ;
      RECT 42.42 2.572 42.43 3.143 ;
      RECT 42.4 2.582 42.42 3.126 ;
      RECT 42.395 2.591 42.4 3.113 ;
      RECT 42.39 2.595 42.395 3.063 ;
      RECT 42.38 2.601 42.39 2.98 ;
      RECT 42.375 2.605 42.38 2.894 ;
      RECT 42.37 2.625 42.375 2.831 ;
      RECT 42.365 2.648 42.37 2.778 ;
      RECT 42.36 2.666 42.365 2.723 ;
      RECT 42.97 2.485 43.14 2.745 ;
      RECT 43.14 2.45 43.185 2.731 ;
      RECT 43.101 2.452 43.19 2.714 ;
      RECT 42.99 2.469 43.276 2.685 ;
      RECT 42.99 2.484 43.28 2.657 ;
      RECT 42.99 2.465 43.19 2.714 ;
      RECT 43.015 2.453 43.14 2.745 ;
      RECT 43.101 2.451 43.185 2.731 ;
      RECT 42.155 1.84 42.325 2.33 ;
      RECT 42.155 1.84 42.36 2.31 ;
      RECT 42.29 1.76 42.4 2.27 ;
      RECT 42.271 1.764 42.42 2.24 ;
      RECT 42.185 1.772 42.44 2.223 ;
      RECT 42.185 1.778 42.445 2.213 ;
      RECT 42.185 1.787 42.465 2.201 ;
      RECT 42.16 1.812 42.495 2.179 ;
      RECT 42.16 1.832 42.5 2.159 ;
      RECT 42.155 1.845 42.51 2.139 ;
      RECT 42.155 1.912 42.515 2.12 ;
      RECT 42.155 2.045 42.52 2.107 ;
      RECT 42.15 1.85 42.51 1.94 ;
      RECT 42.16 1.807 42.465 2.201 ;
      RECT 42.271 1.762 42.4 2.27 ;
      RECT 42.145 3.515 42.445 3.77 ;
      RECT 42.23 3.481 42.445 3.77 ;
      RECT 42.23 3.484 42.45 3.63 ;
      RECT 42.165 3.505 42.45 3.63 ;
      RECT 42.2 3.495 42.445 3.77 ;
      RECT 42.195 3.5 42.45 3.63 ;
      RECT 42.23 3.479 42.431 3.77 ;
      RECT 42.316 3.47 42.431 3.77 ;
      RECT 42.316 3.464 42.345 3.77 ;
      RECT 41.805 3.105 41.815 3.595 ;
      RECT 41.465 3.04 41.475 3.34 ;
      RECT 41.98 3.212 41.985 3.431 ;
      RECT 41.97 3.192 41.98 3.448 ;
      RECT 41.96 3.172 41.97 3.478 ;
      RECT 41.955 3.162 41.96 3.493 ;
      RECT 41.95 3.158 41.955 3.498 ;
      RECT 41.935 3.15 41.95 3.505 ;
      RECT 41.895 3.13 41.935 3.53 ;
      RECT 41.87 3.112 41.895 3.563 ;
      RECT 41.865 3.11 41.87 3.576 ;
      RECT 41.845 3.107 41.865 3.58 ;
      RECT 41.815 3.105 41.845 3.59 ;
      RECT 41.745 3.107 41.805 3.591 ;
      RECT 41.725 3.107 41.745 3.585 ;
      RECT 41.7 3.105 41.725 3.582 ;
      RECT 41.665 3.1 41.7 3.578 ;
      RECT 41.645 3.094 41.665 3.565 ;
      RECT 41.635 3.091 41.645 3.553 ;
      RECT 41.615 3.088 41.635 3.538 ;
      RECT 41.595 3.084 41.615 3.52 ;
      RECT 41.59 3.081 41.595 3.51 ;
      RECT 41.585 3.08 41.59 3.508 ;
      RECT 41.575 3.077 41.585 3.5 ;
      RECT 41.565 3.071 41.575 3.483 ;
      RECT 41.555 3.065 41.565 3.465 ;
      RECT 41.545 3.059 41.555 3.453 ;
      RECT 41.535 3.053 41.545 3.433 ;
      RECT 41.53 3.049 41.535 3.418 ;
      RECT 41.525 3.047 41.53 3.41 ;
      RECT 41.52 3.045 41.525 3.403 ;
      RECT 41.515 3.043 41.52 3.393 ;
      RECT 41.51 3.041 41.515 3.387 ;
      RECT 41.5 3.04 41.51 3.377 ;
      RECT 41.49 3.04 41.5 3.368 ;
      RECT 41.475 3.04 41.49 3.353 ;
      RECT 41.435 3.04 41.465 3.337 ;
      RECT 41.415 3.042 41.435 3.332 ;
      RECT 41.41 3.047 41.415 3.33 ;
      RECT 41.38 3.055 41.41 3.328 ;
      RECT 41.35 3.07 41.38 3.327 ;
      RECT 41.305 3.092 41.35 3.332 ;
      RECT 41.3 3.107 41.305 3.336 ;
      RECT 41.285 3.112 41.3 3.338 ;
      RECT 41.28 3.116 41.285 3.34 ;
      RECT 41.22 3.139 41.28 3.349 ;
      RECT 41.2 3.165 41.22 3.362 ;
      RECT 41.19 3.172 41.2 3.366 ;
      RECT 41.175 3.179 41.19 3.369 ;
      RECT 41.155 3.189 41.175 3.372 ;
      RECT 41.15 3.197 41.155 3.375 ;
      RECT 41.105 3.202 41.15 3.382 ;
      RECT 41.095 3.205 41.105 3.389 ;
      RECT 41.085 3.205 41.095 3.393 ;
      RECT 41.05 3.207 41.085 3.405 ;
      RECT 41.03 3.21 41.05 3.418 ;
      RECT 40.99 3.213 41.03 3.429 ;
      RECT 40.975 3.215 40.99 3.442 ;
      RECT 40.965 3.215 40.975 3.447 ;
      RECT 40.94 3.216 40.965 3.455 ;
      RECT 40.93 3.218 40.94 3.46 ;
      RECT 40.925 3.219 40.93 3.463 ;
      RECT 40.9 3.217 40.925 3.466 ;
      RECT 40.885 3.215 40.9 3.467 ;
      RECT 40.865 3.212 40.885 3.469 ;
      RECT 40.845 3.207 40.865 3.469 ;
      RECT 40.785 3.202 40.845 3.466 ;
      RECT 40.75 3.177 40.785 3.462 ;
      RECT 40.74 3.154 40.75 3.46 ;
      RECT 40.71 3.131 40.74 3.46 ;
      RECT 40.7 3.11 40.71 3.46 ;
      RECT 40.675 3.092 40.7 3.458 ;
      RECT 40.66 3.07 40.675 3.455 ;
      RECT 40.645 3.052 40.66 3.453 ;
      RECT 40.625 3.042 40.645 3.451 ;
      RECT 40.61 3.037 40.625 3.45 ;
      RECT 40.595 3.035 40.61 3.449 ;
      RECT 40.565 3.036 40.595 3.447 ;
      RECT 40.545 3.039 40.565 3.445 ;
      RECT 40.488 3.043 40.545 3.445 ;
      RECT 40.402 3.052 40.488 3.445 ;
      RECT 40.316 3.063 40.402 3.445 ;
      RECT 40.23 3.074 40.316 3.445 ;
      RECT 40.21 3.081 40.23 3.453 ;
      RECT 40.2 3.084 40.21 3.46 ;
      RECT 40.135 3.089 40.2 3.478 ;
      RECT 40.105 3.096 40.135 3.503 ;
      RECT 40.095 3.099 40.105 3.51 ;
      RECT 40.05 3.103 40.095 3.515 ;
      RECT 40.02 3.108 40.05 3.52 ;
      RECT 40.019 3.11 40.02 3.52 ;
      RECT 39.933 3.116 40.019 3.52 ;
      RECT 39.847 3.127 39.933 3.52 ;
      RECT 39.761 3.139 39.847 3.52 ;
      RECT 39.675 3.15 39.761 3.52 ;
      RECT 39.66 3.157 39.675 3.515 ;
      RECT 39.655 3.159 39.66 3.509 ;
      RECT 39.635 3.17 39.655 3.504 ;
      RECT 39.625 3.188 39.635 3.498 ;
      RECT 39.62 3.2 39.625 3.298 ;
      RECT 41.915 1.953 41.935 2.04 ;
      RECT 41.91 1.888 41.915 2.072 ;
      RECT 41.9 1.855 41.91 2.077 ;
      RECT 41.895 1.835 41.9 2.083 ;
      RECT 41.865 1.835 41.895 2.1 ;
      RECT 41.816 1.835 41.865 2.136 ;
      RECT 41.73 1.835 41.816 2.194 ;
      RECT 41.701 1.845 41.73 2.243 ;
      RECT 41.615 1.887 41.701 2.296 ;
      RECT 41.595 1.925 41.615 2.343 ;
      RECT 41.57 1.942 41.595 2.363 ;
      RECT 41.56 1.956 41.57 2.383 ;
      RECT 41.555 1.962 41.56 2.393 ;
      RECT 41.55 1.966 41.555 2.4 ;
      RECT 41.5 1.986 41.55 2.405 ;
      RECT 41.435 2.03 41.5 2.405 ;
      RECT 41.41 2.08 41.435 2.405 ;
      RECT 41.4 2.11 41.41 2.405 ;
      RECT 41.395 2.137 41.4 2.405 ;
      RECT 41.39 2.155 41.395 2.405 ;
      RECT 41.38 2.197 41.39 2.405 ;
      RECT 41.73 2.755 41.9 2.93 ;
      RECT 41.67 2.583 41.73 2.918 ;
      RECT 41.66 2.576 41.67 2.901 ;
      RECT 41.615 2.755 41.9 2.881 ;
      RECT 41.596 2.755 41.9 2.859 ;
      RECT 41.51 2.755 41.9 2.824 ;
      RECT 41.49 2.575 41.66 2.78 ;
      RECT 41.49 2.722 41.895 2.78 ;
      RECT 41.49 2.67 41.87 2.78 ;
      RECT 41.49 2.625 41.835 2.78 ;
      RECT 41.49 2.607 41.8 2.78 ;
      RECT 41.49 2.597 41.795 2.78 ;
      RECT 41.66 7.855 41.83 8.305 ;
      RECT 41.715 6.075 41.885 8.025 ;
      RECT 41.66 5.015 41.83 6.245 ;
      RECT 41.14 5.015 41.31 8.305 ;
      RECT 41.14 7.315 41.545 7.645 ;
      RECT 41.14 6.475 41.545 6.805 ;
      RECT 41.21 3.555 41.4 3.78 ;
      RECT 41.2 3.556 41.405 3.775 ;
      RECT 41.2 3.558 41.415 3.755 ;
      RECT 41.2 3.562 41.42 3.74 ;
      RECT 41.2 3.549 41.37 3.775 ;
      RECT 41.2 3.552 41.395 3.775 ;
      RECT 41.21 3.548 41.37 3.78 ;
      RECT 41.296 3.546 41.37 3.78 ;
      RECT 40.92 2.797 41.09 3.035 ;
      RECT 40.92 2.797 41.176 2.949 ;
      RECT 40.92 2.797 41.18 2.859 ;
      RECT 40.97 2.57 41.19 2.838 ;
      RECT 40.965 2.587 41.195 2.811 ;
      RECT 40.93 2.745 41.195 2.811 ;
      RECT 40.95 2.595 41.09 3.035 ;
      RECT 40.94 2.677 41.2 2.794 ;
      RECT 40.935 2.725 41.2 2.794 ;
      RECT 40.94 2.635 41.195 2.811 ;
      RECT 40.965 2.572 41.19 2.838 ;
      RECT 40.53 2.547 40.7 2.745 ;
      RECT 40.53 2.547 40.745 2.72 ;
      RECT 40.6 2.49 40.77 2.678 ;
      RECT 40.575 2.505 40.77 2.678 ;
      RECT 40.19 2.551 40.22 2.745 ;
      RECT 40.185 2.523 40.19 2.745 ;
      RECT 40.155 2.497 40.185 2.747 ;
      RECT 40.13 2.455 40.155 2.75 ;
      RECT 40.12 2.427 40.13 2.752 ;
      RECT 40.085 2.407 40.12 2.754 ;
      RECT 40.02 2.392 40.085 2.76 ;
      RECT 39.97 2.39 40.02 2.766 ;
      RECT 39.947 2.392 39.97 2.771 ;
      RECT 39.861 2.403 39.947 2.777 ;
      RECT 39.775 2.421 39.861 2.787 ;
      RECT 39.76 2.432 39.775 2.793 ;
      RECT 39.69 2.455 39.76 2.799 ;
      RECT 39.635 2.487 39.69 2.807 ;
      RECT 39.595 2.51 39.635 2.813 ;
      RECT 39.581 2.523 39.595 2.816 ;
      RECT 39.495 2.545 39.581 2.822 ;
      RECT 39.48 2.57 39.495 2.828 ;
      RECT 39.44 2.585 39.48 2.832 ;
      RECT 39.39 2.6 39.44 2.837 ;
      RECT 39.365 2.607 39.39 2.841 ;
      RECT 39.305 2.602 39.365 2.845 ;
      RECT 39.29 2.593 39.305 2.849 ;
      RECT 39.22 2.583 39.29 2.845 ;
      RECT 39.195 2.575 39.215 2.835 ;
      RECT 39.136 2.575 39.195 2.813 ;
      RECT 39.05 2.575 39.136 2.77 ;
      RECT 39.215 2.575 39.22 2.84 ;
      RECT 39.91 1.806 40.08 2.14 ;
      RECT 39.88 1.806 40.08 2.135 ;
      RECT 39.82 1.773 39.88 2.123 ;
      RECT 39.82 1.829 40.09 2.118 ;
      RECT 39.795 1.829 40.09 2.112 ;
      RECT 39.79 1.77 39.82 2.109 ;
      RECT 39.775 1.776 39.91 2.107 ;
      RECT 39.77 1.784 39.995 2.095 ;
      RECT 39.77 1.836 40.105 2.048 ;
      RECT 39.755 1.792 39.995 2.043 ;
      RECT 39.755 1.862 40.115 1.984 ;
      RECT 39.725 1.812 40.08 1.945 ;
      RECT 39.725 1.902 40.125 1.941 ;
      RECT 39.775 1.781 39.995 2.107 ;
      RECT 39.115 2.111 39.17 2.375 ;
      RECT 39.115 2.111 39.235 2.374 ;
      RECT 39.115 2.111 39.26 2.373 ;
      RECT 39.115 2.111 39.325 2.372 ;
      RECT 39.26 2.077 39.34 2.371 ;
      RECT 39.075 2.121 39.485 2.37 ;
      RECT 39.115 2.118 39.485 2.37 ;
      RECT 39.075 2.126 39.49 2.363 ;
      RECT 39.06 2.128 39.49 2.362 ;
      RECT 39.06 2.135 39.495 2.358 ;
      RECT 39.04 2.134 39.49 2.354 ;
      RECT 39.04 2.142 39.5 2.353 ;
      RECT 39.035 2.139 39.495 2.349 ;
      RECT 39.035 2.152 39.51 2.348 ;
      RECT 39.02 2.142 39.5 2.347 ;
      RECT 38.985 2.155 39.51 2.34 ;
      RECT 39.17 2.11 39.48 2.37 ;
      RECT 39.17 2.095 39.43 2.37 ;
      RECT 39.235 2.082 39.365 2.37 ;
      RECT 38.78 3.171 38.795 3.564 ;
      RECT 38.745 3.176 38.795 3.563 ;
      RECT 38.78 3.175 38.84 3.562 ;
      RECT 38.725 3.186 38.84 3.561 ;
      RECT 38.74 3.182 38.84 3.561 ;
      RECT 38.705 3.192 38.915 3.558 ;
      RECT 38.705 3.211 38.96 3.556 ;
      RECT 38.705 3.218 38.965 3.553 ;
      RECT 38.69 3.195 38.915 3.55 ;
      RECT 38.67 3.2 38.915 3.543 ;
      RECT 38.665 3.204 38.915 3.539 ;
      RECT 38.665 3.221 38.975 3.538 ;
      RECT 38.645 3.215 38.96 3.534 ;
      RECT 38.645 3.224 38.98 3.528 ;
      RECT 38.64 3.23 38.98 3.3 ;
      RECT 38.705 3.19 38.84 3.558 ;
      RECT 38.58 2.553 38.78 2.865 ;
      RECT 38.655 2.531 38.78 2.865 ;
      RECT 38.595 2.55 38.785 2.85 ;
      RECT 38.565 2.561 38.785 2.848 ;
      RECT 38.58 2.556 38.79 2.814 ;
      RECT 38.565 2.66 38.795 2.781 ;
      RECT 38.595 2.532 38.78 2.865 ;
      RECT 38.655 2.51 38.755 2.865 ;
      RECT 38.68 2.507 38.755 2.865 ;
      RECT 38.68 2.502 38.7 2.865 ;
      RECT 38.085 2.57 38.26 2.745 ;
      RECT 38.08 2.57 38.26 2.743 ;
      RECT 38.055 2.57 38.26 2.738 ;
      RECT 38 2.55 38.17 2.728 ;
      RECT 38 2.557 38.235 2.728 ;
      RECT 38.085 3.237 38.1 3.42 ;
      RECT 38.075 3.215 38.085 3.42 ;
      RECT 38.06 3.195 38.075 3.42 ;
      RECT 38.05 3.17 38.06 3.42 ;
      RECT 38.02 3.135 38.05 3.42 ;
      RECT 37.985 3.075 38.02 3.42 ;
      RECT 37.98 3.037 37.985 3.42 ;
      RECT 37.93 2.988 37.98 3.42 ;
      RECT 37.92 2.938 37.93 3.408 ;
      RECT 37.905 2.917 37.92 3.368 ;
      RECT 37.885 2.885 37.905 3.318 ;
      RECT 37.86 2.841 37.885 3.258 ;
      RECT 37.855 2.813 37.86 3.213 ;
      RECT 37.85 2.804 37.855 3.199 ;
      RECT 37.845 2.797 37.85 3.186 ;
      RECT 37.84 2.792 37.845 3.175 ;
      RECT 37.835 2.777 37.84 3.165 ;
      RECT 37.83 2.755 37.835 3.152 ;
      RECT 37.82 2.715 37.83 3.127 ;
      RECT 37.795 2.645 37.82 3.083 ;
      RECT 37.79 2.585 37.795 3.048 ;
      RECT 37.775 2.565 37.79 3.015 ;
      RECT 37.77 2.565 37.775 2.99 ;
      RECT 37.74 2.565 37.77 2.945 ;
      RECT 37.695 2.565 37.74 2.885 ;
      RECT 37.62 2.565 37.695 2.833 ;
      RECT 37.615 2.565 37.62 2.798 ;
      RECT 37.61 2.565 37.615 2.788 ;
      RECT 37.605 2.565 37.61 2.768 ;
      RECT 37.87 1.785 38.04 2.255 ;
      RECT 37.815 1.778 38.01 2.239 ;
      RECT 37.815 1.792 38.045 2.238 ;
      RECT 37.8 1.793 38.045 2.219 ;
      RECT 37.795 1.811 38.045 2.205 ;
      RECT 37.8 1.794 38.05 2.203 ;
      RECT 37.785 1.825 38.05 2.188 ;
      RECT 37.8 1.8 38.055 2.173 ;
      RECT 37.78 1.84 38.055 2.17 ;
      RECT 37.795 1.812 38.06 2.155 ;
      RECT 37.795 1.824 38.065 2.135 ;
      RECT 37.78 1.84 38.07 2.118 ;
      RECT 37.78 1.85 38.075 1.973 ;
      RECT 37.775 1.85 38.075 1.93 ;
      RECT 37.775 1.865 38.08 1.908 ;
      RECT 37.87 1.775 38.01 2.255 ;
      RECT 37.87 1.773 37.98 2.255 ;
      RECT 37.956 1.77 37.98 2.255 ;
      RECT 37.615 3.437 37.62 3.483 ;
      RECT 37.605 3.285 37.615 3.507 ;
      RECT 37.6 3.13 37.605 3.532 ;
      RECT 37.585 3.092 37.6 3.543 ;
      RECT 37.58 3.075 37.585 3.55 ;
      RECT 37.57 3.063 37.58 3.557 ;
      RECT 37.565 3.054 37.57 3.559 ;
      RECT 37.56 3.052 37.565 3.563 ;
      RECT 37.515 3.043 37.56 3.578 ;
      RECT 37.51 3.035 37.515 3.592 ;
      RECT 37.505 3.032 37.51 3.596 ;
      RECT 37.49 3.027 37.505 3.604 ;
      RECT 37.435 3.017 37.49 3.615 ;
      RECT 37.4 3.005 37.435 3.616 ;
      RECT 37.391 3 37.4 3.61 ;
      RECT 37.305 3 37.391 3.6 ;
      RECT 37.275 3 37.305 3.578 ;
      RECT 37.265 3 37.27 3.558 ;
      RECT 37.26 3 37.265 3.52 ;
      RECT 37.255 3 37.26 3.478 ;
      RECT 37.25 3 37.255 3.438 ;
      RECT 37.245 3 37.25 3.368 ;
      RECT 37.235 3 37.245 3.29 ;
      RECT 37.23 3 37.235 3.19 ;
      RECT 37.27 3 37.275 3.56 ;
      RECT 36.765 3.082 36.855 3.56 ;
      RECT 36.75 3.085 36.87 3.558 ;
      RECT 36.765 3.084 36.87 3.558 ;
      RECT 36.73 3.091 36.895 3.548 ;
      RECT 36.75 3.085 36.895 3.548 ;
      RECT 36.715 3.097 36.895 3.536 ;
      RECT 36.75 3.088 36.945 3.529 ;
      RECT 36.701 3.105 36.945 3.527 ;
      RECT 36.73 3.095 36.955 3.515 ;
      RECT 36.701 3.116 36.985 3.506 ;
      RECT 36.615 3.14 36.985 3.5 ;
      RECT 36.615 3.153 37.025 3.483 ;
      RECT 36.61 3.175 37.025 3.476 ;
      RECT 36.58 3.19 37.025 3.466 ;
      RECT 36.575 3.201 37.025 3.456 ;
      RECT 36.545 3.214 37.025 3.447 ;
      RECT 36.53 3.232 37.025 3.436 ;
      RECT 36.505 3.245 37.025 3.426 ;
      RECT 36.765 3.081 36.775 3.56 ;
      RECT 36.811 2.505 36.85 2.75 ;
      RECT 36.725 2.505 36.86 2.748 ;
      RECT 36.61 2.53 36.86 2.745 ;
      RECT 36.61 2.53 36.865 2.743 ;
      RECT 36.61 2.53 36.88 2.738 ;
      RECT 36.716 2.505 36.895 2.718 ;
      RECT 36.63 2.513 36.895 2.718 ;
      RECT 36.3 1.865 36.47 2.3 ;
      RECT 36.29 1.899 36.47 2.283 ;
      RECT 36.37 1.835 36.54 2.27 ;
      RECT 36.275 1.91 36.54 2.248 ;
      RECT 36.37 1.845 36.545 2.238 ;
      RECT 36.3 1.897 36.575 2.223 ;
      RECT 36.26 1.923 36.575 2.208 ;
      RECT 36.26 1.965 36.585 2.188 ;
      RECT 36.255 1.99 36.59 2.17 ;
      RECT 36.255 2 36.595 2.155 ;
      RECT 36.25 1.937 36.575 2.153 ;
      RECT 36.25 2.01 36.6 2.138 ;
      RECT 36.245 1.947 36.575 2.135 ;
      RECT 36.24 2.031 36.605 2.118 ;
      RECT 36.24 2.063 36.61 2.098 ;
      RECT 36.235 1.977 36.585 2.09 ;
      RECT 36.24 1.962 36.575 2.118 ;
      RECT 36.255 1.932 36.575 2.17 ;
      RECT 36.1 2.519 36.325 2.775 ;
      RECT 36.1 2.552 36.345 2.765 ;
      RECT 36.065 2.552 36.345 2.763 ;
      RECT 36.065 2.565 36.35 2.753 ;
      RECT 36.065 2.585 36.36 2.745 ;
      RECT 36.065 2.682 36.365 2.738 ;
      RECT 36.045 2.43 36.175 2.728 ;
      RECT 36 2.585 36.36 2.67 ;
      RECT 35.99 2.43 36.175 2.615 ;
      RECT 35.99 2.462 36.261 2.615 ;
      RECT 35.955 2.992 35.975 3.17 ;
      RECT 35.92 2.945 35.955 3.17 ;
      RECT 35.905 2.885 35.92 3.17 ;
      RECT 35.88 2.832 35.905 3.17 ;
      RECT 35.865 2.785 35.88 3.17 ;
      RECT 35.845 2.762 35.865 3.17 ;
      RECT 35.82 2.727 35.845 3.17 ;
      RECT 35.81 2.573 35.82 3.17 ;
      RECT 35.78 2.568 35.81 3.161 ;
      RECT 35.775 2.565 35.78 3.151 ;
      RECT 35.76 2.565 35.775 3.125 ;
      RECT 35.755 2.565 35.76 3.088 ;
      RECT 35.73 2.565 35.755 3.04 ;
      RECT 35.71 2.565 35.73 2.965 ;
      RECT 35.7 2.565 35.71 2.925 ;
      RECT 35.695 2.565 35.7 2.9 ;
      RECT 35.69 2.565 35.695 2.883 ;
      RECT 35.685 2.565 35.69 2.865 ;
      RECT 35.68 2.566 35.685 2.855 ;
      RECT 35.67 2.568 35.68 2.823 ;
      RECT 35.66 2.57 35.67 2.79 ;
      RECT 35.65 2.573 35.66 2.763 ;
      RECT 35.975 3 36.2 3.17 ;
      RECT 35.305 1.812 35.475 2.265 ;
      RECT 35.305 1.812 35.565 2.231 ;
      RECT 35.305 1.812 35.595 2.215 ;
      RECT 35.305 1.812 35.625 2.188 ;
      RECT 35.561 1.79 35.64 2.17 ;
      RECT 35.34 1.797 35.645 2.155 ;
      RECT 35.34 1.805 35.655 2.118 ;
      RECT 35.3 1.832 35.655 2.09 ;
      RECT 35.285 1.845 35.655 2.055 ;
      RECT 35.305 1.82 35.675 2.045 ;
      RECT 35.28 1.885 35.675 2.015 ;
      RECT 35.28 1.915 35.68 1.998 ;
      RECT 35.275 1.945 35.68 1.985 ;
      RECT 35.34 1.794 35.64 2.17 ;
      RECT 35.475 1.791 35.561 2.249 ;
      RECT 35.426 1.792 35.64 2.17 ;
      RECT 35.57 3.452 35.615 3.645 ;
      RECT 35.56 3.422 35.57 3.645 ;
      RECT 35.555 3.407 35.56 3.645 ;
      RECT 35.515 3.317 35.555 3.645 ;
      RECT 35.51 3.23 35.515 3.645 ;
      RECT 35.5 3.2 35.51 3.645 ;
      RECT 35.495 3.16 35.5 3.645 ;
      RECT 35.485 3.122 35.495 3.645 ;
      RECT 35.48 3.087 35.485 3.645 ;
      RECT 35.46 3.04 35.48 3.645 ;
      RECT 35.445 2.965 35.46 3.645 ;
      RECT 35.44 2.92 35.445 3.64 ;
      RECT 35.435 2.9 35.44 3.613 ;
      RECT 35.43 2.88 35.435 3.598 ;
      RECT 35.425 2.855 35.43 3.578 ;
      RECT 35.42 2.833 35.425 3.563 ;
      RECT 35.415 2.811 35.42 3.545 ;
      RECT 35.41 2.79 35.415 3.535 ;
      RECT 35.4 2.762 35.41 3.505 ;
      RECT 35.39 2.725 35.4 3.473 ;
      RECT 35.38 2.685 35.39 3.44 ;
      RECT 35.37 2.663 35.38 3.41 ;
      RECT 35.34 2.615 35.37 3.342 ;
      RECT 35.325 2.575 35.34 3.269 ;
      RECT 35.315 2.575 35.325 3.235 ;
      RECT 35.31 2.575 35.315 3.21 ;
      RECT 35.305 2.575 35.31 3.195 ;
      RECT 35.3 2.575 35.305 3.173 ;
      RECT 35.295 2.575 35.3 3.16 ;
      RECT 35.28 2.575 35.295 3.125 ;
      RECT 35.26 2.575 35.28 3.065 ;
      RECT 35.25 2.575 35.26 3.015 ;
      RECT 35.23 2.575 35.25 2.963 ;
      RECT 35.21 2.575 35.23 2.92 ;
      RECT 35.2 2.575 35.21 2.908 ;
      RECT 35.17 2.575 35.2 2.895 ;
      RECT 35.14 2.596 35.17 2.875 ;
      RECT 35.13 2.624 35.14 2.855 ;
      RECT 35.115 2.641 35.13 2.823 ;
      RECT 35.11 2.655 35.115 2.79 ;
      RECT 35.105 2.663 35.11 2.763 ;
      RECT 35.1 2.671 35.105 2.725 ;
      RECT 35.105 3.195 35.11 3.53 ;
      RECT 35.07 3.182 35.105 3.529 ;
      RECT 35 3.122 35.07 3.528 ;
      RECT 34.92 3.065 35 3.527 ;
      RECT 34.785 3.025 34.92 3.526 ;
      RECT 34.785 3.212 35.12 3.515 ;
      RECT 34.745 3.212 35.12 3.505 ;
      RECT 34.745 3.23 35.125 3.5 ;
      RECT 34.745 3.32 35.13 3.49 ;
      RECT 34.74 3.015 34.905 3.47 ;
      RECT 34.735 3.015 34.905 3.213 ;
      RECT 34.735 3.172 35.1 3.213 ;
      RECT 34.735 3.16 35.095 3.213 ;
      RECT 33.875 5.02 34.045 6.49 ;
      RECT 33.875 6.315 34.05 6.485 ;
      RECT 33.505 1.74 33.675 2.93 ;
      RECT 33.505 1.74 33.975 1.91 ;
      RECT 33.505 6.97 33.975 7.14 ;
      RECT 33.505 5.95 33.675 7.14 ;
      RECT 32.515 1.74 32.685 2.93 ;
      RECT 32.515 1.74 32.985 1.91 ;
      RECT 32.515 6.97 32.985 7.14 ;
      RECT 32.515 5.95 32.685 7.14 ;
      RECT 30.665 2.635 30.835 3.865 ;
      RECT 30.72 0.855 30.89 2.805 ;
      RECT 30.665 0.575 30.835 1.025 ;
      RECT 30.665 7.855 30.835 8.305 ;
      RECT 30.72 6.075 30.89 8.025 ;
      RECT 30.665 5.015 30.835 6.245 ;
      RECT 30.145 0.575 30.315 3.865 ;
      RECT 30.145 2.075 30.55 2.405 ;
      RECT 30.145 1.235 30.55 1.565 ;
      RECT 30.145 5.015 30.315 8.305 ;
      RECT 30.145 7.315 30.55 7.645 ;
      RECT 30.145 6.475 30.55 6.805 ;
      RECT 27.48 1.975 28.21 2.215 ;
      RECT 28.022 1.77 28.21 2.215 ;
      RECT 27.85 1.782 28.225 2.209 ;
      RECT 27.765 1.797 28.245 2.194 ;
      RECT 27.765 1.812 28.25 2.184 ;
      RECT 27.72 1.832 28.265 2.176 ;
      RECT 27.697 1.867 28.28 2.13 ;
      RECT 27.611 1.89 28.285 2.09 ;
      RECT 27.611 1.908 28.295 2.06 ;
      RECT 27.48 1.977 28.3 2.023 ;
      RECT 27.525 1.92 28.295 2.06 ;
      RECT 27.611 1.872 28.28 2.13 ;
      RECT 27.697 1.841 28.265 2.176 ;
      RECT 27.72 1.822 28.25 2.184 ;
      RECT 27.765 1.795 28.225 2.209 ;
      RECT 27.85 1.777 28.21 2.215 ;
      RECT 27.936 1.771 28.21 2.215 ;
      RECT 28.022 1.766 28.155 2.215 ;
      RECT 28.108 1.761 28.155 2.215 ;
      RECT 27.8 2.659 27.97 3.045 ;
      RECT 27.795 2.659 27.97 3.04 ;
      RECT 27.77 2.659 27.97 3.005 ;
      RECT 27.77 2.687 27.98 2.995 ;
      RECT 27.75 2.687 27.98 2.955 ;
      RECT 27.745 2.687 27.98 2.928 ;
      RECT 27.745 2.705 27.985 2.92 ;
      RECT 27.69 2.705 27.985 2.855 ;
      RECT 27.69 2.722 27.995 2.838 ;
      RECT 27.68 2.722 27.995 2.778 ;
      RECT 27.68 2.739 28 2.775 ;
      RECT 27.675 2.575 27.845 2.753 ;
      RECT 27.675 2.609 27.931 2.753 ;
      RECT 27.67 3.375 27.675 3.388 ;
      RECT 27.665 3.27 27.67 3.393 ;
      RECT 27.64 3.13 27.665 3.408 ;
      RECT 27.605 3.081 27.64 3.44 ;
      RECT 27.6 3.049 27.605 3.46 ;
      RECT 27.595 3.04 27.6 3.46 ;
      RECT 27.515 3.005 27.595 3.46 ;
      RECT 27.452 2.975 27.515 3.46 ;
      RECT 27.366 2.963 27.452 3.46 ;
      RECT 27.28 2.949 27.366 3.46 ;
      RECT 27.2 2.936 27.28 3.446 ;
      RECT 27.165 2.928 27.2 3.426 ;
      RECT 27.155 2.925 27.165 3.417 ;
      RECT 27.125 2.92 27.155 3.404 ;
      RECT 27.075 2.895 27.125 3.38 ;
      RECT 27.061 2.869 27.075 3.362 ;
      RECT 26.975 2.829 27.061 3.338 ;
      RECT 26.93 2.777 26.975 3.307 ;
      RECT 26.92 2.752 26.93 3.294 ;
      RECT 26.915 2.533 26.92 2.555 ;
      RECT 26.91 2.735 26.92 3.29 ;
      RECT 26.91 2.531 26.915 2.645 ;
      RECT 26.9 2.527 26.91 3.286 ;
      RECT 26.856 2.525 26.9 3.274 ;
      RECT 26.77 2.525 26.856 3.245 ;
      RECT 26.74 2.525 26.77 3.218 ;
      RECT 26.725 2.525 26.74 3.206 ;
      RECT 26.685 2.537 26.725 3.191 ;
      RECT 26.665 2.556 26.685 3.17 ;
      RECT 26.655 2.566 26.665 3.154 ;
      RECT 26.645 2.572 26.655 3.143 ;
      RECT 26.625 2.582 26.645 3.126 ;
      RECT 26.62 2.591 26.625 3.113 ;
      RECT 26.615 2.595 26.62 3.063 ;
      RECT 26.605 2.601 26.615 2.98 ;
      RECT 26.6 2.605 26.605 2.894 ;
      RECT 26.595 2.625 26.6 2.831 ;
      RECT 26.59 2.648 26.595 2.778 ;
      RECT 26.585 2.666 26.59 2.723 ;
      RECT 27.195 2.485 27.365 2.745 ;
      RECT 27.365 2.45 27.41 2.731 ;
      RECT 27.326 2.452 27.415 2.714 ;
      RECT 27.215 2.469 27.501 2.685 ;
      RECT 27.215 2.484 27.505 2.657 ;
      RECT 27.215 2.465 27.415 2.714 ;
      RECT 27.24 2.453 27.365 2.745 ;
      RECT 27.326 2.451 27.41 2.731 ;
      RECT 26.38 1.84 26.55 2.33 ;
      RECT 26.38 1.84 26.585 2.31 ;
      RECT 26.515 1.76 26.625 2.27 ;
      RECT 26.496 1.764 26.645 2.24 ;
      RECT 26.41 1.772 26.665 2.223 ;
      RECT 26.41 1.778 26.67 2.213 ;
      RECT 26.41 1.787 26.69 2.201 ;
      RECT 26.385 1.812 26.72 2.179 ;
      RECT 26.385 1.832 26.725 2.159 ;
      RECT 26.38 1.845 26.735 2.139 ;
      RECT 26.38 1.912 26.74 2.12 ;
      RECT 26.38 2.045 26.745 2.107 ;
      RECT 26.375 1.85 26.735 1.94 ;
      RECT 26.385 1.807 26.69 2.201 ;
      RECT 26.496 1.762 26.625 2.27 ;
      RECT 26.37 3.515 26.67 3.77 ;
      RECT 26.455 3.481 26.67 3.77 ;
      RECT 26.455 3.484 26.675 3.63 ;
      RECT 26.39 3.505 26.675 3.63 ;
      RECT 26.425 3.495 26.67 3.77 ;
      RECT 26.42 3.5 26.675 3.63 ;
      RECT 26.455 3.479 26.656 3.77 ;
      RECT 26.541 3.47 26.656 3.77 ;
      RECT 26.541 3.464 26.57 3.77 ;
      RECT 26.03 3.105 26.04 3.595 ;
      RECT 25.69 3.04 25.7 3.34 ;
      RECT 26.205 3.212 26.21 3.431 ;
      RECT 26.195 3.192 26.205 3.448 ;
      RECT 26.185 3.172 26.195 3.478 ;
      RECT 26.18 3.162 26.185 3.493 ;
      RECT 26.175 3.158 26.18 3.498 ;
      RECT 26.16 3.15 26.175 3.505 ;
      RECT 26.12 3.13 26.16 3.53 ;
      RECT 26.095 3.112 26.12 3.563 ;
      RECT 26.09 3.11 26.095 3.576 ;
      RECT 26.07 3.107 26.09 3.58 ;
      RECT 26.04 3.105 26.07 3.59 ;
      RECT 25.97 3.107 26.03 3.591 ;
      RECT 25.95 3.107 25.97 3.585 ;
      RECT 25.925 3.105 25.95 3.582 ;
      RECT 25.89 3.1 25.925 3.578 ;
      RECT 25.87 3.094 25.89 3.565 ;
      RECT 25.86 3.091 25.87 3.553 ;
      RECT 25.84 3.088 25.86 3.538 ;
      RECT 25.82 3.084 25.84 3.52 ;
      RECT 25.815 3.081 25.82 3.51 ;
      RECT 25.81 3.08 25.815 3.508 ;
      RECT 25.8 3.077 25.81 3.5 ;
      RECT 25.79 3.071 25.8 3.483 ;
      RECT 25.78 3.065 25.79 3.465 ;
      RECT 25.77 3.059 25.78 3.453 ;
      RECT 25.76 3.053 25.77 3.433 ;
      RECT 25.755 3.049 25.76 3.418 ;
      RECT 25.75 3.047 25.755 3.41 ;
      RECT 25.745 3.045 25.75 3.403 ;
      RECT 25.74 3.043 25.745 3.393 ;
      RECT 25.735 3.041 25.74 3.387 ;
      RECT 25.725 3.04 25.735 3.377 ;
      RECT 25.715 3.04 25.725 3.368 ;
      RECT 25.7 3.04 25.715 3.353 ;
      RECT 25.66 3.04 25.69 3.337 ;
      RECT 25.64 3.042 25.66 3.332 ;
      RECT 25.635 3.047 25.64 3.33 ;
      RECT 25.605 3.055 25.635 3.328 ;
      RECT 25.575 3.07 25.605 3.327 ;
      RECT 25.53 3.092 25.575 3.332 ;
      RECT 25.525 3.107 25.53 3.336 ;
      RECT 25.51 3.112 25.525 3.338 ;
      RECT 25.505 3.116 25.51 3.34 ;
      RECT 25.445 3.139 25.505 3.349 ;
      RECT 25.425 3.165 25.445 3.362 ;
      RECT 25.415 3.172 25.425 3.366 ;
      RECT 25.4 3.179 25.415 3.369 ;
      RECT 25.38 3.189 25.4 3.372 ;
      RECT 25.375 3.197 25.38 3.375 ;
      RECT 25.33 3.202 25.375 3.382 ;
      RECT 25.32 3.205 25.33 3.389 ;
      RECT 25.31 3.205 25.32 3.393 ;
      RECT 25.275 3.207 25.31 3.405 ;
      RECT 25.255 3.21 25.275 3.418 ;
      RECT 25.215 3.213 25.255 3.429 ;
      RECT 25.2 3.215 25.215 3.442 ;
      RECT 25.19 3.215 25.2 3.447 ;
      RECT 25.165 3.216 25.19 3.455 ;
      RECT 25.155 3.218 25.165 3.46 ;
      RECT 25.15 3.219 25.155 3.463 ;
      RECT 25.125 3.217 25.15 3.466 ;
      RECT 25.11 3.215 25.125 3.467 ;
      RECT 25.09 3.212 25.11 3.469 ;
      RECT 25.07 3.207 25.09 3.469 ;
      RECT 25.01 3.202 25.07 3.466 ;
      RECT 24.975 3.177 25.01 3.462 ;
      RECT 24.965 3.154 24.975 3.46 ;
      RECT 24.935 3.131 24.965 3.46 ;
      RECT 24.925 3.11 24.935 3.46 ;
      RECT 24.9 3.092 24.925 3.458 ;
      RECT 24.885 3.07 24.9 3.455 ;
      RECT 24.87 3.052 24.885 3.453 ;
      RECT 24.85 3.042 24.87 3.451 ;
      RECT 24.835 3.037 24.85 3.45 ;
      RECT 24.82 3.035 24.835 3.449 ;
      RECT 24.79 3.036 24.82 3.447 ;
      RECT 24.77 3.039 24.79 3.445 ;
      RECT 24.713 3.043 24.77 3.445 ;
      RECT 24.627 3.052 24.713 3.445 ;
      RECT 24.541 3.063 24.627 3.445 ;
      RECT 24.455 3.074 24.541 3.445 ;
      RECT 24.435 3.081 24.455 3.453 ;
      RECT 24.425 3.084 24.435 3.46 ;
      RECT 24.36 3.089 24.425 3.478 ;
      RECT 24.33 3.096 24.36 3.503 ;
      RECT 24.32 3.099 24.33 3.51 ;
      RECT 24.275 3.103 24.32 3.515 ;
      RECT 24.245 3.108 24.275 3.52 ;
      RECT 24.244 3.11 24.245 3.52 ;
      RECT 24.158 3.116 24.244 3.52 ;
      RECT 24.072 3.127 24.158 3.52 ;
      RECT 23.986 3.139 24.072 3.52 ;
      RECT 23.9 3.15 23.986 3.52 ;
      RECT 23.885 3.157 23.9 3.515 ;
      RECT 23.88 3.159 23.885 3.509 ;
      RECT 23.86 3.17 23.88 3.504 ;
      RECT 23.85 3.188 23.86 3.498 ;
      RECT 23.845 3.2 23.85 3.298 ;
      RECT 26.14 1.953 26.16 2.04 ;
      RECT 26.135 1.888 26.14 2.072 ;
      RECT 26.125 1.855 26.135 2.077 ;
      RECT 26.12 1.835 26.125 2.083 ;
      RECT 26.09 1.835 26.12 2.1 ;
      RECT 26.041 1.835 26.09 2.136 ;
      RECT 25.955 1.835 26.041 2.194 ;
      RECT 25.926 1.845 25.955 2.243 ;
      RECT 25.84 1.887 25.926 2.296 ;
      RECT 25.82 1.925 25.84 2.343 ;
      RECT 25.795 1.942 25.82 2.363 ;
      RECT 25.785 1.956 25.795 2.383 ;
      RECT 25.78 1.962 25.785 2.393 ;
      RECT 25.775 1.966 25.78 2.4 ;
      RECT 25.725 1.986 25.775 2.405 ;
      RECT 25.66 2.03 25.725 2.405 ;
      RECT 25.635 2.08 25.66 2.405 ;
      RECT 25.625 2.11 25.635 2.405 ;
      RECT 25.62 2.137 25.625 2.405 ;
      RECT 25.615 2.155 25.62 2.405 ;
      RECT 25.605 2.197 25.615 2.405 ;
      RECT 25.955 2.755 26.125 2.93 ;
      RECT 25.895 2.583 25.955 2.918 ;
      RECT 25.885 2.576 25.895 2.901 ;
      RECT 25.84 2.755 26.125 2.881 ;
      RECT 25.821 2.755 26.125 2.859 ;
      RECT 25.735 2.755 26.125 2.824 ;
      RECT 25.715 2.575 25.885 2.78 ;
      RECT 25.715 2.722 26.12 2.78 ;
      RECT 25.715 2.67 26.095 2.78 ;
      RECT 25.715 2.625 26.06 2.78 ;
      RECT 25.715 2.607 26.025 2.78 ;
      RECT 25.715 2.597 26.02 2.78 ;
      RECT 25.885 7.855 26.055 8.305 ;
      RECT 25.94 6.075 26.11 8.025 ;
      RECT 25.885 5.015 26.055 6.245 ;
      RECT 25.365 5.015 25.535 8.305 ;
      RECT 25.365 7.315 25.77 7.645 ;
      RECT 25.365 6.475 25.77 6.805 ;
      RECT 25.435 3.555 25.625 3.78 ;
      RECT 25.425 3.556 25.63 3.775 ;
      RECT 25.425 3.558 25.64 3.755 ;
      RECT 25.425 3.562 25.645 3.74 ;
      RECT 25.425 3.549 25.595 3.775 ;
      RECT 25.425 3.552 25.62 3.775 ;
      RECT 25.435 3.548 25.595 3.78 ;
      RECT 25.521 3.546 25.595 3.78 ;
      RECT 25.145 2.797 25.315 3.035 ;
      RECT 25.145 2.797 25.401 2.949 ;
      RECT 25.145 2.797 25.405 2.859 ;
      RECT 25.195 2.57 25.415 2.838 ;
      RECT 25.19 2.587 25.42 2.811 ;
      RECT 25.155 2.745 25.42 2.811 ;
      RECT 25.175 2.595 25.315 3.035 ;
      RECT 25.165 2.677 25.425 2.794 ;
      RECT 25.16 2.725 25.425 2.794 ;
      RECT 25.165 2.635 25.42 2.811 ;
      RECT 25.19 2.572 25.415 2.838 ;
      RECT 24.755 2.547 24.925 2.745 ;
      RECT 24.755 2.547 24.97 2.72 ;
      RECT 24.825 2.49 24.995 2.678 ;
      RECT 24.8 2.505 24.995 2.678 ;
      RECT 24.415 2.551 24.445 2.745 ;
      RECT 24.41 2.523 24.415 2.745 ;
      RECT 24.38 2.497 24.41 2.747 ;
      RECT 24.355 2.455 24.38 2.75 ;
      RECT 24.345 2.427 24.355 2.752 ;
      RECT 24.31 2.407 24.345 2.754 ;
      RECT 24.245 2.392 24.31 2.76 ;
      RECT 24.195 2.39 24.245 2.766 ;
      RECT 24.172 2.392 24.195 2.771 ;
      RECT 24.086 2.403 24.172 2.777 ;
      RECT 24 2.421 24.086 2.787 ;
      RECT 23.985 2.432 24 2.793 ;
      RECT 23.915 2.455 23.985 2.799 ;
      RECT 23.86 2.487 23.915 2.807 ;
      RECT 23.82 2.51 23.86 2.813 ;
      RECT 23.806 2.523 23.82 2.816 ;
      RECT 23.72 2.545 23.806 2.822 ;
      RECT 23.705 2.57 23.72 2.828 ;
      RECT 23.665 2.585 23.705 2.832 ;
      RECT 23.615 2.6 23.665 2.837 ;
      RECT 23.59 2.607 23.615 2.841 ;
      RECT 23.53 2.602 23.59 2.845 ;
      RECT 23.515 2.593 23.53 2.849 ;
      RECT 23.445 2.583 23.515 2.845 ;
      RECT 23.42 2.575 23.44 2.835 ;
      RECT 23.361 2.575 23.42 2.813 ;
      RECT 23.275 2.575 23.361 2.77 ;
      RECT 23.44 2.575 23.445 2.84 ;
      RECT 24.135 1.806 24.305 2.14 ;
      RECT 24.105 1.806 24.305 2.135 ;
      RECT 24.045 1.773 24.105 2.123 ;
      RECT 24.045 1.829 24.315 2.118 ;
      RECT 24.02 1.829 24.315 2.112 ;
      RECT 24.015 1.77 24.045 2.109 ;
      RECT 24 1.776 24.135 2.107 ;
      RECT 23.995 1.784 24.22 2.095 ;
      RECT 23.995 1.836 24.33 2.048 ;
      RECT 23.98 1.792 24.22 2.043 ;
      RECT 23.98 1.862 24.34 1.984 ;
      RECT 23.95 1.812 24.305 1.945 ;
      RECT 23.95 1.902 24.35 1.941 ;
      RECT 24 1.781 24.22 2.107 ;
      RECT 23.34 2.111 23.395 2.375 ;
      RECT 23.34 2.111 23.46 2.374 ;
      RECT 23.34 2.111 23.485 2.373 ;
      RECT 23.34 2.111 23.55 2.372 ;
      RECT 23.485 2.077 23.565 2.371 ;
      RECT 23.3 2.121 23.71 2.37 ;
      RECT 23.34 2.118 23.71 2.37 ;
      RECT 23.3 2.126 23.715 2.363 ;
      RECT 23.285 2.128 23.715 2.362 ;
      RECT 23.285 2.135 23.72 2.358 ;
      RECT 23.265 2.134 23.715 2.354 ;
      RECT 23.265 2.142 23.725 2.353 ;
      RECT 23.26 2.139 23.72 2.349 ;
      RECT 23.26 2.152 23.735 2.348 ;
      RECT 23.245 2.142 23.725 2.347 ;
      RECT 23.21 2.155 23.735 2.34 ;
      RECT 23.395 2.11 23.705 2.37 ;
      RECT 23.395 2.095 23.655 2.37 ;
      RECT 23.46 2.082 23.59 2.37 ;
      RECT 23.005 3.171 23.02 3.564 ;
      RECT 22.97 3.176 23.02 3.563 ;
      RECT 23.005 3.175 23.065 3.562 ;
      RECT 22.95 3.186 23.065 3.561 ;
      RECT 22.965 3.182 23.065 3.561 ;
      RECT 22.93 3.192 23.14 3.558 ;
      RECT 22.93 3.211 23.185 3.556 ;
      RECT 22.93 3.218 23.19 3.553 ;
      RECT 22.915 3.195 23.14 3.55 ;
      RECT 22.895 3.2 23.14 3.543 ;
      RECT 22.89 3.204 23.14 3.539 ;
      RECT 22.89 3.221 23.2 3.538 ;
      RECT 22.87 3.215 23.185 3.534 ;
      RECT 22.87 3.224 23.205 3.528 ;
      RECT 22.865 3.23 23.205 3.3 ;
      RECT 22.93 3.19 23.065 3.558 ;
      RECT 22.805 2.553 23.005 2.865 ;
      RECT 22.88 2.531 23.005 2.865 ;
      RECT 22.82 2.55 23.01 2.85 ;
      RECT 22.79 2.561 23.01 2.848 ;
      RECT 22.805 2.556 23.015 2.814 ;
      RECT 22.79 2.66 23.02 2.781 ;
      RECT 22.82 2.532 23.005 2.865 ;
      RECT 22.88 2.51 22.98 2.865 ;
      RECT 22.905 2.507 22.98 2.865 ;
      RECT 22.905 2.502 22.925 2.865 ;
      RECT 22.31 2.57 22.485 2.745 ;
      RECT 22.305 2.57 22.485 2.743 ;
      RECT 22.28 2.57 22.485 2.738 ;
      RECT 22.225 2.55 22.395 2.728 ;
      RECT 22.225 2.557 22.46 2.728 ;
      RECT 22.31 3.237 22.325 3.42 ;
      RECT 22.3 3.215 22.31 3.42 ;
      RECT 22.285 3.195 22.3 3.42 ;
      RECT 22.275 3.17 22.285 3.42 ;
      RECT 22.245 3.135 22.275 3.42 ;
      RECT 22.21 3.075 22.245 3.42 ;
      RECT 22.205 3.037 22.21 3.42 ;
      RECT 22.155 2.988 22.205 3.42 ;
      RECT 22.145 2.938 22.155 3.408 ;
      RECT 22.13 2.917 22.145 3.368 ;
      RECT 22.11 2.885 22.13 3.318 ;
      RECT 22.085 2.841 22.11 3.258 ;
      RECT 22.08 2.813 22.085 3.213 ;
      RECT 22.075 2.804 22.08 3.199 ;
      RECT 22.07 2.797 22.075 3.186 ;
      RECT 22.065 2.792 22.07 3.175 ;
      RECT 22.06 2.777 22.065 3.165 ;
      RECT 22.055 2.755 22.06 3.152 ;
      RECT 22.045 2.715 22.055 3.127 ;
      RECT 22.02 2.645 22.045 3.083 ;
      RECT 22.015 2.585 22.02 3.048 ;
      RECT 22 2.565 22.015 3.015 ;
      RECT 21.995 2.565 22 2.99 ;
      RECT 21.965 2.565 21.995 2.945 ;
      RECT 21.92 2.565 21.965 2.885 ;
      RECT 21.845 2.565 21.92 2.833 ;
      RECT 21.84 2.565 21.845 2.798 ;
      RECT 21.835 2.565 21.84 2.788 ;
      RECT 21.83 2.565 21.835 2.768 ;
      RECT 22.095 1.785 22.265 2.255 ;
      RECT 22.04 1.778 22.235 2.239 ;
      RECT 22.04 1.792 22.27 2.238 ;
      RECT 22.025 1.793 22.27 2.219 ;
      RECT 22.02 1.811 22.27 2.205 ;
      RECT 22.025 1.794 22.275 2.203 ;
      RECT 22.01 1.825 22.275 2.188 ;
      RECT 22.025 1.8 22.28 2.173 ;
      RECT 22.005 1.84 22.28 2.17 ;
      RECT 22.02 1.812 22.285 2.155 ;
      RECT 22.02 1.824 22.29 2.135 ;
      RECT 22.005 1.84 22.295 2.118 ;
      RECT 22.005 1.85 22.3 1.973 ;
      RECT 22 1.85 22.3 1.93 ;
      RECT 22 1.865 22.305 1.908 ;
      RECT 22.095 1.775 22.235 2.255 ;
      RECT 22.095 1.773 22.205 2.255 ;
      RECT 22.181 1.77 22.205 2.255 ;
      RECT 21.84 3.437 21.845 3.483 ;
      RECT 21.83 3.285 21.84 3.507 ;
      RECT 21.825 3.13 21.83 3.532 ;
      RECT 21.81 3.092 21.825 3.543 ;
      RECT 21.805 3.075 21.81 3.55 ;
      RECT 21.795 3.063 21.805 3.557 ;
      RECT 21.79 3.054 21.795 3.559 ;
      RECT 21.785 3.052 21.79 3.563 ;
      RECT 21.74 3.043 21.785 3.578 ;
      RECT 21.735 3.035 21.74 3.592 ;
      RECT 21.73 3.032 21.735 3.596 ;
      RECT 21.715 3.027 21.73 3.604 ;
      RECT 21.66 3.017 21.715 3.615 ;
      RECT 21.625 3.005 21.66 3.616 ;
      RECT 21.616 3 21.625 3.61 ;
      RECT 21.53 3 21.616 3.6 ;
      RECT 21.5 3 21.53 3.578 ;
      RECT 21.49 3 21.495 3.558 ;
      RECT 21.485 3 21.49 3.52 ;
      RECT 21.48 3 21.485 3.478 ;
      RECT 21.475 3 21.48 3.438 ;
      RECT 21.47 3 21.475 3.368 ;
      RECT 21.46 3 21.47 3.29 ;
      RECT 21.455 3 21.46 3.19 ;
      RECT 21.495 3 21.5 3.56 ;
      RECT 20.99 3.082 21.08 3.56 ;
      RECT 20.975 3.085 21.095 3.558 ;
      RECT 20.99 3.084 21.095 3.558 ;
      RECT 20.955 3.091 21.12 3.548 ;
      RECT 20.975 3.085 21.12 3.548 ;
      RECT 20.94 3.097 21.12 3.536 ;
      RECT 20.975 3.088 21.17 3.529 ;
      RECT 20.926 3.105 21.17 3.527 ;
      RECT 20.955 3.095 21.18 3.515 ;
      RECT 20.926 3.116 21.21 3.506 ;
      RECT 20.84 3.14 21.21 3.5 ;
      RECT 20.84 3.153 21.25 3.483 ;
      RECT 20.835 3.175 21.25 3.476 ;
      RECT 20.805 3.19 21.25 3.466 ;
      RECT 20.8 3.201 21.25 3.456 ;
      RECT 20.77 3.214 21.25 3.447 ;
      RECT 20.755 3.232 21.25 3.436 ;
      RECT 20.73 3.245 21.25 3.426 ;
      RECT 20.99 3.081 21 3.56 ;
      RECT 21.036 2.505 21.075 2.75 ;
      RECT 20.95 2.505 21.085 2.748 ;
      RECT 20.835 2.53 21.085 2.745 ;
      RECT 20.835 2.53 21.09 2.743 ;
      RECT 20.835 2.53 21.105 2.738 ;
      RECT 20.941 2.505 21.12 2.718 ;
      RECT 20.855 2.513 21.12 2.718 ;
      RECT 20.525 1.865 20.695 2.3 ;
      RECT 20.515 1.899 20.695 2.283 ;
      RECT 20.595 1.835 20.765 2.27 ;
      RECT 20.5 1.91 20.765 2.248 ;
      RECT 20.595 1.845 20.77 2.238 ;
      RECT 20.525 1.897 20.8 2.223 ;
      RECT 20.485 1.923 20.8 2.208 ;
      RECT 20.485 1.965 20.81 2.188 ;
      RECT 20.48 1.99 20.815 2.17 ;
      RECT 20.48 2 20.82 2.155 ;
      RECT 20.475 1.937 20.8 2.153 ;
      RECT 20.475 2.01 20.825 2.138 ;
      RECT 20.47 1.947 20.8 2.135 ;
      RECT 20.465 2.031 20.83 2.118 ;
      RECT 20.465 2.063 20.835 2.098 ;
      RECT 20.46 1.977 20.81 2.09 ;
      RECT 20.465 1.962 20.8 2.118 ;
      RECT 20.48 1.932 20.8 2.17 ;
      RECT 20.325 2.519 20.55 2.775 ;
      RECT 20.325 2.552 20.57 2.765 ;
      RECT 20.29 2.552 20.57 2.763 ;
      RECT 20.29 2.565 20.575 2.753 ;
      RECT 20.29 2.585 20.585 2.745 ;
      RECT 20.29 2.682 20.59 2.738 ;
      RECT 20.27 2.43 20.4 2.728 ;
      RECT 20.225 2.585 20.585 2.67 ;
      RECT 20.215 2.43 20.4 2.615 ;
      RECT 20.215 2.462 20.486 2.615 ;
      RECT 20.18 2.992 20.2 3.17 ;
      RECT 20.145 2.945 20.18 3.17 ;
      RECT 20.13 2.885 20.145 3.17 ;
      RECT 20.105 2.832 20.13 3.17 ;
      RECT 20.09 2.785 20.105 3.17 ;
      RECT 20.07 2.762 20.09 3.17 ;
      RECT 20.045 2.727 20.07 3.17 ;
      RECT 20.035 2.573 20.045 3.17 ;
      RECT 20.005 2.568 20.035 3.161 ;
      RECT 20 2.565 20.005 3.151 ;
      RECT 19.985 2.565 20 3.125 ;
      RECT 19.98 2.565 19.985 3.088 ;
      RECT 19.955 2.565 19.98 3.04 ;
      RECT 19.935 2.565 19.955 2.965 ;
      RECT 19.925 2.565 19.935 2.925 ;
      RECT 19.92 2.565 19.925 2.9 ;
      RECT 19.915 2.565 19.92 2.883 ;
      RECT 19.91 2.565 19.915 2.865 ;
      RECT 19.905 2.566 19.91 2.855 ;
      RECT 19.895 2.568 19.905 2.823 ;
      RECT 19.885 2.57 19.895 2.79 ;
      RECT 19.875 2.573 19.885 2.763 ;
      RECT 20.2 3 20.425 3.17 ;
      RECT 19.53 1.812 19.7 2.265 ;
      RECT 19.53 1.812 19.79 2.231 ;
      RECT 19.53 1.812 19.82 2.215 ;
      RECT 19.53 1.812 19.85 2.188 ;
      RECT 19.786 1.79 19.865 2.17 ;
      RECT 19.565 1.797 19.87 2.155 ;
      RECT 19.565 1.805 19.88 2.118 ;
      RECT 19.525 1.832 19.88 2.09 ;
      RECT 19.51 1.845 19.88 2.055 ;
      RECT 19.53 1.82 19.9 2.045 ;
      RECT 19.505 1.885 19.9 2.015 ;
      RECT 19.505 1.915 19.905 1.998 ;
      RECT 19.5 1.945 19.905 1.985 ;
      RECT 19.565 1.794 19.865 2.17 ;
      RECT 19.7 1.791 19.786 2.249 ;
      RECT 19.651 1.792 19.865 2.17 ;
      RECT 19.795 3.452 19.84 3.645 ;
      RECT 19.785 3.422 19.795 3.645 ;
      RECT 19.78 3.407 19.785 3.645 ;
      RECT 19.74 3.317 19.78 3.645 ;
      RECT 19.735 3.23 19.74 3.645 ;
      RECT 19.725 3.2 19.735 3.645 ;
      RECT 19.72 3.16 19.725 3.645 ;
      RECT 19.71 3.122 19.72 3.645 ;
      RECT 19.705 3.087 19.71 3.645 ;
      RECT 19.685 3.04 19.705 3.645 ;
      RECT 19.67 2.965 19.685 3.645 ;
      RECT 19.665 2.92 19.67 3.64 ;
      RECT 19.66 2.9 19.665 3.613 ;
      RECT 19.655 2.88 19.66 3.598 ;
      RECT 19.65 2.855 19.655 3.578 ;
      RECT 19.645 2.833 19.65 3.563 ;
      RECT 19.64 2.811 19.645 3.545 ;
      RECT 19.635 2.79 19.64 3.535 ;
      RECT 19.625 2.762 19.635 3.505 ;
      RECT 19.615 2.725 19.625 3.473 ;
      RECT 19.605 2.685 19.615 3.44 ;
      RECT 19.595 2.663 19.605 3.41 ;
      RECT 19.565 2.615 19.595 3.342 ;
      RECT 19.55 2.575 19.565 3.269 ;
      RECT 19.54 2.575 19.55 3.235 ;
      RECT 19.535 2.575 19.54 3.21 ;
      RECT 19.53 2.575 19.535 3.195 ;
      RECT 19.525 2.575 19.53 3.173 ;
      RECT 19.52 2.575 19.525 3.16 ;
      RECT 19.505 2.575 19.52 3.125 ;
      RECT 19.485 2.575 19.505 3.065 ;
      RECT 19.475 2.575 19.485 3.015 ;
      RECT 19.455 2.575 19.475 2.963 ;
      RECT 19.435 2.575 19.455 2.92 ;
      RECT 19.425 2.575 19.435 2.908 ;
      RECT 19.395 2.575 19.425 2.895 ;
      RECT 19.365 2.596 19.395 2.875 ;
      RECT 19.355 2.624 19.365 2.855 ;
      RECT 19.34 2.641 19.355 2.823 ;
      RECT 19.335 2.655 19.34 2.79 ;
      RECT 19.33 2.663 19.335 2.763 ;
      RECT 19.325 2.671 19.33 2.725 ;
      RECT 19.33 3.195 19.335 3.53 ;
      RECT 19.295 3.182 19.33 3.529 ;
      RECT 19.225 3.122 19.295 3.528 ;
      RECT 19.145 3.065 19.225 3.527 ;
      RECT 19.01 3.025 19.145 3.526 ;
      RECT 19.01 3.212 19.345 3.515 ;
      RECT 18.97 3.212 19.345 3.505 ;
      RECT 18.97 3.23 19.35 3.5 ;
      RECT 18.97 3.32 19.355 3.49 ;
      RECT 18.965 3.015 19.13 3.47 ;
      RECT 18.96 3.015 19.13 3.213 ;
      RECT 18.96 3.172 19.325 3.213 ;
      RECT 18.96 3.16 19.32 3.213 ;
      RECT 18.095 5.02 18.265 6.49 ;
      RECT 18.095 6.315 18.27 6.485 ;
      RECT 17.725 1.74 17.895 2.93 ;
      RECT 17.725 1.74 18.195 1.91 ;
      RECT 17.725 6.97 18.195 7.14 ;
      RECT 17.725 5.95 17.895 7.14 ;
      RECT 16.735 1.74 16.905 2.93 ;
      RECT 16.735 1.74 17.205 1.91 ;
      RECT 16.735 6.97 17.205 7.14 ;
      RECT 16.735 5.95 16.905 7.14 ;
      RECT 14.885 2.635 15.055 3.865 ;
      RECT 14.94 0.855 15.11 2.805 ;
      RECT 14.885 0.575 15.055 1.025 ;
      RECT 14.885 7.855 15.055 8.305 ;
      RECT 14.94 6.075 15.11 8.025 ;
      RECT 14.885 5.015 15.055 6.245 ;
      RECT 14.365 0.575 14.535 3.865 ;
      RECT 14.365 2.075 14.77 2.405 ;
      RECT 14.365 1.235 14.77 1.565 ;
      RECT 14.365 5.015 14.535 8.305 ;
      RECT 14.365 7.315 14.77 7.645 ;
      RECT 14.365 6.475 14.77 6.805 ;
      RECT 11.7 1.975 12.43 2.215 ;
      RECT 12.242 1.77 12.43 2.215 ;
      RECT 12.07 1.782 12.445 2.209 ;
      RECT 11.985 1.797 12.465 2.194 ;
      RECT 11.985 1.812 12.47 2.184 ;
      RECT 11.94 1.832 12.485 2.176 ;
      RECT 11.917 1.867 12.5 2.13 ;
      RECT 11.831 1.89 12.505 2.09 ;
      RECT 11.831 1.908 12.515 2.06 ;
      RECT 11.7 1.977 12.52 2.023 ;
      RECT 11.745 1.92 12.515 2.06 ;
      RECT 11.831 1.872 12.5 2.13 ;
      RECT 11.917 1.841 12.485 2.176 ;
      RECT 11.94 1.822 12.47 2.184 ;
      RECT 11.985 1.795 12.445 2.209 ;
      RECT 12.07 1.777 12.43 2.215 ;
      RECT 12.156 1.771 12.43 2.215 ;
      RECT 12.242 1.766 12.375 2.215 ;
      RECT 12.328 1.761 12.375 2.215 ;
      RECT 12.02 2.659 12.19 3.045 ;
      RECT 12.015 2.659 12.19 3.04 ;
      RECT 11.99 2.659 12.19 3.005 ;
      RECT 11.99 2.687 12.2 2.995 ;
      RECT 11.97 2.687 12.2 2.955 ;
      RECT 11.965 2.687 12.2 2.928 ;
      RECT 11.965 2.705 12.205 2.92 ;
      RECT 11.91 2.705 12.205 2.855 ;
      RECT 11.91 2.722 12.215 2.838 ;
      RECT 11.9 2.722 12.215 2.778 ;
      RECT 11.9 2.739 12.22 2.775 ;
      RECT 11.895 2.575 12.065 2.753 ;
      RECT 11.895 2.609 12.151 2.753 ;
      RECT 11.89 3.375 11.895 3.388 ;
      RECT 11.885 3.27 11.89 3.393 ;
      RECT 11.86 3.13 11.885 3.408 ;
      RECT 11.825 3.081 11.86 3.44 ;
      RECT 11.82 3.049 11.825 3.46 ;
      RECT 11.815 3.04 11.82 3.46 ;
      RECT 11.735 3.005 11.815 3.46 ;
      RECT 11.672 2.975 11.735 3.46 ;
      RECT 11.586 2.963 11.672 3.46 ;
      RECT 11.5 2.949 11.586 3.46 ;
      RECT 11.42 2.936 11.5 3.446 ;
      RECT 11.385 2.928 11.42 3.426 ;
      RECT 11.375 2.925 11.385 3.417 ;
      RECT 11.345 2.92 11.375 3.404 ;
      RECT 11.295 2.895 11.345 3.38 ;
      RECT 11.281 2.869 11.295 3.362 ;
      RECT 11.195 2.829 11.281 3.338 ;
      RECT 11.15 2.777 11.195 3.307 ;
      RECT 11.14 2.752 11.15 3.294 ;
      RECT 11.135 2.533 11.14 2.555 ;
      RECT 11.13 2.735 11.14 3.29 ;
      RECT 11.13 2.531 11.135 2.645 ;
      RECT 11.12 2.527 11.13 3.286 ;
      RECT 11.076 2.525 11.12 3.274 ;
      RECT 10.99 2.525 11.076 3.245 ;
      RECT 10.96 2.525 10.99 3.218 ;
      RECT 10.945 2.525 10.96 3.206 ;
      RECT 10.905 2.537 10.945 3.191 ;
      RECT 10.885 2.556 10.905 3.17 ;
      RECT 10.875 2.566 10.885 3.154 ;
      RECT 10.865 2.572 10.875 3.143 ;
      RECT 10.845 2.582 10.865 3.126 ;
      RECT 10.84 2.591 10.845 3.113 ;
      RECT 10.835 2.595 10.84 3.063 ;
      RECT 10.825 2.601 10.835 2.98 ;
      RECT 10.82 2.605 10.825 2.894 ;
      RECT 10.815 2.625 10.82 2.831 ;
      RECT 10.81 2.648 10.815 2.778 ;
      RECT 10.805 2.666 10.81 2.723 ;
      RECT 11.415 2.485 11.585 2.745 ;
      RECT 11.585 2.45 11.63 2.731 ;
      RECT 11.546 2.452 11.635 2.714 ;
      RECT 11.435 2.469 11.721 2.685 ;
      RECT 11.435 2.484 11.725 2.657 ;
      RECT 11.435 2.465 11.635 2.714 ;
      RECT 11.46 2.453 11.585 2.745 ;
      RECT 11.546 2.451 11.63 2.731 ;
      RECT 10.6 1.84 10.77 2.33 ;
      RECT 10.6 1.84 10.805 2.31 ;
      RECT 10.735 1.76 10.845 2.27 ;
      RECT 10.716 1.764 10.865 2.24 ;
      RECT 10.63 1.772 10.885 2.223 ;
      RECT 10.63 1.778 10.89 2.213 ;
      RECT 10.63 1.787 10.91 2.201 ;
      RECT 10.605 1.812 10.94 2.179 ;
      RECT 10.605 1.832 10.945 2.159 ;
      RECT 10.6 1.845 10.955 2.139 ;
      RECT 10.6 1.912 10.96 2.12 ;
      RECT 10.6 2.045 10.965 2.107 ;
      RECT 10.595 1.85 10.955 1.94 ;
      RECT 10.605 1.807 10.91 2.201 ;
      RECT 10.716 1.762 10.845 2.27 ;
      RECT 10.59 3.515 10.89 3.77 ;
      RECT 10.675 3.481 10.89 3.77 ;
      RECT 10.675 3.484 10.895 3.63 ;
      RECT 10.61 3.505 10.895 3.63 ;
      RECT 10.645 3.495 10.89 3.77 ;
      RECT 10.64 3.5 10.895 3.63 ;
      RECT 10.675 3.479 10.876 3.77 ;
      RECT 10.761 3.47 10.876 3.77 ;
      RECT 10.761 3.464 10.79 3.77 ;
      RECT 10.25 3.105 10.26 3.595 ;
      RECT 9.91 3.04 9.92 3.34 ;
      RECT 10.425 3.212 10.43 3.431 ;
      RECT 10.415 3.192 10.425 3.448 ;
      RECT 10.405 3.172 10.415 3.478 ;
      RECT 10.4 3.162 10.405 3.493 ;
      RECT 10.395 3.158 10.4 3.498 ;
      RECT 10.38 3.15 10.395 3.505 ;
      RECT 10.34 3.13 10.38 3.53 ;
      RECT 10.315 3.112 10.34 3.563 ;
      RECT 10.31 3.11 10.315 3.576 ;
      RECT 10.29 3.107 10.31 3.58 ;
      RECT 10.26 3.105 10.29 3.59 ;
      RECT 10.19 3.107 10.25 3.591 ;
      RECT 10.17 3.107 10.19 3.585 ;
      RECT 10.145 3.105 10.17 3.582 ;
      RECT 10.11 3.1 10.145 3.578 ;
      RECT 10.09 3.094 10.11 3.565 ;
      RECT 10.08 3.091 10.09 3.553 ;
      RECT 10.06 3.088 10.08 3.538 ;
      RECT 10.04 3.084 10.06 3.52 ;
      RECT 10.035 3.081 10.04 3.51 ;
      RECT 10.03 3.08 10.035 3.508 ;
      RECT 10.02 3.077 10.03 3.5 ;
      RECT 10.01 3.071 10.02 3.483 ;
      RECT 10 3.065 10.01 3.465 ;
      RECT 9.99 3.059 10 3.453 ;
      RECT 9.98 3.053 9.99 3.433 ;
      RECT 9.975 3.049 9.98 3.418 ;
      RECT 9.97 3.047 9.975 3.41 ;
      RECT 9.965 3.045 9.97 3.403 ;
      RECT 9.96 3.043 9.965 3.393 ;
      RECT 9.955 3.041 9.96 3.387 ;
      RECT 9.945 3.04 9.955 3.377 ;
      RECT 9.935 3.04 9.945 3.368 ;
      RECT 9.92 3.04 9.935 3.353 ;
      RECT 9.88 3.04 9.91 3.337 ;
      RECT 9.86 3.042 9.88 3.332 ;
      RECT 9.855 3.047 9.86 3.33 ;
      RECT 9.825 3.055 9.855 3.328 ;
      RECT 9.795 3.07 9.825 3.327 ;
      RECT 9.75 3.092 9.795 3.332 ;
      RECT 9.745 3.107 9.75 3.336 ;
      RECT 9.73 3.112 9.745 3.338 ;
      RECT 9.725 3.116 9.73 3.34 ;
      RECT 9.665 3.139 9.725 3.349 ;
      RECT 9.645 3.165 9.665 3.362 ;
      RECT 9.635 3.172 9.645 3.366 ;
      RECT 9.62 3.179 9.635 3.369 ;
      RECT 9.6 3.189 9.62 3.372 ;
      RECT 9.595 3.197 9.6 3.375 ;
      RECT 9.55 3.202 9.595 3.382 ;
      RECT 9.54 3.205 9.55 3.389 ;
      RECT 9.53 3.205 9.54 3.393 ;
      RECT 9.495 3.207 9.53 3.405 ;
      RECT 9.475 3.21 9.495 3.418 ;
      RECT 9.435 3.213 9.475 3.429 ;
      RECT 9.42 3.215 9.435 3.442 ;
      RECT 9.41 3.215 9.42 3.447 ;
      RECT 9.385 3.216 9.41 3.455 ;
      RECT 9.375 3.218 9.385 3.46 ;
      RECT 9.37 3.219 9.375 3.463 ;
      RECT 9.345 3.217 9.37 3.466 ;
      RECT 9.33 3.215 9.345 3.467 ;
      RECT 9.31 3.212 9.33 3.469 ;
      RECT 9.29 3.207 9.31 3.469 ;
      RECT 9.23 3.202 9.29 3.466 ;
      RECT 9.195 3.177 9.23 3.462 ;
      RECT 9.185 3.154 9.195 3.46 ;
      RECT 9.155 3.131 9.185 3.46 ;
      RECT 9.145 3.11 9.155 3.46 ;
      RECT 9.12 3.092 9.145 3.458 ;
      RECT 9.105 3.07 9.12 3.455 ;
      RECT 9.09 3.052 9.105 3.453 ;
      RECT 9.07 3.042 9.09 3.451 ;
      RECT 9.055 3.037 9.07 3.45 ;
      RECT 9.04 3.035 9.055 3.449 ;
      RECT 9.01 3.036 9.04 3.447 ;
      RECT 8.99 3.039 9.01 3.445 ;
      RECT 8.933 3.043 8.99 3.445 ;
      RECT 8.847 3.052 8.933 3.445 ;
      RECT 8.761 3.063 8.847 3.445 ;
      RECT 8.675 3.074 8.761 3.445 ;
      RECT 8.655 3.081 8.675 3.453 ;
      RECT 8.645 3.084 8.655 3.46 ;
      RECT 8.58 3.089 8.645 3.478 ;
      RECT 8.55 3.096 8.58 3.503 ;
      RECT 8.54 3.099 8.55 3.51 ;
      RECT 8.495 3.103 8.54 3.515 ;
      RECT 8.465 3.108 8.495 3.52 ;
      RECT 8.464 3.11 8.465 3.52 ;
      RECT 8.378 3.116 8.464 3.52 ;
      RECT 8.292 3.127 8.378 3.52 ;
      RECT 8.206 3.139 8.292 3.52 ;
      RECT 8.12 3.15 8.206 3.52 ;
      RECT 8.105 3.157 8.12 3.515 ;
      RECT 8.1 3.159 8.105 3.509 ;
      RECT 8.08 3.17 8.1 3.504 ;
      RECT 8.07 3.188 8.08 3.498 ;
      RECT 8.065 3.2 8.07 3.298 ;
      RECT 10.36 1.953 10.38 2.04 ;
      RECT 10.355 1.888 10.36 2.072 ;
      RECT 10.345 1.855 10.355 2.077 ;
      RECT 10.34 1.835 10.345 2.083 ;
      RECT 10.31 1.835 10.34 2.1 ;
      RECT 10.261 1.835 10.31 2.136 ;
      RECT 10.175 1.835 10.261 2.194 ;
      RECT 10.146 1.845 10.175 2.243 ;
      RECT 10.06 1.887 10.146 2.296 ;
      RECT 10.04 1.925 10.06 2.343 ;
      RECT 10.015 1.942 10.04 2.363 ;
      RECT 10.005 1.956 10.015 2.383 ;
      RECT 10 1.962 10.005 2.393 ;
      RECT 9.995 1.966 10 2.4 ;
      RECT 9.945 1.986 9.995 2.405 ;
      RECT 9.88 2.03 9.945 2.405 ;
      RECT 9.855 2.08 9.88 2.405 ;
      RECT 9.845 2.11 9.855 2.405 ;
      RECT 9.84 2.137 9.845 2.405 ;
      RECT 9.835 2.155 9.84 2.405 ;
      RECT 9.825 2.197 9.835 2.405 ;
      RECT 10.175 2.755 10.345 2.93 ;
      RECT 10.115 2.583 10.175 2.918 ;
      RECT 10.105 2.576 10.115 2.901 ;
      RECT 10.06 2.755 10.345 2.881 ;
      RECT 10.041 2.755 10.345 2.859 ;
      RECT 9.955 2.755 10.345 2.824 ;
      RECT 9.935 2.575 10.105 2.78 ;
      RECT 9.935 2.722 10.34 2.78 ;
      RECT 9.935 2.67 10.315 2.78 ;
      RECT 9.935 2.625 10.28 2.78 ;
      RECT 9.935 2.607 10.245 2.78 ;
      RECT 9.935 2.597 10.24 2.78 ;
      RECT 10.105 7.855 10.275 8.305 ;
      RECT 10.16 6.075 10.33 8.025 ;
      RECT 10.105 5.015 10.275 6.245 ;
      RECT 9.585 5.015 9.755 8.305 ;
      RECT 9.585 7.315 9.99 7.645 ;
      RECT 9.585 6.475 9.99 6.805 ;
      RECT 9.655 3.555 9.845 3.78 ;
      RECT 9.645 3.556 9.85 3.775 ;
      RECT 9.645 3.558 9.86 3.755 ;
      RECT 9.645 3.562 9.865 3.74 ;
      RECT 9.645 3.549 9.815 3.775 ;
      RECT 9.645 3.552 9.84 3.775 ;
      RECT 9.655 3.548 9.815 3.78 ;
      RECT 9.741 3.546 9.815 3.78 ;
      RECT 9.365 2.797 9.535 3.035 ;
      RECT 9.365 2.797 9.621 2.949 ;
      RECT 9.365 2.797 9.625 2.859 ;
      RECT 9.415 2.57 9.635 2.838 ;
      RECT 9.41 2.587 9.64 2.811 ;
      RECT 9.375 2.745 9.64 2.811 ;
      RECT 9.395 2.595 9.535 3.035 ;
      RECT 9.385 2.677 9.645 2.794 ;
      RECT 9.38 2.725 9.645 2.794 ;
      RECT 9.385 2.635 9.64 2.811 ;
      RECT 9.41 2.572 9.635 2.838 ;
      RECT 8.975 2.547 9.145 2.745 ;
      RECT 8.975 2.547 9.19 2.72 ;
      RECT 9.045 2.49 9.215 2.678 ;
      RECT 9.02 2.505 9.215 2.678 ;
      RECT 8.635 2.551 8.665 2.745 ;
      RECT 8.63 2.523 8.635 2.745 ;
      RECT 8.6 2.497 8.63 2.747 ;
      RECT 8.575 2.455 8.6 2.75 ;
      RECT 8.565 2.427 8.575 2.752 ;
      RECT 8.53 2.407 8.565 2.754 ;
      RECT 8.465 2.392 8.53 2.76 ;
      RECT 8.415 2.39 8.465 2.766 ;
      RECT 8.392 2.392 8.415 2.771 ;
      RECT 8.306 2.403 8.392 2.777 ;
      RECT 8.22 2.421 8.306 2.787 ;
      RECT 8.205 2.432 8.22 2.793 ;
      RECT 8.135 2.455 8.205 2.799 ;
      RECT 8.08 2.487 8.135 2.807 ;
      RECT 8.04 2.51 8.08 2.813 ;
      RECT 8.026 2.523 8.04 2.816 ;
      RECT 7.94 2.545 8.026 2.822 ;
      RECT 7.925 2.57 7.94 2.828 ;
      RECT 7.885 2.585 7.925 2.832 ;
      RECT 7.835 2.6 7.885 2.837 ;
      RECT 7.81 2.607 7.835 2.841 ;
      RECT 7.75 2.602 7.81 2.845 ;
      RECT 7.735 2.593 7.75 2.849 ;
      RECT 7.665 2.583 7.735 2.845 ;
      RECT 7.64 2.575 7.66 2.835 ;
      RECT 7.581 2.575 7.64 2.813 ;
      RECT 7.495 2.575 7.581 2.77 ;
      RECT 7.66 2.575 7.665 2.84 ;
      RECT 8.355 1.806 8.525 2.14 ;
      RECT 8.325 1.806 8.525 2.135 ;
      RECT 8.265 1.773 8.325 2.123 ;
      RECT 8.265 1.829 8.535 2.118 ;
      RECT 8.24 1.829 8.535 2.112 ;
      RECT 8.235 1.77 8.265 2.109 ;
      RECT 8.22 1.776 8.355 2.107 ;
      RECT 8.215 1.784 8.44 2.095 ;
      RECT 8.215 1.836 8.55 2.048 ;
      RECT 8.2 1.792 8.44 2.043 ;
      RECT 8.2 1.862 8.56 1.984 ;
      RECT 8.17 1.812 8.525 1.945 ;
      RECT 8.17 1.902 8.57 1.941 ;
      RECT 8.22 1.781 8.44 2.107 ;
      RECT 7.56 2.111 7.615 2.375 ;
      RECT 7.56 2.111 7.68 2.374 ;
      RECT 7.56 2.111 7.705 2.373 ;
      RECT 7.56 2.111 7.77 2.372 ;
      RECT 7.705 2.077 7.785 2.371 ;
      RECT 7.52 2.121 7.93 2.37 ;
      RECT 7.56 2.118 7.93 2.37 ;
      RECT 7.52 2.126 7.935 2.363 ;
      RECT 7.505 2.128 7.935 2.362 ;
      RECT 7.505 2.135 7.94 2.358 ;
      RECT 7.485 2.134 7.935 2.354 ;
      RECT 7.485 2.142 7.945 2.353 ;
      RECT 7.48 2.139 7.94 2.349 ;
      RECT 7.48 2.152 7.955 2.348 ;
      RECT 7.465 2.142 7.945 2.347 ;
      RECT 7.43 2.155 7.955 2.34 ;
      RECT 7.615 2.11 7.925 2.37 ;
      RECT 7.615 2.095 7.875 2.37 ;
      RECT 7.68 2.082 7.81 2.37 ;
      RECT 7.225 3.171 7.24 3.564 ;
      RECT 7.19 3.176 7.24 3.563 ;
      RECT 7.225 3.175 7.285 3.562 ;
      RECT 7.17 3.186 7.285 3.561 ;
      RECT 7.185 3.182 7.285 3.561 ;
      RECT 7.15 3.192 7.36 3.558 ;
      RECT 7.15 3.211 7.405 3.556 ;
      RECT 7.15 3.218 7.41 3.553 ;
      RECT 7.135 3.195 7.36 3.55 ;
      RECT 7.115 3.2 7.36 3.543 ;
      RECT 7.11 3.204 7.36 3.539 ;
      RECT 7.11 3.221 7.42 3.538 ;
      RECT 7.09 3.215 7.405 3.534 ;
      RECT 7.09 3.224 7.425 3.528 ;
      RECT 7.085 3.23 7.425 3.3 ;
      RECT 7.15 3.19 7.285 3.558 ;
      RECT 7.025 2.553 7.225 2.865 ;
      RECT 7.1 2.531 7.225 2.865 ;
      RECT 7.04 2.55 7.23 2.85 ;
      RECT 7.01 2.561 7.23 2.848 ;
      RECT 7.025 2.556 7.235 2.814 ;
      RECT 7.01 2.66 7.24 2.781 ;
      RECT 7.04 2.532 7.225 2.865 ;
      RECT 7.1 2.51 7.2 2.865 ;
      RECT 7.125 2.507 7.2 2.865 ;
      RECT 7.125 2.502 7.145 2.865 ;
      RECT 6.53 2.57 6.705 2.745 ;
      RECT 6.525 2.57 6.705 2.743 ;
      RECT 6.5 2.57 6.705 2.738 ;
      RECT 6.445 2.55 6.615 2.728 ;
      RECT 6.445 2.557 6.68 2.728 ;
      RECT 6.53 3.237 6.545 3.42 ;
      RECT 6.52 3.215 6.53 3.42 ;
      RECT 6.505 3.195 6.52 3.42 ;
      RECT 6.495 3.17 6.505 3.42 ;
      RECT 6.465 3.135 6.495 3.42 ;
      RECT 6.43 3.075 6.465 3.42 ;
      RECT 6.425 3.037 6.43 3.42 ;
      RECT 6.375 2.988 6.425 3.42 ;
      RECT 6.365 2.938 6.375 3.408 ;
      RECT 6.35 2.917 6.365 3.368 ;
      RECT 6.33 2.885 6.35 3.318 ;
      RECT 6.305 2.841 6.33 3.258 ;
      RECT 6.3 2.813 6.305 3.213 ;
      RECT 6.295 2.804 6.3 3.199 ;
      RECT 6.29 2.797 6.295 3.186 ;
      RECT 6.285 2.792 6.29 3.175 ;
      RECT 6.28 2.777 6.285 3.165 ;
      RECT 6.275 2.755 6.28 3.152 ;
      RECT 6.265 2.715 6.275 3.127 ;
      RECT 6.24 2.645 6.265 3.083 ;
      RECT 6.235 2.585 6.24 3.048 ;
      RECT 6.22 2.565 6.235 3.015 ;
      RECT 6.215 2.565 6.22 2.99 ;
      RECT 6.185 2.565 6.215 2.945 ;
      RECT 6.14 2.565 6.185 2.885 ;
      RECT 6.065 2.565 6.14 2.833 ;
      RECT 6.06 2.565 6.065 2.798 ;
      RECT 6.055 2.565 6.06 2.788 ;
      RECT 6.05 2.565 6.055 2.768 ;
      RECT 6.315 1.785 6.485 2.255 ;
      RECT 6.26 1.778 6.455 2.239 ;
      RECT 6.26 1.792 6.49 2.238 ;
      RECT 6.245 1.793 6.49 2.219 ;
      RECT 6.24 1.811 6.49 2.205 ;
      RECT 6.245 1.794 6.495 2.203 ;
      RECT 6.23 1.825 6.495 2.188 ;
      RECT 6.245 1.8 6.5 2.173 ;
      RECT 6.225 1.84 6.5 2.17 ;
      RECT 6.24 1.812 6.505 2.155 ;
      RECT 6.24 1.824 6.51 2.135 ;
      RECT 6.225 1.84 6.515 2.118 ;
      RECT 6.225 1.85 6.52 1.973 ;
      RECT 6.22 1.85 6.52 1.93 ;
      RECT 6.22 1.865 6.525 1.908 ;
      RECT 6.315 1.775 6.455 2.255 ;
      RECT 6.315 1.773 6.425 2.255 ;
      RECT 6.401 1.77 6.425 2.255 ;
      RECT 6.06 3.437 6.065 3.483 ;
      RECT 6.05 3.285 6.06 3.507 ;
      RECT 6.045 3.13 6.05 3.532 ;
      RECT 6.03 3.092 6.045 3.543 ;
      RECT 6.025 3.075 6.03 3.55 ;
      RECT 6.015 3.063 6.025 3.557 ;
      RECT 6.01 3.054 6.015 3.559 ;
      RECT 6.005 3.052 6.01 3.563 ;
      RECT 5.96 3.043 6.005 3.578 ;
      RECT 5.955 3.035 5.96 3.592 ;
      RECT 5.95 3.032 5.955 3.596 ;
      RECT 5.935 3.027 5.95 3.604 ;
      RECT 5.88 3.017 5.935 3.615 ;
      RECT 5.845 3.005 5.88 3.616 ;
      RECT 5.836 3 5.845 3.61 ;
      RECT 5.75 3 5.836 3.6 ;
      RECT 5.72 3 5.75 3.578 ;
      RECT 5.71 3 5.715 3.558 ;
      RECT 5.705 3 5.71 3.52 ;
      RECT 5.7 3 5.705 3.478 ;
      RECT 5.695 3 5.7 3.438 ;
      RECT 5.69 3 5.695 3.368 ;
      RECT 5.68 3 5.69 3.29 ;
      RECT 5.675 3 5.68 3.19 ;
      RECT 5.715 3 5.72 3.56 ;
      RECT 5.21 3.082 5.3 3.56 ;
      RECT 5.195 3.085 5.315 3.558 ;
      RECT 5.21 3.084 5.315 3.558 ;
      RECT 5.175 3.091 5.34 3.548 ;
      RECT 5.195 3.085 5.34 3.548 ;
      RECT 5.16 3.097 5.34 3.536 ;
      RECT 5.195 3.088 5.39 3.529 ;
      RECT 5.146 3.105 5.39 3.527 ;
      RECT 5.175 3.095 5.4 3.515 ;
      RECT 5.146 3.116 5.43 3.506 ;
      RECT 5.06 3.14 5.43 3.5 ;
      RECT 5.06 3.153 5.47 3.483 ;
      RECT 5.055 3.175 5.47 3.476 ;
      RECT 5.025 3.19 5.47 3.466 ;
      RECT 5.02 3.201 5.47 3.456 ;
      RECT 4.99 3.214 5.47 3.447 ;
      RECT 4.975 3.232 5.47 3.436 ;
      RECT 4.95 3.245 5.47 3.426 ;
      RECT 5.21 3.081 5.22 3.56 ;
      RECT 5.256 2.505 5.295 2.75 ;
      RECT 5.17 2.505 5.305 2.748 ;
      RECT 5.055 2.53 5.305 2.745 ;
      RECT 5.055 2.53 5.31 2.743 ;
      RECT 5.055 2.53 5.325 2.738 ;
      RECT 5.161 2.505 5.34 2.718 ;
      RECT 5.075 2.513 5.34 2.718 ;
      RECT 4.745 1.865 4.915 2.3 ;
      RECT 4.735 1.899 4.915 2.283 ;
      RECT 4.815 1.835 4.985 2.27 ;
      RECT 4.72 1.91 4.985 2.248 ;
      RECT 4.815 1.845 4.99 2.238 ;
      RECT 4.745 1.897 5.02 2.223 ;
      RECT 4.705 1.923 5.02 2.208 ;
      RECT 4.705 1.965 5.03 2.188 ;
      RECT 4.7 1.99 5.035 2.17 ;
      RECT 4.7 2 5.04 2.155 ;
      RECT 4.695 1.937 5.02 2.153 ;
      RECT 4.695 2.01 5.045 2.138 ;
      RECT 4.69 1.947 5.02 2.135 ;
      RECT 4.685 2.031 5.05 2.118 ;
      RECT 4.685 2.063 5.055 2.098 ;
      RECT 4.68 1.977 5.03 2.09 ;
      RECT 4.685 1.962 5.02 2.118 ;
      RECT 4.7 1.932 5.02 2.17 ;
      RECT 4.545 2.519 4.77 2.775 ;
      RECT 4.545 2.552 4.79 2.765 ;
      RECT 4.51 2.552 4.79 2.763 ;
      RECT 4.51 2.565 4.795 2.753 ;
      RECT 4.51 2.585 4.805 2.745 ;
      RECT 4.51 2.682 4.81 2.738 ;
      RECT 4.49 2.43 4.62 2.728 ;
      RECT 4.445 2.585 4.805 2.67 ;
      RECT 4.435 2.43 4.62 2.615 ;
      RECT 4.435 2.462 4.706 2.615 ;
      RECT 4.4 2.992 4.42 3.17 ;
      RECT 4.365 2.945 4.4 3.17 ;
      RECT 4.35 2.885 4.365 3.17 ;
      RECT 4.325 2.832 4.35 3.17 ;
      RECT 4.31 2.785 4.325 3.17 ;
      RECT 4.29 2.762 4.31 3.17 ;
      RECT 4.265 2.727 4.29 3.17 ;
      RECT 4.255 2.573 4.265 3.17 ;
      RECT 4.225 2.568 4.255 3.161 ;
      RECT 4.22 2.565 4.225 3.151 ;
      RECT 4.205 2.565 4.22 3.125 ;
      RECT 4.2 2.565 4.205 3.088 ;
      RECT 4.175 2.565 4.2 3.04 ;
      RECT 4.155 2.565 4.175 2.965 ;
      RECT 4.145 2.565 4.155 2.925 ;
      RECT 4.14 2.565 4.145 2.9 ;
      RECT 4.135 2.565 4.14 2.883 ;
      RECT 4.13 2.565 4.135 2.865 ;
      RECT 4.125 2.566 4.13 2.855 ;
      RECT 4.115 2.568 4.125 2.823 ;
      RECT 4.105 2.57 4.115 2.79 ;
      RECT 4.095 2.573 4.105 2.763 ;
      RECT 4.42 3 4.645 3.17 ;
      RECT 3.75 1.812 3.92 2.265 ;
      RECT 3.75 1.812 4.01 2.231 ;
      RECT 3.75 1.812 4.04 2.215 ;
      RECT 3.75 1.812 4.07 2.188 ;
      RECT 4.006 1.79 4.085 2.17 ;
      RECT 3.785 1.797 4.09 2.155 ;
      RECT 3.785 1.805 4.1 2.118 ;
      RECT 3.745 1.832 4.1 2.09 ;
      RECT 3.73 1.845 4.1 2.055 ;
      RECT 3.75 1.82 4.12 2.045 ;
      RECT 3.725 1.885 4.12 2.015 ;
      RECT 3.725 1.915 4.125 1.998 ;
      RECT 3.72 1.945 4.125 1.985 ;
      RECT 3.785 1.794 4.085 2.17 ;
      RECT 3.92 1.791 4.006 2.249 ;
      RECT 3.871 1.792 4.085 2.17 ;
      RECT 4.015 3.452 4.06 3.645 ;
      RECT 4.005 3.422 4.015 3.645 ;
      RECT 4 3.407 4.005 3.645 ;
      RECT 3.96 3.317 4 3.645 ;
      RECT 3.955 3.23 3.96 3.645 ;
      RECT 3.945 3.2 3.955 3.645 ;
      RECT 3.94 3.16 3.945 3.645 ;
      RECT 3.93 3.122 3.94 3.645 ;
      RECT 3.925 3.087 3.93 3.645 ;
      RECT 3.905 3.04 3.925 3.645 ;
      RECT 3.89 2.965 3.905 3.645 ;
      RECT 3.885 2.92 3.89 3.64 ;
      RECT 3.88 2.9 3.885 3.613 ;
      RECT 3.875 2.88 3.88 3.598 ;
      RECT 3.87 2.855 3.875 3.578 ;
      RECT 3.865 2.833 3.87 3.563 ;
      RECT 3.86 2.811 3.865 3.545 ;
      RECT 3.855 2.79 3.86 3.535 ;
      RECT 3.845 2.762 3.855 3.505 ;
      RECT 3.835 2.725 3.845 3.473 ;
      RECT 3.825 2.685 3.835 3.44 ;
      RECT 3.815 2.663 3.825 3.41 ;
      RECT 3.785 2.615 3.815 3.342 ;
      RECT 3.77 2.575 3.785 3.269 ;
      RECT 3.76 2.575 3.77 3.235 ;
      RECT 3.755 2.575 3.76 3.21 ;
      RECT 3.75 2.575 3.755 3.195 ;
      RECT 3.745 2.575 3.75 3.173 ;
      RECT 3.74 2.575 3.745 3.16 ;
      RECT 3.725 2.575 3.74 3.125 ;
      RECT 3.705 2.575 3.725 3.065 ;
      RECT 3.695 2.575 3.705 3.015 ;
      RECT 3.675 2.575 3.695 2.963 ;
      RECT 3.655 2.575 3.675 2.92 ;
      RECT 3.645 2.575 3.655 2.908 ;
      RECT 3.615 2.575 3.645 2.895 ;
      RECT 3.585 2.596 3.615 2.875 ;
      RECT 3.575 2.624 3.585 2.855 ;
      RECT 3.56 2.641 3.575 2.823 ;
      RECT 3.555 2.655 3.56 2.79 ;
      RECT 3.55 2.663 3.555 2.763 ;
      RECT 3.545 2.671 3.55 2.725 ;
      RECT 3.55 3.195 3.555 3.53 ;
      RECT 3.515 3.182 3.55 3.529 ;
      RECT 3.445 3.122 3.515 3.528 ;
      RECT 3.365 3.065 3.445 3.527 ;
      RECT 3.23 3.025 3.365 3.526 ;
      RECT 3.23 3.212 3.565 3.515 ;
      RECT 3.19 3.212 3.565 3.505 ;
      RECT 3.19 3.23 3.57 3.5 ;
      RECT 3.19 3.32 3.575 3.49 ;
      RECT 3.185 3.015 3.35 3.47 ;
      RECT 3.18 3.015 3.35 3.213 ;
      RECT 3.18 3.172 3.545 3.213 ;
      RECT 3.18 3.16 3.54 3.213 ;
      RECT 1.17 7.855 1.34 8.305 ;
      RECT 1.225 6.075 1.395 8.025 ;
      RECT 1.17 5.015 1.34 6.245 ;
      RECT 0.65 5.015 0.82 8.305 ;
      RECT 0.65 7.315 1.055 7.645 ;
      RECT 0.65 6.475 1.055 6.805 ;
      RECT 81.22 7.8 81.39 8.31 ;
      RECT 80.23 0.57 80.4 1.08 ;
      RECT 80.23 2.39 80.4 3.86 ;
      RECT 80.23 5.02 80.4 6.49 ;
      RECT 80.23 7.8 80.4 8.31 ;
      RECT 78.87 0.575 79.04 3.865 ;
      RECT 78.87 5.015 79.04 8.305 ;
      RECT 78.44 0.575 78.61 1.085 ;
      RECT 78.44 1.655 78.61 3.865 ;
      RECT 78.44 5.015 78.61 7.225 ;
      RECT 78.44 7.795 78.61 8.305 ;
      RECT 76.05 2.85 76.42 3.22 ;
      RECT 74.09 5.015 74.26 8.305 ;
      RECT 73.66 5.015 73.83 7.225 ;
      RECT 73.66 7.795 73.83 8.305 ;
      RECT 65.435 7.8 65.605 8.31 ;
      RECT 64.445 0.57 64.615 1.08 ;
      RECT 64.445 2.39 64.615 3.86 ;
      RECT 64.445 5.02 64.615 6.49 ;
      RECT 64.445 7.8 64.615 8.31 ;
      RECT 63.085 0.575 63.255 3.865 ;
      RECT 63.085 5.015 63.255 8.305 ;
      RECT 62.655 0.575 62.825 1.085 ;
      RECT 62.655 1.655 62.825 3.865 ;
      RECT 62.655 5.015 62.825 7.225 ;
      RECT 62.655 7.795 62.825 8.305 ;
      RECT 60.265 2.85 60.635 3.22 ;
      RECT 58.305 5.015 58.475 8.305 ;
      RECT 57.875 5.015 58.045 7.225 ;
      RECT 57.875 7.795 58.045 8.305 ;
      RECT 49.65 7.8 49.82 8.31 ;
      RECT 48.66 0.57 48.83 1.08 ;
      RECT 48.66 2.39 48.83 3.86 ;
      RECT 48.66 5.02 48.83 6.49 ;
      RECT 48.66 7.8 48.83 8.31 ;
      RECT 47.3 0.575 47.47 3.865 ;
      RECT 47.3 5.015 47.47 8.305 ;
      RECT 46.87 0.575 47.04 1.085 ;
      RECT 46.87 1.655 47.04 3.865 ;
      RECT 46.87 5.015 47.04 7.225 ;
      RECT 46.87 7.795 47.04 8.305 ;
      RECT 44.48 2.85 44.85 3.22 ;
      RECT 42.52 5.015 42.69 8.305 ;
      RECT 42.09 5.015 42.26 7.225 ;
      RECT 42.09 7.795 42.26 8.305 ;
      RECT 33.875 7.8 34.045 8.31 ;
      RECT 32.885 0.57 33.055 1.08 ;
      RECT 32.885 2.39 33.055 3.86 ;
      RECT 32.885 5.02 33.055 6.49 ;
      RECT 32.885 7.8 33.055 8.31 ;
      RECT 31.525 0.575 31.695 3.865 ;
      RECT 31.525 5.015 31.695 8.305 ;
      RECT 31.095 0.575 31.265 1.085 ;
      RECT 31.095 1.655 31.265 3.865 ;
      RECT 31.095 5.015 31.265 7.225 ;
      RECT 31.095 7.795 31.265 8.305 ;
      RECT 28.705 2.85 29.075 3.22 ;
      RECT 26.745 5.015 26.915 8.305 ;
      RECT 26.315 5.015 26.485 7.225 ;
      RECT 26.315 7.795 26.485 8.305 ;
      RECT 18.095 7.8 18.265 8.31 ;
      RECT 17.105 0.57 17.275 1.08 ;
      RECT 17.105 2.39 17.275 3.86 ;
      RECT 17.105 5.02 17.275 6.49 ;
      RECT 17.105 7.8 17.275 8.31 ;
      RECT 15.745 0.575 15.915 3.865 ;
      RECT 15.745 5.015 15.915 8.305 ;
      RECT 15.315 0.575 15.485 1.085 ;
      RECT 15.315 1.655 15.485 3.865 ;
      RECT 15.315 5.015 15.485 7.225 ;
      RECT 15.315 7.795 15.485 8.305 ;
      RECT 12.925 2.85 13.295 3.22 ;
      RECT 10.965 5.015 11.135 8.305 ;
      RECT 10.535 5.015 10.705 7.225 ;
      RECT 10.535 7.795 10.705 8.305 ;
      RECT 1.6 5.015 1.77 7.225 ;
      RECT 1.6 7.795 1.77 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r1
  CLASS BLOCK ;
  ORIGIN -1.46 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8_b0r1 ;
  SIZE 92.435 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 21.655 0.915 21.825 1.085 ;
        RECT 21.65 0.91 21.82 1.08 ;
        RECT 21.65 2.39 21.82 2.56 ;
      LAYER li1 ;
        RECT 21.655 0.915 21.825 1.085 ;
        RECT 21.65 0.57 21.82 1.08 ;
        RECT 21.65 2.39 21.82 3.86 ;
      LAYER met1 ;
        RECT 21.59 2.36 21.88 2.59 ;
        RECT 21.59 0.88 21.88 1.11 ;
        RECT 21.65 0.88 21.82 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 39.58 0.915 39.75 1.085 ;
        RECT 39.575 0.91 39.745 1.08 ;
        RECT 39.575 2.39 39.745 2.56 ;
      LAYER li1 ;
        RECT 39.58 0.915 39.75 1.085 ;
        RECT 39.575 0.57 39.745 1.08 ;
        RECT 39.575 2.39 39.745 3.86 ;
      LAYER met1 ;
        RECT 39.515 2.36 39.805 2.59 ;
        RECT 39.515 0.88 39.805 1.11 ;
        RECT 39.575 0.88 39.745 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 57.505 0.915 57.675 1.085 ;
        RECT 57.5 0.91 57.67 1.08 ;
        RECT 57.5 2.39 57.67 2.56 ;
      LAYER li1 ;
        RECT 57.505 0.915 57.675 1.085 ;
        RECT 57.5 0.57 57.67 1.08 ;
        RECT 57.5 2.39 57.67 3.86 ;
      LAYER met1 ;
        RECT 57.44 2.36 57.73 2.59 ;
        RECT 57.44 0.88 57.73 1.11 ;
        RECT 57.5 0.88 57.67 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 75.43 0.915 75.6 1.085 ;
        RECT 75.425 0.91 75.595 1.08 ;
        RECT 75.425 2.39 75.595 2.56 ;
      LAYER li1 ;
        RECT 75.43 0.915 75.6 1.085 ;
        RECT 75.425 0.57 75.595 1.08 ;
        RECT 75.425 2.39 75.595 3.86 ;
      LAYER met1 ;
        RECT 75.365 2.36 75.655 2.59 ;
        RECT 75.365 0.88 75.655 1.11 ;
        RECT 75.425 0.88 75.595 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 93.355 0.915 93.525 1.085 ;
        RECT 93.35 0.91 93.52 1.08 ;
        RECT 93.35 2.39 93.52 2.56 ;
      LAYER li1 ;
        RECT 93.355 0.915 93.525 1.085 ;
        RECT 93.35 0.57 93.52 1.08 ;
        RECT 93.35 2.39 93.52 3.86 ;
      LAYER met1 ;
        RECT 93.29 2.36 93.58 2.59 ;
        RECT 93.29 0.88 93.58 1.11 ;
        RECT 93.35 0.88 93.52 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 17.5 1.66 17.67 2.935 ;
        RECT 17.5 5.945 17.67 7.22 ;
        RECT 12.74 5.945 12.91 7.22 ;
      LAYER met2 ;
        RECT 17.42 2.705 17.77 3.055 ;
        RECT 17.41 5.84 17.76 6.19 ;
        RECT 17.485 2.705 17.66 6.19 ;
      LAYER met1 ;
        RECT 17.42 2.765 17.9 2.935 ;
        RECT 17.42 2.705 17.77 3.055 ;
        RECT 12.68 5.945 17.9 6.115 ;
        RECT 17.41 5.84 17.76 6.19 ;
        RECT 12.68 5.915 12.97 6.145 ;
      LAYER mcon ;
        RECT 12.74 5.945 12.91 6.115 ;
        RECT 17.5 5.945 17.67 6.115 ;
        RECT 17.5 2.765 17.67 2.935 ;
      LAYER via1 ;
        RECT 17.51 5.94 17.66 6.09 ;
        RECT 17.52 2.805 17.67 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 35.425 1.66 35.595 2.935 ;
        RECT 35.425 5.945 35.595 7.22 ;
        RECT 30.665 5.945 30.835 7.22 ;
      LAYER met2 ;
        RECT 35.345 2.705 35.695 3.055 ;
        RECT 35.335 5.84 35.685 6.19 ;
        RECT 35.41 2.705 35.585 6.19 ;
      LAYER met1 ;
        RECT 35.345 2.765 35.825 2.935 ;
        RECT 35.345 2.705 35.695 3.055 ;
        RECT 30.605 5.945 35.825 6.115 ;
        RECT 35.335 5.84 35.685 6.19 ;
        RECT 30.605 5.915 30.895 6.145 ;
      LAYER mcon ;
        RECT 30.665 5.945 30.835 6.115 ;
        RECT 35.425 5.945 35.595 6.115 ;
        RECT 35.425 2.765 35.595 2.935 ;
      LAYER via1 ;
        RECT 35.435 5.94 35.585 6.09 ;
        RECT 35.445 2.805 35.595 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 53.35 1.66 53.52 2.935 ;
        RECT 53.35 5.945 53.52 7.22 ;
        RECT 48.59 5.945 48.76 7.22 ;
      LAYER met2 ;
        RECT 53.27 2.705 53.62 3.055 ;
        RECT 53.26 5.84 53.61 6.19 ;
        RECT 53.335 2.705 53.51 6.19 ;
      LAYER met1 ;
        RECT 53.27 2.765 53.75 2.935 ;
        RECT 53.27 2.705 53.62 3.055 ;
        RECT 48.53 5.945 53.75 6.115 ;
        RECT 53.26 5.84 53.61 6.19 ;
        RECT 48.53 5.915 48.82 6.145 ;
      LAYER mcon ;
        RECT 48.59 5.945 48.76 6.115 ;
        RECT 53.35 5.945 53.52 6.115 ;
        RECT 53.35 2.765 53.52 2.935 ;
      LAYER via1 ;
        RECT 53.36 5.94 53.51 6.09 ;
        RECT 53.37 2.805 53.52 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 71.275 1.66 71.445 2.935 ;
        RECT 71.275 5.945 71.445 7.22 ;
        RECT 66.515 5.945 66.685 7.22 ;
      LAYER met2 ;
        RECT 71.195 2.705 71.545 3.055 ;
        RECT 71.185 5.84 71.535 6.19 ;
        RECT 71.26 2.705 71.435 6.19 ;
      LAYER met1 ;
        RECT 71.195 2.765 71.675 2.935 ;
        RECT 71.195 2.705 71.545 3.055 ;
        RECT 66.455 5.945 71.675 6.115 ;
        RECT 71.185 5.84 71.535 6.19 ;
        RECT 66.455 5.915 66.745 6.145 ;
      LAYER mcon ;
        RECT 66.515 5.945 66.685 6.115 ;
        RECT 71.275 5.945 71.445 6.115 ;
        RECT 71.275 2.765 71.445 2.935 ;
      LAYER via1 ;
        RECT 71.285 5.94 71.435 6.09 ;
        RECT 71.295 2.805 71.445 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 89.2 1.66 89.37 2.935 ;
        RECT 89.2 5.945 89.37 7.22 ;
        RECT 84.44 5.945 84.61 7.22 ;
      LAYER met2 ;
        RECT 89.12 2.705 89.47 3.055 ;
        RECT 89.11 5.84 89.46 6.19 ;
        RECT 89.185 2.705 89.36 6.19 ;
      LAYER met1 ;
        RECT 89.12 2.765 89.6 2.935 ;
        RECT 89.12 2.705 89.47 3.055 ;
        RECT 84.38 5.945 89.6 6.115 ;
        RECT 89.11 5.84 89.46 6.19 ;
        RECT 84.38 5.915 84.67 6.145 ;
      LAYER mcon ;
        RECT 84.44 5.945 84.61 6.115 ;
        RECT 89.2 5.945 89.37 6.115 ;
        RECT 89.2 2.765 89.37 2.935 ;
      LAYER via1 ;
        RECT 89.21 5.94 89.36 6.09 ;
        RECT 89.22 2.805 89.37 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 1.71 5.945 1.88 7.22 ;
      LAYER met1 ;
        RECT 1.65 5.945 2.11 6.115 ;
        RECT 1.65 5.915 1.94 6.145 ;
      LAYER mcon ;
        RECT 1.71 5.945 1.88 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 2.74 4.33 3.545 4.71 ;
      LAYER li1 ;
        RECT 1.48 4.44 93.895 4.745 ;
        RECT 87.935 4.135 93.895 4.745 ;
        RECT 91.76 4.13 93.74 4.75 ;
        RECT 92.92 3.4 93.09 5.48 ;
        RECT 91.93 3.4 92.1 5.48 ;
        RECT 89.19 3.405 89.36 5.475 ;
        RECT 3.205 4.285 93.895 4.745 ;
        RECT 86.435 3.785 86.605 4.745 ;
        RECT 84.43 4.285 84.6 5.475 ;
        RECT 83.995 3.785 84.165 4.745 ;
        RECT 82.035 3.785 82.205 4.745 ;
        RECT 81.075 3.785 81.245 4.745 ;
        RECT 79.115 3.785 79.285 4.745 ;
        RECT 78.115 3.785 78.285 4.745 ;
        RECT 77.155 3.785 77.325 4.745 ;
        RECT 70.01 4.135 75.97 4.745 ;
        RECT 73.835 4.13 75.815 4.75 ;
        RECT 74.995 3.4 75.165 5.48 ;
        RECT 74.005 3.4 74.175 5.48 ;
        RECT 71.265 3.405 71.435 5.475 ;
        RECT 68.51 3.785 68.68 4.745 ;
        RECT 66.505 4.285 66.675 5.475 ;
        RECT 66.07 3.785 66.24 4.745 ;
        RECT 64.11 3.785 64.28 4.745 ;
        RECT 63.15 3.785 63.32 4.745 ;
        RECT 61.19 3.785 61.36 4.745 ;
        RECT 60.19 3.785 60.36 4.745 ;
        RECT 59.23 3.785 59.4 4.745 ;
        RECT 52.085 4.135 58.045 4.745 ;
        RECT 55.91 4.13 57.89 4.75 ;
        RECT 57.07 3.4 57.24 5.48 ;
        RECT 56.08 3.4 56.25 5.48 ;
        RECT 53.34 3.405 53.51 5.475 ;
        RECT 50.585 3.785 50.755 4.745 ;
        RECT 48.58 4.285 48.75 5.475 ;
        RECT 48.145 3.785 48.315 4.745 ;
        RECT 46.185 3.785 46.355 4.745 ;
        RECT 45.225 3.785 45.395 4.745 ;
        RECT 43.265 3.785 43.435 4.745 ;
        RECT 42.265 3.785 42.435 4.745 ;
        RECT 41.305 3.785 41.475 4.745 ;
        RECT 34.16 4.135 40.12 4.745 ;
        RECT 37.985 4.13 39.965 4.75 ;
        RECT 39.145 3.4 39.315 5.48 ;
        RECT 38.155 3.4 38.325 5.48 ;
        RECT 35.415 3.405 35.585 5.475 ;
        RECT 32.66 3.785 32.83 4.745 ;
        RECT 30.655 4.285 30.825 5.475 ;
        RECT 30.22 3.785 30.39 4.745 ;
        RECT 28.26 3.785 28.43 4.745 ;
        RECT 27.3 3.785 27.47 4.745 ;
        RECT 25.34 3.785 25.51 4.745 ;
        RECT 24.34 3.785 24.51 4.745 ;
        RECT 23.38 3.785 23.55 4.745 ;
        RECT 16.235 4.135 22.195 4.745 ;
        RECT 20.06 4.13 22.04 4.75 ;
        RECT 21.22 3.4 21.39 5.48 ;
        RECT 20.23 3.4 20.4 5.48 ;
        RECT 17.49 3.405 17.66 5.475 ;
        RECT 14.735 3.785 14.905 4.745 ;
        RECT 12.73 4.285 12.9 5.475 ;
        RECT 12.295 3.785 12.465 4.745 ;
        RECT 10.335 3.785 10.505 4.745 ;
        RECT 9.375 3.785 9.545 4.745 ;
        RECT 7.415 3.785 7.585 4.745 ;
        RECT 6.415 3.785 6.585 4.745 ;
        RECT 5.455 3.785 5.625 4.745 ;
        RECT 3.51 4.285 3.68 8.305 ;
        RECT 1.48 4.285 93.895 4.405 ;
        RECT 1.48 4.285 3.035 4.745 ;
        RECT 1.7 4.285 1.87 5.475 ;
      LAYER met2 ;
        RECT 2.93 4.33 3.31 4.71 ;
      LAYER met1 ;
        RECT 1.48 4.285 93.895 4.745 ;
        RECT 76.345 4.135 93.895 4.745 ;
        RECT 91.76 4.13 93.74 4.75 ;
        RECT 76.345 4.125 88.305 4.745 ;
        RECT 58.42 4.135 75.97 4.745 ;
        RECT 73.835 4.13 75.815 4.75 ;
        RECT 58.42 4.125 70.38 4.745 ;
        RECT 40.495 4.135 58.045 4.745 ;
        RECT 55.91 4.13 57.89 4.75 ;
        RECT 40.495 4.125 52.455 4.745 ;
        RECT 22.57 4.135 40.12 4.745 ;
        RECT 37.985 4.13 39.965 4.75 ;
        RECT 22.57 4.125 34.53 4.745 ;
        RECT 4.645 4.135 22.195 4.745 ;
        RECT 20.06 4.13 22.04 4.75 ;
        RECT 4.645 4.125 16.605 4.745 ;
        RECT 3.45 6.655 3.74 6.885 ;
        RECT 3.28 6.685 3.74 6.855 ;
      LAYER via2 ;
        RECT 3.02 4.42 3.22 4.62 ;
      LAYER mcon ;
        RECT 3.51 6.685 3.68 6.855 ;
        RECT 3.82 4.545 3.99 4.715 ;
        RECT 4.785 4.285 4.955 4.455 ;
        RECT 5.245 4.285 5.415 4.455 ;
        RECT 5.705 4.285 5.875 4.455 ;
        RECT 6.165 4.285 6.335 4.455 ;
        RECT 6.625 4.285 6.795 4.455 ;
        RECT 7.085 4.285 7.255 4.455 ;
        RECT 7.545 4.285 7.715 4.455 ;
        RECT 8.005 4.285 8.175 4.455 ;
        RECT 8.465 4.285 8.635 4.455 ;
        RECT 8.925 4.285 9.095 4.455 ;
        RECT 9.385 4.285 9.555 4.455 ;
        RECT 9.845 4.285 10.015 4.455 ;
        RECT 10.305 4.285 10.475 4.455 ;
        RECT 10.765 4.285 10.935 4.455 ;
        RECT 11.225 4.285 11.395 4.455 ;
        RECT 11.685 4.285 11.855 4.455 ;
        RECT 12.145 4.285 12.315 4.455 ;
        RECT 12.605 4.285 12.775 4.455 ;
        RECT 13.065 4.285 13.235 4.455 ;
        RECT 13.525 4.285 13.695 4.455 ;
        RECT 13.985 4.285 14.155 4.455 ;
        RECT 14.445 4.285 14.615 4.455 ;
        RECT 14.85 4.545 15.02 4.715 ;
        RECT 14.905 4.285 15.075 4.455 ;
        RECT 15.365 4.285 15.535 4.455 ;
        RECT 15.825 4.285 15.995 4.455 ;
        RECT 16.285 4.285 16.455 4.455 ;
        RECT 19.61 4.545 19.78 4.715 ;
        RECT 19.61 4.165 19.78 4.335 ;
        RECT 20.31 4.55 20.48 4.72 ;
        RECT 20.31 4.16 20.48 4.33 ;
        RECT 21.3 4.55 21.47 4.72 ;
        RECT 21.3 4.16 21.47 4.33 ;
        RECT 22.71 4.285 22.88 4.455 ;
        RECT 23.17 4.285 23.34 4.455 ;
        RECT 23.63 4.285 23.8 4.455 ;
        RECT 24.09 4.285 24.26 4.455 ;
        RECT 24.55 4.285 24.72 4.455 ;
        RECT 25.01 4.285 25.18 4.455 ;
        RECT 25.47 4.285 25.64 4.455 ;
        RECT 25.93 4.285 26.1 4.455 ;
        RECT 26.39 4.285 26.56 4.455 ;
        RECT 26.85 4.285 27.02 4.455 ;
        RECT 27.31 4.285 27.48 4.455 ;
        RECT 27.77 4.285 27.94 4.455 ;
        RECT 28.23 4.285 28.4 4.455 ;
        RECT 28.69 4.285 28.86 4.455 ;
        RECT 29.15 4.285 29.32 4.455 ;
        RECT 29.61 4.285 29.78 4.455 ;
        RECT 30.07 4.285 30.24 4.455 ;
        RECT 30.53 4.285 30.7 4.455 ;
        RECT 30.99 4.285 31.16 4.455 ;
        RECT 31.45 4.285 31.62 4.455 ;
        RECT 31.91 4.285 32.08 4.455 ;
        RECT 32.37 4.285 32.54 4.455 ;
        RECT 32.775 4.545 32.945 4.715 ;
        RECT 32.83 4.285 33 4.455 ;
        RECT 33.29 4.285 33.46 4.455 ;
        RECT 33.75 4.285 33.92 4.455 ;
        RECT 34.21 4.285 34.38 4.455 ;
        RECT 37.535 4.545 37.705 4.715 ;
        RECT 37.535 4.165 37.705 4.335 ;
        RECT 38.235 4.55 38.405 4.72 ;
        RECT 38.235 4.16 38.405 4.33 ;
        RECT 39.225 4.55 39.395 4.72 ;
        RECT 39.225 4.16 39.395 4.33 ;
        RECT 40.635 4.285 40.805 4.455 ;
        RECT 41.095 4.285 41.265 4.455 ;
        RECT 41.555 4.285 41.725 4.455 ;
        RECT 42.015 4.285 42.185 4.455 ;
        RECT 42.475 4.285 42.645 4.455 ;
        RECT 42.935 4.285 43.105 4.455 ;
        RECT 43.395 4.285 43.565 4.455 ;
        RECT 43.855 4.285 44.025 4.455 ;
        RECT 44.315 4.285 44.485 4.455 ;
        RECT 44.775 4.285 44.945 4.455 ;
        RECT 45.235 4.285 45.405 4.455 ;
        RECT 45.695 4.285 45.865 4.455 ;
        RECT 46.155 4.285 46.325 4.455 ;
        RECT 46.615 4.285 46.785 4.455 ;
        RECT 47.075 4.285 47.245 4.455 ;
        RECT 47.535 4.285 47.705 4.455 ;
        RECT 47.995 4.285 48.165 4.455 ;
        RECT 48.455 4.285 48.625 4.455 ;
        RECT 48.915 4.285 49.085 4.455 ;
        RECT 49.375 4.285 49.545 4.455 ;
        RECT 49.835 4.285 50.005 4.455 ;
        RECT 50.295 4.285 50.465 4.455 ;
        RECT 50.7 4.545 50.87 4.715 ;
        RECT 50.755 4.285 50.925 4.455 ;
        RECT 51.215 4.285 51.385 4.455 ;
        RECT 51.675 4.285 51.845 4.455 ;
        RECT 52.135 4.285 52.305 4.455 ;
        RECT 55.46 4.545 55.63 4.715 ;
        RECT 55.46 4.165 55.63 4.335 ;
        RECT 56.16 4.55 56.33 4.72 ;
        RECT 56.16 4.16 56.33 4.33 ;
        RECT 57.15 4.55 57.32 4.72 ;
        RECT 57.15 4.16 57.32 4.33 ;
        RECT 58.56 4.285 58.73 4.455 ;
        RECT 59.02 4.285 59.19 4.455 ;
        RECT 59.48 4.285 59.65 4.455 ;
        RECT 59.94 4.285 60.11 4.455 ;
        RECT 60.4 4.285 60.57 4.455 ;
        RECT 60.86 4.285 61.03 4.455 ;
        RECT 61.32 4.285 61.49 4.455 ;
        RECT 61.78 4.285 61.95 4.455 ;
        RECT 62.24 4.285 62.41 4.455 ;
        RECT 62.7 4.285 62.87 4.455 ;
        RECT 63.16 4.285 63.33 4.455 ;
        RECT 63.62 4.285 63.79 4.455 ;
        RECT 64.08 4.285 64.25 4.455 ;
        RECT 64.54 4.285 64.71 4.455 ;
        RECT 65 4.285 65.17 4.455 ;
        RECT 65.46 4.285 65.63 4.455 ;
        RECT 65.92 4.285 66.09 4.455 ;
        RECT 66.38 4.285 66.55 4.455 ;
        RECT 66.84 4.285 67.01 4.455 ;
        RECT 67.3 4.285 67.47 4.455 ;
        RECT 67.76 4.285 67.93 4.455 ;
        RECT 68.22 4.285 68.39 4.455 ;
        RECT 68.625 4.545 68.795 4.715 ;
        RECT 68.68 4.285 68.85 4.455 ;
        RECT 69.14 4.285 69.31 4.455 ;
        RECT 69.6 4.285 69.77 4.455 ;
        RECT 70.06 4.285 70.23 4.455 ;
        RECT 73.385 4.545 73.555 4.715 ;
        RECT 73.385 4.165 73.555 4.335 ;
        RECT 74.085 4.55 74.255 4.72 ;
        RECT 74.085 4.16 74.255 4.33 ;
        RECT 75.075 4.55 75.245 4.72 ;
        RECT 75.075 4.16 75.245 4.33 ;
        RECT 76.485 4.285 76.655 4.455 ;
        RECT 76.945 4.285 77.115 4.455 ;
        RECT 77.405 4.285 77.575 4.455 ;
        RECT 77.865 4.285 78.035 4.455 ;
        RECT 78.325 4.285 78.495 4.455 ;
        RECT 78.785 4.285 78.955 4.455 ;
        RECT 79.245 4.285 79.415 4.455 ;
        RECT 79.705 4.285 79.875 4.455 ;
        RECT 80.165 4.285 80.335 4.455 ;
        RECT 80.625 4.285 80.795 4.455 ;
        RECT 81.085 4.285 81.255 4.455 ;
        RECT 81.545 4.285 81.715 4.455 ;
        RECT 82.005 4.285 82.175 4.455 ;
        RECT 82.465 4.285 82.635 4.455 ;
        RECT 82.925 4.285 83.095 4.455 ;
        RECT 83.385 4.285 83.555 4.455 ;
        RECT 83.845 4.285 84.015 4.455 ;
        RECT 84.305 4.285 84.475 4.455 ;
        RECT 84.765 4.285 84.935 4.455 ;
        RECT 85.225 4.285 85.395 4.455 ;
        RECT 85.685 4.285 85.855 4.455 ;
        RECT 86.145 4.285 86.315 4.455 ;
        RECT 86.55 4.545 86.72 4.715 ;
        RECT 86.605 4.285 86.775 4.455 ;
        RECT 87.065 4.285 87.235 4.455 ;
        RECT 87.525 4.285 87.695 4.455 ;
        RECT 87.985 4.285 88.155 4.455 ;
        RECT 91.31 4.545 91.48 4.715 ;
        RECT 91.31 4.165 91.48 4.335 ;
        RECT 92.01 4.55 92.18 4.72 ;
        RECT 92.01 4.16 92.18 4.33 ;
        RECT 93 4.55 93.17 4.72 ;
        RECT 93 4.16 93.17 4.33 ;
      LAYER via1 ;
        RECT 3.045 4.445 3.195 4.595 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 85.7 7.055 86.075 7.425 ;
      RECT 85.735 4.925 86.045 7.425 ;
      RECT 85.735 4.925 88.83 5.235 ;
      RECT 88.52 1.125 88.83 5.235 ;
      RECT 88.52 1.14 88.895 1.51 ;
      RECT 85.645 3.685 86.205 4.015 ;
      RECT 85.645 2.015 85.945 4.015 ;
      RECT 81.715 3.125 82.265 3.455 ;
      RECT 81.965 2.015 82.265 3.455 ;
      RECT 82.765 1.885 82.915 2.535 ;
      RECT 81.965 2.015 85.945 2.315 ;
      RECT 80.485 0.96 80.785 3.91 ;
      RECT 80.475 2.565 81.205 2.895 ;
      RECT 80.44 0.96 80.815 1.33 ;
      RECT 79.035 3.125 79.765 3.455 ;
      RECT 79.05 0.96 79.35 3.455 ;
      RECT 76.925 2.565 77.655 2.895 ;
      RECT 77.08 0.93 77.38 2.895 ;
      RECT 79.005 0.96 79.38 1.33 ;
      RECT 77.035 0.93 77.41 1.3 ;
      RECT 77.035 0.97 79.38 1.27 ;
      RECT 67.775 7.055 68.15 7.425 ;
      RECT 67.81 4.925 68.12 7.425 ;
      RECT 67.81 4.925 70.905 5.235 ;
      RECT 70.595 1.125 70.905 5.235 ;
      RECT 70.595 1.14 70.97 1.51 ;
      RECT 67.72 3.685 68.28 4.015 ;
      RECT 67.72 2.015 68.02 4.015 ;
      RECT 63.79 3.125 64.34 3.455 ;
      RECT 64.04 2.015 64.34 3.455 ;
      RECT 64.84 1.885 64.99 2.535 ;
      RECT 64.04 2.015 68.02 2.315 ;
      RECT 62.56 0.96 62.86 3.91 ;
      RECT 62.55 2.565 63.28 2.895 ;
      RECT 62.515 0.96 62.89 1.33 ;
      RECT 61.11 3.125 61.84 3.455 ;
      RECT 61.125 0.96 61.425 3.455 ;
      RECT 59 2.565 59.73 2.895 ;
      RECT 59.155 0.93 59.455 2.895 ;
      RECT 61.08 0.96 61.455 1.33 ;
      RECT 59.11 0.93 59.485 1.3 ;
      RECT 59.11 0.97 61.455 1.27 ;
      RECT 49.85 7.055 50.225 7.425 ;
      RECT 49.885 4.925 50.195 7.425 ;
      RECT 49.885 4.925 52.98 5.235 ;
      RECT 52.67 1.125 52.98 5.235 ;
      RECT 52.67 1.14 53.045 1.51 ;
      RECT 49.795 3.685 50.355 4.015 ;
      RECT 49.795 2.015 50.095 4.015 ;
      RECT 45.865 3.125 46.415 3.455 ;
      RECT 46.115 2.015 46.415 3.455 ;
      RECT 46.915 1.885 47.065 2.535 ;
      RECT 46.115 2.015 50.095 2.315 ;
      RECT 44.635 0.96 44.935 3.91 ;
      RECT 44.625 2.565 45.355 2.895 ;
      RECT 44.59 0.96 44.965 1.33 ;
      RECT 43.185 3.125 43.915 3.455 ;
      RECT 43.2 0.96 43.5 3.455 ;
      RECT 41.075 2.565 41.805 2.895 ;
      RECT 41.23 0.93 41.53 2.895 ;
      RECT 43.155 0.96 43.53 1.33 ;
      RECT 41.185 0.93 41.56 1.3 ;
      RECT 41.185 0.97 43.53 1.27 ;
      RECT 31.925 7.055 32.3 7.425 ;
      RECT 31.96 4.925 32.27 7.425 ;
      RECT 31.96 4.925 35.055 5.235 ;
      RECT 34.745 1.125 35.055 5.235 ;
      RECT 34.745 1.14 35.12 1.51 ;
      RECT 31.87 3.685 32.43 4.015 ;
      RECT 31.87 2.015 32.17 4.015 ;
      RECT 27.94 3.125 28.49 3.455 ;
      RECT 28.19 2.015 28.49 3.455 ;
      RECT 28.99 1.885 29.14 2.535 ;
      RECT 28.19 2.015 32.17 2.315 ;
      RECT 26.71 0.96 27.01 3.91 ;
      RECT 26.7 2.565 27.43 2.895 ;
      RECT 26.665 0.96 27.04 1.33 ;
      RECT 25.26 3.125 25.99 3.455 ;
      RECT 25.275 0.96 25.575 3.455 ;
      RECT 23.15 2.565 23.88 2.895 ;
      RECT 23.305 0.93 23.605 2.895 ;
      RECT 25.23 0.96 25.605 1.33 ;
      RECT 23.26 0.93 23.635 1.3 ;
      RECT 23.26 0.97 25.605 1.27 ;
      RECT 14 7.055 14.375 7.425 ;
      RECT 14.035 4.925 14.345 7.425 ;
      RECT 14.035 4.925 17.13 5.235 ;
      RECT 16.82 1.125 17.13 5.235 ;
      RECT 16.82 1.14 17.195 1.51 ;
      RECT 13.945 3.685 14.505 4.015 ;
      RECT 13.945 2.015 14.245 4.015 ;
      RECT 10.015 3.125 10.565 3.455 ;
      RECT 10.265 2.015 10.565 3.455 ;
      RECT 11.065 1.885 11.215 2.535 ;
      RECT 10.265 2.015 14.245 2.315 ;
      RECT 8.785 0.96 9.085 3.91 ;
      RECT 8.775 2.565 9.505 2.895 ;
      RECT 8.74 0.96 9.115 1.33 ;
      RECT 7.335 3.125 8.065 3.455 ;
      RECT 7.35 0.96 7.65 3.455 ;
      RECT 5.225 2.565 5.955 2.895 ;
      RECT 5.38 0.93 5.68 2.895 ;
      RECT 7.305 0.96 7.68 1.33 ;
      RECT 5.335 0.93 5.71 1.3 ;
      RECT 5.335 0.97 7.68 1.27 ;
      RECT 86.835 2.005 87.565 2.335 ;
      RECT 84.615 3.685 85.345 4.015 ;
      RECT 82.915 3.685 83.645 4.015 ;
      RECT 77.955 2.565 78.685 2.895 ;
      RECT 76.595 3.685 77.325 4.015 ;
      RECT 68.91 2.005 69.64 2.335 ;
      RECT 66.69 3.685 67.42 4.015 ;
      RECT 64.99 3.685 65.72 4.015 ;
      RECT 60.03 2.565 60.76 2.895 ;
      RECT 58.67 3.685 59.4 4.015 ;
      RECT 50.985 2.005 51.715 2.335 ;
      RECT 48.765 3.685 49.495 4.015 ;
      RECT 47.065 3.685 47.795 4.015 ;
      RECT 42.105 2.565 42.835 2.895 ;
      RECT 40.745 3.685 41.475 4.015 ;
      RECT 33.06 2.005 33.79 2.335 ;
      RECT 30.84 3.685 31.57 4.015 ;
      RECT 29.14 3.685 29.87 4.015 ;
      RECT 24.18 2.565 24.91 2.895 ;
      RECT 22.82 3.685 23.55 4.015 ;
      RECT 15.135 2.005 15.865 2.335 ;
      RECT 12.915 3.685 13.645 4.015 ;
      RECT 11.215 3.685 11.945 4.015 ;
      RECT 6.255 2.565 6.985 2.895 ;
      RECT 4.895 3.685 5.625 4.015 ;
      RECT 1.46 8.5 2.265 8.88 ;
    LAYER via2 ;
      RECT 78.36 2.63 78.56 2.83 ;
      RECT 78.355 2.625 78.555 2.825 ;
      RECT 60.435 2.63 60.635 2.83 ;
      RECT 60.43 2.625 60.63 2.825 ;
      RECT 42.51 2.63 42.71 2.83 ;
      RECT 42.505 2.625 42.705 2.825 ;
      RECT 24.585 2.63 24.785 2.83 ;
      RECT 24.58 2.625 24.78 2.825 ;
      RECT 6.66 2.63 6.86 2.83 ;
      RECT 6.655 2.625 6.855 2.825 ;
      RECT 88.61 1.225 88.81 1.425 ;
      RECT 86.895 2.065 87.095 2.265 ;
      RECT 85.935 3.745 86.135 3.945 ;
      RECT 85.79 7.14 85.99 7.34 ;
      RECT 84.935 3.745 85.135 3.945 ;
      RECT 82.975 3.745 83.175 3.945 ;
      RECT 81.775 3.185 81.975 3.385 ;
      RECT 80.535 2.625 80.735 2.825 ;
      RECT 80.53 1.045 80.73 1.245 ;
      RECT 79.095 1.04 79.295 1.24 ;
      RECT 79.095 3.185 79.295 3.385 ;
      RECT 77.135 2.625 77.335 2.825 ;
      RECT 77.125 1.015 77.325 1.215 ;
      RECT 76.655 3.745 76.855 3.945 ;
      RECT 70.685 1.225 70.885 1.425 ;
      RECT 68.97 2.065 69.17 2.265 ;
      RECT 68.01 3.745 68.21 3.945 ;
      RECT 67.865 7.14 68.065 7.34 ;
      RECT 67.01 3.745 67.21 3.945 ;
      RECT 65.05 3.745 65.25 3.945 ;
      RECT 63.85 3.185 64.05 3.385 ;
      RECT 62.61 2.625 62.81 2.825 ;
      RECT 62.605 1.045 62.805 1.245 ;
      RECT 61.17 1.04 61.37 1.24 ;
      RECT 61.17 3.185 61.37 3.385 ;
      RECT 59.21 2.625 59.41 2.825 ;
      RECT 59.2 1.015 59.4 1.215 ;
      RECT 58.73 3.745 58.93 3.945 ;
      RECT 52.76 1.225 52.96 1.425 ;
      RECT 51.045 2.065 51.245 2.265 ;
      RECT 50.085 3.745 50.285 3.945 ;
      RECT 49.94 7.14 50.14 7.34 ;
      RECT 49.085 3.745 49.285 3.945 ;
      RECT 47.125 3.745 47.325 3.945 ;
      RECT 45.925 3.185 46.125 3.385 ;
      RECT 44.685 2.625 44.885 2.825 ;
      RECT 44.68 1.045 44.88 1.245 ;
      RECT 43.245 1.04 43.445 1.24 ;
      RECT 43.245 3.185 43.445 3.385 ;
      RECT 41.285 2.625 41.485 2.825 ;
      RECT 41.275 1.015 41.475 1.215 ;
      RECT 40.805 3.745 41.005 3.945 ;
      RECT 34.835 1.225 35.035 1.425 ;
      RECT 33.12 2.065 33.32 2.265 ;
      RECT 32.16 3.745 32.36 3.945 ;
      RECT 32.015 7.14 32.215 7.34 ;
      RECT 31.16 3.745 31.36 3.945 ;
      RECT 29.2 3.745 29.4 3.945 ;
      RECT 28 3.185 28.2 3.385 ;
      RECT 26.76 2.625 26.96 2.825 ;
      RECT 26.755 1.045 26.955 1.245 ;
      RECT 25.32 1.04 25.52 1.24 ;
      RECT 25.32 3.185 25.52 3.385 ;
      RECT 23.36 2.625 23.56 2.825 ;
      RECT 23.35 1.015 23.55 1.215 ;
      RECT 22.88 3.745 23.08 3.945 ;
      RECT 16.91 1.225 17.11 1.425 ;
      RECT 15.195 2.065 15.395 2.265 ;
      RECT 14.235 3.745 14.435 3.945 ;
      RECT 14.09 7.14 14.29 7.34 ;
      RECT 13.235 3.745 13.435 3.945 ;
      RECT 11.275 3.745 11.475 3.945 ;
      RECT 10.075 3.185 10.275 3.385 ;
      RECT 8.835 2.625 9.035 2.825 ;
      RECT 8.83 1.045 9.03 1.245 ;
      RECT 7.395 1.04 7.595 1.24 ;
      RECT 7.395 3.185 7.595 3.385 ;
      RECT 5.435 2.625 5.635 2.825 ;
      RECT 5.425 1.015 5.625 1.215 ;
      RECT 4.955 3.745 5.155 3.945 ;
      RECT 1.74 8.59 1.94 8.79 ;
    LAYER met2 ;
      RECT 2.7 8.4 93.52 8.57 ;
      RECT 93.35 7.275 93.52 8.57 ;
      RECT 2.7 6.255 2.87 8.57 ;
      RECT 93.32 7.275 93.67 7.625 ;
      RECT 2.645 6.255 2.935 6.605 ;
      RECT 90.165 6.225 90.485 6.545 ;
      RECT 90.195 5.695 90.365 6.545 ;
      RECT 90.195 5.695 90.37 6.045 ;
      RECT 90.195 5.695 91.17 5.87 ;
      RECT 90.995 1.965 91.17 5.87 ;
      RECT 90.94 1.965 91.29 2.315 ;
      RECT 90.965 6.655 91.29 6.98 ;
      RECT 89.85 6.745 91.29 6.915 ;
      RECT 89.85 2.395 90.01 6.915 ;
      RECT 90.165 2.365 90.485 2.685 ;
      RECT 89.85 2.395 90.485 2.565 ;
      RECT 88.52 1.14 88.895 1.51 ;
      RECT 80.44 0.96 80.815 1.33 ;
      RECT 79.005 0.96 79.38 1.33 ;
      RECT 79.005 1.08 88.825 1.25 ;
      RECT 84.95 4.36 88.805 4.53 ;
      RECT 88.635 3.425 88.805 4.53 ;
      RECT 84.95 3.665 85.12 4.53 ;
      RECT 84.895 3.705 85.175 3.985 ;
      RECT 84.915 3.665 85.175 3.985 ;
      RECT 84.555 3.625 84.665 3.885 ;
      RECT 88.545 3.43 88.895 3.78 ;
      RECT 84.415 2.115 84.505 2.375 ;
      RECT 84.945 3.17 84.955 3.3 ;
      RECT 84.935 3.135 84.945 3.454 ;
      RECT 84.855 3.067 84.935 3.534 ;
      RECT 84.885 3.71 84.895 3.93 ;
      RECT 84.865 3.705 84.885 3.919 ;
      RECT 84.835 3.7 84.865 3.904 ;
      RECT 84.845 3.002 84.855 3.61 ;
      RECT 84.825 2.946 84.845 3.625 ;
      RECT 84.815 3.685 84.835 3.89 ;
      RECT 84.815 2.874 84.825 3.645 ;
      RECT 84.785 2.777 84.815 3.885 ;
      RECT 84.765 2.66 84.785 3.885 ;
      RECT 84.735 2.54 84.765 3.885 ;
      RECT 84.725 2.455 84.735 3.885 ;
      RECT 84.715 2.4 84.725 3.885 ;
      RECT 84.705 2.355 84.715 3.104 ;
      RECT 84.695 3.315 84.715 3.885 ;
      RECT 84.695 2.285 84.705 3.061 ;
      RECT 84.675 2.235 84.695 2.996 ;
      RECT 84.685 3.395 84.695 3.885 ;
      RECT 84.665 3.495 84.685 3.885 ;
      RECT 84.615 2.115 84.675 2.824 ;
      RECT 84.605 2.115 84.615 2.66 ;
      RECT 84.595 2.115 84.605 2.61 ;
      RECT 84.545 2.115 84.595 2.54 ;
      RECT 84.525 2.115 84.545 2.455 ;
      RECT 84.505 2.115 84.525 2.41 ;
      RECT 86.895 2.155 87.155 2.415 ;
      RECT 86.885 2.155 87.155 2.365 ;
      RECT 86.855 2.025 87.135 2.305 ;
      RECT 75.375 6.655 75.725 7.005 ;
      RECT 86.62 6.61 86.97 6.96 ;
      RECT 75.375 6.685 86.97 6.885 ;
      RECT 85.895 3.705 86.175 3.985 ;
      RECT 85.935 3.665 86.205 3.925 ;
      RECT 85.925 3.7 86.205 3.925 ;
      RECT 85.935 3.66 86.145 3.985 ;
      RECT 85.935 3.655 86.135 3.985 ;
      RECT 85.975 3.645 86.135 3.985 ;
      RECT 85.945 3.65 86.135 3.985 ;
      RECT 85.985 3.64 86.075 3.985 ;
      RECT 86.005 3.635 86.075 3.985 ;
      RECT 85.315 3.155 85.575 3.415 ;
      RECT 85.365 3.065 85.555 3.415 ;
      RECT 85.395 2.85 85.555 3.415 ;
      RECT 85.485 2.455 85.555 3.415 ;
      RECT 85.505 2.165 85.641 2.893 ;
      RECT 85.445 2.66 85.641 2.893 ;
      RECT 85.465 2.54 85.555 3.415 ;
      RECT 85.505 2.165 85.665 2.558 ;
      RECT 85.505 2.165 85.675 2.455 ;
      RECT 85.495 2.165 85.755 2.425 ;
      RECT 83.825 3.565 83.875 3.825 ;
      RECT 83.735 2.095 83.875 2.355 ;
      RECT 84.235 2.72 84.245 2.808 ;
      RECT 84.225 2.655 84.235 2.854 ;
      RECT 84.215 2.605 84.225 2.9 ;
      RECT 84.165 2.552 84.215 3.039 ;
      RECT 84.155 2.501 84.165 3.23 ;
      RECT 84.115 2.459 84.155 3.335 ;
      RECT 84.095 2.405 84.115 3.472 ;
      RECT 84.085 2.38 84.095 2.688 ;
      RECT 84.085 2.77 84.095 3.542 ;
      RECT 84.075 2.366 84.085 2.673 ;
      RECT 84.075 2.825 84.085 3.825 ;
      RECT 84.055 2.341 84.075 2.655 ;
      RECT 84.035 3 84.075 3.825 ;
      RECT 84.045 2.315 84.055 2.635 ;
      RECT 84.015 2.28 84.045 2.589 ;
      RECT 84.025 3.125 84.035 3.825 ;
      RECT 84.015 3.205 84.025 3.825 ;
      RECT 84.005 2.245 84.015 2.554 ;
      RECT 83.965 3.275 84.015 3.825 ;
      RECT 83.995 2.225 84.005 2.53 ;
      RECT 83.965 2.095 83.995 2.495 ;
      RECT 83.955 2.095 83.965 2.46 ;
      RECT 83.935 3.375 83.965 3.825 ;
      RECT 83.935 2.095 83.955 2.435 ;
      RECT 83.925 2.095 83.935 2.41 ;
      RECT 83.885 3.475 83.935 3.825 ;
      RECT 83.905 2.095 83.925 2.38 ;
      RECT 83.875 2.095 83.905 2.365 ;
      RECT 83.875 3.55 83.885 3.825 ;
      RECT 83.795 2.635 83.835 2.895 ;
      RECT 79.525 2.055 79.785 2.315 ;
      RECT 79.525 2.085 79.805 2.295 ;
      RECT 81.735 1.905 81.915 2.055 ;
      RECT 83.785 2.63 83.795 2.895 ;
      RECT 83.765 2.62 83.785 2.895 ;
      RECT 83.747 2.613 83.765 2.895 ;
      RECT 83.661 2.602 83.747 2.895 ;
      RECT 83.575 2.585 83.661 2.895 ;
      RECT 83.525 2.572 83.575 2.82 ;
      RECT 83.491 2.564 83.525 2.795 ;
      RECT 83.405 2.553 83.491 2.76 ;
      RECT 83.365 2.53 83.405 2.723 ;
      RECT 83.355 2.495 83.365 2.708 ;
      RECT 83.345 2.455 83.355 2.703 ;
      RECT 83.335 2.435 83.345 2.698 ;
      RECT 83.32 2.395 83.335 2.693 ;
      RECT 83.305 2.347 83.32 2.689 ;
      RECT 83.295 2.306 83.305 2.686 ;
      RECT 83.285 2.268 83.295 2.675 ;
      RECT 83.265 2.212 83.285 2.655 ;
      RECT 83.245 2.16 83.265 2.591 ;
      RECT 83.225 2.11 83.245 2.543 ;
      RECT 83.215 2.08 83.225 2.507 ;
      RECT 83.21 2.062 83.215 2.493 ;
      RECT 83.195 2.053 83.21 2.475 ;
      RECT 83.165 2.034 83.195 2.415 ;
      RECT 83.155 2.017 83.165 2.37 ;
      RECT 83.145 2.009 83.155 2.34 ;
      RECT 83.115 1.997 83.145 2.29 ;
      RECT 83.095 1.985 83.115 2.225 ;
      RECT 83.085 1.977 83.095 2.185 ;
      RECT 83.065 1.974 83.085 2.175 ;
      RECT 83.05 1.972 83.065 2.17 ;
      RECT 83.03 1.971 83.05 2.16 ;
      RECT 83.015 1.97 83.03 2.15 ;
      RECT 82.995 1.969 83.015 2.145 ;
      RECT 82.993 1.969 82.995 2.145 ;
      RECT 82.907 1.966 82.993 2.142 ;
      RECT 82.821 1.961 82.907 2.135 ;
      RECT 82.735 1.956 82.821 2.129 ;
      RECT 82.685 1.953 82.735 2.12 ;
      RECT 82.641 1.951 82.685 2.114 ;
      RECT 82.555 1.947 82.641 2.109 ;
      RECT 82.551 1.945 82.555 2.105 ;
      RECT 82.465 1.942 82.551 2.1 ;
      RECT 82.411 1.938 82.465 2.093 ;
      RECT 82.325 1.935 82.411 2.088 ;
      RECT 82.301 1.932 82.325 2.084 ;
      RECT 82.215 1.93 82.301 2.079 ;
      RECT 82.155 1.926 82.215 2.073 ;
      RECT 82.147 1.924 82.155 2.07 ;
      RECT 82.061 1.92 82.147 2.066 ;
      RECT 81.975 1.913 82.061 2.059 ;
      RECT 81.915 1.907 81.975 2.055 ;
      RECT 81.715 1.905 81.735 2.058 ;
      RECT 81.665 1.915 81.715 2.068 ;
      RECT 81.635 1.925 81.665 2.08 ;
      RECT 81.611 1.927 81.635 2.086 ;
      RECT 81.525 1.93 81.611 2.091 ;
      RECT 81.455 1.935 81.525 2.1 ;
      RECT 81.441 1.937 81.455 2.106 ;
      RECT 81.355 1.941 81.441 2.111 ;
      RECT 81.315 1.945 81.355 2.12 ;
      RECT 81.301 1.947 81.315 2.126 ;
      RECT 81.215 1.951 81.301 2.131 ;
      RECT 81.131 1.957 81.215 2.138 ;
      RECT 81.045 1.963 81.131 2.143 ;
      RECT 81.021 1.967 81.045 2.146 ;
      RECT 80.935 1.971 81.021 2.151 ;
      RECT 80.885 1.976 80.935 2.16 ;
      RECT 80.805 1.981 80.885 2.17 ;
      RECT 80.725 1.987 80.805 2.185 ;
      RECT 80.705 1.991 80.725 2.195 ;
      RECT 80.635 1.994 80.705 2.205 ;
      RECT 80.585 1.999 80.635 2.22 ;
      RECT 80.555 2.002 80.585 2.24 ;
      RECT 80.545 2.004 80.555 2.256 ;
      RECT 80.485 2.016 80.545 2.266 ;
      RECT 80.465 2.031 80.485 2.275 ;
      RECT 80.455 2.05 80.465 2.275 ;
      RECT 80.445 2.07 80.455 2.275 ;
      RECT 80.425 2.08 80.445 2.275 ;
      RECT 80.375 2.09 80.425 2.275 ;
      RECT 80.345 2.096 80.375 2.275 ;
      RECT 80.275 2.101 80.345 2.277 ;
      RECT 80.195 2.102 80.275 2.282 ;
      RECT 80.191 2.1 80.195 2.285 ;
      RECT 80.105 2.097 80.191 2.286 ;
      RECT 80.063 2.094 80.105 2.288 ;
      RECT 79.977 2.092 80.063 2.289 ;
      RECT 79.891 2.089 79.977 2.292 ;
      RECT 79.805 2.086 79.891 2.294 ;
      RECT 83.185 3.705 83.215 3.985 ;
      RECT 82.935 3.595 82.955 3.985 ;
      RECT 82.895 3.595 82.955 3.855 ;
      RECT 82.725 2.225 82.755 2.485 ;
      RECT 82.495 2.225 82.555 2.485 ;
      RECT 83.175 3.685 83.185 3.985 ;
      RECT 83.155 3.605 83.175 3.985 ;
      RECT 83.145 3.545 83.155 3.985 ;
      RECT 83.095 3.435 83.145 3.985 ;
      RECT 83.085 3.305 83.095 3.985 ;
      RECT 83.045 3.245 83.085 3.985 ;
      RECT 83.041 3.214 83.045 3.985 ;
      RECT 82.955 3.205 83.041 3.985 ;
      RECT 82.945 3.196 82.955 3.55 ;
      RECT 82.915 3.175 82.945 3.517 ;
      RECT 82.905 3.125 82.915 3.493 ;
      RECT 82.895 3.09 82.905 3.481 ;
      RECT 82.855 3.015 82.895 3.45 ;
      RECT 82.835 2.925 82.855 3.415 ;
      RECT 82.825 2.866 82.835 3.4 ;
      RECT 82.775 2.756 82.825 3.36 ;
      RECT 82.765 2.65 82.775 3.315 ;
      RECT 82.735 2.579 82.765 3.235 ;
      RECT 82.725 2.511 82.735 3.16 ;
      RECT 82.715 2.225 82.725 3.125 ;
      RECT 82.685 2.225 82.715 3.055 ;
      RECT 82.675 2.225 82.685 2.95 ;
      RECT 82.665 2.225 82.675 2.915 ;
      RECT 82.595 2.225 82.665 2.775 ;
      RECT 82.565 2.225 82.595 2.575 ;
      RECT 82.555 2.225 82.565 2.5 ;
      RECT 81.735 3.145 82.015 3.425 ;
      RECT 81.765 3.125 82.035 3.385 ;
      RECT 81.765 3.075 81.995 3.425 ;
      RECT 81.835 3.065 81.995 3.425 ;
      RECT 81.835 2.775 81.985 3.425 ;
      RECT 81.825 2.455 81.975 2.825 ;
      RECT 81.815 2.455 81.975 2.695 ;
      RECT 81.795 2.165 81.965 2.5 ;
      RECT 81.775 2.165 81.965 2.45 ;
      RECT 81.735 2.165 81.995 2.425 ;
      RECT 81.645 3.635 81.725 3.895 ;
      RECT 80.935 2.355 81.055 2.615 ;
      RECT 81.62 3.615 81.645 3.895 ;
      RECT 81.605 3.577 81.62 3.895 ;
      RECT 81.565 3.52 81.605 3.895 ;
      RECT 81.535 3.43 81.565 3.895 ;
      RECT 81.495 3.33 81.535 3.895 ;
      RECT 81.465 3.23 81.495 3.895 ;
      RECT 81.46 3.177 81.465 3.718 ;
      RECT 81.445 3.147 81.46 3.684 ;
      RECT 81.435 3.108 81.445 3.649 ;
      RECT 81.425 3.075 81.435 3.605 ;
      RECT 81.415 3.042 81.425 3.57 ;
      RECT 81.385 2.976 81.415 3.505 ;
      RECT 81.375 2.911 81.385 3.43 ;
      RECT 81.365 2.881 81.375 3.4 ;
      RECT 81.325 2.811 81.365 3.33 ;
      RECT 81.315 2.746 81.325 3.245 ;
      RECT 81.305 2.728 81.315 3.23 ;
      RECT 81.295 2.711 81.305 3.195 ;
      RECT 81.285 2.694 81.295 3.165 ;
      RECT 81.275 2.677 81.285 3.135 ;
      RECT 81.255 2.652 81.275 3.075 ;
      RECT 81.245 2.626 81.255 3.02 ;
      RECT 81.225 2.601 81.245 2.98 ;
      RECT 81.215 2.57 81.225 2.945 ;
      RECT 81.205 2.557 81.215 2.9 ;
      RECT 81.195 2.542 81.205 2.875 ;
      RECT 81.185 2.355 81.195 2.835 ;
      RECT 81.175 2.355 81.185 2.805 ;
      RECT 81.17 2.355 81.175 2.788 ;
      RECT 81.165 2.355 81.17 2.77 ;
      RECT 81.095 2.355 81.165 2.71 ;
      RECT 81.055 2.355 81.095 2.645 ;
      RECT 80.885 3.225 81.145 3.485 ;
      RECT 79.055 3.145 79.135 3.465 ;
      RECT 78.875 3.205 79.025 3.465 ;
      RECT 79.055 3.145 79.165 3.425 ;
      RECT 80.875 3.317 80.885 3.48 ;
      RECT 80.845 3.327 80.875 3.488 ;
      RECT 80.825 3.335 80.845 3.493 ;
      RECT 80.757 3.343 80.825 3.503 ;
      RECT 80.671 3.363 80.757 3.52 ;
      RECT 80.585 3.384 80.671 3.539 ;
      RECT 80.575 3.4 80.585 3.55 ;
      RECT 80.535 3.41 80.575 3.556 ;
      RECT 80.515 3.415 80.535 3.563 ;
      RECT 80.477 3.416 80.515 3.566 ;
      RECT 80.391 3.419 80.477 3.567 ;
      RECT 80.305 3.423 80.391 3.568 ;
      RECT 80.251 3.425 80.305 3.57 ;
      RECT 80.165 3.425 80.251 3.572 ;
      RECT 80.125 3.42 80.165 3.574 ;
      RECT 80.115 3.414 80.125 3.575 ;
      RECT 80.075 3.409 80.115 3.571 ;
      RECT 80.065 3.4 80.075 3.567 ;
      RECT 80.033 3.391 80.065 3.564 ;
      RECT 79.947 3.379 80.033 3.554 ;
      RECT 79.861 3.362 79.947 3.539 ;
      RECT 79.775 3.344 79.861 3.525 ;
      RECT 79.755 3.335 79.775 3.516 ;
      RECT 79.685 3.325 79.755 3.509 ;
      RECT 79.635 3.31 79.685 3.499 ;
      RECT 79.575 3.3 79.635 3.49 ;
      RECT 79.535 3.29 79.575 3.485 ;
      RECT 79.485 3.28 79.535 3.479 ;
      RECT 79.445 3.268 79.485 3.469 ;
      RECT 79.425 3.258 79.445 3.465 ;
      RECT 79.405 3.248 79.425 3.465 ;
      RECT 79.395 3.238 79.405 3.464 ;
      RECT 79.375 3.23 79.395 3.46 ;
      RECT 79.335 3.205 79.375 3.454 ;
      RECT 79.315 3.145 79.335 3.447 ;
      RECT 79.291 3.145 79.315 3.444 ;
      RECT 79.205 3.145 79.291 3.439 ;
      RECT 79.165 3.145 79.205 3.43 ;
      RECT 79.025 3.195 79.055 3.465 ;
      RECT 80.705 2.775 80.965 3.035 ;
      RECT 80.665 2.775 80.965 2.915 ;
      RECT 80.635 2.775 80.965 2.9 ;
      RECT 80.575 2.775 80.965 2.88 ;
      RECT 80.495 2.585 80.775 2.865 ;
      RECT 80.495 2.77 80.845 2.865 ;
      RECT 80.495 2.71 80.835 2.865 ;
      RECT 80.495 2.66 80.785 2.865 ;
      RECT 78.265 3.115 78.525 3.375 ;
      RECT 78.41 1.205 78.525 3.375 ;
      RECT 78.325 2.585 78.525 3.375 ;
      RECT 79.635 2.635 79.895 2.895 ;
      RECT 78.32 2.585 78.525 2.87 ;
      RECT 78.315 2.585 78.525 2.865 ;
      RECT 79.615 2.645 79.895 2.825 ;
      RECT 79.205 2.615 79.345 2.765 ;
      RECT 78.58 1.205 78.66 1.55 ;
      RECT 78.315 1.205 78.525 1.55 ;
      RECT 79.605 2.644 79.615 2.825 ;
      RECT 79.601 2.644 79.605 2.825 ;
      RECT 79.515 2.639 79.601 2.814 ;
      RECT 79.441 2.63 79.515 2.794 ;
      RECT 79.355 2.621 79.441 2.775 ;
      RECT 79.345 2.615 79.355 2.765 ;
      RECT 79.165 2.615 79.205 2.768 ;
      RECT 79.079 2.615 79.165 2.776 ;
      RECT 78.993 2.615 79.079 2.787 ;
      RECT 78.907 2.615 78.993 2.798 ;
      RECT 78.821 2.615 78.907 2.809 ;
      RECT 78.735 2.615 78.821 2.82 ;
      RECT 78.705 2.615 78.735 2.86 ;
      RECT 78.675 2.615 78.705 2.91 ;
      RECT 78.6 2.615 78.675 2.93 ;
      RECT 78.595 2.59 78.6 2.935 ;
      RECT 78.58 2.585 78.595 2.943 ;
      RECT 78.575 1.205 78.58 2.953 ;
      RECT 78.545 1.205 78.575 2.995 ;
      RECT 78.525 1.205 78.545 3.075 ;
      RECT 77.655 2.965 77.675 3.404 ;
      RECT 77.655 2.965 77.761 3.401 ;
      RECT 77.645 3.08 77.761 3.4 ;
      RECT 77.675 2.115 77.805 3.397 ;
      RECT 77.655 2.985 77.815 3.395 ;
      RECT 77.655 3.07 77.825 3.39 ;
      RECT 77.625 3.115 77.825 3.385 ;
      RECT 77.625 3.115 77.835 3.38 ;
      RECT 77.605 3.115 77.865 3.375 ;
      RECT 77.675 2.115 77.835 2.765 ;
      RECT 77.665 2.115 77.835 2.74 ;
      RECT 77.665 2.115 77.855 2.505 ;
      RECT 77.615 2.115 77.875 2.375 ;
      RECT 77.085 2.605 77.375 2.865 ;
      RECT 77.095 2.585 77.375 2.865 ;
      RECT 77.045 2.665 77.375 2.86 ;
      RECT 77.115 2.578 77.285 2.865 ;
      RECT 77.115 2.565 77.241 2.865 ;
      RECT 77.155 2.558 77.241 2.865 ;
      RECT 76.615 3.705 76.895 3.985 ;
      RECT 76.575 3.67 76.875 3.78 ;
      RECT 76.565 3.62 76.855 3.675 ;
      RECT 76.505 3.385 76.765 3.645 ;
      RECT 76.505 3.525 76.845 3.645 ;
      RECT 76.505 3.475 76.825 3.645 ;
      RECT 76.505 3.43 76.815 3.645 ;
      RECT 76.505 3.415 76.785 3.645 ;
      RECT 72.24 6.225 72.56 6.545 ;
      RECT 72.27 5.695 72.44 6.545 ;
      RECT 72.27 5.695 72.445 6.045 ;
      RECT 72.27 5.695 73.245 5.87 ;
      RECT 73.07 1.965 73.245 5.87 ;
      RECT 73.015 1.965 73.365 2.315 ;
      RECT 73.04 6.655 73.365 6.98 ;
      RECT 71.925 6.745 73.365 6.915 ;
      RECT 71.925 2.395 72.085 6.915 ;
      RECT 72.24 2.365 72.56 2.685 ;
      RECT 71.925 2.395 72.56 2.565 ;
      RECT 70.595 1.14 70.97 1.51 ;
      RECT 62.515 0.96 62.89 1.33 ;
      RECT 61.08 0.96 61.455 1.33 ;
      RECT 61.08 1.08 70.9 1.25 ;
      RECT 67.025 4.36 70.88 4.53 ;
      RECT 70.71 3.425 70.88 4.53 ;
      RECT 67.025 3.665 67.195 4.53 ;
      RECT 66.97 3.705 67.25 3.985 ;
      RECT 66.99 3.665 67.25 3.985 ;
      RECT 66.63 3.625 66.74 3.885 ;
      RECT 70.62 3.43 70.97 3.78 ;
      RECT 66.49 2.115 66.58 2.375 ;
      RECT 67.02 3.17 67.03 3.3 ;
      RECT 67.01 3.135 67.02 3.454 ;
      RECT 66.93 3.067 67.01 3.534 ;
      RECT 66.96 3.71 66.97 3.93 ;
      RECT 66.94 3.705 66.96 3.919 ;
      RECT 66.91 3.7 66.94 3.904 ;
      RECT 66.92 3.002 66.93 3.61 ;
      RECT 66.9 2.946 66.92 3.625 ;
      RECT 66.89 3.685 66.91 3.89 ;
      RECT 66.89 2.874 66.9 3.645 ;
      RECT 66.86 2.777 66.89 3.885 ;
      RECT 66.84 2.66 66.86 3.885 ;
      RECT 66.81 2.54 66.84 3.885 ;
      RECT 66.8 2.455 66.81 3.885 ;
      RECT 66.79 2.4 66.8 3.885 ;
      RECT 66.78 2.355 66.79 3.104 ;
      RECT 66.77 3.315 66.79 3.885 ;
      RECT 66.77 2.285 66.78 3.061 ;
      RECT 66.75 2.235 66.77 2.996 ;
      RECT 66.76 3.395 66.77 3.885 ;
      RECT 66.74 3.495 66.76 3.885 ;
      RECT 66.69 2.115 66.75 2.824 ;
      RECT 66.68 2.115 66.69 2.66 ;
      RECT 66.67 2.115 66.68 2.61 ;
      RECT 66.62 2.115 66.67 2.54 ;
      RECT 66.6 2.115 66.62 2.455 ;
      RECT 66.58 2.115 66.6 2.41 ;
      RECT 68.97 2.155 69.23 2.415 ;
      RECT 68.96 2.155 69.23 2.365 ;
      RECT 68.93 2.025 69.21 2.305 ;
      RECT 57.45 6.655 57.8 7.005 ;
      RECT 68.415 6.61 68.765 6.96 ;
      RECT 57.45 6.685 68.765 6.885 ;
      RECT 67.97 3.705 68.25 3.985 ;
      RECT 68.01 3.665 68.28 3.925 ;
      RECT 68 3.7 68.28 3.925 ;
      RECT 68.01 3.66 68.22 3.985 ;
      RECT 68.01 3.655 68.21 3.985 ;
      RECT 68.05 3.645 68.21 3.985 ;
      RECT 68.02 3.65 68.21 3.985 ;
      RECT 68.06 3.64 68.15 3.985 ;
      RECT 68.08 3.635 68.15 3.985 ;
      RECT 67.39 3.155 67.65 3.415 ;
      RECT 67.44 3.065 67.63 3.415 ;
      RECT 67.47 2.85 67.63 3.415 ;
      RECT 67.56 2.455 67.63 3.415 ;
      RECT 67.58 2.165 67.716 2.893 ;
      RECT 67.52 2.66 67.716 2.893 ;
      RECT 67.54 2.54 67.63 3.415 ;
      RECT 67.58 2.165 67.74 2.558 ;
      RECT 67.58 2.165 67.75 2.455 ;
      RECT 67.57 2.165 67.83 2.425 ;
      RECT 65.9 3.565 65.95 3.825 ;
      RECT 65.81 2.095 65.95 2.355 ;
      RECT 66.31 2.72 66.32 2.808 ;
      RECT 66.3 2.655 66.31 2.854 ;
      RECT 66.29 2.605 66.3 2.9 ;
      RECT 66.24 2.552 66.29 3.039 ;
      RECT 66.23 2.501 66.24 3.23 ;
      RECT 66.19 2.459 66.23 3.335 ;
      RECT 66.17 2.405 66.19 3.472 ;
      RECT 66.16 2.38 66.17 2.688 ;
      RECT 66.16 2.77 66.17 3.542 ;
      RECT 66.15 2.366 66.16 2.673 ;
      RECT 66.15 2.825 66.16 3.825 ;
      RECT 66.13 2.341 66.15 2.655 ;
      RECT 66.11 3 66.15 3.825 ;
      RECT 66.12 2.315 66.13 2.635 ;
      RECT 66.09 2.28 66.12 2.589 ;
      RECT 66.1 3.125 66.11 3.825 ;
      RECT 66.09 3.205 66.1 3.825 ;
      RECT 66.08 2.245 66.09 2.554 ;
      RECT 66.04 3.275 66.09 3.825 ;
      RECT 66.07 2.225 66.08 2.53 ;
      RECT 66.04 2.095 66.07 2.495 ;
      RECT 66.03 2.095 66.04 2.46 ;
      RECT 66.01 3.375 66.04 3.825 ;
      RECT 66.01 2.095 66.03 2.435 ;
      RECT 66 2.095 66.01 2.41 ;
      RECT 65.96 3.475 66.01 3.825 ;
      RECT 65.98 2.095 66 2.38 ;
      RECT 65.95 2.095 65.98 2.365 ;
      RECT 65.95 3.55 65.96 3.825 ;
      RECT 65.87 2.635 65.91 2.895 ;
      RECT 61.6 2.055 61.86 2.315 ;
      RECT 61.6 2.085 61.88 2.295 ;
      RECT 63.81 1.905 63.99 2.055 ;
      RECT 65.86 2.63 65.87 2.895 ;
      RECT 65.84 2.62 65.86 2.895 ;
      RECT 65.822 2.613 65.84 2.895 ;
      RECT 65.736 2.602 65.822 2.895 ;
      RECT 65.65 2.585 65.736 2.895 ;
      RECT 65.6 2.572 65.65 2.82 ;
      RECT 65.566 2.564 65.6 2.795 ;
      RECT 65.48 2.553 65.566 2.76 ;
      RECT 65.44 2.53 65.48 2.723 ;
      RECT 65.43 2.495 65.44 2.708 ;
      RECT 65.42 2.455 65.43 2.703 ;
      RECT 65.41 2.435 65.42 2.698 ;
      RECT 65.395 2.395 65.41 2.693 ;
      RECT 65.38 2.347 65.395 2.689 ;
      RECT 65.37 2.306 65.38 2.686 ;
      RECT 65.36 2.268 65.37 2.675 ;
      RECT 65.34 2.212 65.36 2.655 ;
      RECT 65.32 2.16 65.34 2.591 ;
      RECT 65.3 2.11 65.32 2.543 ;
      RECT 65.29 2.08 65.3 2.507 ;
      RECT 65.285 2.062 65.29 2.493 ;
      RECT 65.27 2.053 65.285 2.475 ;
      RECT 65.24 2.034 65.27 2.415 ;
      RECT 65.23 2.017 65.24 2.37 ;
      RECT 65.22 2.009 65.23 2.34 ;
      RECT 65.19 1.997 65.22 2.29 ;
      RECT 65.17 1.985 65.19 2.225 ;
      RECT 65.16 1.977 65.17 2.185 ;
      RECT 65.14 1.974 65.16 2.175 ;
      RECT 65.125 1.972 65.14 2.17 ;
      RECT 65.105 1.971 65.125 2.16 ;
      RECT 65.09 1.97 65.105 2.15 ;
      RECT 65.07 1.969 65.09 2.145 ;
      RECT 65.068 1.969 65.07 2.145 ;
      RECT 64.982 1.966 65.068 2.142 ;
      RECT 64.896 1.961 64.982 2.135 ;
      RECT 64.81 1.956 64.896 2.129 ;
      RECT 64.76 1.953 64.81 2.12 ;
      RECT 64.716 1.951 64.76 2.114 ;
      RECT 64.63 1.947 64.716 2.109 ;
      RECT 64.626 1.945 64.63 2.105 ;
      RECT 64.54 1.942 64.626 2.1 ;
      RECT 64.486 1.938 64.54 2.093 ;
      RECT 64.4 1.935 64.486 2.088 ;
      RECT 64.376 1.932 64.4 2.084 ;
      RECT 64.29 1.93 64.376 2.079 ;
      RECT 64.23 1.926 64.29 2.073 ;
      RECT 64.222 1.924 64.23 2.07 ;
      RECT 64.136 1.92 64.222 2.066 ;
      RECT 64.05 1.913 64.136 2.059 ;
      RECT 63.99 1.907 64.05 2.055 ;
      RECT 63.79 1.905 63.81 2.058 ;
      RECT 63.74 1.915 63.79 2.068 ;
      RECT 63.71 1.925 63.74 2.08 ;
      RECT 63.686 1.927 63.71 2.086 ;
      RECT 63.6 1.93 63.686 2.091 ;
      RECT 63.53 1.935 63.6 2.1 ;
      RECT 63.516 1.937 63.53 2.106 ;
      RECT 63.43 1.941 63.516 2.111 ;
      RECT 63.39 1.945 63.43 2.12 ;
      RECT 63.376 1.947 63.39 2.126 ;
      RECT 63.29 1.951 63.376 2.131 ;
      RECT 63.206 1.957 63.29 2.138 ;
      RECT 63.12 1.963 63.206 2.143 ;
      RECT 63.096 1.967 63.12 2.146 ;
      RECT 63.01 1.971 63.096 2.151 ;
      RECT 62.96 1.976 63.01 2.16 ;
      RECT 62.88 1.981 62.96 2.17 ;
      RECT 62.8 1.987 62.88 2.185 ;
      RECT 62.78 1.991 62.8 2.195 ;
      RECT 62.71 1.994 62.78 2.205 ;
      RECT 62.66 1.999 62.71 2.22 ;
      RECT 62.63 2.002 62.66 2.24 ;
      RECT 62.62 2.004 62.63 2.256 ;
      RECT 62.56 2.016 62.62 2.266 ;
      RECT 62.54 2.031 62.56 2.275 ;
      RECT 62.53 2.05 62.54 2.275 ;
      RECT 62.52 2.07 62.53 2.275 ;
      RECT 62.5 2.08 62.52 2.275 ;
      RECT 62.45 2.09 62.5 2.275 ;
      RECT 62.42 2.096 62.45 2.275 ;
      RECT 62.35 2.101 62.42 2.277 ;
      RECT 62.27 2.102 62.35 2.282 ;
      RECT 62.266 2.1 62.27 2.285 ;
      RECT 62.18 2.097 62.266 2.286 ;
      RECT 62.138 2.094 62.18 2.288 ;
      RECT 62.052 2.092 62.138 2.289 ;
      RECT 61.966 2.089 62.052 2.292 ;
      RECT 61.88 2.086 61.966 2.294 ;
      RECT 65.26 3.705 65.29 3.985 ;
      RECT 65.01 3.595 65.03 3.985 ;
      RECT 64.97 3.595 65.03 3.855 ;
      RECT 64.8 2.225 64.83 2.485 ;
      RECT 64.57 2.225 64.63 2.485 ;
      RECT 65.25 3.685 65.26 3.985 ;
      RECT 65.23 3.605 65.25 3.985 ;
      RECT 65.22 3.545 65.23 3.985 ;
      RECT 65.17 3.435 65.22 3.985 ;
      RECT 65.16 3.305 65.17 3.985 ;
      RECT 65.12 3.245 65.16 3.985 ;
      RECT 65.116 3.214 65.12 3.985 ;
      RECT 65.03 3.205 65.116 3.985 ;
      RECT 65.02 3.196 65.03 3.55 ;
      RECT 64.99 3.175 65.02 3.517 ;
      RECT 64.98 3.125 64.99 3.493 ;
      RECT 64.97 3.09 64.98 3.481 ;
      RECT 64.93 3.015 64.97 3.45 ;
      RECT 64.91 2.925 64.93 3.415 ;
      RECT 64.9 2.866 64.91 3.4 ;
      RECT 64.85 2.756 64.9 3.36 ;
      RECT 64.84 2.65 64.85 3.315 ;
      RECT 64.81 2.579 64.84 3.235 ;
      RECT 64.8 2.511 64.81 3.16 ;
      RECT 64.79 2.225 64.8 3.125 ;
      RECT 64.76 2.225 64.79 3.055 ;
      RECT 64.75 2.225 64.76 2.95 ;
      RECT 64.74 2.225 64.75 2.915 ;
      RECT 64.67 2.225 64.74 2.775 ;
      RECT 64.64 2.225 64.67 2.575 ;
      RECT 64.63 2.225 64.64 2.5 ;
      RECT 63.81 3.145 64.09 3.425 ;
      RECT 63.84 3.125 64.11 3.385 ;
      RECT 63.84 3.075 64.07 3.425 ;
      RECT 63.91 3.065 64.07 3.425 ;
      RECT 63.91 2.775 64.06 3.425 ;
      RECT 63.9 2.455 64.05 2.825 ;
      RECT 63.89 2.455 64.05 2.695 ;
      RECT 63.87 2.165 64.04 2.5 ;
      RECT 63.85 2.165 64.04 2.45 ;
      RECT 63.81 2.165 64.07 2.425 ;
      RECT 63.72 3.635 63.8 3.895 ;
      RECT 63.01 2.355 63.13 2.615 ;
      RECT 63.695 3.615 63.72 3.895 ;
      RECT 63.68 3.577 63.695 3.895 ;
      RECT 63.64 3.52 63.68 3.895 ;
      RECT 63.61 3.43 63.64 3.895 ;
      RECT 63.57 3.33 63.61 3.895 ;
      RECT 63.54 3.23 63.57 3.895 ;
      RECT 63.535 3.177 63.54 3.718 ;
      RECT 63.52 3.147 63.535 3.684 ;
      RECT 63.51 3.108 63.52 3.649 ;
      RECT 63.5 3.075 63.51 3.605 ;
      RECT 63.49 3.042 63.5 3.57 ;
      RECT 63.46 2.976 63.49 3.505 ;
      RECT 63.45 2.911 63.46 3.43 ;
      RECT 63.44 2.881 63.45 3.4 ;
      RECT 63.4 2.811 63.44 3.33 ;
      RECT 63.39 2.746 63.4 3.245 ;
      RECT 63.38 2.728 63.39 3.23 ;
      RECT 63.37 2.711 63.38 3.195 ;
      RECT 63.36 2.694 63.37 3.165 ;
      RECT 63.35 2.677 63.36 3.135 ;
      RECT 63.33 2.652 63.35 3.075 ;
      RECT 63.32 2.626 63.33 3.02 ;
      RECT 63.3 2.601 63.32 2.98 ;
      RECT 63.29 2.57 63.3 2.945 ;
      RECT 63.28 2.557 63.29 2.9 ;
      RECT 63.27 2.542 63.28 2.875 ;
      RECT 63.26 2.355 63.27 2.835 ;
      RECT 63.25 2.355 63.26 2.805 ;
      RECT 63.245 2.355 63.25 2.788 ;
      RECT 63.24 2.355 63.245 2.77 ;
      RECT 63.17 2.355 63.24 2.71 ;
      RECT 63.13 2.355 63.17 2.645 ;
      RECT 62.96 3.225 63.22 3.485 ;
      RECT 61.13 3.145 61.21 3.465 ;
      RECT 60.95 3.205 61.1 3.465 ;
      RECT 61.13 3.145 61.24 3.425 ;
      RECT 62.95 3.317 62.96 3.48 ;
      RECT 62.92 3.327 62.95 3.488 ;
      RECT 62.9 3.335 62.92 3.493 ;
      RECT 62.832 3.343 62.9 3.503 ;
      RECT 62.746 3.363 62.832 3.52 ;
      RECT 62.66 3.384 62.746 3.539 ;
      RECT 62.65 3.4 62.66 3.55 ;
      RECT 62.61 3.41 62.65 3.556 ;
      RECT 62.59 3.415 62.61 3.563 ;
      RECT 62.552 3.416 62.59 3.566 ;
      RECT 62.466 3.419 62.552 3.567 ;
      RECT 62.38 3.423 62.466 3.568 ;
      RECT 62.326 3.425 62.38 3.57 ;
      RECT 62.24 3.425 62.326 3.572 ;
      RECT 62.2 3.42 62.24 3.574 ;
      RECT 62.19 3.414 62.2 3.575 ;
      RECT 62.15 3.409 62.19 3.571 ;
      RECT 62.14 3.4 62.15 3.567 ;
      RECT 62.108 3.391 62.14 3.564 ;
      RECT 62.022 3.379 62.108 3.554 ;
      RECT 61.936 3.362 62.022 3.539 ;
      RECT 61.85 3.344 61.936 3.525 ;
      RECT 61.83 3.335 61.85 3.516 ;
      RECT 61.76 3.325 61.83 3.509 ;
      RECT 61.71 3.31 61.76 3.499 ;
      RECT 61.65 3.3 61.71 3.49 ;
      RECT 61.61 3.29 61.65 3.485 ;
      RECT 61.56 3.28 61.61 3.479 ;
      RECT 61.52 3.268 61.56 3.469 ;
      RECT 61.5 3.258 61.52 3.465 ;
      RECT 61.48 3.248 61.5 3.465 ;
      RECT 61.47 3.238 61.48 3.464 ;
      RECT 61.45 3.23 61.47 3.46 ;
      RECT 61.41 3.205 61.45 3.454 ;
      RECT 61.39 3.145 61.41 3.447 ;
      RECT 61.366 3.145 61.39 3.444 ;
      RECT 61.28 3.145 61.366 3.439 ;
      RECT 61.24 3.145 61.28 3.43 ;
      RECT 61.1 3.195 61.13 3.465 ;
      RECT 62.78 2.775 63.04 3.035 ;
      RECT 62.74 2.775 63.04 2.915 ;
      RECT 62.71 2.775 63.04 2.9 ;
      RECT 62.65 2.775 63.04 2.88 ;
      RECT 62.57 2.585 62.85 2.865 ;
      RECT 62.57 2.77 62.92 2.865 ;
      RECT 62.57 2.71 62.91 2.865 ;
      RECT 62.57 2.66 62.86 2.865 ;
      RECT 60.34 3.115 60.6 3.375 ;
      RECT 60.485 1.205 60.6 3.375 ;
      RECT 60.4 2.585 60.6 3.375 ;
      RECT 61.71 2.635 61.97 2.895 ;
      RECT 60.395 2.585 60.6 2.87 ;
      RECT 60.39 2.585 60.6 2.865 ;
      RECT 61.69 2.645 61.97 2.825 ;
      RECT 61.28 2.615 61.42 2.765 ;
      RECT 60.655 1.205 60.735 1.55 ;
      RECT 60.39 1.205 60.6 1.55 ;
      RECT 61.68 2.644 61.69 2.825 ;
      RECT 61.676 2.644 61.68 2.825 ;
      RECT 61.59 2.639 61.676 2.814 ;
      RECT 61.516 2.63 61.59 2.794 ;
      RECT 61.43 2.621 61.516 2.775 ;
      RECT 61.42 2.615 61.43 2.765 ;
      RECT 61.24 2.615 61.28 2.768 ;
      RECT 61.154 2.615 61.24 2.776 ;
      RECT 61.068 2.615 61.154 2.787 ;
      RECT 60.982 2.615 61.068 2.798 ;
      RECT 60.896 2.615 60.982 2.809 ;
      RECT 60.81 2.615 60.896 2.82 ;
      RECT 60.78 2.615 60.81 2.86 ;
      RECT 60.75 2.615 60.78 2.91 ;
      RECT 60.675 2.615 60.75 2.93 ;
      RECT 60.67 2.59 60.675 2.935 ;
      RECT 60.655 2.585 60.67 2.943 ;
      RECT 60.65 1.205 60.655 2.953 ;
      RECT 60.62 1.205 60.65 2.995 ;
      RECT 60.6 1.205 60.62 3.075 ;
      RECT 59.73 2.965 59.75 3.404 ;
      RECT 59.73 2.965 59.836 3.401 ;
      RECT 59.72 3.08 59.836 3.4 ;
      RECT 59.75 2.115 59.88 3.397 ;
      RECT 59.73 2.985 59.89 3.395 ;
      RECT 59.73 3.07 59.9 3.39 ;
      RECT 59.7 3.115 59.9 3.385 ;
      RECT 59.7 3.115 59.91 3.38 ;
      RECT 59.68 3.115 59.94 3.375 ;
      RECT 59.75 2.115 59.91 2.765 ;
      RECT 59.74 2.115 59.91 2.74 ;
      RECT 59.74 2.115 59.93 2.505 ;
      RECT 59.69 2.115 59.95 2.375 ;
      RECT 59.16 2.605 59.45 2.865 ;
      RECT 59.17 2.585 59.45 2.865 ;
      RECT 59.12 2.665 59.45 2.86 ;
      RECT 59.19 2.578 59.36 2.865 ;
      RECT 59.19 2.565 59.316 2.865 ;
      RECT 59.23 2.558 59.316 2.865 ;
      RECT 58.69 3.705 58.97 3.985 ;
      RECT 58.65 3.67 58.95 3.78 ;
      RECT 58.64 3.62 58.93 3.675 ;
      RECT 58.58 3.385 58.84 3.645 ;
      RECT 58.58 3.525 58.92 3.645 ;
      RECT 58.58 3.475 58.9 3.645 ;
      RECT 58.58 3.43 58.89 3.645 ;
      RECT 58.58 3.415 58.86 3.645 ;
      RECT 54.315 6.225 54.635 6.545 ;
      RECT 54.345 5.695 54.515 6.545 ;
      RECT 54.345 5.695 54.52 6.045 ;
      RECT 54.345 5.695 55.32 5.87 ;
      RECT 55.145 1.965 55.32 5.87 ;
      RECT 55.09 1.965 55.44 2.315 ;
      RECT 55.115 6.655 55.44 6.98 ;
      RECT 54 6.745 55.44 6.915 ;
      RECT 54 2.395 54.16 6.915 ;
      RECT 54.315 2.365 54.635 2.685 ;
      RECT 54 2.395 54.635 2.565 ;
      RECT 52.67 1.14 53.045 1.51 ;
      RECT 44.59 0.96 44.965 1.33 ;
      RECT 43.155 0.96 43.53 1.33 ;
      RECT 43.155 1.08 52.975 1.25 ;
      RECT 49.1 4.36 52.955 4.53 ;
      RECT 52.785 3.425 52.955 4.53 ;
      RECT 49.1 3.665 49.27 4.53 ;
      RECT 49.045 3.705 49.325 3.985 ;
      RECT 49.065 3.665 49.325 3.985 ;
      RECT 48.705 3.625 48.815 3.885 ;
      RECT 52.695 3.43 53.045 3.78 ;
      RECT 48.565 2.115 48.655 2.375 ;
      RECT 49.095 3.17 49.105 3.3 ;
      RECT 49.085 3.135 49.095 3.454 ;
      RECT 49.005 3.067 49.085 3.534 ;
      RECT 49.035 3.71 49.045 3.93 ;
      RECT 49.015 3.705 49.035 3.919 ;
      RECT 48.985 3.7 49.015 3.904 ;
      RECT 48.995 3.002 49.005 3.61 ;
      RECT 48.975 2.946 48.995 3.625 ;
      RECT 48.965 3.685 48.985 3.89 ;
      RECT 48.965 2.874 48.975 3.645 ;
      RECT 48.935 2.777 48.965 3.885 ;
      RECT 48.915 2.66 48.935 3.885 ;
      RECT 48.885 2.54 48.915 3.885 ;
      RECT 48.875 2.455 48.885 3.885 ;
      RECT 48.865 2.4 48.875 3.885 ;
      RECT 48.855 2.355 48.865 3.104 ;
      RECT 48.845 3.315 48.865 3.885 ;
      RECT 48.845 2.285 48.855 3.061 ;
      RECT 48.825 2.235 48.845 2.996 ;
      RECT 48.835 3.395 48.845 3.885 ;
      RECT 48.815 3.495 48.835 3.885 ;
      RECT 48.765 2.115 48.825 2.824 ;
      RECT 48.755 2.115 48.765 2.66 ;
      RECT 48.745 2.115 48.755 2.61 ;
      RECT 48.695 2.115 48.745 2.54 ;
      RECT 48.675 2.115 48.695 2.455 ;
      RECT 48.655 2.115 48.675 2.41 ;
      RECT 51.045 2.155 51.305 2.415 ;
      RECT 51.035 2.155 51.305 2.365 ;
      RECT 51.005 2.025 51.285 2.305 ;
      RECT 39.57 6.66 39.92 7.01 ;
      RECT 50.545 6.615 50.895 6.965 ;
      RECT 39.57 6.69 50.895 6.89 ;
      RECT 50.045 3.705 50.325 3.985 ;
      RECT 50.085 3.665 50.355 3.925 ;
      RECT 50.075 3.7 50.355 3.925 ;
      RECT 50.085 3.66 50.295 3.985 ;
      RECT 50.085 3.655 50.285 3.985 ;
      RECT 50.125 3.645 50.285 3.985 ;
      RECT 50.095 3.65 50.285 3.985 ;
      RECT 50.135 3.64 50.225 3.985 ;
      RECT 50.155 3.635 50.225 3.985 ;
      RECT 49.465 3.155 49.725 3.415 ;
      RECT 49.515 3.065 49.705 3.415 ;
      RECT 49.545 2.85 49.705 3.415 ;
      RECT 49.635 2.455 49.705 3.415 ;
      RECT 49.655 2.165 49.791 2.893 ;
      RECT 49.595 2.66 49.791 2.893 ;
      RECT 49.615 2.54 49.705 3.415 ;
      RECT 49.655 2.165 49.815 2.558 ;
      RECT 49.655 2.165 49.825 2.455 ;
      RECT 49.645 2.165 49.905 2.425 ;
      RECT 47.975 3.565 48.025 3.825 ;
      RECT 47.885 2.095 48.025 2.355 ;
      RECT 48.385 2.72 48.395 2.808 ;
      RECT 48.375 2.655 48.385 2.854 ;
      RECT 48.365 2.605 48.375 2.9 ;
      RECT 48.315 2.552 48.365 3.039 ;
      RECT 48.305 2.501 48.315 3.23 ;
      RECT 48.265 2.459 48.305 3.335 ;
      RECT 48.245 2.405 48.265 3.472 ;
      RECT 48.235 2.38 48.245 2.688 ;
      RECT 48.235 2.77 48.245 3.542 ;
      RECT 48.225 2.366 48.235 2.673 ;
      RECT 48.225 2.825 48.235 3.825 ;
      RECT 48.205 2.341 48.225 2.655 ;
      RECT 48.185 3 48.225 3.825 ;
      RECT 48.195 2.315 48.205 2.635 ;
      RECT 48.165 2.28 48.195 2.589 ;
      RECT 48.175 3.125 48.185 3.825 ;
      RECT 48.165 3.205 48.175 3.825 ;
      RECT 48.155 2.245 48.165 2.554 ;
      RECT 48.115 3.275 48.165 3.825 ;
      RECT 48.145 2.225 48.155 2.53 ;
      RECT 48.115 2.095 48.145 2.495 ;
      RECT 48.105 2.095 48.115 2.46 ;
      RECT 48.085 3.375 48.115 3.825 ;
      RECT 48.085 2.095 48.105 2.435 ;
      RECT 48.075 2.095 48.085 2.41 ;
      RECT 48.035 3.475 48.085 3.825 ;
      RECT 48.055 2.095 48.075 2.38 ;
      RECT 48.025 2.095 48.055 2.365 ;
      RECT 48.025 3.55 48.035 3.825 ;
      RECT 47.945 2.635 47.985 2.895 ;
      RECT 43.675 2.055 43.935 2.315 ;
      RECT 43.675 2.085 43.955 2.295 ;
      RECT 45.885 1.905 46.065 2.055 ;
      RECT 47.935 2.63 47.945 2.895 ;
      RECT 47.915 2.62 47.935 2.895 ;
      RECT 47.897 2.613 47.915 2.895 ;
      RECT 47.811 2.602 47.897 2.895 ;
      RECT 47.725 2.585 47.811 2.895 ;
      RECT 47.675 2.572 47.725 2.82 ;
      RECT 47.641 2.564 47.675 2.795 ;
      RECT 47.555 2.553 47.641 2.76 ;
      RECT 47.515 2.53 47.555 2.723 ;
      RECT 47.505 2.495 47.515 2.708 ;
      RECT 47.495 2.455 47.505 2.703 ;
      RECT 47.485 2.435 47.495 2.698 ;
      RECT 47.47 2.395 47.485 2.693 ;
      RECT 47.455 2.347 47.47 2.689 ;
      RECT 47.445 2.306 47.455 2.686 ;
      RECT 47.435 2.268 47.445 2.675 ;
      RECT 47.415 2.212 47.435 2.655 ;
      RECT 47.395 2.16 47.415 2.591 ;
      RECT 47.375 2.11 47.395 2.543 ;
      RECT 47.365 2.08 47.375 2.507 ;
      RECT 47.36 2.062 47.365 2.493 ;
      RECT 47.345 2.053 47.36 2.475 ;
      RECT 47.315 2.034 47.345 2.415 ;
      RECT 47.305 2.017 47.315 2.37 ;
      RECT 47.295 2.009 47.305 2.34 ;
      RECT 47.265 1.997 47.295 2.29 ;
      RECT 47.245 1.985 47.265 2.225 ;
      RECT 47.235 1.977 47.245 2.185 ;
      RECT 47.215 1.974 47.235 2.175 ;
      RECT 47.2 1.972 47.215 2.17 ;
      RECT 47.18 1.971 47.2 2.16 ;
      RECT 47.165 1.97 47.18 2.15 ;
      RECT 47.145 1.969 47.165 2.145 ;
      RECT 47.143 1.969 47.145 2.145 ;
      RECT 47.057 1.966 47.143 2.142 ;
      RECT 46.971 1.961 47.057 2.135 ;
      RECT 46.885 1.956 46.971 2.129 ;
      RECT 46.835 1.953 46.885 2.12 ;
      RECT 46.791 1.951 46.835 2.114 ;
      RECT 46.705 1.947 46.791 2.109 ;
      RECT 46.701 1.945 46.705 2.105 ;
      RECT 46.615 1.942 46.701 2.1 ;
      RECT 46.561 1.938 46.615 2.093 ;
      RECT 46.475 1.935 46.561 2.088 ;
      RECT 46.451 1.932 46.475 2.084 ;
      RECT 46.365 1.93 46.451 2.079 ;
      RECT 46.305 1.926 46.365 2.073 ;
      RECT 46.297 1.924 46.305 2.07 ;
      RECT 46.211 1.92 46.297 2.066 ;
      RECT 46.125 1.913 46.211 2.059 ;
      RECT 46.065 1.907 46.125 2.055 ;
      RECT 45.865 1.905 45.885 2.058 ;
      RECT 45.815 1.915 45.865 2.068 ;
      RECT 45.785 1.925 45.815 2.08 ;
      RECT 45.761 1.927 45.785 2.086 ;
      RECT 45.675 1.93 45.761 2.091 ;
      RECT 45.605 1.935 45.675 2.1 ;
      RECT 45.591 1.937 45.605 2.106 ;
      RECT 45.505 1.941 45.591 2.111 ;
      RECT 45.465 1.945 45.505 2.12 ;
      RECT 45.451 1.947 45.465 2.126 ;
      RECT 45.365 1.951 45.451 2.131 ;
      RECT 45.281 1.957 45.365 2.138 ;
      RECT 45.195 1.963 45.281 2.143 ;
      RECT 45.171 1.967 45.195 2.146 ;
      RECT 45.085 1.971 45.171 2.151 ;
      RECT 45.035 1.976 45.085 2.16 ;
      RECT 44.955 1.981 45.035 2.17 ;
      RECT 44.875 1.987 44.955 2.185 ;
      RECT 44.855 1.991 44.875 2.195 ;
      RECT 44.785 1.994 44.855 2.205 ;
      RECT 44.735 1.999 44.785 2.22 ;
      RECT 44.705 2.002 44.735 2.24 ;
      RECT 44.695 2.004 44.705 2.256 ;
      RECT 44.635 2.016 44.695 2.266 ;
      RECT 44.615 2.031 44.635 2.275 ;
      RECT 44.605 2.05 44.615 2.275 ;
      RECT 44.595 2.07 44.605 2.275 ;
      RECT 44.575 2.08 44.595 2.275 ;
      RECT 44.525 2.09 44.575 2.275 ;
      RECT 44.495 2.096 44.525 2.275 ;
      RECT 44.425 2.101 44.495 2.277 ;
      RECT 44.345 2.102 44.425 2.282 ;
      RECT 44.341 2.1 44.345 2.285 ;
      RECT 44.255 2.097 44.341 2.286 ;
      RECT 44.213 2.094 44.255 2.288 ;
      RECT 44.127 2.092 44.213 2.289 ;
      RECT 44.041 2.089 44.127 2.292 ;
      RECT 43.955 2.086 44.041 2.294 ;
      RECT 47.335 3.705 47.365 3.985 ;
      RECT 47.085 3.595 47.105 3.985 ;
      RECT 47.045 3.595 47.105 3.855 ;
      RECT 46.875 2.225 46.905 2.485 ;
      RECT 46.645 2.225 46.705 2.485 ;
      RECT 47.325 3.685 47.335 3.985 ;
      RECT 47.305 3.605 47.325 3.985 ;
      RECT 47.295 3.545 47.305 3.985 ;
      RECT 47.245 3.435 47.295 3.985 ;
      RECT 47.235 3.305 47.245 3.985 ;
      RECT 47.195 3.245 47.235 3.985 ;
      RECT 47.191 3.214 47.195 3.985 ;
      RECT 47.105 3.205 47.191 3.985 ;
      RECT 47.095 3.196 47.105 3.55 ;
      RECT 47.065 3.175 47.095 3.517 ;
      RECT 47.055 3.125 47.065 3.493 ;
      RECT 47.045 3.09 47.055 3.481 ;
      RECT 47.005 3.015 47.045 3.45 ;
      RECT 46.985 2.925 47.005 3.415 ;
      RECT 46.975 2.866 46.985 3.4 ;
      RECT 46.925 2.756 46.975 3.36 ;
      RECT 46.915 2.65 46.925 3.315 ;
      RECT 46.885 2.579 46.915 3.235 ;
      RECT 46.875 2.511 46.885 3.16 ;
      RECT 46.865 2.225 46.875 3.125 ;
      RECT 46.835 2.225 46.865 3.055 ;
      RECT 46.825 2.225 46.835 2.95 ;
      RECT 46.815 2.225 46.825 2.915 ;
      RECT 46.745 2.225 46.815 2.775 ;
      RECT 46.715 2.225 46.745 2.575 ;
      RECT 46.705 2.225 46.715 2.5 ;
      RECT 45.885 3.145 46.165 3.425 ;
      RECT 45.915 3.125 46.185 3.385 ;
      RECT 45.915 3.075 46.145 3.425 ;
      RECT 45.985 3.065 46.145 3.425 ;
      RECT 45.985 2.775 46.135 3.425 ;
      RECT 45.975 2.455 46.125 2.825 ;
      RECT 45.965 2.455 46.125 2.695 ;
      RECT 45.945 2.165 46.115 2.5 ;
      RECT 45.925 2.165 46.115 2.45 ;
      RECT 45.885 2.165 46.145 2.425 ;
      RECT 45.795 3.635 45.875 3.895 ;
      RECT 45.085 2.355 45.205 2.615 ;
      RECT 45.77 3.615 45.795 3.895 ;
      RECT 45.755 3.577 45.77 3.895 ;
      RECT 45.715 3.52 45.755 3.895 ;
      RECT 45.685 3.43 45.715 3.895 ;
      RECT 45.645 3.33 45.685 3.895 ;
      RECT 45.615 3.23 45.645 3.895 ;
      RECT 45.61 3.177 45.615 3.718 ;
      RECT 45.595 3.147 45.61 3.684 ;
      RECT 45.585 3.108 45.595 3.649 ;
      RECT 45.575 3.075 45.585 3.605 ;
      RECT 45.565 3.042 45.575 3.57 ;
      RECT 45.535 2.976 45.565 3.505 ;
      RECT 45.525 2.911 45.535 3.43 ;
      RECT 45.515 2.881 45.525 3.4 ;
      RECT 45.475 2.811 45.515 3.33 ;
      RECT 45.465 2.746 45.475 3.245 ;
      RECT 45.455 2.728 45.465 3.23 ;
      RECT 45.445 2.711 45.455 3.195 ;
      RECT 45.435 2.694 45.445 3.165 ;
      RECT 45.425 2.677 45.435 3.135 ;
      RECT 45.405 2.652 45.425 3.075 ;
      RECT 45.395 2.626 45.405 3.02 ;
      RECT 45.375 2.601 45.395 2.98 ;
      RECT 45.365 2.57 45.375 2.945 ;
      RECT 45.355 2.557 45.365 2.9 ;
      RECT 45.345 2.542 45.355 2.875 ;
      RECT 45.335 2.355 45.345 2.835 ;
      RECT 45.325 2.355 45.335 2.805 ;
      RECT 45.32 2.355 45.325 2.788 ;
      RECT 45.315 2.355 45.32 2.77 ;
      RECT 45.245 2.355 45.315 2.71 ;
      RECT 45.205 2.355 45.245 2.645 ;
      RECT 45.035 3.225 45.295 3.485 ;
      RECT 43.205 3.145 43.285 3.465 ;
      RECT 43.025 3.205 43.175 3.465 ;
      RECT 43.205 3.145 43.315 3.425 ;
      RECT 45.025 3.317 45.035 3.48 ;
      RECT 44.995 3.327 45.025 3.488 ;
      RECT 44.975 3.335 44.995 3.493 ;
      RECT 44.907 3.343 44.975 3.503 ;
      RECT 44.821 3.363 44.907 3.52 ;
      RECT 44.735 3.384 44.821 3.539 ;
      RECT 44.725 3.4 44.735 3.55 ;
      RECT 44.685 3.41 44.725 3.556 ;
      RECT 44.665 3.415 44.685 3.563 ;
      RECT 44.627 3.416 44.665 3.566 ;
      RECT 44.541 3.419 44.627 3.567 ;
      RECT 44.455 3.423 44.541 3.568 ;
      RECT 44.401 3.425 44.455 3.57 ;
      RECT 44.315 3.425 44.401 3.572 ;
      RECT 44.275 3.42 44.315 3.574 ;
      RECT 44.265 3.414 44.275 3.575 ;
      RECT 44.225 3.409 44.265 3.571 ;
      RECT 44.215 3.4 44.225 3.567 ;
      RECT 44.183 3.391 44.215 3.564 ;
      RECT 44.097 3.379 44.183 3.554 ;
      RECT 44.011 3.362 44.097 3.539 ;
      RECT 43.925 3.344 44.011 3.525 ;
      RECT 43.905 3.335 43.925 3.516 ;
      RECT 43.835 3.325 43.905 3.509 ;
      RECT 43.785 3.31 43.835 3.499 ;
      RECT 43.725 3.3 43.785 3.49 ;
      RECT 43.685 3.29 43.725 3.485 ;
      RECT 43.635 3.28 43.685 3.479 ;
      RECT 43.595 3.268 43.635 3.469 ;
      RECT 43.575 3.258 43.595 3.465 ;
      RECT 43.555 3.248 43.575 3.465 ;
      RECT 43.545 3.238 43.555 3.464 ;
      RECT 43.525 3.23 43.545 3.46 ;
      RECT 43.485 3.205 43.525 3.454 ;
      RECT 43.465 3.145 43.485 3.447 ;
      RECT 43.441 3.145 43.465 3.444 ;
      RECT 43.355 3.145 43.441 3.439 ;
      RECT 43.315 3.145 43.355 3.43 ;
      RECT 43.175 3.195 43.205 3.465 ;
      RECT 44.855 2.775 45.115 3.035 ;
      RECT 44.815 2.775 45.115 2.915 ;
      RECT 44.785 2.775 45.115 2.9 ;
      RECT 44.725 2.775 45.115 2.88 ;
      RECT 44.645 2.585 44.925 2.865 ;
      RECT 44.645 2.77 44.995 2.865 ;
      RECT 44.645 2.71 44.985 2.865 ;
      RECT 44.645 2.66 44.935 2.865 ;
      RECT 42.415 3.115 42.675 3.375 ;
      RECT 42.56 1.205 42.675 3.375 ;
      RECT 42.475 2.585 42.675 3.375 ;
      RECT 43.785 2.635 44.045 2.895 ;
      RECT 42.47 2.585 42.675 2.87 ;
      RECT 42.465 2.585 42.675 2.865 ;
      RECT 43.765 2.645 44.045 2.825 ;
      RECT 43.355 2.615 43.495 2.765 ;
      RECT 42.73 1.205 42.81 1.55 ;
      RECT 42.465 1.205 42.675 1.55 ;
      RECT 43.755 2.644 43.765 2.825 ;
      RECT 43.751 2.644 43.755 2.825 ;
      RECT 43.665 2.639 43.751 2.814 ;
      RECT 43.591 2.63 43.665 2.794 ;
      RECT 43.505 2.621 43.591 2.775 ;
      RECT 43.495 2.615 43.505 2.765 ;
      RECT 43.315 2.615 43.355 2.768 ;
      RECT 43.229 2.615 43.315 2.776 ;
      RECT 43.143 2.615 43.229 2.787 ;
      RECT 43.057 2.615 43.143 2.798 ;
      RECT 42.971 2.615 43.057 2.809 ;
      RECT 42.885 2.615 42.971 2.82 ;
      RECT 42.855 2.615 42.885 2.86 ;
      RECT 42.825 2.615 42.855 2.91 ;
      RECT 42.75 2.615 42.825 2.93 ;
      RECT 42.745 2.59 42.75 2.935 ;
      RECT 42.73 2.585 42.745 2.943 ;
      RECT 42.725 1.205 42.73 2.953 ;
      RECT 42.695 1.205 42.725 2.995 ;
      RECT 42.675 1.205 42.695 3.075 ;
      RECT 41.805 2.965 41.825 3.404 ;
      RECT 41.805 2.965 41.911 3.401 ;
      RECT 41.795 3.08 41.911 3.4 ;
      RECT 41.825 2.115 41.955 3.397 ;
      RECT 41.805 2.985 41.965 3.395 ;
      RECT 41.805 3.07 41.975 3.39 ;
      RECT 41.775 3.115 41.975 3.385 ;
      RECT 41.775 3.115 41.985 3.38 ;
      RECT 41.755 3.115 42.015 3.375 ;
      RECT 41.825 2.115 41.985 2.765 ;
      RECT 41.815 2.115 41.985 2.74 ;
      RECT 41.815 2.115 42.005 2.505 ;
      RECT 41.765 2.115 42.025 2.375 ;
      RECT 41.235 2.605 41.525 2.865 ;
      RECT 41.245 2.585 41.525 2.865 ;
      RECT 41.195 2.665 41.525 2.86 ;
      RECT 41.265 2.578 41.435 2.865 ;
      RECT 41.265 2.565 41.391 2.865 ;
      RECT 41.305 2.558 41.391 2.865 ;
      RECT 40.765 3.705 41.045 3.985 ;
      RECT 40.725 3.67 41.025 3.78 ;
      RECT 40.715 3.62 41.005 3.675 ;
      RECT 40.655 3.385 40.915 3.645 ;
      RECT 40.655 3.525 40.995 3.645 ;
      RECT 40.655 3.475 40.975 3.645 ;
      RECT 40.655 3.43 40.965 3.645 ;
      RECT 40.655 3.415 40.935 3.645 ;
      RECT 36.39 6.225 36.71 6.545 ;
      RECT 36.42 5.695 36.59 6.545 ;
      RECT 36.42 5.695 36.595 6.045 ;
      RECT 36.42 5.695 37.395 5.87 ;
      RECT 37.22 1.965 37.395 5.87 ;
      RECT 37.165 1.965 37.515 2.315 ;
      RECT 37.19 6.655 37.515 6.98 ;
      RECT 36.075 6.745 37.515 6.915 ;
      RECT 36.075 2.395 36.235 6.915 ;
      RECT 36.39 2.365 36.71 2.685 ;
      RECT 36.075 2.395 36.71 2.565 ;
      RECT 34.745 1.14 35.12 1.51 ;
      RECT 26.665 0.96 27.04 1.33 ;
      RECT 25.23 0.96 25.605 1.33 ;
      RECT 25.23 1.08 35.05 1.25 ;
      RECT 31.175 4.36 35.03 4.53 ;
      RECT 34.86 3.425 35.03 4.53 ;
      RECT 31.175 3.665 31.345 4.53 ;
      RECT 31.12 3.705 31.4 3.985 ;
      RECT 31.14 3.665 31.4 3.985 ;
      RECT 30.78 3.625 30.89 3.885 ;
      RECT 34.77 3.43 35.12 3.78 ;
      RECT 30.64 2.115 30.73 2.375 ;
      RECT 31.17 3.17 31.18 3.3 ;
      RECT 31.16 3.135 31.17 3.454 ;
      RECT 31.08 3.067 31.16 3.534 ;
      RECT 31.11 3.71 31.12 3.93 ;
      RECT 31.09 3.705 31.11 3.919 ;
      RECT 31.06 3.7 31.09 3.904 ;
      RECT 31.07 3.002 31.08 3.61 ;
      RECT 31.05 2.946 31.07 3.625 ;
      RECT 31.04 3.685 31.06 3.89 ;
      RECT 31.04 2.874 31.05 3.645 ;
      RECT 31.01 2.777 31.04 3.885 ;
      RECT 30.99 2.66 31.01 3.885 ;
      RECT 30.96 2.54 30.99 3.885 ;
      RECT 30.95 2.455 30.96 3.885 ;
      RECT 30.94 2.4 30.95 3.885 ;
      RECT 30.93 2.355 30.94 3.104 ;
      RECT 30.92 3.315 30.94 3.885 ;
      RECT 30.92 2.285 30.93 3.061 ;
      RECT 30.9 2.235 30.92 2.996 ;
      RECT 30.91 3.395 30.92 3.885 ;
      RECT 30.89 3.495 30.91 3.885 ;
      RECT 30.84 2.115 30.9 2.824 ;
      RECT 30.83 2.115 30.84 2.66 ;
      RECT 30.82 2.115 30.83 2.61 ;
      RECT 30.77 2.115 30.82 2.54 ;
      RECT 30.75 2.115 30.77 2.455 ;
      RECT 30.73 2.115 30.75 2.41 ;
      RECT 33.12 2.155 33.38 2.415 ;
      RECT 33.11 2.155 33.38 2.365 ;
      RECT 33.08 2.025 33.36 2.305 ;
      RECT 21.645 6.655 21.995 7.005 ;
      RECT 32.615 6.61 32.965 6.96 ;
      RECT 21.645 6.685 32.965 6.885 ;
      RECT 32.12 3.705 32.4 3.985 ;
      RECT 32.16 3.665 32.43 3.925 ;
      RECT 32.15 3.7 32.43 3.925 ;
      RECT 32.16 3.66 32.37 3.985 ;
      RECT 32.16 3.655 32.36 3.985 ;
      RECT 32.2 3.645 32.36 3.985 ;
      RECT 32.17 3.65 32.36 3.985 ;
      RECT 32.21 3.64 32.3 3.985 ;
      RECT 32.23 3.635 32.3 3.985 ;
      RECT 31.54 3.155 31.8 3.415 ;
      RECT 31.59 3.065 31.78 3.415 ;
      RECT 31.62 2.85 31.78 3.415 ;
      RECT 31.71 2.455 31.78 3.415 ;
      RECT 31.73 2.165 31.866 2.893 ;
      RECT 31.67 2.66 31.866 2.893 ;
      RECT 31.69 2.54 31.78 3.415 ;
      RECT 31.73 2.165 31.89 2.558 ;
      RECT 31.73 2.165 31.9 2.455 ;
      RECT 31.72 2.165 31.98 2.425 ;
      RECT 30.05 3.565 30.1 3.825 ;
      RECT 29.96 2.095 30.1 2.355 ;
      RECT 30.46 2.72 30.47 2.808 ;
      RECT 30.45 2.655 30.46 2.854 ;
      RECT 30.44 2.605 30.45 2.9 ;
      RECT 30.39 2.552 30.44 3.039 ;
      RECT 30.38 2.501 30.39 3.23 ;
      RECT 30.34 2.459 30.38 3.335 ;
      RECT 30.32 2.405 30.34 3.472 ;
      RECT 30.31 2.38 30.32 2.688 ;
      RECT 30.31 2.77 30.32 3.542 ;
      RECT 30.3 2.366 30.31 2.673 ;
      RECT 30.3 2.825 30.31 3.825 ;
      RECT 30.28 2.341 30.3 2.655 ;
      RECT 30.26 3 30.3 3.825 ;
      RECT 30.27 2.315 30.28 2.635 ;
      RECT 30.24 2.28 30.27 2.589 ;
      RECT 30.25 3.125 30.26 3.825 ;
      RECT 30.24 3.205 30.25 3.825 ;
      RECT 30.23 2.245 30.24 2.554 ;
      RECT 30.19 3.275 30.24 3.825 ;
      RECT 30.22 2.225 30.23 2.53 ;
      RECT 30.19 2.095 30.22 2.495 ;
      RECT 30.18 2.095 30.19 2.46 ;
      RECT 30.16 3.375 30.19 3.825 ;
      RECT 30.16 2.095 30.18 2.435 ;
      RECT 30.15 2.095 30.16 2.41 ;
      RECT 30.11 3.475 30.16 3.825 ;
      RECT 30.13 2.095 30.15 2.38 ;
      RECT 30.1 2.095 30.13 2.365 ;
      RECT 30.1 3.55 30.11 3.825 ;
      RECT 30.02 2.635 30.06 2.895 ;
      RECT 25.75 2.055 26.01 2.315 ;
      RECT 25.75 2.085 26.03 2.295 ;
      RECT 27.96 1.905 28.14 2.055 ;
      RECT 30.01 2.63 30.02 2.895 ;
      RECT 29.99 2.62 30.01 2.895 ;
      RECT 29.972 2.613 29.99 2.895 ;
      RECT 29.886 2.602 29.972 2.895 ;
      RECT 29.8 2.585 29.886 2.895 ;
      RECT 29.75 2.572 29.8 2.82 ;
      RECT 29.716 2.564 29.75 2.795 ;
      RECT 29.63 2.553 29.716 2.76 ;
      RECT 29.59 2.53 29.63 2.723 ;
      RECT 29.58 2.495 29.59 2.708 ;
      RECT 29.57 2.455 29.58 2.703 ;
      RECT 29.56 2.435 29.57 2.698 ;
      RECT 29.545 2.395 29.56 2.693 ;
      RECT 29.53 2.347 29.545 2.689 ;
      RECT 29.52 2.306 29.53 2.686 ;
      RECT 29.51 2.268 29.52 2.675 ;
      RECT 29.49 2.212 29.51 2.655 ;
      RECT 29.47 2.16 29.49 2.591 ;
      RECT 29.45 2.11 29.47 2.543 ;
      RECT 29.44 2.08 29.45 2.507 ;
      RECT 29.435 2.062 29.44 2.493 ;
      RECT 29.42 2.053 29.435 2.475 ;
      RECT 29.39 2.034 29.42 2.415 ;
      RECT 29.38 2.017 29.39 2.37 ;
      RECT 29.37 2.009 29.38 2.34 ;
      RECT 29.34 1.997 29.37 2.29 ;
      RECT 29.32 1.985 29.34 2.225 ;
      RECT 29.31 1.977 29.32 2.185 ;
      RECT 29.29 1.974 29.31 2.175 ;
      RECT 29.275 1.972 29.29 2.17 ;
      RECT 29.255 1.971 29.275 2.16 ;
      RECT 29.24 1.97 29.255 2.15 ;
      RECT 29.22 1.969 29.24 2.145 ;
      RECT 29.218 1.969 29.22 2.145 ;
      RECT 29.132 1.966 29.218 2.142 ;
      RECT 29.046 1.961 29.132 2.135 ;
      RECT 28.96 1.956 29.046 2.129 ;
      RECT 28.91 1.953 28.96 2.12 ;
      RECT 28.866 1.951 28.91 2.114 ;
      RECT 28.78 1.947 28.866 2.109 ;
      RECT 28.776 1.945 28.78 2.105 ;
      RECT 28.69 1.942 28.776 2.1 ;
      RECT 28.636 1.938 28.69 2.093 ;
      RECT 28.55 1.935 28.636 2.088 ;
      RECT 28.526 1.932 28.55 2.084 ;
      RECT 28.44 1.93 28.526 2.079 ;
      RECT 28.38 1.926 28.44 2.073 ;
      RECT 28.372 1.924 28.38 2.07 ;
      RECT 28.286 1.92 28.372 2.066 ;
      RECT 28.2 1.913 28.286 2.059 ;
      RECT 28.14 1.907 28.2 2.055 ;
      RECT 27.94 1.905 27.96 2.058 ;
      RECT 27.89 1.915 27.94 2.068 ;
      RECT 27.86 1.925 27.89 2.08 ;
      RECT 27.836 1.927 27.86 2.086 ;
      RECT 27.75 1.93 27.836 2.091 ;
      RECT 27.68 1.935 27.75 2.1 ;
      RECT 27.666 1.937 27.68 2.106 ;
      RECT 27.58 1.941 27.666 2.111 ;
      RECT 27.54 1.945 27.58 2.12 ;
      RECT 27.526 1.947 27.54 2.126 ;
      RECT 27.44 1.951 27.526 2.131 ;
      RECT 27.356 1.957 27.44 2.138 ;
      RECT 27.27 1.963 27.356 2.143 ;
      RECT 27.246 1.967 27.27 2.146 ;
      RECT 27.16 1.971 27.246 2.151 ;
      RECT 27.11 1.976 27.16 2.16 ;
      RECT 27.03 1.981 27.11 2.17 ;
      RECT 26.95 1.987 27.03 2.185 ;
      RECT 26.93 1.991 26.95 2.195 ;
      RECT 26.86 1.994 26.93 2.205 ;
      RECT 26.81 1.999 26.86 2.22 ;
      RECT 26.78 2.002 26.81 2.24 ;
      RECT 26.77 2.004 26.78 2.256 ;
      RECT 26.71 2.016 26.77 2.266 ;
      RECT 26.69 2.031 26.71 2.275 ;
      RECT 26.68 2.05 26.69 2.275 ;
      RECT 26.67 2.07 26.68 2.275 ;
      RECT 26.65 2.08 26.67 2.275 ;
      RECT 26.6 2.09 26.65 2.275 ;
      RECT 26.57 2.096 26.6 2.275 ;
      RECT 26.5 2.101 26.57 2.277 ;
      RECT 26.42 2.102 26.5 2.282 ;
      RECT 26.416 2.1 26.42 2.285 ;
      RECT 26.33 2.097 26.416 2.286 ;
      RECT 26.288 2.094 26.33 2.288 ;
      RECT 26.202 2.092 26.288 2.289 ;
      RECT 26.116 2.089 26.202 2.292 ;
      RECT 26.03 2.086 26.116 2.294 ;
      RECT 29.41 3.705 29.44 3.985 ;
      RECT 29.16 3.595 29.18 3.985 ;
      RECT 29.12 3.595 29.18 3.855 ;
      RECT 28.95 2.225 28.98 2.485 ;
      RECT 28.72 2.225 28.78 2.485 ;
      RECT 29.4 3.685 29.41 3.985 ;
      RECT 29.38 3.605 29.4 3.985 ;
      RECT 29.37 3.545 29.38 3.985 ;
      RECT 29.32 3.435 29.37 3.985 ;
      RECT 29.31 3.305 29.32 3.985 ;
      RECT 29.27 3.245 29.31 3.985 ;
      RECT 29.266 3.214 29.27 3.985 ;
      RECT 29.18 3.205 29.266 3.985 ;
      RECT 29.17 3.196 29.18 3.55 ;
      RECT 29.14 3.175 29.17 3.517 ;
      RECT 29.13 3.125 29.14 3.493 ;
      RECT 29.12 3.09 29.13 3.481 ;
      RECT 29.08 3.015 29.12 3.45 ;
      RECT 29.06 2.925 29.08 3.415 ;
      RECT 29.05 2.866 29.06 3.4 ;
      RECT 29 2.756 29.05 3.36 ;
      RECT 28.99 2.65 29 3.315 ;
      RECT 28.96 2.579 28.99 3.235 ;
      RECT 28.95 2.511 28.96 3.16 ;
      RECT 28.94 2.225 28.95 3.125 ;
      RECT 28.91 2.225 28.94 3.055 ;
      RECT 28.9 2.225 28.91 2.95 ;
      RECT 28.89 2.225 28.9 2.915 ;
      RECT 28.82 2.225 28.89 2.775 ;
      RECT 28.79 2.225 28.82 2.575 ;
      RECT 28.78 2.225 28.79 2.5 ;
      RECT 27.96 3.145 28.24 3.425 ;
      RECT 27.99 3.125 28.26 3.385 ;
      RECT 27.99 3.075 28.22 3.425 ;
      RECT 28.06 3.065 28.22 3.425 ;
      RECT 28.06 2.775 28.21 3.425 ;
      RECT 28.05 2.455 28.2 2.825 ;
      RECT 28.04 2.455 28.2 2.695 ;
      RECT 28.02 2.165 28.19 2.5 ;
      RECT 28 2.165 28.19 2.45 ;
      RECT 27.96 2.165 28.22 2.425 ;
      RECT 27.87 3.635 27.95 3.895 ;
      RECT 27.16 2.355 27.28 2.615 ;
      RECT 27.845 3.615 27.87 3.895 ;
      RECT 27.83 3.577 27.845 3.895 ;
      RECT 27.79 3.52 27.83 3.895 ;
      RECT 27.76 3.43 27.79 3.895 ;
      RECT 27.72 3.33 27.76 3.895 ;
      RECT 27.69 3.23 27.72 3.895 ;
      RECT 27.685 3.177 27.69 3.718 ;
      RECT 27.67 3.147 27.685 3.684 ;
      RECT 27.66 3.108 27.67 3.649 ;
      RECT 27.65 3.075 27.66 3.605 ;
      RECT 27.64 3.042 27.65 3.57 ;
      RECT 27.61 2.976 27.64 3.505 ;
      RECT 27.6 2.911 27.61 3.43 ;
      RECT 27.59 2.881 27.6 3.4 ;
      RECT 27.55 2.811 27.59 3.33 ;
      RECT 27.54 2.746 27.55 3.245 ;
      RECT 27.53 2.728 27.54 3.23 ;
      RECT 27.52 2.711 27.53 3.195 ;
      RECT 27.51 2.694 27.52 3.165 ;
      RECT 27.5 2.677 27.51 3.135 ;
      RECT 27.48 2.652 27.5 3.075 ;
      RECT 27.47 2.626 27.48 3.02 ;
      RECT 27.45 2.601 27.47 2.98 ;
      RECT 27.44 2.57 27.45 2.945 ;
      RECT 27.43 2.557 27.44 2.9 ;
      RECT 27.42 2.542 27.43 2.875 ;
      RECT 27.41 2.355 27.42 2.835 ;
      RECT 27.4 2.355 27.41 2.805 ;
      RECT 27.395 2.355 27.4 2.788 ;
      RECT 27.39 2.355 27.395 2.77 ;
      RECT 27.32 2.355 27.39 2.71 ;
      RECT 27.28 2.355 27.32 2.645 ;
      RECT 27.11 3.225 27.37 3.485 ;
      RECT 25.28 3.145 25.36 3.465 ;
      RECT 25.1 3.205 25.25 3.465 ;
      RECT 25.28 3.145 25.39 3.425 ;
      RECT 27.1 3.317 27.11 3.48 ;
      RECT 27.07 3.327 27.1 3.488 ;
      RECT 27.05 3.335 27.07 3.493 ;
      RECT 26.982 3.343 27.05 3.503 ;
      RECT 26.896 3.363 26.982 3.52 ;
      RECT 26.81 3.384 26.896 3.539 ;
      RECT 26.8 3.4 26.81 3.55 ;
      RECT 26.76 3.41 26.8 3.556 ;
      RECT 26.74 3.415 26.76 3.563 ;
      RECT 26.702 3.416 26.74 3.566 ;
      RECT 26.616 3.419 26.702 3.567 ;
      RECT 26.53 3.423 26.616 3.568 ;
      RECT 26.476 3.425 26.53 3.57 ;
      RECT 26.39 3.425 26.476 3.572 ;
      RECT 26.35 3.42 26.39 3.574 ;
      RECT 26.34 3.414 26.35 3.575 ;
      RECT 26.3 3.409 26.34 3.571 ;
      RECT 26.29 3.4 26.3 3.567 ;
      RECT 26.258 3.391 26.29 3.564 ;
      RECT 26.172 3.379 26.258 3.554 ;
      RECT 26.086 3.362 26.172 3.539 ;
      RECT 26 3.344 26.086 3.525 ;
      RECT 25.98 3.335 26 3.516 ;
      RECT 25.91 3.325 25.98 3.509 ;
      RECT 25.86 3.31 25.91 3.499 ;
      RECT 25.8 3.3 25.86 3.49 ;
      RECT 25.76 3.29 25.8 3.485 ;
      RECT 25.71 3.28 25.76 3.479 ;
      RECT 25.67 3.268 25.71 3.469 ;
      RECT 25.65 3.258 25.67 3.465 ;
      RECT 25.63 3.248 25.65 3.465 ;
      RECT 25.62 3.238 25.63 3.464 ;
      RECT 25.6 3.23 25.62 3.46 ;
      RECT 25.56 3.205 25.6 3.454 ;
      RECT 25.54 3.145 25.56 3.447 ;
      RECT 25.516 3.145 25.54 3.444 ;
      RECT 25.43 3.145 25.516 3.439 ;
      RECT 25.39 3.145 25.43 3.43 ;
      RECT 25.25 3.195 25.28 3.465 ;
      RECT 26.93 2.775 27.19 3.035 ;
      RECT 26.89 2.775 27.19 2.915 ;
      RECT 26.86 2.775 27.19 2.9 ;
      RECT 26.8 2.775 27.19 2.88 ;
      RECT 26.72 2.585 27 2.865 ;
      RECT 26.72 2.77 27.07 2.865 ;
      RECT 26.72 2.71 27.06 2.865 ;
      RECT 26.72 2.66 27.01 2.865 ;
      RECT 24.49 3.115 24.75 3.375 ;
      RECT 24.635 1.205 24.75 3.375 ;
      RECT 24.55 2.585 24.75 3.375 ;
      RECT 25.86 2.635 26.12 2.895 ;
      RECT 24.545 2.585 24.75 2.87 ;
      RECT 24.54 2.585 24.75 2.865 ;
      RECT 25.84 2.645 26.12 2.825 ;
      RECT 25.43 2.615 25.57 2.765 ;
      RECT 24.805 1.205 24.885 1.55 ;
      RECT 24.54 1.205 24.75 1.55 ;
      RECT 25.83 2.644 25.84 2.825 ;
      RECT 25.826 2.644 25.83 2.825 ;
      RECT 25.74 2.639 25.826 2.814 ;
      RECT 25.666 2.63 25.74 2.794 ;
      RECT 25.58 2.621 25.666 2.775 ;
      RECT 25.57 2.615 25.58 2.765 ;
      RECT 25.39 2.615 25.43 2.768 ;
      RECT 25.304 2.615 25.39 2.776 ;
      RECT 25.218 2.615 25.304 2.787 ;
      RECT 25.132 2.615 25.218 2.798 ;
      RECT 25.046 2.615 25.132 2.809 ;
      RECT 24.96 2.615 25.046 2.82 ;
      RECT 24.93 2.615 24.96 2.86 ;
      RECT 24.9 2.615 24.93 2.91 ;
      RECT 24.825 2.615 24.9 2.93 ;
      RECT 24.82 2.59 24.825 2.935 ;
      RECT 24.805 2.585 24.82 2.943 ;
      RECT 24.8 1.205 24.805 2.953 ;
      RECT 24.77 1.205 24.8 2.995 ;
      RECT 24.75 1.205 24.77 3.075 ;
      RECT 23.88 2.965 23.9 3.404 ;
      RECT 23.88 2.965 23.986 3.401 ;
      RECT 23.87 3.08 23.986 3.4 ;
      RECT 23.9 2.115 24.03 3.397 ;
      RECT 23.88 2.985 24.04 3.395 ;
      RECT 23.88 3.07 24.05 3.39 ;
      RECT 23.85 3.115 24.05 3.385 ;
      RECT 23.85 3.115 24.06 3.38 ;
      RECT 23.83 3.115 24.09 3.375 ;
      RECT 23.9 2.115 24.06 2.765 ;
      RECT 23.89 2.115 24.06 2.74 ;
      RECT 23.89 2.115 24.08 2.505 ;
      RECT 23.84 2.115 24.1 2.375 ;
      RECT 23.31 2.605 23.6 2.865 ;
      RECT 23.32 2.585 23.6 2.865 ;
      RECT 23.27 2.665 23.6 2.86 ;
      RECT 23.34 2.578 23.51 2.865 ;
      RECT 23.34 2.565 23.466 2.865 ;
      RECT 23.38 2.558 23.466 2.865 ;
      RECT 22.84 3.705 23.12 3.985 ;
      RECT 22.8 3.67 23.1 3.78 ;
      RECT 22.79 3.62 23.08 3.675 ;
      RECT 22.73 3.385 22.99 3.645 ;
      RECT 22.73 3.525 23.07 3.645 ;
      RECT 22.73 3.475 23.05 3.645 ;
      RECT 22.73 3.43 23.04 3.645 ;
      RECT 22.73 3.415 23.01 3.645 ;
      RECT 18.465 6.225 18.785 6.545 ;
      RECT 18.495 5.695 18.665 6.545 ;
      RECT 18.495 5.695 18.67 6.045 ;
      RECT 18.495 5.695 19.47 5.87 ;
      RECT 19.295 1.965 19.47 5.87 ;
      RECT 19.24 1.965 19.59 2.315 ;
      RECT 19.265 6.655 19.59 6.98 ;
      RECT 18.15 6.745 19.59 6.915 ;
      RECT 18.15 2.395 18.31 6.915 ;
      RECT 18.465 2.365 18.785 2.685 ;
      RECT 18.15 2.395 18.785 2.565 ;
      RECT 16.82 1.14 17.195 1.51 ;
      RECT 8.74 0.96 9.115 1.33 ;
      RECT 7.305 0.96 7.68 1.33 ;
      RECT 7.305 1.08 17.125 1.25 ;
      RECT 13.25 4.36 17.105 4.53 ;
      RECT 16.935 3.425 17.105 4.53 ;
      RECT 13.25 3.665 13.42 4.53 ;
      RECT 13.195 3.705 13.475 3.985 ;
      RECT 13.215 3.665 13.475 3.985 ;
      RECT 12.855 3.625 12.965 3.885 ;
      RECT 16.845 3.43 17.195 3.78 ;
      RECT 12.715 2.115 12.805 2.375 ;
      RECT 13.245 3.17 13.255 3.3 ;
      RECT 13.235 3.135 13.245 3.454 ;
      RECT 13.155 3.067 13.235 3.534 ;
      RECT 13.185 3.71 13.195 3.93 ;
      RECT 13.165 3.705 13.185 3.919 ;
      RECT 13.135 3.7 13.165 3.904 ;
      RECT 13.145 3.002 13.155 3.61 ;
      RECT 13.125 2.946 13.145 3.625 ;
      RECT 13.115 3.685 13.135 3.89 ;
      RECT 13.115 2.874 13.125 3.645 ;
      RECT 13.085 2.777 13.115 3.885 ;
      RECT 13.065 2.66 13.085 3.885 ;
      RECT 13.035 2.54 13.065 3.885 ;
      RECT 13.025 2.455 13.035 3.885 ;
      RECT 13.015 2.4 13.025 3.885 ;
      RECT 13.005 2.355 13.015 3.104 ;
      RECT 12.995 3.315 13.015 3.885 ;
      RECT 12.995 2.285 13.005 3.061 ;
      RECT 12.975 2.235 12.995 2.996 ;
      RECT 12.985 3.395 12.995 3.885 ;
      RECT 12.965 3.495 12.985 3.885 ;
      RECT 12.915 2.115 12.975 2.824 ;
      RECT 12.905 2.115 12.915 2.66 ;
      RECT 12.895 2.115 12.905 2.61 ;
      RECT 12.845 2.115 12.895 2.54 ;
      RECT 12.825 2.115 12.845 2.455 ;
      RECT 12.805 2.115 12.825 2.41 ;
      RECT 15.195 2.155 15.455 2.415 ;
      RECT 15.185 2.155 15.455 2.365 ;
      RECT 15.155 2.025 15.435 2.305 ;
      RECT 3.02 6.995 3.31 7.345 ;
      RECT 3.02 7.055 4.155 7.225 ;
      RECT 3.985 6.685 4.155 7.225 ;
      RECT 14.71 6.605 14.88 6.96 ;
      RECT 14.66 6.605 15.01 6.955 ;
      RECT 3.985 6.685 15.01 6.855 ;
      RECT 14.195 3.705 14.475 3.985 ;
      RECT 14.235 3.665 14.505 3.925 ;
      RECT 14.225 3.7 14.505 3.925 ;
      RECT 14.235 3.66 14.445 3.985 ;
      RECT 14.235 3.655 14.435 3.985 ;
      RECT 14.275 3.645 14.435 3.985 ;
      RECT 14.245 3.65 14.435 3.985 ;
      RECT 14.285 3.64 14.375 3.985 ;
      RECT 14.305 3.635 14.375 3.985 ;
      RECT 13.615 3.155 13.875 3.415 ;
      RECT 13.665 3.065 13.855 3.415 ;
      RECT 13.695 2.85 13.855 3.415 ;
      RECT 13.785 2.455 13.855 3.415 ;
      RECT 13.805 2.165 13.941 2.893 ;
      RECT 13.745 2.66 13.941 2.893 ;
      RECT 13.765 2.54 13.855 3.415 ;
      RECT 13.805 2.165 13.965 2.558 ;
      RECT 13.805 2.165 13.975 2.455 ;
      RECT 13.795 2.165 14.055 2.425 ;
      RECT 12.125 3.565 12.175 3.825 ;
      RECT 12.035 2.095 12.175 2.355 ;
      RECT 12.535 2.72 12.545 2.808 ;
      RECT 12.525 2.655 12.535 2.854 ;
      RECT 12.515 2.605 12.525 2.9 ;
      RECT 12.465 2.552 12.515 3.039 ;
      RECT 12.455 2.501 12.465 3.23 ;
      RECT 12.415 2.459 12.455 3.335 ;
      RECT 12.395 2.405 12.415 3.472 ;
      RECT 12.385 2.38 12.395 2.688 ;
      RECT 12.385 2.77 12.395 3.542 ;
      RECT 12.375 2.366 12.385 2.673 ;
      RECT 12.375 2.825 12.385 3.825 ;
      RECT 12.355 2.341 12.375 2.655 ;
      RECT 12.335 3 12.375 3.825 ;
      RECT 12.345 2.315 12.355 2.635 ;
      RECT 12.315 2.28 12.345 2.589 ;
      RECT 12.325 3.125 12.335 3.825 ;
      RECT 12.315 3.205 12.325 3.825 ;
      RECT 12.305 2.245 12.315 2.554 ;
      RECT 12.265 3.275 12.315 3.825 ;
      RECT 12.295 2.225 12.305 2.53 ;
      RECT 12.265 2.095 12.295 2.495 ;
      RECT 12.255 2.095 12.265 2.46 ;
      RECT 12.235 3.375 12.265 3.825 ;
      RECT 12.235 2.095 12.255 2.435 ;
      RECT 12.225 2.095 12.235 2.41 ;
      RECT 12.185 3.475 12.235 3.825 ;
      RECT 12.205 2.095 12.225 2.38 ;
      RECT 12.175 2.095 12.205 2.365 ;
      RECT 12.175 3.55 12.185 3.825 ;
      RECT 12.095 2.635 12.135 2.895 ;
      RECT 7.825 2.055 8.085 2.315 ;
      RECT 7.825 2.085 8.105 2.295 ;
      RECT 10.035 1.905 10.215 2.055 ;
      RECT 12.085 2.63 12.095 2.895 ;
      RECT 12.065 2.62 12.085 2.895 ;
      RECT 12.047 2.613 12.065 2.895 ;
      RECT 11.961 2.602 12.047 2.895 ;
      RECT 11.875 2.585 11.961 2.895 ;
      RECT 11.825 2.572 11.875 2.82 ;
      RECT 11.791 2.564 11.825 2.795 ;
      RECT 11.705 2.553 11.791 2.76 ;
      RECT 11.665 2.53 11.705 2.723 ;
      RECT 11.655 2.495 11.665 2.708 ;
      RECT 11.645 2.455 11.655 2.703 ;
      RECT 11.635 2.435 11.645 2.698 ;
      RECT 11.62 2.395 11.635 2.693 ;
      RECT 11.605 2.347 11.62 2.689 ;
      RECT 11.595 2.306 11.605 2.686 ;
      RECT 11.585 2.268 11.595 2.675 ;
      RECT 11.565 2.212 11.585 2.655 ;
      RECT 11.545 2.16 11.565 2.591 ;
      RECT 11.525 2.11 11.545 2.543 ;
      RECT 11.515 2.08 11.525 2.507 ;
      RECT 11.51 2.062 11.515 2.493 ;
      RECT 11.495 2.053 11.51 2.475 ;
      RECT 11.465 2.034 11.495 2.415 ;
      RECT 11.455 2.017 11.465 2.37 ;
      RECT 11.445 2.009 11.455 2.34 ;
      RECT 11.415 1.997 11.445 2.29 ;
      RECT 11.395 1.985 11.415 2.225 ;
      RECT 11.385 1.977 11.395 2.185 ;
      RECT 11.365 1.974 11.385 2.175 ;
      RECT 11.35 1.972 11.365 2.17 ;
      RECT 11.33 1.971 11.35 2.16 ;
      RECT 11.315 1.97 11.33 2.15 ;
      RECT 11.295 1.969 11.315 2.145 ;
      RECT 11.293 1.969 11.295 2.145 ;
      RECT 11.207 1.966 11.293 2.142 ;
      RECT 11.121 1.961 11.207 2.135 ;
      RECT 11.035 1.956 11.121 2.129 ;
      RECT 10.985 1.953 11.035 2.12 ;
      RECT 10.941 1.951 10.985 2.114 ;
      RECT 10.855 1.947 10.941 2.109 ;
      RECT 10.851 1.945 10.855 2.105 ;
      RECT 10.765 1.942 10.851 2.1 ;
      RECT 10.711 1.938 10.765 2.093 ;
      RECT 10.625 1.935 10.711 2.088 ;
      RECT 10.601 1.932 10.625 2.084 ;
      RECT 10.515 1.93 10.601 2.079 ;
      RECT 10.455 1.926 10.515 2.073 ;
      RECT 10.447 1.924 10.455 2.07 ;
      RECT 10.361 1.92 10.447 2.066 ;
      RECT 10.275 1.913 10.361 2.059 ;
      RECT 10.215 1.907 10.275 2.055 ;
      RECT 10.015 1.905 10.035 2.058 ;
      RECT 9.965 1.915 10.015 2.068 ;
      RECT 9.935 1.925 9.965 2.08 ;
      RECT 9.911 1.927 9.935 2.086 ;
      RECT 9.825 1.93 9.911 2.091 ;
      RECT 9.755 1.935 9.825 2.1 ;
      RECT 9.741 1.937 9.755 2.106 ;
      RECT 9.655 1.941 9.741 2.111 ;
      RECT 9.615 1.945 9.655 2.12 ;
      RECT 9.601 1.947 9.615 2.126 ;
      RECT 9.515 1.951 9.601 2.131 ;
      RECT 9.431 1.957 9.515 2.138 ;
      RECT 9.345 1.963 9.431 2.143 ;
      RECT 9.321 1.967 9.345 2.146 ;
      RECT 9.235 1.971 9.321 2.151 ;
      RECT 9.185 1.976 9.235 2.16 ;
      RECT 9.105 1.981 9.185 2.17 ;
      RECT 9.025 1.987 9.105 2.185 ;
      RECT 9.005 1.991 9.025 2.195 ;
      RECT 8.935 1.994 9.005 2.205 ;
      RECT 8.885 1.999 8.935 2.22 ;
      RECT 8.855 2.002 8.885 2.24 ;
      RECT 8.845 2.004 8.855 2.256 ;
      RECT 8.785 2.016 8.845 2.266 ;
      RECT 8.765 2.031 8.785 2.275 ;
      RECT 8.755 2.05 8.765 2.275 ;
      RECT 8.745 2.07 8.755 2.275 ;
      RECT 8.725 2.08 8.745 2.275 ;
      RECT 8.675 2.09 8.725 2.275 ;
      RECT 8.645 2.096 8.675 2.275 ;
      RECT 8.575 2.101 8.645 2.277 ;
      RECT 8.495 2.102 8.575 2.282 ;
      RECT 8.491 2.1 8.495 2.285 ;
      RECT 8.405 2.097 8.491 2.286 ;
      RECT 8.363 2.094 8.405 2.288 ;
      RECT 8.277 2.092 8.363 2.289 ;
      RECT 8.191 2.089 8.277 2.292 ;
      RECT 8.105 2.086 8.191 2.294 ;
      RECT 11.485 3.705 11.515 3.985 ;
      RECT 11.235 3.595 11.255 3.985 ;
      RECT 11.195 3.595 11.255 3.855 ;
      RECT 11.025 2.225 11.055 2.485 ;
      RECT 10.795 2.225 10.855 2.485 ;
      RECT 11.475 3.685 11.485 3.985 ;
      RECT 11.455 3.605 11.475 3.985 ;
      RECT 11.445 3.545 11.455 3.985 ;
      RECT 11.395 3.435 11.445 3.985 ;
      RECT 11.385 3.305 11.395 3.985 ;
      RECT 11.345 3.245 11.385 3.985 ;
      RECT 11.341 3.214 11.345 3.985 ;
      RECT 11.255 3.205 11.341 3.985 ;
      RECT 11.245 3.196 11.255 3.55 ;
      RECT 11.215 3.175 11.245 3.517 ;
      RECT 11.205 3.125 11.215 3.493 ;
      RECT 11.195 3.09 11.205 3.481 ;
      RECT 11.155 3.015 11.195 3.45 ;
      RECT 11.135 2.925 11.155 3.415 ;
      RECT 11.125 2.866 11.135 3.4 ;
      RECT 11.075 2.756 11.125 3.36 ;
      RECT 11.065 2.65 11.075 3.315 ;
      RECT 11.035 2.579 11.065 3.235 ;
      RECT 11.025 2.511 11.035 3.16 ;
      RECT 11.015 2.225 11.025 3.125 ;
      RECT 10.985 2.225 11.015 3.055 ;
      RECT 10.975 2.225 10.985 2.95 ;
      RECT 10.965 2.225 10.975 2.915 ;
      RECT 10.895 2.225 10.965 2.775 ;
      RECT 10.865 2.225 10.895 2.575 ;
      RECT 10.855 2.225 10.865 2.5 ;
      RECT 10.035 3.145 10.315 3.425 ;
      RECT 10.065 3.125 10.335 3.385 ;
      RECT 10.065 3.075 10.295 3.425 ;
      RECT 10.135 3.065 10.295 3.425 ;
      RECT 10.135 2.775 10.285 3.425 ;
      RECT 10.125 2.455 10.275 2.825 ;
      RECT 10.115 2.455 10.275 2.695 ;
      RECT 10.095 2.165 10.265 2.5 ;
      RECT 10.075 2.165 10.265 2.45 ;
      RECT 10.035 2.165 10.295 2.425 ;
      RECT 9.945 3.635 10.025 3.895 ;
      RECT 9.235 2.355 9.355 2.615 ;
      RECT 9.92 3.615 9.945 3.895 ;
      RECT 9.905 3.577 9.92 3.895 ;
      RECT 9.865 3.52 9.905 3.895 ;
      RECT 9.835 3.43 9.865 3.895 ;
      RECT 9.795 3.33 9.835 3.895 ;
      RECT 9.765 3.23 9.795 3.895 ;
      RECT 9.76 3.177 9.765 3.718 ;
      RECT 9.745 3.147 9.76 3.684 ;
      RECT 9.735 3.108 9.745 3.649 ;
      RECT 9.725 3.075 9.735 3.605 ;
      RECT 9.715 3.042 9.725 3.57 ;
      RECT 9.685 2.976 9.715 3.505 ;
      RECT 9.675 2.911 9.685 3.43 ;
      RECT 9.665 2.881 9.675 3.4 ;
      RECT 9.625 2.811 9.665 3.33 ;
      RECT 9.615 2.746 9.625 3.245 ;
      RECT 9.605 2.728 9.615 3.23 ;
      RECT 9.595 2.711 9.605 3.195 ;
      RECT 9.585 2.694 9.595 3.165 ;
      RECT 9.575 2.677 9.585 3.135 ;
      RECT 9.555 2.652 9.575 3.075 ;
      RECT 9.545 2.626 9.555 3.02 ;
      RECT 9.525 2.601 9.545 2.98 ;
      RECT 9.515 2.57 9.525 2.945 ;
      RECT 9.505 2.557 9.515 2.9 ;
      RECT 9.495 2.542 9.505 2.875 ;
      RECT 9.485 2.355 9.495 2.835 ;
      RECT 9.475 2.355 9.485 2.805 ;
      RECT 9.47 2.355 9.475 2.788 ;
      RECT 9.465 2.355 9.47 2.77 ;
      RECT 9.395 2.355 9.465 2.71 ;
      RECT 9.355 2.355 9.395 2.645 ;
      RECT 9.185 3.225 9.445 3.485 ;
      RECT 7.355 3.145 7.435 3.465 ;
      RECT 7.175 3.205 7.325 3.465 ;
      RECT 7.355 3.145 7.465 3.425 ;
      RECT 9.175 3.317 9.185 3.48 ;
      RECT 9.145 3.327 9.175 3.488 ;
      RECT 9.125 3.335 9.145 3.493 ;
      RECT 9.057 3.343 9.125 3.503 ;
      RECT 8.971 3.363 9.057 3.52 ;
      RECT 8.885 3.384 8.971 3.539 ;
      RECT 8.875 3.4 8.885 3.55 ;
      RECT 8.835 3.41 8.875 3.556 ;
      RECT 8.815 3.415 8.835 3.563 ;
      RECT 8.777 3.416 8.815 3.566 ;
      RECT 8.691 3.419 8.777 3.567 ;
      RECT 8.605 3.423 8.691 3.568 ;
      RECT 8.551 3.425 8.605 3.57 ;
      RECT 8.465 3.425 8.551 3.572 ;
      RECT 8.425 3.42 8.465 3.574 ;
      RECT 8.415 3.414 8.425 3.575 ;
      RECT 8.375 3.409 8.415 3.571 ;
      RECT 8.365 3.4 8.375 3.567 ;
      RECT 8.333 3.391 8.365 3.564 ;
      RECT 8.247 3.379 8.333 3.554 ;
      RECT 8.161 3.362 8.247 3.539 ;
      RECT 8.075 3.344 8.161 3.525 ;
      RECT 8.055 3.335 8.075 3.516 ;
      RECT 7.985 3.325 8.055 3.509 ;
      RECT 7.935 3.31 7.985 3.499 ;
      RECT 7.875 3.3 7.935 3.49 ;
      RECT 7.835 3.29 7.875 3.485 ;
      RECT 7.785 3.28 7.835 3.479 ;
      RECT 7.745 3.268 7.785 3.469 ;
      RECT 7.725 3.258 7.745 3.465 ;
      RECT 7.705 3.248 7.725 3.465 ;
      RECT 7.695 3.238 7.705 3.464 ;
      RECT 7.675 3.23 7.695 3.46 ;
      RECT 7.635 3.205 7.675 3.454 ;
      RECT 7.615 3.145 7.635 3.447 ;
      RECT 7.591 3.145 7.615 3.444 ;
      RECT 7.505 3.145 7.591 3.439 ;
      RECT 7.465 3.145 7.505 3.43 ;
      RECT 7.325 3.195 7.355 3.465 ;
      RECT 9.005 2.775 9.265 3.035 ;
      RECT 8.965 2.775 9.265 2.915 ;
      RECT 8.935 2.775 9.265 2.9 ;
      RECT 8.875 2.775 9.265 2.88 ;
      RECT 8.795 2.585 9.075 2.865 ;
      RECT 8.795 2.77 9.145 2.865 ;
      RECT 8.795 2.71 9.135 2.865 ;
      RECT 8.795 2.66 9.085 2.865 ;
      RECT 6.565 3.115 6.825 3.375 ;
      RECT 6.71 1.205 6.825 3.375 ;
      RECT 6.625 2.585 6.825 3.375 ;
      RECT 7.935 2.635 8.195 2.895 ;
      RECT 6.62 2.585 6.825 2.87 ;
      RECT 6.615 2.585 6.825 2.865 ;
      RECT 7.915 2.645 8.195 2.825 ;
      RECT 7.505 2.615 7.645 2.765 ;
      RECT 6.88 1.205 6.96 1.55 ;
      RECT 6.615 1.205 6.825 1.55 ;
      RECT 7.905 2.644 7.915 2.825 ;
      RECT 7.901 2.644 7.905 2.825 ;
      RECT 7.815 2.639 7.901 2.814 ;
      RECT 7.741 2.63 7.815 2.794 ;
      RECT 7.655 2.621 7.741 2.775 ;
      RECT 7.645 2.615 7.655 2.765 ;
      RECT 7.465 2.615 7.505 2.768 ;
      RECT 7.379 2.615 7.465 2.776 ;
      RECT 7.293 2.615 7.379 2.787 ;
      RECT 7.207 2.615 7.293 2.798 ;
      RECT 7.121 2.615 7.207 2.809 ;
      RECT 7.035 2.615 7.121 2.82 ;
      RECT 7.005 2.615 7.035 2.86 ;
      RECT 6.975 2.615 7.005 2.91 ;
      RECT 6.9 2.615 6.975 2.93 ;
      RECT 6.895 2.59 6.9 2.935 ;
      RECT 6.88 2.585 6.895 2.943 ;
      RECT 6.875 1.205 6.88 2.953 ;
      RECT 6.845 1.205 6.875 2.995 ;
      RECT 6.825 1.205 6.845 3.075 ;
      RECT 5.955 2.965 5.975 3.404 ;
      RECT 5.955 2.965 6.061 3.401 ;
      RECT 5.945 3.08 6.061 3.4 ;
      RECT 5.975 2.115 6.105 3.397 ;
      RECT 5.955 2.985 6.115 3.395 ;
      RECT 5.955 3.07 6.125 3.39 ;
      RECT 5.925 3.115 6.125 3.385 ;
      RECT 5.925 3.115 6.135 3.38 ;
      RECT 5.905 3.115 6.165 3.375 ;
      RECT 5.975 2.115 6.135 2.765 ;
      RECT 5.965 2.115 6.135 2.74 ;
      RECT 5.965 2.115 6.155 2.505 ;
      RECT 5.915 2.115 6.175 2.375 ;
      RECT 5.385 2.605 5.675 2.865 ;
      RECT 5.395 2.585 5.675 2.865 ;
      RECT 5.345 2.665 5.675 2.86 ;
      RECT 5.415 2.578 5.585 2.865 ;
      RECT 5.415 2.565 5.541 2.865 ;
      RECT 5.455 2.558 5.541 2.865 ;
      RECT 4.915 3.705 5.195 3.985 ;
      RECT 4.875 3.67 5.175 3.78 ;
      RECT 4.865 3.62 5.155 3.675 ;
      RECT 4.805 3.385 5.065 3.645 ;
      RECT 4.805 3.525 5.145 3.645 ;
      RECT 4.805 3.475 5.125 3.645 ;
      RECT 4.805 3.43 5.115 3.645 ;
      RECT 4.805 3.415 5.085 3.645 ;
      RECT 1.65 8.5 2.03 8.88 ;
      RECT 1.715 8.485 1.855 8.88 ;
      RECT 85.7 7.055 86.075 7.425 ;
      RECT 77.035 0.93 77.41 1.3 ;
      RECT 67.775 7.055 68.15 7.425 ;
      RECT 59.11 0.93 59.485 1.3 ;
      RECT 49.85 7.055 50.225 7.425 ;
      RECT 41.185 0.93 41.56 1.3 ;
      RECT 31.925 7.055 32.3 7.425 ;
      RECT 23.26 0.93 23.635 1.3 ;
      RECT 14 7.055 14.375 7.425 ;
      RECT 5.335 0.93 5.71 1.3 ;
    LAYER via1 ;
      RECT 93.42 7.375 93.57 7.525 ;
      RECT 91.055 6.74 91.205 6.89 ;
      RECT 91.04 2.065 91.19 2.215 ;
      RECT 90.25 2.45 90.4 2.6 ;
      RECT 90.25 6.325 90.4 6.475 ;
      RECT 88.645 3.53 88.795 3.68 ;
      RECT 88.635 1.25 88.785 1.4 ;
      RECT 86.95 2.21 87.1 2.36 ;
      RECT 86.72 6.71 86.87 6.86 ;
      RECT 86 3.72 86.15 3.87 ;
      RECT 85.815 7.165 85.965 7.315 ;
      RECT 85.55 2.22 85.7 2.37 ;
      RECT 85.37 3.21 85.52 3.36 ;
      RECT 84.97 3.72 85.12 3.87 ;
      RECT 84.61 3.68 84.76 3.83 ;
      RECT 84.47 2.17 84.62 2.32 ;
      RECT 83.88 3.62 84.03 3.77 ;
      RECT 83.79 2.15 83.94 2.3 ;
      RECT 83.63 2.69 83.78 2.84 ;
      RECT 82.95 3.65 83.1 3.8 ;
      RECT 82.55 2.28 82.7 2.43 ;
      RECT 81.83 3.18 81.98 3.33 ;
      RECT 81.79 2.22 81.94 2.37 ;
      RECT 81.52 3.69 81.67 3.84 ;
      RECT 80.99 2.41 81.14 2.56 ;
      RECT 80.94 3.28 81.09 3.43 ;
      RECT 80.76 2.83 80.91 2.98 ;
      RECT 79.69 2.69 79.84 2.84 ;
      RECT 79.58 2.11 79.73 2.26 ;
      RECT 78.93 3.26 79.08 3.41 ;
      RECT 78.41 1.3 78.56 1.45 ;
      RECT 78.32 3.17 78.47 3.32 ;
      RECT 77.67 2.17 77.82 2.32 ;
      RECT 77.66 3.17 77.81 3.32 ;
      RECT 77.14 2.66 77.29 2.81 ;
      RECT 76.56 3.44 76.71 3.59 ;
      RECT 75.475 6.755 75.625 6.905 ;
      RECT 73.13 6.74 73.28 6.89 ;
      RECT 73.115 2.065 73.265 2.215 ;
      RECT 72.325 2.45 72.475 2.6 ;
      RECT 72.325 6.325 72.475 6.475 ;
      RECT 70.72 3.53 70.87 3.68 ;
      RECT 70.71 1.25 70.86 1.4 ;
      RECT 69.025 2.21 69.175 2.36 ;
      RECT 68.515 6.71 68.665 6.86 ;
      RECT 68.075 3.72 68.225 3.87 ;
      RECT 67.89 7.165 68.04 7.315 ;
      RECT 67.625 2.22 67.775 2.37 ;
      RECT 67.445 3.21 67.595 3.36 ;
      RECT 67.045 3.72 67.195 3.87 ;
      RECT 66.685 3.68 66.835 3.83 ;
      RECT 66.545 2.17 66.695 2.32 ;
      RECT 65.955 3.62 66.105 3.77 ;
      RECT 65.865 2.15 66.015 2.3 ;
      RECT 65.705 2.69 65.855 2.84 ;
      RECT 65.025 3.65 65.175 3.8 ;
      RECT 64.625 2.28 64.775 2.43 ;
      RECT 63.905 3.18 64.055 3.33 ;
      RECT 63.865 2.22 64.015 2.37 ;
      RECT 63.595 3.69 63.745 3.84 ;
      RECT 63.065 2.41 63.215 2.56 ;
      RECT 63.015 3.28 63.165 3.43 ;
      RECT 62.835 2.83 62.985 2.98 ;
      RECT 61.765 2.69 61.915 2.84 ;
      RECT 61.655 2.11 61.805 2.26 ;
      RECT 61.005 3.26 61.155 3.41 ;
      RECT 60.485 1.3 60.635 1.45 ;
      RECT 60.395 3.17 60.545 3.32 ;
      RECT 59.745 2.17 59.895 2.32 ;
      RECT 59.735 3.17 59.885 3.32 ;
      RECT 59.215 2.66 59.365 2.81 ;
      RECT 58.635 3.44 58.785 3.59 ;
      RECT 57.55 6.755 57.7 6.905 ;
      RECT 55.205 6.74 55.355 6.89 ;
      RECT 55.19 2.065 55.34 2.215 ;
      RECT 54.4 2.45 54.55 2.6 ;
      RECT 54.4 6.325 54.55 6.475 ;
      RECT 52.795 3.53 52.945 3.68 ;
      RECT 52.785 1.25 52.935 1.4 ;
      RECT 51.1 2.21 51.25 2.36 ;
      RECT 50.645 6.715 50.795 6.865 ;
      RECT 50.15 3.72 50.3 3.87 ;
      RECT 49.965 7.165 50.115 7.315 ;
      RECT 49.7 2.22 49.85 2.37 ;
      RECT 49.52 3.21 49.67 3.36 ;
      RECT 49.12 3.72 49.27 3.87 ;
      RECT 48.76 3.68 48.91 3.83 ;
      RECT 48.62 2.17 48.77 2.32 ;
      RECT 48.03 3.62 48.18 3.77 ;
      RECT 47.94 2.15 48.09 2.3 ;
      RECT 47.78 2.69 47.93 2.84 ;
      RECT 47.1 3.65 47.25 3.8 ;
      RECT 46.7 2.28 46.85 2.43 ;
      RECT 45.98 3.18 46.13 3.33 ;
      RECT 45.94 2.22 46.09 2.37 ;
      RECT 45.67 3.69 45.82 3.84 ;
      RECT 45.14 2.41 45.29 2.56 ;
      RECT 45.09 3.28 45.24 3.43 ;
      RECT 44.91 2.83 45.06 2.98 ;
      RECT 43.84 2.69 43.99 2.84 ;
      RECT 43.73 2.11 43.88 2.26 ;
      RECT 43.08 3.26 43.23 3.41 ;
      RECT 42.56 1.3 42.71 1.45 ;
      RECT 42.47 3.17 42.62 3.32 ;
      RECT 41.82 2.17 41.97 2.32 ;
      RECT 41.81 3.17 41.96 3.32 ;
      RECT 41.29 2.66 41.44 2.81 ;
      RECT 40.71 3.44 40.86 3.59 ;
      RECT 39.67 6.76 39.82 6.91 ;
      RECT 37.28 6.74 37.43 6.89 ;
      RECT 37.265 2.065 37.415 2.215 ;
      RECT 36.475 2.45 36.625 2.6 ;
      RECT 36.475 6.325 36.625 6.475 ;
      RECT 34.87 3.53 35.02 3.68 ;
      RECT 34.86 1.25 35.01 1.4 ;
      RECT 33.175 2.21 33.325 2.36 ;
      RECT 32.715 6.71 32.865 6.86 ;
      RECT 32.225 3.72 32.375 3.87 ;
      RECT 32.04 7.165 32.19 7.315 ;
      RECT 31.775 2.22 31.925 2.37 ;
      RECT 31.595 3.21 31.745 3.36 ;
      RECT 31.195 3.72 31.345 3.87 ;
      RECT 30.835 3.68 30.985 3.83 ;
      RECT 30.695 2.17 30.845 2.32 ;
      RECT 30.105 3.62 30.255 3.77 ;
      RECT 30.015 2.15 30.165 2.3 ;
      RECT 29.855 2.69 30.005 2.84 ;
      RECT 29.175 3.65 29.325 3.8 ;
      RECT 28.775 2.28 28.925 2.43 ;
      RECT 28.055 3.18 28.205 3.33 ;
      RECT 28.015 2.22 28.165 2.37 ;
      RECT 27.745 3.69 27.895 3.84 ;
      RECT 27.215 2.41 27.365 2.56 ;
      RECT 27.165 3.28 27.315 3.43 ;
      RECT 26.985 2.83 27.135 2.98 ;
      RECT 25.915 2.69 26.065 2.84 ;
      RECT 25.805 2.11 25.955 2.26 ;
      RECT 25.155 3.26 25.305 3.41 ;
      RECT 24.635 1.3 24.785 1.45 ;
      RECT 24.545 3.17 24.695 3.32 ;
      RECT 23.895 2.17 24.045 2.32 ;
      RECT 23.885 3.17 24.035 3.32 ;
      RECT 23.365 2.66 23.515 2.81 ;
      RECT 22.785 3.44 22.935 3.59 ;
      RECT 21.745 6.755 21.895 6.905 ;
      RECT 19.355 6.74 19.505 6.89 ;
      RECT 19.34 2.065 19.49 2.215 ;
      RECT 18.55 2.45 18.7 2.6 ;
      RECT 18.55 6.325 18.7 6.475 ;
      RECT 16.945 3.53 17.095 3.68 ;
      RECT 16.935 1.25 17.085 1.4 ;
      RECT 15.25 2.21 15.4 2.36 ;
      RECT 14.76 6.705 14.91 6.855 ;
      RECT 14.3 3.72 14.45 3.87 ;
      RECT 14.115 7.165 14.265 7.315 ;
      RECT 13.85 2.22 14 2.37 ;
      RECT 13.67 3.21 13.82 3.36 ;
      RECT 13.27 3.72 13.42 3.87 ;
      RECT 12.91 3.68 13.06 3.83 ;
      RECT 12.77 2.17 12.92 2.32 ;
      RECT 12.18 3.62 12.33 3.77 ;
      RECT 12.09 2.15 12.24 2.3 ;
      RECT 11.93 2.69 12.08 2.84 ;
      RECT 11.25 3.65 11.4 3.8 ;
      RECT 10.85 2.28 11 2.43 ;
      RECT 10.13 3.18 10.28 3.33 ;
      RECT 10.09 2.22 10.24 2.37 ;
      RECT 9.82 3.69 9.97 3.84 ;
      RECT 9.29 2.41 9.44 2.56 ;
      RECT 9.24 3.28 9.39 3.43 ;
      RECT 9.06 2.83 9.21 2.98 ;
      RECT 7.99 2.69 8.14 2.84 ;
      RECT 7.88 2.11 8.03 2.26 ;
      RECT 7.23 3.26 7.38 3.41 ;
      RECT 6.71 1.3 6.86 1.45 ;
      RECT 6.62 3.17 6.77 3.32 ;
      RECT 5.97 2.17 6.12 2.32 ;
      RECT 5.96 3.17 6.11 3.32 ;
      RECT 5.44 2.66 5.59 2.81 ;
      RECT 4.86 3.44 5.01 3.59 ;
      RECT 3.09 7.095 3.24 7.245 ;
      RECT 2.715 6.355 2.865 6.505 ;
      RECT 1.765 8.615 1.915 8.765 ;
    LAYER met1 ;
      RECT 76.345 1.285 88.305 1.885 ;
      RECT 80.77 0 88.305 1.885 ;
      RECT 58.42 1.285 70.38 1.885 ;
      RECT 62.845 0 70.38 1.885 ;
      RECT 40.495 1.285 52.455 1.885 ;
      RECT 44.92 0 52.455 1.885 ;
      RECT 22.57 1.285 34.53 1.885 ;
      RECT 26.995 0 34.53 1.885 ;
      RECT 4.645 1.285 16.605 1.885 ;
      RECT 9.07 0 16.605 1.885 ;
      RECT 76.34 0 77.085 1.68 ;
      RECT 58.415 0 59.16 1.68 ;
      RECT 40.49 0 41.235 1.68 ;
      RECT 22.565 0 23.31 1.68 ;
      RECT 4.64 0 5.385 1.68 ;
      RECT 79.335 0 80.49 1.885 ;
      RECT 76.34 1.255 79.055 1.68 ;
      RECT 77.365 0 79.055 1.885 ;
      RECT 61.41 0 62.565 1.885 ;
      RECT 58.415 1.255 61.13 1.68 ;
      RECT 59.44 0 61.13 1.885 ;
      RECT 43.485 0 44.64 1.885 ;
      RECT 40.49 1.255 43.205 1.68 ;
      RECT 41.515 0 43.205 1.885 ;
      RECT 25.56 0 26.715 1.885 ;
      RECT 22.565 1.255 25.28 1.68 ;
      RECT 23.59 0 25.28 1.885 ;
      RECT 7.635 0 8.79 1.885 ;
      RECT 4.64 1.255 7.355 1.68 ;
      RECT 5.665 0 7.355 1.885 ;
      RECT 77.365 0 88.305 1.005 ;
      RECT 59.44 0 70.38 1.005 ;
      RECT 41.515 0 52.455 1.005 ;
      RECT 23.59 0 34.53 1.005 ;
      RECT 5.665 0 16.605 1.005 ;
      RECT 76.34 0 88.305 0.975 ;
      RECT 58.415 0 70.38 0.975 ;
      RECT 40.49 0 52.455 0.975 ;
      RECT 22.565 0 34.53 0.975 ;
      RECT 4.64 0 16.605 0.975 ;
      RECT 93.715 0 93.895 0.305 ;
      RECT 75.79 0 91.765 0.305 ;
      RECT 57.865 0 73.84 0.305 ;
      RECT 39.94 0 55.915 0.305 ;
      RECT 22.015 0 37.99 0.305 ;
      RECT 1.48 0 20.065 0.305 ;
      RECT 1.48 0 93.895 0.3 ;
      RECT 1.46 8.58 93.895 8.88 ;
      RECT 93.715 8.575 93.895 8.88 ;
      RECT 75.79 8.575 91.765 8.88 ;
      RECT 57.865 8.575 73.84 8.88 ;
      RECT 39.94 8.575 55.915 8.88 ;
      RECT 22.015 8.575 37.99 8.88 ;
      RECT 1.46 8.575 20.065 8.88 ;
      RECT 85.04 6.315 85.21 8.88 ;
      RECT 67.115 6.315 67.285 8.88 ;
      RECT 49.19 6.315 49.36 8.88 ;
      RECT 31.265 6.315 31.435 8.88 ;
      RECT 13.34 6.315 13.51 8.88 ;
      RECT 1.46 8.565 2.265 8.88 ;
      RECT 1.665 8.545 2.015 8.88 ;
      RECT 85.375 6.285 85.665 6.515 ;
      RECT 67.45 6.285 67.74 6.515 ;
      RECT 49.525 6.285 49.815 6.515 ;
      RECT 31.6 6.285 31.89 6.515 ;
      RECT 13.675 6.285 13.965 6.515 ;
      RECT 85.04 6.315 85.665 6.485 ;
      RECT 67.115 6.315 67.74 6.485 ;
      RECT 49.19 6.315 49.815 6.485 ;
      RECT 31.265 6.315 31.89 6.485 ;
      RECT 13.34 6.315 13.965 6.485 ;
      RECT 93.29 7.77 93.58 8 ;
      RECT 93.35 6.29 93.52 8 ;
      RECT 93.32 7.275 93.67 7.625 ;
      RECT 93.29 6.29 93.58 6.52 ;
      RECT 92.885 2.395 92.99 2.965 ;
      RECT 92.885 2.73 93.21 2.96 ;
      RECT 92.885 2.76 93.38 2.93 ;
      RECT 92.885 2.395 93.075 2.96 ;
      RECT 92.3 2.36 92.59 2.59 ;
      RECT 92.3 2.395 93.075 2.565 ;
      RECT 92.36 0.88 92.53 2.59 ;
      RECT 92.3 0.88 92.59 1.11 ;
      RECT 92.3 7.77 92.59 8 ;
      RECT 92.36 6.29 92.53 8 ;
      RECT 92.3 6.29 92.59 6.52 ;
      RECT 92.3 6.325 93.155 6.485 ;
      RECT 92.985 5.92 93.155 6.485 ;
      RECT 92.3 6.32 92.695 6.485 ;
      RECT 92.92 5.92 93.21 6.15 ;
      RECT 92.92 5.95 93.38 6.12 ;
      RECT 91.93 2.73 92.22 2.96 ;
      RECT 91.93 2.76 92.39 2.93 ;
      RECT 91.995 1.655 92.16 2.96 ;
      RECT 90.51 1.625 90.8 1.855 ;
      RECT 90.51 1.655 92.16 1.825 ;
      RECT 90.57 0.885 90.74 1.855 ;
      RECT 90.51 0.885 90.8 1.115 ;
      RECT 90.51 7.765 90.8 7.995 ;
      RECT 90.57 7.025 90.74 7.995 ;
      RECT 90.57 7.12 92.16 7.29 ;
      RECT 91.99 5.92 92.16 7.29 ;
      RECT 90.51 7.025 90.8 7.255 ;
      RECT 91.93 5.92 92.22 6.15 ;
      RECT 91.93 5.95 92.39 6.12 ;
      RECT 88.545 3.43 88.895 3.78 ;
      RECT 88.635 2.025 88.805 3.78 ;
      RECT 90.94 1.965 91.29 2.315 ;
      RECT 88.635 2.025 90.255 2.2 ;
      RECT 88.635 2.025 91.29 2.195 ;
      RECT 90.965 6.655 91.29 6.98 ;
      RECT 86.62 6.61 86.97 6.96 ;
      RECT 90.94 6.655 91.29 6.885 ;
      RECT 86.18 6.655 86.47 6.885 ;
      RECT 86.01 6.685 91.29 6.855 ;
      RECT 90.165 2.365 90.485 2.685 ;
      RECT 90.135 2.365 90.485 2.595 ;
      RECT 89.965 2.395 90.485 2.565 ;
      RECT 90.165 6.225 90.485 6.545 ;
      RECT 90.135 6.285 90.485 6.515 ;
      RECT 89.965 6.315 90.485 6.485 ;
      RECT 86.005 3.255 86.195 3.925 ;
      RECT 85.945 3.665 85.985 3.925 ;
      RECT 87.315 2.89 87.325 3.111 ;
      RECT 87.245 2.885 87.315 3.236 ;
      RECT 87.235 2.885 87.245 3.36 ;
      RECT 87.205 2.885 87.235 3.41 ;
      RECT 87.185 2.885 87.205 3.485 ;
      RECT 87.165 2.885 87.185 3.555 ;
      RECT 87.135 2.885 87.165 3.595 ;
      RECT 87.125 2.885 87.135 3.615 ;
      RECT 87.115 2.885 87.125 3.626 ;
      RECT 87.105 3.135 87.115 3.628 ;
      RECT 87.095 3.2 87.105 3.63 ;
      RECT 87.085 3.295 87.095 3.632 ;
      RECT 87.075 3.37 87.085 3.634 ;
      RECT 87.025 3.394 87.075 3.64 ;
      RECT 86.985 3.429 87.025 3.649 ;
      RECT 86.975 3.445 86.985 3.654 ;
      RECT 86.961 3.45 86.975 3.657 ;
      RECT 86.875 3.49 86.961 3.668 ;
      RECT 86.795 3.533 86.875 3.686 ;
      RECT 86.775 3.543 86.795 3.697 ;
      RECT 86.745 3.551 86.775 3.702 ;
      RECT 86.725 3.561 86.745 3.707 ;
      RECT 86.701 3.567 86.725 3.712 ;
      RECT 86.615 3.577 86.701 3.725 ;
      RECT 86.537 3.583 86.615 3.745 ;
      RECT 86.451 3.578 86.537 3.764 ;
      RECT 86.365 3.574 86.451 3.785 ;
      RECT 86.285 3.57 86.365 3.8 ;
      RECT 86.215 3.566 86.285 3.831 ;
      RECT 86.205 3.277 86.215 3.345 ;
      RECT 86.205 3.555 86.215 3.861 ;
      RECT 86.195 3.262 86.205 3.49 ;
      RECT 86.195 3.535 86.205 3.925 ;
      RECT 85.985 3.285 86.005 3.925 ;
      RECT 86.785 2.605 86.795 3.345 ;
      RECT 86.605 3.125 86.625 3.345 ;
      RECT 86.615 3.115 86.625 3.345 ;
      RECT 87.115 2.155 87.155 2.415 ;
      RECT 87.105 2.155 87.115 2.425 ;
      RECT 87.071 2.155 87.105 2.452 ;
      RECT 86.985 2.155 87.071 2.512 ;
      RECT 86.965 2.155 86.985 2.575 ;
      RECT 86.905 2.155 86.965 2.74 ;
      RECT 86.895 2.155 86.905 2.9 ;
      RECT 86.865 2.346 86.895 2.995 ;
      RECT 86.855 2.401 86.865 3.095 ;
      RECT 86.845 2.43 86.855 3.14 ;
      RECT 86.835 2.455 86.845 3.173 ;
      RECT 86.825 2.49 86.835 3.228 ;
      RECT 86.805 2.535 86.825 3.29 ;
      RECT 86.795 2.58 86.805 3.34 ;
      RECT 86.775 2.64 86.785 3.345 ;
      RECT 86.765 2.67 86.775 3.345 ;
      RECT 86.745 2.7 86.765 3.345 ;
      RECT 86.695 2.805 86.745 3.345 ;
      RECT 86.685 2.9 86.695 3.345 ;
      RECT 86.675 2.93 86.685 3.345 ;
      RECT 86.65 2.98 86.675 3.345 ;
      RECT 86.645 3.035 86.65 3.345 ;
      RECT 86.625 3.06 86.645 3.345 ;
      RECT 86.585 3.14 86.605 3.335 ;
      RECT 86.335 2.725 86.405 2.935 ;
      RECT 83.575 2.635 83.835 2.895 ;
      RECT 86.405 2.73 86.415 2.93 ;
      RECT 86.291 2.723 86.335 2.935 ;
      RECT 86.205 2.716 86.291 2.935 ;
      RECT 86.185 2.711 86.205 2.925 ;
      RECT 86.175 2.709 86.185 2.905 ;
      RECT 86.125 2.706 86.175 2.9 ;
      RECT 86.095 2.702 86.125 2.895 ;
      RECT 86.075 2.7 86.095 2.89 ;
      RECT 86.035 2.697 86.075 2.885 ;
      RECT 85.965 2.691 86.035 2.88 ;
      RECT 85.935 2.686 85.965 2.875 ;
      RECT 85.915 2.684 85.935 2.87 ;
      RECT 85.885 2.681 85.915 2.865 ;
      RECT 85.825 2.677 85.885 2.86 ;
      RECT 85.755 2.675 85.825 2.85 ;
      RECT 85.721 2.673 85.755 2.843 ;
      RECT 85.635 2.668 85.721 2.835 ;
      RECT 85.601 2.662 85.635 2.827 ;
      RECT 85.515 2.652 85.601 2.819 ;
      RECT 85.481 2.643 85.515 2.811 ;
      RECT 85.395 2.638 85.481 2.803 ;
      RECT 85.325 2.635 85.395 2.793 ;
      RECT 85.305 2.63 85.325 2.787 ;
      RECT 85.301 2.625 85.305 2.786 ;
      RECT 85.215 2.621 85.301 2.781 ;
      RECT 85.175 2.616 85.215 2.774 ;
      RECT 85.095 2.615 85.175 2.769 ;
      RECT 85.075 2.615 85.095 2.766 ;
      RECT 85.049 2.615 85.075 2.766 ;
      RECT 84.963 2.617 85.049 2.77 ;
      RECT 84.877 2.619 84.963 2.777 ;
      RECT 84.791 2.621 84.877 2.783 ;
      RECT 84.705 2.624 84.791 2.79 ;
      RECT 84.671 2.626 84.705 2.795 ;
      RECT 84.585 2.631 84.671 2.8 ;
      RECT 84.561 2.626 84.585 2.804 ;
      RECT 84.475 2.631 84.561 2.809 ;
      RECT 84.437 2.636 84.475 2.814 ;
      RECT 84.351 2.639 84.437 2.819 ;
      RECT 84.265 2.643 84.351 2.826 ;
      RECT 84.201 2.645 84.265 2.832 ;
      RECT 84.115 2.645 84.201 2.838 ;
      RECT 84.031 2.646 84.115 2.845 ;
      RECT 83.945 2.649 84.031 2.852 ;
      RECT 83.921 2.651 83.945 2.856 ;
      RECT 83.835 2.653 83.921 2.861 ;
      RECT 83.565 2.67 83.575 2.865 ;
      RECT 85.75 7.765 86.04 7.995 ;
      RECT 85.81 7.025 85.98 7.995 ;
      RECT 85.7 7.055 86.075 7.425 ;
      RECT 85.75 7.025 86.04 7.425 ;
      RECT 85.805 2.247 85.995 2.455 ;
      RECT 85.795 2.252 86.005 2.45 ;
      RECT 85.785 2.233 85.795 2.445 ;
      RECT 85.755 2.228 85.785 2.44 ;
      RECT 85.715 2.252 86.005 2.43 ;
      RECT 85.495 2.165 85.755 2.425 ;
      RECT 85.795 2.236 85.805 2.45 ;
      RECT 85.495 2.245 85.985 2.425 ;
      RECT 85.495 2.241 85.845 2.425 ;
      RECT 85.445 3.155 85.495 3.435 ;
      RECT 85.375 3.125 85.405 3.435 ;
      RECT 85.515 3.155 85.575 3.415 ;
      RECT 85.375 3.115 85.395 3.435 ;
      RECT 85.495 3.155 85.515 3.425 ;
      RECT 85.415 3.145 85.445 3.435 ;
      RECT 85.405 3.13 85.415 3.435 ;
      RECT 85.355 3.105 85.375 3.435 ;
      RECT 85.325 3.09 85.355 3.435 ;
      RECT 85.315 3.08 85.325 3.435 ;
      RECT 85.295 3.069 85.315 3.43 ;
      RECT 85.275 3.057 85.295 3.4 ;
      RECT 85.265 3.048 85.275 3.383 ;
      RECT 85.235 3.03 85.265 3.375 ;
      RECT 85.225 2.995 85.235 3.367 ;
      RECT 85.215 2.975 85.225 3.36 ;
      RECT 85.205 2.955 85.215 3.353 ;
      RECT 85.195 2.94 85.205 3.348 ;
      RECT 85.185 2.92 85.195 3.343 ;
      RECT 85.175 2.915 85.185 3.338 ;
      RECT 85.171 2.905 85.175 3.334 ;
      RECT 85.085 2.905 85.171 3.309 ;
      RECT 85.055 2.905 85.085 3.275 ;
      RECT 85.045 2.905 85.055 3.255 ;
      RECT 84.985 2.905 85.045 3.2 ;
      RECT 84.975 2.92 84.985 3.145 ;
      RECT 84.965 2.93 84.975 3.125 ;
      RECT 84.915 3.665 85.175 3.925 ;
      RECT 84.835 3.685 85.175 3.901 ;
      RECT 84.815 3.685 85.175 3.896 ;
      RECT 84.791 3.685 85.175 3.894 ;
      RECT 84.705 3.685 85.175 3.889 ;
      RECT 84.555 3.625 84.815 3.885 ;
      RECT 84.515 3.68 84.835 3.88 ;
      RECT 84.505 3.69 85.175 3.875 ;
      RECT 84.525 3.675 84.815 3.885 ;
      RECT 84.415 2.115 84.675 2.375 ;
      RECT 84.415 2.2 84.685 2.3 ;
      RECT 83.585 3.63 83.605 3.874 ;
      RECT 83.585 3.63 83.655 3.869 ;
      RECT 83.565 3.635 83.655 3.868 ;
      RECT 83.555 3.65 83.741 3.858 ;
      RECT 83.555 3.65 83.815 3.855 ;
      RECT 83.55 3.687 83.825 3.845 ;
      RECT 83.55 3.687 83.911 3.841 ;
      RECT 83.55 3.687 83.925 3.827 ;
      RECT 83.825 3.565 84.085 3.825 ;
      RECT 83.545 3.692 84.085 3.82 ;
      RECT 83.535 3.74 84.085 3.795 ;
      RECT 83.805 3.605 83.825 3.854 ;
      RECT 83.741 3.609 83.805 3.857 ;
      RECT 83.605 3.622 84.085 3.825 ;
      RECT 83.655 3.616 83.741 3.862 ;
      RECT 83.055 2.475 83.065 2.645 ;
      RECT 83.115 2.435 83.125 2.615 ;
      RECT 83.415 2.245 83.425 2.455 ;
      RECT 83.745 2.095 83.995 2.355 ;
      RECT 83.735 2.095 83.745 2.357 ;
      RECT 83.725 2.155 83.735 2.361 ;
      RECT 83.695 2.157 83.725 2.369 ;
      RECT 83.665 2.162 83.695 2.383 ;
      RECT 83.655 2.166 83.665 2.393 ;
      RECT 83.625 2.171 83.655 2.405 ;
      RECT 83.595 2.18 83.625 2.406 ;
      RECT 83.525 2.19 83.595 2.41 ;
      RECT 83.485 2.195 83.525 2.414 ;
      RECT 83.465 2.195 83.485 2.425 ;
      RECT 83.455 2.2 83.465 2.435 ;
      RECT 83.445 2.21 83.455 2.438 ;
      RECT 83.435 2.23 83.445 2.443 ;
      RECT 83.425 2.24 83.435 2.445 ;
      RECT 83.395 2.255 83.415 2.462 ;
      RECT 83.385 2.267 83.395 2.472 ;
      RECT 83.375 2.273 83.385 2.475 ;
      RECT 83.341 2.286 83.375 2.485 ;
      RECT 83.255 2.32 83.341 2.518 ;
      RECT 83.235 2.355 83.255 2.547 ;
      RECT 83.215 2.37 83.235 2.559 ;
      RECT 83.195 2.38 83.215 2.571 ;
      RECT 83.145 2.399 83.195 2.591 ;
      RECT 83.135 2.416 83.145 2.605 ;
      RECT 83.125 2.422 83.135 2.61 ;
      RECT 83.105 2.44 83.115 2.618 ;
      RECT 83.095 2.445 83.105 2.625 ;
      RECT 83.085 2.456 83.095 2.632 ;
      RECT 83.065 2.461 83.085 2.64 ;
      RECT 83.045 2.475 83.055 2.65 ;
      RECT 83.035 2.48 83.045 2.66 ;
      RECT 83.005 2.494 83.035 2.67 ;
      RECT 82.995 2.507 83.005 2.68 ;
      RECT 82.915 2.538 82.995 2.705 ;
      RECT 82.895 2.568 82.915 2.73 ;
      RECT 82.885 2.573 82.895 2.737 ;
      RECT 82.855 2.585 82.885 2.743 ;
      RECT 82.845 2.6 82.855 2.749 ;
      RECT 82.835 2.605 82.845 2.752 ;
      RECT 82.815 2.615 82.835 2.756 ;
      RECT 82.795 2.62 82.815 2.762 ;
      RECT 82.765 2.625 82.795 2.77 ;
      RECT 82.735 2.63 82.765 2.78 ;
      RECT 82.705 2.64 82.735 2.789 ;
      RECT 82.665 2.645 82.705 2.797 ;
      RECT 82.615 2.638 82.665 2.809 ;
      RECT 82.595 2.629 82.615 2.82 ;
      RECT 82.585 2.626 82.595 2.825 ;
      RECT 82.545 2.625 82.585 2.826 ;
      RECT 82.535 2.61 82.545 2.827 ;
      RECT 82.507 2.595 82.535 2.828 ;
      RECT 82.421 2.595 82.507 2.83 ;
      RECT 82.335 2.595 82.421 2.834 ;
      RECT 82.315 2.595 82.335 2.83 ;
      RECT 82.305 2.605 82.315 2.823 ;
      RECT 82.295 2.62 82.305 2.818 ;
      RECT 82.285 2.625 82.295 2.795 ;
      RECT 83.765 3.13 83.775 3.33 ;
      RECT 83.715 3.125 83.765 3.35 ;
      RECT 83.705 3.125 83.715 3.37 ;
      RECT 83.661 3.125 83.705 3.374 ;
      RECT 83.575 3.125 83.661 3.371 ;
      RECT 83.515 3.135 83.575 3.368 ;
      RECT 83.455 3.149 83.515 3.366 ;
      RECT 83.445 3.154 83.455 3.364 ;
      RECT 83.435 3.16 83.445 3.363 ;
      RECT 83.365 3.173 83.435 3.359 ;
      RECT 83.317 3.187 83.365 3.36 ;
      RECT 83.231 3.203 83.317 3.372 ;
      RECT 83.145 3.224 83.231 3.388 ;
      RECT 83.125 3.235 83.145 3.398 ;
      RECT 83.045 3.245 83.125 3.408 ;
      RECT 83.011 3.259 83.045 3.42 ;
      RECT 82.925 3.274 83.011 3.435 ;
      RECT 82.895 3.29 82.925 3.445 ;
      RECT 82.84 3.305 82.895 3.456 ;
      RECT 82.795 3.323 82.84 3.476 ;
      RECT 82.741 3.342 82.795 3.496 ;
      RECT 82.655 3.368 82.741 3.523 ;
      RECT 82.635 3.39 82.655 3.543 ;
      RECT 82.575 3.405 82.635 3.559 ;
      RECT 82.565 3.42 82.575 3.573 ;
      RECT 82.545 3.425 82.565 3.579 ;
      RECT 82.515 3.438 82.545 3.589 ;
      RECT 82.495 3.443 82.515 3.598 ;
      RECT 82.485 3.45 82.495 3.603 ;
      RECT 82.475 3.455 82.485 3.606 ;
      RECT 82.435 3.465 82.475 3.615 ;
      RECT 82.41 3.48 82.435 3.627 ;
      RECT 82.365 3.495 82.41 3.639 ;
      RECT 82.345 3.507 82.365 3.651 ;
      RECT 82.315 3.512 82.345 3.661 ;
      RECT 82.295 3.519 82.315 3.671 ;
      RECT 82.285 3.525 82.295 3.68 ;
      RECT 82.261 3.532 82.285 3.69 ;
      RECT 82.175 3.554 82.261 3.71 ;
      RECT 82.165 3.573 82.175 3.725 ;
      RECT 82.141 3.58 82.165 3.731 ;
      RECT 82.055 3.602 82.141 3.756 ;
      RECT 82.015 3.627 82.055 3.783 ;
      RECT 82.005 3.636 82.015 3.793 ;
      RECT 81.955 3.646 82.005 3.802 ;
      RECT 81.935 3.66 81.955 3.812 ;
      RECT 81.905 3.67 81.935 3.817 ;
      RECT 81.895 3.675 81.905 3.82 ;
      RECT 81.821 3.677 81.895 3.827 ;
      RECT 81.735 3.681 81.821 3.839 ;
      RECT 81.725 3.684 81.735 3.845 ;
      RECT 81.465 3.635 81.725 3.895 ;
      RECT 82.995 3.705 83.185 3.915 ;
      RECT 82.985 3.71 83.195 3.91 ;
      RECT 82.975 3.71 83.195 3.875 ;
      RECT 82.895 3.595 83.155 3.855 ;
      RECT 81.805 3.125 81.995 3.425 ;
      RECT 81.795 3.125 81.995 3.42 ;
      RECT 81.785 3.125 82.005 3.415 ;
      RECT 81.775 3.125 82.005 3.41 ;
      RECT 81.775 3.125 82.035 3.385 ;
      RECT 81.735 2.165 81.995 2.425 ;
      RECT 81.545 2.09 81.631 2.423 ;
      RECT 81.545 2.09 81.675 2.419 ;
      RECT 81.525 2.094 81.685 2.418 ;
      RECT 81.675 2.085 81.685 2.418 ;
      RECT 81.545 2.09 81.695 2.417 ;
      RECT 81.525 2.1 81.735 2.416 ;
      RECT 81.515 2.095 81.695 2.408 ;
      RECT 81.505 2.11 81.735 2.315 ;
      RECT 81.505 2.16 81.935 2.315 ;
      RECT 81.505 2.15 81.915 2.315 ;
      RECT 81.505 2.14 81.885 2.315 ;
      RECT 81.505 2.13 81.825 2.315 ;
      RECT 81.505 2.115 81.805 2.315 ;
      RECT 81.631 2.086 81.685 2.418 ;
      RECT 80.705 2.745 80.845 3.035 ;
      RECT 80.965 2.768 80.975 2.955 ;
      RECT 81.665 2.665 81.845 2.895 ;
      RECT 81.665 2.665 81.855 2.885 ;
      RECT 81.875 2.67 81.885 2.875 ;
      RECT 81.855 2.665 81.875 2.88 ;
      RECT 81.615 2.669 81.665 2.895 ;
      RECT 81.605 2.674 81.615 2.895 ;
      RECT 81.571 2.679 81.605 2.896 ;
      RECT 81.485 2.694 81.571 2.898 ;
      RECT 81.471 2.706 81.485 2.901 ;
      RECT 81.385 2.716 81.471 2.903 ;
      RECT 81.361 2.726 81.385 2.905 ;
      RECT 81.275 2.737 81.361 2.905 ;
      RECT 81.245 2.747 81.275 2.905 ;
      RECT 81.215 2.752 81.245 2.908 ;
      RECT 81.195 2.757 81.215 2.913 ;
      RECT 81.175 2.762 81.195 2.915 ;
      RECT 81.125 2.77 81.175 2.915 ;
      RECT 81.105 2.774 81.125 2.915 ;
      RECT 81.085 2.773 81.105 2.92 ;
      RECT 81.025 2.771 81.085 2.935 ;
      RECT 80.975 2.769 81.025 2.95 ;
      RECT 80.885 2.766 80.965 3.035 ;
      RECT 80.855 2.76 80.885 3.035 ;
      RECT 80.845 2.75 80.855 3.035 ;
      RECT 80.655 2.745 80.705 2.96 ;
      RECT 80.645 2.75 80.655 2.95 ;
      RECT 80.885 3.225 81.145 3.485 ;
      RECT 80.885 3.225 81.175 3.375 ;
      RECT 80.885 3.225 81.215 3.36 ;
      RECT 81.145 3.145 81.335 3.355 ;
      RECT 81.145 3.15 81.345 3.345 ;
      RECT 81.095 3.22 81.345 3.345 ;
      RECT 81.125 3.155 81.145 3.485 ;
      RECT 81.115 3.18 81.345 3.345 ;
      RECT 80.295 3.125 80.305 3.355 ;
      RECT 80.195 2.245 80.265 3.355 ;
      RECT 80.935 2.355 81.195 2.615 ;
      RECT 80.635 2.405 80.765 2.565 ;
      RECT 80.851 2.412 80.935 2.565 ;
      RECT 80.765 2.407 80.851 2.565 ;
      RECT 80.575 2.405 80.635 2.575 ;
      RECT 80.545 2.403 80.575 2.59 ;
      RECT 80.525 2.401 80.545 2.6 ;
      RECT 80.515 2.399 80.525 2.605 ;
      RECT 80.495 2.398 80.515 2.615 ;
      RECT 80.485 2.396 80.495 2.62 ;
      RECT 80.465 2.395 80.485 2.625 ;
      RECT 80.445 2.39 80.465 2.63 ;
      RECT 80.415 2.376 80.445 2.64 ;
      RECT 80.375 2.355 80.415 2.655 ;
      RECT 80.365 2.34 80.375 2.665 ;
      RECT 80.345 2.331 80.365 2.675 ;
      RECT 80.335 2.322 80.345 2.695 ;
      RECT 80.325 2.317 80.335 2.755 ;
      RECT 80.305 2.311 80.325 2.84 ;
      RECT 80.305 3.15 80.315 3.35 ;
      RECT 80.295 2.306 80.305 3.07 ;
      RECT 80.285 2.28 80.295 3.355 ;
      RECT 80.265 2.25 80.285 3.355 ;
      RECT 80.175 2.245 80.195 2.58 ;
      RECT 80.185 2.68 80.195 3.355 ;
      RECT 80.175 2.72 80.185 3.355 ;
      RECT 80.145 2.245 80.175 2.525 ;
      RECT 80.155 2.81 80.175 3.355 ;
      RECT 80.14 2.915 80.155 3.355 ;
      RECT 80.115 2.245 80.145 2.48 ;
      RECT 80.135 2.947 80.14 3.355 ;
      RECT 80.115 3.05 80.135 3.355 ;
      RECT 80.105 2.245 80.115 2.47 ;
      RECT 80.105 3.12 80.115 3.35 ;
      RECT 80.085 2.245 80.105 2.46 ;
      RECT 80.075 2.25 80.085 2.45 ;
      RECT 80.285 3.525 80.305 3.765 ;
      RECT 79.605 3.455 79.685 3.725 ;
      RECT 79.515 3.455 79.525 3.665 ;
      RECT 80.795 3.525 80.805 3.725 ;
      RECT 80.715 3.515 80.795 3.75 ;
      RECT 80.711 3.515 80.715 3.776 ;
      RECT 80.625 3.515 80.711 3.786 ;
      RECT 80.605 3.515 80.625 3.794 ;
      RECT 80.581 3.516 80.605 3.792 ;
      RECT 80.495 3.521 80.581 3.787 ;
      RECT 80.477 3.525 80.495 3.781 ;
      RECT 80.391 3.525 80.477 3.777 ;
      RECT 80.305 3.525 80.391 3.769 ;
      RECT 80.201 3.525 80.285 3.762 ;
      RECT 80.115 3.525 80.201 3.756 ;
      RECT 80.055 3.52 80.115 3.75 ;
      RECT 80.027 3.514 80.055 3.747 ;
      RECT 79.941 3.511 80.027 3.744 ;
      RECT 79.855 3.507 79.941 3.738 ;
      RECT 79.81 3.495 79.855 3.734 ;
      RECT 79.785 3.48 79.81 3.732 ;
      RECT 79.745 3.465 79.785 3.73 ;
      RECT 79.685 3.455 79.745 3.727 ;
      RECT 79.595 3.455 79.605 3.72 ;
      RECT 79.58 3.455 79.595 3.71 ;
      RECT 79.525 3.455 79.58 3.685 ;
      RECT 79.505 3.47 79.515 3.66 ;
      RECT 79.635 2.635 79.895 2.895 ;
      RECT 79.635 2.645 79.915 2.855 ;
      RECT 79.635 2.65 79.925 2.85 ;
      RECT 77.615 2.115 77.875 2.375 ;
      RECT 77.605 2.145 77.875 2.355 ;
      RECT 79.535 2.055 79.785 2.315 ;
      RECT 79.525 2.055 79.535 2.316 ;
      RECT 79.495 2.14 79.525 2.318 ;
      RECT 79.485 2.145 79.495 2.32 ;
      RECT 79.425 2.16 79.485 2.326 ;
      RECT 79.395 2.18 79.425 2.333 ;
      RECT 79.365 2.191 79.395 2.34 ;
      RECT 79.345 2.201 79.365 2.345 ;
      RECT 79.327 2.204 79.345 2.344 ;
      RECT 79.241 2.203 79.327 2.344 ;
      RECT 79.155 2.2 79.241 2.343 ;
      RECT 79.069 2.197 79.155 2.342 ;
      RECT 78.983 2.194 79.069 2.342 ;
      RECT 78.897 2.192 78.983 2.341 ;
      RECT 78.811 2.189 78.897 2.34 ;
      RECT 78.725 2.186 78.811 2.34 ;
      RECT 78.707 2.185 78.725 2.339 ;
      RECT 78.621 2.184 78.707 2.339 ;
      RECT 78.535 2.182 78.621 2.338 ;
      RECT 78.449 2.181 78.535 2.338 ;
      RECT 78.363 2.18 78.449 2.337 ;
      RECT 78.277 2.178 78.363 2.337 ;
      RECT 78.191 2.177 78.277 2.336 ;
      RECT 78.105 2.175 78.191 2.336 ;
      RECT 78.081 2.174 78.105 2.335 ;
      RECT 77.995 2.169 78.081 2.335 ;
      RECT 77.961 2.162 77.995 2.335 ;
      RECT 77.875 2.152 77.961 2.335 ;
      RECT 77.595 2.15 77.605 2.35 ;
      RECT 78.875 3.205 79.135 3.465 ;
      RECT 78.875 3.205 79.215 3.251 ;
      RECT 79.015 3.185 79.225 3.24 ;
      RECT 79.075 3.16 79.285 3.2 ;
      RECT 79.085 3.155 79.285 3.2 ;
      RECT 79.095 3.13 79.285 3.2 ;
      RECT 79.155 2.96 79.205 3.29 ;
      RECT 79.105 3.09 79.295 3.15 ;
      RECT 79.145 3.016 79.155 3.329 ;
      RECT 79.105 3.09 79.325 3.125 ;
      RECT 79.105 3.09 79.345 3.1 ;
      RECT 79.215 2.89 79.405 3.095 ;
      RECT 79.205 2.9 79.415 3.09 ;
      RECT 79.125 3.063 79.415 3.09 ;
      RECT 79.135 3.039 79.145 3.345 ;
      RECT 79.225 2.885 79.395 3.095 ;
      RECT 78.515 2.675 78.705 2.885 ;
      RECT 77.085 2.605 77.345 2.865 ;
      RECT 77.435 2.595 77.535 2.805 ;
      RECT 77.385 2.615 77.425 2.805 ;
      RECT 78.705 2.685 78.715 2.88 ;
      RECT 78.505 2.685 78.515 2.88 ;
      RECT 78.485 2.7 78.505 2.87 ;
      RECT 78.475 2.71 78.485 2.865 ;
      RECT 78.435 2.71 78.475 2.863 ;
      RECT 78.411 2.704 78.435 2.86 ;
      RECT 78.325 2.699 78.411 2.857 ;
      RECT 78.265 2.695 78.325 2.852 ;
      RECT 78.231 2.692 78.265 2.849 ;
      RECT 78.145 2.682 78.231 2.845 ;
      RECT 78.141 2.675 78.145 2.842 ;
      RECT 78.055 2.67 78.141 2.84 ;
      RECT 78.027 2.663 78.055 2.836 ;
      RECT 77.941 2.658 78.027 2.833 ;
      RECT 77.855 2.649 77.941 2.828 ;
      RECT 77.845 2.644 77.855 2.825 ;
      RECT 77.831 2.643 77.845 2.825 ;
      RECT 77.745 2.639 77.831 2.82 ;
      RECT 77.725 2.633 77.745 2.816 ;
      RECT 77.665 2.628 77.725 2.815 ;
      RECT 77.635 2.62 77.665 2.815 ;
      RECT 77.625 2.605 77.635 2.815 ;
      RECT 77.621 2.595 77.625 2.814 ;
      RECT 77.535 2.595 77.621 2.81 ;
      RECT 77.425 2.605 77.435 2.805 ;
      RECT 77.355 2.615 77.385 2.8 ;
      RECT 77.345 2.615 77.355 2.8 ;
      RECT 78.265 3.115 78.525 3.375 ;
      RECT 78.195 3.125 78.525 3.335 ;
      RECT 78.185 3.13 78.525 3.33 ;
      RECT 77.605 3.115 77.865 3.375 ;
      RECT 77.605 3.16 77.975 3.365 ;
      RECT 77.605 3.155 77.965 3.365 ;
      RECT 76.515 3.322 76.695 3.765 ;
      RECT 76.505 3.322 76.695 3.763 ;
      RECT 76.505 3.337 76.705 3.76 ;
      RECT 76.495 2.26 76.625 3.758 ;
      RECT 76.495 3.385 76.765 3.645 ;
      RECT 76.495 3.36 76.715 3.645 ;
      RECT 76.495 3.295 76.685 3.758 ;
      RECT 76.495 3.255 76.655 3.758 ;
      RECT 76.495 3.21 76.645 3.758 ;
      RECT 76.495 3.15 76.635 3.758 ;
      RECT 76.485 2.545 76.625 3.2 ;
      RECT 76.525 2.245 76.635 3.065 ;
      RECT 76.495 2.26 76.675 2.52 ;
      RECT 76.495 2.26 76.685 2.47 ;
      RECT 76.525 2.245 76.695 2.463 ;
      RECT 76.515 2.247 76.705 2.458 ;
      RECT 76.505 2.252 76.715 2.45 ;
      RECT 75.365 7.77 75.655 8 ;
      RECT 75.425 6.29 75.595 8 ;
      RECT 75.375 6.655 75.725 7.005 ;
      RECT 75.365 6.29 75.655 6.52 ;
      RECT 74.96 2.395 75.065 2.965 ;
      RECT 74.96 2.73 75.285 2.96 ;
      RECT 74.96 2.76 75.455 2.93 ;
      RECT 74.96 2.395 75.15 2.96 ;
      RECT 74.375 2.36 74.665 2.59 ;
      RECT 74.375 2.395 75.15 2.565 ;
      RECT 74.435 0.88 74.605 2.59 ;
      RECT 74.375 0.88 74.665 1.11 ;
      RECT 74.375 7.77 74.665 8 ;
      RECT 74.435 6.29 74.605 8 ;
      RECT 74.375 6.29 74.665 6.52 ;
      RECT 74.375 6.325 75.23 6.485 ;
      RECT 75.06 5.92 75.23 6.485 ;
      RECT 74.375 6.32 74.77 6.485 ;
      RECT 74.995 5.92 75.285 6.15 ;
      RECT 74.995 5.95 75.455 6.12 ;
      RECT 74.005 2.73 74.295 2.96 ;
      RECT 74.005 2.76 74.465 2.93 ;
      RECT 74.07 1.655 74.235 2.96 ;
      RECT 72.585 1.625 72.875 1.855 ;
      RECT 72.585 1.655 74.235 1.825 ;
      RECT 72.645 0.885 72.815 1.855 ;
      RECT 72.585 0.885 72.875 1.115 ;
      RECT 72.585 7.765 72.875 7.995 ;
      RECT 72.645 7.025 72.815 7.995 ;
      RECT 72.645 7.12 74.235 7.29 ;
      RECT 74.065 5.92 74.235 7.29 ;
      RECT 72.585 7.025 72.875 7.255 ;
      RECT 74.005 5.92 74.295 6.15 ;
      RECT 74.005 5.95 74.465 6.12 ;
      RECT 70.62 3.43 70.97 3.78 ;
      RECT 70.71 2.025 70.88 3.78 ;
      RECT 73.015 1.965 73.365 2.315 ;
      RECT 70.71 2.025 72.33 2.2 ;
      RECT 70.71 2.025 73.365 2.195 ;
      RECT 73.04 6.655 73.365 6.98 ;
      RECT 68.415 6.61 68.765 6.96 ;
      RECT 73.015 6.655 73.365 6.885 ;
      RECT 68.255 6.655 68.765 6.885 ;
      RECT 68.085 6.685 73.365 6.855 ;
      RECT 72.24 2.365 72.56 2.685 ;
      RECT 72.21 2.365 72.56 2.595 ;
      RECT 72.04 2.395 72.56 2.565 ;
      RECT 72.24 6.225 72.56 6.545 ;
      RECT 72.21 6.285 72.56 6.515 ;
      RECT 72.04 6.315 72.56 6.485 ;
      RECT 68.08 3.255 68.27 3.925 ;
      RECT 68.02 3.665 68.06 3.925 ;
      RECT 69.39 2.89 69.4 3.111 ;
      RECT 69.32 2.885 69.39 3.236 ;
      RECT 69.31 2.885 69.32 3.36 ;
      RECT 69.28 2.885 69.31 3.41 ;
      RECT 69.26 2.885 69.28 3.485 ;
      RECT 69.24 2.885 69.26 3.555 ;
      RECT 69.21 2.885 69.24 3.595 ;
      RECT 69.2 2.885 69.21 3.615 ;
      RECT 69.19 2.885 69.2 3.626 ;
      RECT 69.18 3.135 69.19 3.628 ;
      RECT 69.17 3.2 69.18 3.63 ;
      RECT 69.16 3.295 69.17 3.632 ;
      RECT 69.15 3.37 69.16 3.634 ;
      RECT 69.1 3.394 69.15 3.64 ;
      RECT 69.06 3.429 69.1 3.649 ;
      RECT 69.05 3.445 69.06 3.654 ;
      RECT 69.036 3.45 69.05 3.657 ;
      RECT 68.95 3.49 69.036 3.668 ;
      RECT 68.87 3.533 68.95 3.686 ;
      RECT 68.85 3.543 68.87 3.697 ;
      RECT 68.82 3.551 68.85 3.702 ;
      RECT 68.8 3.561 68.82 3.707 ;
      RECT 68.776 3.567 68.8 3.712 ;
      RECT 68.69 3.577 68.776 3.725 ;
      RECT 68.612 3.583 68.69 3.745 ;
      RECT 68.526 3.578 68.612 3.764 ;
      RECT 68.44 3.574 68.526 3.785 ;
      RECT 68.36 3.57 68.44 3.8 ;
      RECT 68.29 3.566 68.36 3.831 ;
      RECT 68.28 3.277 68.29 3.345 ;
      RECT 68.28 3.555 68.29 3.861 ;
      RECT 68.27 3.262 68.28 3.49 ;
      RECT 68.27 3.535 68.28 3.925 ;
      RECT 68.06 3.285 68.08 3.925 ;
      RECT 68.86 2.605 68.87 3.345 ;
      RECT 68.68 3.125 68.7 3.345 ;
      RECT 68.69 3.115 68.7 3.345 ;
      RECT 69.19 2.155 69.23 2.415 ;
      RECT 69.18 2.155 69.19 2.425 ;
      RECT 69.146 2.155 69.18 2.452 ;
      RECT 69.06 2.155 69.146 2.512 ;
      RECT 69.04 2.155 69.06 2.575 ;
      RECT 68.98 2.155 69.04 2.74 ;
      RECT 68.97 2.155 68.98 2.9 ;
      RECT 68.94 2.346 68.97 2.995 ;
      RECT 68.93 2.401 68.94 3.095 ;
      RECT 68.92 2.43 68.93 3.14 ;
      RECT 68.91 2.455 68.92 3.173 ;
      RECT 68.9 2.49 68.91 3.228 ;
      RECT 68.88 2.535 68.9 3.29 ;
      RECT 68.87 2.58 68.88 3.34 ;
      RECT 68.85 2.64 68.86 3.345 ;
      RECT 68.84 2.67 68.85 3.345 ;
      RECT 68.82 2.7 68.84 3.345 ;
      RECT 68.77 2.805 68.82 3.345 ;
      RECT 68.76 2.9 68.77 3.345 ;
      RECT 68.75 2.93 68.76 3.345 ;
      RECT 68.725 2.98 68.75 3.345 ;
      RECT 68.72 3.035 68.725 3.345 ;
      RECT 68.7 3.06 68.72 3.345 ;
      RECT 68.66 3.14 68.68 3.335 ;
      RECT 68.41 2.725 68.48 2.935 ;
      RECT 65.65 2.635 65.91 2.895 ;
      RECT 68.48 2.73 68.49 2.93 ;
      RECT 68.366 2.723 68.41 2.935 ;
      RECT 68.28 2.716 68.366 2.935 ;
      RECT 68.26 2.711 68.28 2.925 ;
      RECT 68.25 2.709 68.26 2.905 ;
      RECT 68.2 2.706 68.25 2.9 ;
      RECT 68.17 2.702 68.2 2.895 ;
      RECT 68.15 2.7 68.17 2.89 ;
      RECT 68.11 2.697 68.15 2.885 ;
      RECT 68.04 2.691 68.11 2.88 ;
      RECT 68.01 2.686 68.04 2.875 ;
      RECT 67.99 2.684 68.01 2.87 ;
      RECT 67.96 2.681 67.99 2.865 ;
      RECT 67.9 2.677 67.96 2.86 ;
      RECT 67.83 2.675 67.9 2.85 ;
      RECT 67.796 2.673 67.83 2.843 ;
      RECT 67.71 2.668 67.796 2.835 ;
      RECT 67.676 2.662 67.71 2.827 ;
      RECT 67.59 2.652 67.676 2.819 ;
      RECT 67.556 2.643 67.59 2.811 ;
      RECT 67.47 2.638 67.556 2.803 ;
      RECT 67.4 2.635 67.47 2.793 ;
      RECT 67.38 2.63 67.4 2.787 ;
      RECT 67.376 2.625 67.38 2.786 ;
      RECT 67.29 2.621 67.376 2.781 ;
      RECT 67.25 2.616 67.29 2.774 ;
      RECT 67.17 2.615 67.25 2.769 ;
      RECT 67.15 2.615 67.17 2.766 ;
      RECT 67.124 2.615 67.15 2.766 ;
      RECT 67.038 2.617 67.124 2.77 ;
      RECT 66.952 2.619 67.038 2.777 ;
      RECT 66.866 2.621 66.952 2.783 ;
      RECT 66.78 2.624 66.866 2.79 ;
      RECT 66.746 2.626 66.78 2.795 ;
      RECT 66.66 2.631 66.746 2.8 ;
      RECT 66.636 2.626 66.66 2.804 ;
      RECT 66.55 2.631 66.636 2.809 ;
      RECT 66.512 2.636 66.55 2.814 ;
      RECT 66.426 2.639 66.512 2.819 ;
      RECT 66.34 2.643 66.426 2.826 ;
      RECT 66.276 2.645 66.34 2.832 ;
      RECT 66.19 2.645 66.276 2.838 ;
      RECT 66.106 2.646 66.19 2.845 ;
      RECT 66.02 2.649 66.106 2.852 ;
      RECT 65.996 2.651 66.02 2.856 ;
      RECT 65.91 2.653 65.996 2.861 ;
      RECT 65.64 2.67 65.65 2.865 ;
      RECT 67.825 7.765 68.115 7.995 ;
      RECT 67.885 7.025 68.055 7.995 ;
      RECT 67.775 7.055 68.15 7.425 ;
      RECT 67.825 7.025 68.115 7.425 ;
      RECT 67.88 2.247 68.07 2.455 ;
      RECT 67.87 2.252 68.08 2.45 ;
      RECT 67.86 2.233 67.87 2.445 ;
      RECT 67.83 2.228 67.86 2.44 ;
      RECT 67.79 2.252 68.08 2.43 ;
      RECT 67.57 2.165 67.83 2.425 ;
      RECT 67.87 2.236 67.88 2.45 ;
      RECT 67.57 2.245 68.06 2.425 ;
      RECT 67.57 2.241 67.92 2.425 ;
      RECT 67.52 3.155 67.57 3.435 ;
      RECT 67.45 3.125 67.48 3.435 ;
      RECT 67.59 3.155 67.65 3.415 ;
      RECT 67.45 3.115 67.47 3.435 ;
      RECT 67.57 3.155 67.59 3.425 ;
      RECT 67.49 3.145 67.52 3.435 ;
      RECT 67.48 3.13 67.49 3.435 ;
      RECT 67.43 3.105 67.45 3.435 ;
      RECT 67.4 3.09 67.43 3.435 ;
      RECT 67.39 3.08 67.4 3.435 ;
      RECT 67.37 3.069 67.39 3.43 ;
      RECT 67.35 3.057 67.37 3.4 ;
      RECT 67.34 3.048 67.35 3.383 ;
      RECT 67.31 3.03 67.34 3.375 ;
      RECT 67.3 2.995 67.31 3.367 ;
      RECT 67.29 2.975 67.3 3.36 ;
      RECT 67.28 2.955 67.29 3.353 ;
      RECT 67.27 2.94 67.28 3.348 ;
      RECT 67.26 2.92 67.27 3.343 ;
      RECT 67.25 2.915 67.26 3.338 ;
      RECT 67.246 2.905 67.25 3.334 ;
      RECT 67.16 2.905 67.246 3.309 ;
      RECT 67.13 2.905 67.16 3.275 ;
      RECT 67.12 2.905 67.13 3.255 ;
      RECT 67.06 2.905 67.12 3.2 ;
      RECT 67.05 2.92 67.06 3.145 ;
      RECT 67.04 2.93 67.05 3.125 ;
      RECT 66.99 3.665 67.25 3.925 ;
      RECT 66.91 3.685 67.25 3.901 ;
      RECT 66.89 3.685 67.25 3.896 ;
      RECT 66.866 3.685 67.25 3.894 ;
      RECT 66.78 3.685 67.25 3.889 ;
      RECT 66.63 3.625 66.89 3.885 ;
      RECT 66.59 3.68 66.91 3.88 ;
      RECT 66.58 3.69 67.25 3.875 ;
      RECT 66.6 3.675 66.89 3.885 ;
      RECT 66.49 2.115 66.75 2.375 ;
      RECT 66.49 2.2 66.76 2.3 ;
      RECT 65.66 3.63 65.68 3.874 ;
      RECT 65.66 3.63 65.73 3.869 ;
      RECT 65.64 3.635 65.73 3.868 ;
      RECT 65.63 3.65 65.816 3.858 ;
      RECT 65.63 3.65 65.89 3.855 ;
      RECT 65.625 3.687 65.9 3.845 ;
      RECT 65.625 3.687 65.986 3.841 ;
      RECT 65.625 3.687 66 3.827 ;
      RECT 65.9 3.565 66.16 3.825 ;
      RECT 65.62 3.692 66.16 3.82 ;
      RECT 65.61 3.74 66.16 3.795 ;
      RECT 65.88 3.605 65.9 3.854 ;
      RECT 65.816 3.609 65.88 3.857 ;
      RECT 65.68 3.622 66.16 3.825 ;
      RECT 65.73 3.616 65.816 3.862 ;
      RECT 65.13 2.475 65.14 2.645 ;
      RECT 65.19 2.435 65.2 2.615 ;
      RECT 65.49 2.245 65.5 2.455 ;
      RECT 65.82 2.095 66.07 2.355 ;
      RECT 65.81 2.095 65.82 2.357 ;
      RECT 65.8 2.155 65.81 2.361 ;
      RECT 65.77 2.157 65.8 2.369 ;
      RECT 65.74 2.162 65.77 2.383 ;
      RECT 65.73 2.166 65.74 2.393 ;
      RECT 65.7 2.171 65.73 2.405 ;
      RECT 65.67 2.18 65.7 2.406 ;
      RECT 65.6 2.19 65.67 2.41 ;
      RECT 65.56 2.195 65.6 2.414 ;
      RECT 65.54 2.195 65.56 2.425 ;
      RECT 65.53 2.2 65.54 2.435 ;
      RECT 65.52 2.21 65.53 2.438 ;
      RECT 65.51 2.23 65.52 2.443 ;
      RECT 65.5 2.24 65.51 2.445 ;
      RECT 65.47 2.255 65.49 2.462 ;
      RECT 65.46 2.267 65.47 2.472 ;
      RECT 65.45 2.273 65.46 2.475 ;
      RECT 65.416 2.286 65.45 2.485 ;
      RECT 65.33 2.32 65.416 2.518 ;
      RECT 65.31 2.355 65.33 2.547 ;
      RECT 65.29 2.37 65.31 2.559 ;
      RECT 65.27 2.38 65.29 2.571 ;
      RECT 65.22 2.399 65.27 2.591 ;
      RECT 65.21 2.416 65.22 2.605 ;
      RECT 65.2 2.422 65.21 2.61 ;
      RECT 65.18 2.44 65.19 2.618 ;
      RECT 65.17 2.445 65.18 2.625 ;
      RECT 65.16 2.456 65.17 2.632 ;
      RECT 65.14 2.461 65.16 2.64 ;
      RECT 65.12 2.475 65.13 2.65 ;
      RECT 65.11 2.48 65.12 2.66 ;
      RECT 65.08 2.494 65.11 2.67 ;
      RECT 65.07 2.507 65.08 2.68 ;
      RECT 64.99 2.538 65.07 2.705 ;
      RECT 64.97 2.568 64.99 2.73 ;
      RECT 64.96 2.573 64.97 2.737 ;
      RECT 64.93 2.585 64.96 2.743 ;
      RECT 64.92 2.6 64.93 2.749 ;
      RECT 64.91 2.605 64.92 2.752 ;
      RECT 64.89 2.615 64.91 2.756 ;
      RECT 64.87 2.62 64.89 2.762 ;
      RECT 64.84 2.625 64.87 2.77 ;
      RECT 64.81 2.63 64.84 2.78 ;
      RECT 64.78 2.64 64.81 2.789 ;
      RECT 64.74 2.645 64.78 2.797 ;
      RECT 64.69 2.638 64.74 2.809 ;
      RECT 64.67 2.629 64.69 2.82 ;
      RECT 64.66 2.626 64.67 2.825 ;
      RECT 64.62 2.625 64.66 2.826 ;
      RECT 64.61 2.61 64.62 2.827 ;
      RECT 64.582 2.595 64.61 2.828 ;
      RECT 64.496 2.595 64.582 2.83 ;
      RECT 64.41 2.595 64.496 2.834 ;
      RECT 64.39 2.595 64.41 2.83 ;
      RECT 64.38 2.605 64.39 2.823 ;
      RECT 64.37 2.62 64.38 2.818 ;
      RECT 64.36 2.625 64.37 2.795 ;
      RECT 65.84 3.13 65.85 3.33 ;
      RECT 65.79 3.125 65.84 3.35 ;
      RECT 65.78 3.125 65.79 3.37 ;
      RECT 65.736 3.125 65.78 3.374 ;
      RECT 65.65 3.125 65.736 3.371 ;
      RECT 65.59 3.135 65.65 3.368 ;
      RECT 65.53 3.149 65.59 3.366 ;
      RECT 65.52 3.154 65.53 3.364 ;
      RECT 65.51 3.16 65.52 3.363 ;
      RECT 65.44 3.173 65.51 3.359 ;
      RECT 65.392 3.187 65.44 3.36 ;
      RECT 65.306 3.203 65.392 3.372 ;
      RECT 65.22 3.224 65.306 3.388 ;
      RECT 65.2 3.235 65.22 3.398 ;
      RECT 65.12 3.245 65.2 3.408 ;
      RECT 65.086 3.259 65.12 3.42 ;
      RECT 65 3.274 65.086 3.435 ;
      RECT 64.97 3.29 65 3.445 ;
      RECT 64.915 3.305 64.97 3.456 ;
      RECT 64.87 3.323 64.915 3.476 ;
      RECT 64.816 3.342 64.87 3.496 ;
      RECT 64.73 3.368 64.816 3.523 ;
      RECT 64.71 3.39 64.73 3.543 ;
      RECT 64.65 3.405 64.71 3.559 ;
      RECT 64.64 3.42 64.65 3.573 ;
      RECT 64.62 3.425 64.64 3.579 ;
      RECT 64.59 3.438 64.62 3.589 ;
      RECT 64.57 3.443 64.59 3.598 ;
      RECT 64.56 3.45 64.57 3.603 ;
      RECT 64.55 3.455 64.56 3.606 ;
      RECT 64.51 3.465 64.55 3.615 ;
      RECT 64.485 3.48 64.51 3.627 ;
      RECT 64.44 3.495 64.485 3.639 ;
      RECT 64.42 3.507 64.44 3.651 ;
      RECT 64.39 3.512 64.42 3.661 ;
      RECT 64.37 3.519 64.39 3.671 ;
      RECT 64.36 3.525 64.37 3.68 ;
      RECT 64.336 3.532 64.36 3.69 ;
      RECT 64.25 3.554 64.336 3.71 ;
      RECT 64.24 3.573 64.25 3.725 ;
      RECT 64.216 3.58 64.24 3.731 ;
      RECT 64.13 3.602 64.216 3.756 ;
      RECT 64.09 3.627 64.13 3.783 ;
      RECT 64.08 3.636 64.09 3.793 ;
      RECT 64.03 3.646 64.08 3.802 ;
      RECT 64.01 3.66 64.03 3.812 ;
      RECT 63.98 3.67 64.01 3.817 ;
      RECT 63.97 3.675 63.98 3.82 ;
      RECT 63.896 3.677 63.97 3.827 ;
      RECT 63.81 3.681 63.896 3.839 ;
      RECT 63.8 3.684 63.81 3.845 ;
      RECT 63.54 3.635 63.8 3.895 ;
      RECT 65.07 3.705 65.26 3.915 ;
      RECT 65.06 3.71 65.27 3.91 ;
      RECT 65.05 3.71 65.27 3.875 ;
      RECT 64.97 3.595 65.23 3.855 ;
      RECT 63.88 3.125 64.07 3.425 ;
      RECT 63.87 3.125 64.07 3.42 ;
      RECT 63.86 3.125 64.08 3.415 ;
      RECT 63.85 3.125 64.08 3.41 ;
      RECT 63.85 3.125 64.11 3.385 ;
      RECT 63.81 2.165 64.07 2.425 ;
      RECT 63.62 2.09 63.706 2.423 ;
      RECT 63.62 2.09 63.75 2.419 ;
      RECT 63.6 2.094 63.76 2.418 ;
      RECT 63.75 2.085 63.76 2.418 ;
      RECT 63.62 2.09 63.77 2.417 ;
      RECT 63.6 2.1 63.81 2.416 ;
      RECT 63.59 2.095 63.77 2.408 ;
      RECT 63.58 2.11 63.81 2.315 ;
      RECT 63.58 2.16 64.01 2.315 ;
      RECT 63.58 2.15 63.99 2.315 ;
      RECT 63.58 2.14 63.96 2.315 ;
      RECT 63.58 2.13 63.9 2.315 ;
      RECT 63.58 2.115 63.88 2.315 ;
      RECT 63.706 2.086 63.76 2.418 ;
      RECT 62.78 2.745 62.92 3.035 ;
      RECT 63.04 2.768 63.05 2.955 ;
      RECT 63.74 2.665 63.92 2.895 ;
      RECT 63.74 2.665 63.93 2.885 ;
      RECT 63.95 2.67 63.96 2.875 ;
      RECT 63.93 2.665 63.95 2.88 ;
      RECT 63.69 2.669 63.74 2.895 ;
      RECT 63.68 2.674 63.69 2.895 ;
      RECT 63.646 2.679 63.68 2.896 ;
      RECT 63.56 2.694 63.646 2.898 ;
      RECT 63.546 2.706 63.56 2.901 ;
      RECT 63.46 2.716 63.546 2.903 ;
      RECT 63.436 2.726 63.46 2.905 ;
      RECT 63.35 2.737 63.436 2.905 ;
      RECT 63.32 2.747 63.35 2.905 ;
      RECT 63.29 2.752 63.32 2.908 ;
      RECT 63.27 2.757 63.29 2.913 ;
      RECT 63.25 2.762 63.27 2.915 ;
      RECT 63.2 2.77 63.25 2.915 ;
      RECT 63.18 2.774 63.2 2.915 ;
      RECT 63.16 2.773 63.18 2.92 ;
      RECT 63.1 2.771 63.16 2.935 ;
      RECT 63.05 2.769 63.1 2.95 ;
      RECT 62.96 2.766 63.04 3.035 ;
      RECT 62.93 2.76 62.96 3.035 ;
      RECT 62.92 2.75 62.93 3.035 ;
      RECT 62.73 2.745 62.78 2.96 ;
      RECT 62.72 2.75 62.73 2.95 ;
      RECT 62.96 3.225 63.22 3.485 ;
      RECT 62.96 3.225 63.25 3.375 ;
      RECT 62.96 3.225 63.29 3.36 ;
      RECT 63.22 3.145 63.41 3.355 ;
      RECT 63.22 3.15 63.42 3.345 ;
      RECT 63.17 3.22 63.42 3.345 ;
      RECT 63.2 3.155 63.22 3.485 ;
      RECT 63.19 3.18 63.42 3.345 ;
      RECT 62.37 3.125 62.38 3.355 ;
      RECT 62.27 2.245 62.34 3.355 ;
      RECT 63.01 2.355 63.27 2.615 ;
      RECT 62.71 2.405 62.84 2.565 ;
      RECT 62.926 2.412 63.01 2.565 ;
      RECT 62.84 2.407 62.926 2.565 ;
      RECT 62.65 2.405 62.71 2.575 ;
      RECT 62.62 2.403 62.65 2.59 ;
      RECT 62.6 2.401 62.62 2.6 ;
      RECT 62.59 2.399 62.6 2.605 ;
      RECT 62.57 2.398 62.59 2.615 ;
      RECT 62.56 2.396 62.57 2.62 ;
      RECT 62.54 2.395 62.56 2.625 ;
      RECT 62.52 2.39 62.54 2.63 ;
      RECT 62.49 2.376 62.52 2.64 ;
      RECT 62.45 2.355 62.49 2.655 ;
      RECT 62.44 2.34 62.45 2.665 ;
      RECT 62.42 2.331 62.44 2.675 ;
      RECT 62.41 2.322 62.42 2.695 ;
      RECT 62.4 2.317 62.41 2.755 ;
      RECT 62.38 2.311 62.4 2.84 ;
      RECT 62.38 3.15 62.39 3.35 ;
      RECT 62.37 2.306 62.38 3.07 ;
      RECT 62.36 2.28 62.37 3.355 ;
      RECT 62.34 2.25 62.36 3.355 ;
      RECT 62.25 2.245 62.27 2.58 ;
      RECT 62.26 2.68 62.27 3.355 ;
      RECT 62.25 2.72 62.26 3.355 ;
      RECT 62.22 2.245 62.25 2.525 ;
      RECT 62.23 2.81 62.25 3.355 ;
      RECT 62.215 2.915 62.23 3.355 ;
      RECT 62.19 2.245 62.22 2.48 ;
      RECT 62.21 2.947 62.215 3.355 ;
      RECT 62.19 3.05 62.21 3.355 ;
      RECT 62.18 2.245 62.19 2.47 ;
      RECT 62.18 3.12 62.19 3.35 ;
      RECT 62.16 2.245 62.18 2.46 ;
      RECT 62.15 2.25 62.16 2.45 ;
      RECT 62.36 3.525 62.38 3.765 ;
      RECT 61.68 3.455 61.76 3.725 ;
      RECT 61.59 3.455 61.6 3.665 ;
      RECT 62.87 3.525 62.88 3.725 ;
      RECT 62.79 3.515 62.87 3.75 ;
      RECT 62.786 3.515 62.79 3.776 ;
      RECT 62.7 3.515 62.786 3.786 ;
      RECT 62.68 3.515 62.7 3.794 ;
      RECT 62.656 3.516 62.68 3.792 ;
      RECT 62.57 3.521 62.656 3.787 ;
      RECT 62.552 3.525 62.57 3.781 ;
      RECT 62.466 3.525 62.552 3.777 ;
      RECT 62.38 3.525 62.466 3.769 ;
      RECT 62.276 3.525 62.36 3.762 ;
      RECT 62.19 3.525 62.276 3.756 ;
      RECT 62.13 3.52 62.19 3.75 ;
      RECT 62.102 3.514 62.13 3.747 ;
      RECT 62.016 3.511 62.102 3.744 ;
      RECT 61.93 3.507 62.016 3.738 ;
      RECT 61.885 3.495 61.93 3.734 ;
      RECT 61.86 3.48 61.885 3.732 ;
      RECT 61.82 3.465 61.86 3.73 ;
      RECT 61.76 3.455 61.82 3.727 ;
      RECT 61.67 3.455 61.68 3.72 ;
      RECT 61.655 3.455 61.67 3.71 ;
      RECT 61.6 3.455 61.655 3.685 ;
      RECT 61.58 3.47 61.59 3.66 ;
      RECT 61.71 2.635 61.97 2.895 ;
      RECT 61.71 2.645 61.99 2.855 ;
      RECT 61.71 2.65 62 2.85 ;
      RECT 59.69 2.115 59.95 2.375 ;
      RECT 59.68 2.145 59.95 2.355 ;
      RECT 61.61 2.055 61.86 2.315 ;
      RECT 61.6 2.055 61.61 2.316 ;
      RECT 61.57 2.14 61.6 2.318 ;
      RECT 61.56 2.145 61.57 2.32 ;
      RECT 61.5 2.16 61.56 2.326 ;
      RECT 61.47 2.18 61.5 2.333 ;
      RECT 61.44 2.191 61.47 2.34 ;
      RECT 61.42 2.201 61.44 2.345 ;
      RECT 61.402 2.204 61.42 2.344 ;
      RECT 61.316 2.203 61.402 2.344 ;
      RECT 61.23 2.2 61.316 2.343 ;
      RECT 61.144 2.197 61.23 2.342 ;
      RECT 61.058 2.194 61.144 2.342 ;
      RECT 60.972 2.192 61.058 2.341 ;
      RECT 60.886 2.189 60.972 2.34 ;
      RECT 60.8 2.186 60.886 2.34 ;
      RECT 60.782 2.185 60.8 2.339 ;
      RECT 60.696 2.184 60.782 2.339 ;
      RECT 60.61 2.182 60.696 2.338 ;
      RECT 60.524 2.181 60.61 2.338 ;
      RECT 60.438 2.18 60.524 2.337 ;
      RECT 60.352 2.178 60.438 2.337 ;
      RECT 60.266 2.177 60.352 2.336 ;
      RECT 60.18 2.175 60.266 2.336 ;
      RECT 60.156 2.174 60.18 2.335 ;
      RECT 60.07 2.169 60.156 2.335 ;
      RECT 60.036 2.162 60.07 2.335 ;
      RECT 59.95 2.152 60.036 2.335 ;
      RECT 59.67 2.15 59.68 2.35 ;
      RECT 60.95 3.205 61.21 3.465 ;
      RECT 60.95 3.205 61.29 3.251 ;
      RECT 61.09 3.185 61.3 3.24 ;
      RECT 61.15 3.16 61.36 3.2 ;
      RECT 61.16 3.155 61.36 3.2 ;
      RECT 61.17 3.13 61.36 3.2 ;
      RECT 61.23 2.96 61.28 3.29 ;
      RECT 61.18 3.09 61.37 3.15 ;
      RECT 61.22 3.016 61.23 3.329 ;
      RECT 61.18 3.09 61.4 3.125 ;
      RECT 61.18 3.09 61.42 3.1 ;
      RECT 61.29 2.89 61.48 3.095 ;
      RECT 61.28 2.9 61.49 3.09 ;
      RECT 61.2 3.063 61.49 3.09 ;
      RECT 61.21 3.039 61.22 3.345 ;
      RECT 61.3 2.885 61.47 3.095 ;
      RECT 60.59 2.675 60.78 2.885 ;
      RECT 59.16 2.605 59.42 2.865 ;
      RECT 59.51 2.595 59.61 2.805 ;
      RECT 59.46 2.615 59.5 2.805 ;
      RECT 60.78 2.685 60.79 2.88 ;
      RECT 60.58 2.685 60.59 2.88 ;
      RECT 60.56 2.7 60.58 2.87 ;
      RECT 60.55 2.71 60.56 2.865 ;
      RECT 60.51 2.71 60.55 2.863 ;
      RECT 60.486 2.704 60.51 2.86 ;
      RECT 60.4 2.699 60.486 2.857 ;
      RECT 60.34 2.695 60.4 2.852 ;
      RECT 60.306 2.692 60.34 2.849 ;
      RECT 60.22 2.682 60.306 2.845 ;
      RECT 60.216 2.675 60.22 2.842 ;
      RECT 60.13 2.67 60.216 2.84 ;
      RECT 60.102 2.663 60.13 2.836 ;
      RECT 60.016 2.658 60.102 2.833 ;
      RECT 59.93 2.649 60.016 2.828 ;
      RECT 59.92 2.644 59.93 2.825 ;
      RECT 59.906 2.643 59.92 2.825 ;
      RECT 59.82 2.639 59.906 2.82 ;
      RECT 59.8 2.633 59.82 2.816 ;
      RECT 59.74 2.628 59.8 2.815 ;
      RECT 59.71 2.62 59.74 2.815 ;
      RECT 59.7 2.605 59.71 2.815 ;
      RECT 59.696 2.595 59.7 2.814 ;
      RECT 59.61 2.595 59.696 2.81 ;
      RECT 59.5 2.605 59.51 2.805 ;
      RECT 59.43 2.615 59.46 2.8 ;
      RECT 59.42 2.615 59.43 2.8 ;
      RECT 60.34 3.115 60.6 3.375 ;
      RECT 60.27 3.125 60.6 3.335 ;
      RECT 60.26 3.13 60.6 3.33 ;
      RECT 59.68 3.115 59.94 3.375 ;
      RECT 59.68 3.16 60.05 3.365 ;
      RECT 59.68 3.155 60.04 3.365 ;
      RECT 58.59 3.322 58.77 3.765 ;
      RECT 58.58 3.322 58.77 3.763 ;
      RECT 58.58 3.337 58.78 3.76 ;
      RECT 58.57 2.26 58.7 3.758 ;
      RECT 58.57 3.385 58.84 3.645 ;
      RECT 58.57 3.36 58.79 3.645 ;
      RECT 58.57 3.295 58.76 3.758 ;
      RECT 58.57 3.255 58.73 3.758 ;
      RECT 58.57 3.21 58.72 3.758 ;
      RECT 58.57 3.15 58.71 3.758 ;
      RECT 58.56 2.545 58.7 3.2 ;
      RECT 58.6 2.245 58.71 3.065 ;
      RECT 58.57 2.26 58.75 2.52 ;
      RECT 58.57 2.26 58.76 2.47 ;
      RECT 58.6 2.245 58.77 2.463 ;
      RECT 58.59 2.247 58.78 2.458 ;
      RECT 58.58 2.252 58.79 2.45 ;
      RECT 57.44 7.77 57.73 8 ;
      RECT 57.5 6.29 57.67 8 ;
      RECT 57.45 6.655 57.8 7.005 ;
      RECT 57.44 6.29 57.73 6.52 ;
      RECT 57.035 2.395 57.14 2.965 ;
      RECT 57.035 2.73 57.36 2.96 ;
      RECT 57.035 2.76 57.53 2.93 ;
      RECT 57.035 2.395 57.225 2.96 ;
      RECT 56.45 2.36 56.74 2.59 ;
      RECT 56.45 2.395 57.225 2.565 ;
      RECT 56.51 0.88 56.68 2.59 ;
      RECT 56.45 0.88 56.74 1.11 ;
      RECT 56.45 7.77 56.74 8 ;
      RECT 56.51 6.29 56.68 8 ;
      RECT 56.45 6.29 56.74 6.52 ;
      RECT 56.45 6.325 57.305 6.485 ;
      RECT 57.135 5.92 57.305 6.485 ;
      RECT 56.45 6.32 56.845 6.485 ;
      RECT 57.07 5.92 57.36 6.15 ;
      RECT 57.07 5.95 57.53 6.12 ;
      RECT 56.08 2.73 56.37 2.96 ;
      RECT 56.08 2.76 56.54 2.93 ;
      RECT 56.145 1.655 56.31 2.96 ;
      RECT 54.66 1.625 54.95 1.855 ;
      RECT 54.66 1.655 56.31 1.825 ;
      RECT 54.72 0.885 54.89 1.855 ;
      RECT 54.66 0.885 54.95 1.115 ;
      RECT 54.66 7.765 54.95 7.995 ;
      RECT 54.72 7.025 54.89 7.995 ;
      RECT 54.72 7.12 56.31 7.29 ;
      RECT 56.14 5.92 56.31 7.29 ;
      RECT 54.66 7.025 54.95 7.255 ;
      RECT 56.08 5.92 56.37 6.15 ;
      RECT 56.08 5.95 56.54 6.12 ;
      RECT 52.695 3.43 53.045 3.78 ;
      RECT 52.785 2.025 52.955 3.78 ;
      RECT 55.09 1.965 55.44 2.315 ;
      RECT 52.785 2.025 54.405 2.2 ;
      RECT 52.785 2.025 55.44 2.195 ;
      RECT 55.115 6.655 55.44 6.98 ;
      RECT 50.545 6.615 50.895 6.965 ;
      RECT 55.09 6.655 55.44 6.885 ;
      RECT 50.33 6.655 50.895 6.885 ;
      RECT 50.16 6.685 55.44 6.855 ;
      RECT 54.315 2.365 54.635 2.685 ;
      RECT 54.285 2.365 54.635 2.595 ;
      RECT 54.115 2.395 54.635 2.565 ;
      RECT 54.315 6.225 54.635 6.545 ;
      RECT 54.285 6.285 54.635 6.515 ;
      RECT 54.115 6.315 54.635 6.485 ;
      RECT 50.155 3.255 50.345 3.925 ;
      RECT 50.095 3.665 50.135 3.925 ;
      RECT 51.465 2.89 51.475 3.111 ;
      RECT 51.395 2.885 51.465 3.236 ;
      RECT 51.385 2.885 51.395 3.36 ;
      RECT 51.355 2.885 51.385 3.41 ;
      RECT 51.335 2.885 51.355 3.485 ;
      RECT 51.315 2.885 51.335 3.555 ;
      RECT 51.285 2.885 51.315 3.595 ;
      RECT 51.275 2.885 51.285 3.615 ;
      RECT 51.265 2.885 51.275 3.626 ;
      RECT 51.255 3.135 51.265 3.628 ;
      RECT 51.245 3.2 51.255 3.63 ;
      RECT 51.235 3.295 51.245 3.632 ;
      RECT 51.225 3.37 51.235 3.634 ;
      RECT 51.175 3.394 51.225 3.64 ;
      RECT 51.135 3.429 51.175 3.649 ;
      RECT 51.125 3.445 51.135 3.654 ;
      RECT 51.111 3.45 51.125 3.657 ;
      RECT 51.025 3.49 51.111 3.668 ;
      RECT 50.945 3.533 51.025 3.686 ;
      RECT 50.925 3.543 50.945 3.697 ;
      RECT 50.895 3.551 50.925 3.702 ;
      RECT 50.875 3.561 50.895 3.707 ;
      RECT 50.851 3.567 50.875 3.712 ;
      RECT 50.765 3.577 50.851 3.725 ;
      RECT 50.687 3.583 50.765 3.745 ;
      RECT 50.601 3.578 50.687 3.764 ;
      RECT 50.515 3.574 50.601 3.785 ;
      RECT 50.435 3.57 50.515 3.8 ;
      RECT 50.365 3.566 50.435 3.831 ;
      RECT 50.355 3.277 50.365 3.345 ;
      RECT 50.355 3.555 50.365 3.861 ;
      RECT 50.345 3.262 50.355 3.49 ;
      RECT 50.345 3.535 50.355 3.925 ;
      RECT 50.135 3.285 50.155 3.925 ;
      RECT 50.935 2.605 50.945 3.345 ;
      RECT 50.755 3.125 50.775 3.345 ;
      RECT 50.765 3.115 50.775 3.345 ;
      RECT 51.265 2.155 51.305 2.415 ;
      RECT 51.255 2.155 51.265 2.425 ;
      RECT 51.221 2.155 51.255 2.452 ;
      RECT 51.135 2.155 51.221 2.512 ;
      RECT 51.115 2.155 51.135 2.575 ;
      RECT 51.055 2.155 51.115 2.74 ;
      RECT 51.045 2.155 51.055 2.9 ;
      RECT 51.015 2.346 51.045 2.995 ;
      RECT 51.005 2.401 51.015 3.095 ;
      RECT 50.995 2.43 51.005 3.14 ;
      RECT 50.985 2.455 50.995 3.173 ;
      RECT 50.975 2.49 50.985 3.228 ;
      RECT 50.955 2.535 50.975 3.29 ;
      RECT 50.945 2.58 50.955 3.34 ;
      RECT 50.925 2.64 50.935 3.345 ;
      RECT 50.915 2.67 50.925 3.345 ;
      RECT 50.895 2.7 50.915 3.345 ;
      RECT 50.845 2.805 50.895 3.345 ;
      RECT 50.835 2.9 50.845 3.345 ;
      RECT 50.825 2.93 50.835 3.345 ;
      RECT 50.8 2.98 50.825 3.345 ;
      RECT 50.795 3.035 50.8 3.345 ;
      RECT 50.775 3.06 50.795 3.345 ;
      RECT 50.735 3.14 50.755 3.335 ;
      RECT 50.485 2.725 50.555 2.935 ;
      RECT 47.725 2.635 47.985 2.895 ;
      RECT 50.555 2.73 50.565 2.93 ;
      RECT 50.441 2.723 50.485 2.935 ;
      RECT 50.355 2.716 50.441 2.935 ;
      RECT 50.335 2.711 50.355 2.925 ;
      RECT 50.325 2.709 50.335 2.905 ;
      RECT 50.275 2.706 50.325 2.9 ;
      RECT 50.245 2.702 50.275 2.895 ;
      RECT 50.225 2.7 50.245 2.89 ;
      RECT 50.185 2.697 50.225 2.885 ;
      RECT 50.115 2.691 50.185 2.88 ;
      RECT 50.085 2.686 50.115 2.875 ;
      RECT 50.065 2.684 50.085 2.87 ;
      RECT 50.035 2.681 50.065 2.865 ;
      RECT 49.975 2.677 50.035 2.86 ;
      RECT 49.905 2.675 49.975 2.85 ;
      RECT 49.871 2.673 49.905 2.843 ;
      RECT 49.785 2.668 49.871 2.835 ;
      RECT 49.751 2.662 49.785 2.827 ;
      RECT 49.665 2.652 49.751 2.819 ;
      RECT 49.631 2.643 49.665 2.811 ;
      RECT 49.545 2.638 49.631 2.803 ;
      RECT 49.475 2.635 49.545 2.793 ;
      RECT 49.455 2.63 49.475 2.787 ;
      RECT 49.451 2.625 49.455 2.786 ;
      RECT 49.365 2.621 49.451 2.781 ;
      RECT 49.325 2.616 49.365 2.774 ;
      RECT 49.245 2.615 49.325 2.769 ;
      RECT 49.225 2.615 49.245 2.766 ;
      RECT 49.199 2.615 49.225 2.766 ;
      RECT 49.113 2.617 49.199 2.77 ;
      RECT 49.027 2.619 49.113 2.777 ;
      RECT 48.941 2.621 49.027 2.783 ;
      RECT 48.855 2.624 48.941 2.79 ;
      RECT 48.821 2.626 48.855 2.795 ;
      RECT 48.735 2.631 48.821 2.8 ;
      RECT 48.711 2.626 48.735 2.804 ;
      RECT 48.625 2.631 48.711 2.809 ;
      RECT 48.587 2.636 48.625 2.814 ;
      RECT 48.501 2.639 48.587 2.819 ;
      RECT 48.415 2.643 48.501 2.826 ;
      RECT 48.351 2.645 48.415 2.832 ;
      RECT 48.265 2.645 48.351 2.838 ;
      RECT 48.181 2.646 48.265 2.845 ;
      RECT 48.095 2.649 48.181 2.852 ;
      RECT 48.071 2.651 48.095 2.856 ;
      RECT 47.985 2.653 48.071 2.861 ;
      RECT 47.715 2.67 47.725 2.865 ;
      RECT 49.9 7.765 50.19 7.995 ;
      RECT 49.96 7.025 50.13 7.995 ;
      RECT 49.85 7.055 50.225 7.425 ;
      RECT 49.9 7.025 50.19 7.425 ;
      RECT 49.955 2.247 50.145 2.455 ;
      RECT 49.945 2.252 50.155 2.45 ;
      RECT 49.935 2.233 49.945 2.445 ;
      RECT 49.905 2.228 49.935 2.44 ;
      RECT 49.865 2.252 50.155 2.43 ;
      RECT 49.645 2.165 49.905 2.425 ;
      RECT 49.945 2.236 49.955 2.45 ;
      RECT 49.645 2.245 50.135 2.425 ;
      RECT 49.645 2.241 49.995 2.425 ;
      RECT 49.595 3.155 49.645 3.435 ;
      RECT 49.525 3.125 49.555 3.435 ;
      RECT 49.665 3.155 49.725 3.415 ;
      RECT 49.525 3.115 49.545 3.435 ;
      RECT 49.645 3.155 49.665 3.425 ;
      RECT 49.565 3.145 49.595 3.435 ;
      RECT 49.555 3.13 49.565 3.435 ;
      RECT 49.505 3.105 49.525 3.435 ;
      RECT 49.475 3.09 49.505 3.435 ;
      RECT 49.465 3.08 49.475 3.435 ;
      RECT 49.445 3.069 49.465 3.43 ;
      RECT 49.425 3.057 49.445 3.4 ;
      RECT 49.415 3.048 49.425 3.383 ;
      RECT 49.385 3.03 49.415 3.375 ;
      RECT 49.375 2.995 49.385 3.367 ;
      RECT 49.365 2.975 49.375 3.36 ;
      RECT 49.355 2.955 49.365 3.353 ;
      RECT 49.345 2.94 49.355 3.348 ;
      RECT 49.335 2.92 49.345 3.343 ;
      RECT 49.325 2.915 49.335 3.338 ;
      RECT 49.321 2.905 49.325 3.334 ;
      RECT 49.235 2.905 49.321 3.309 ;
      RECT 49.205 2.905 49.235 3.275 ;
      RECT 49.195 2.905 49.205 3.255 ;
      RECT 49.135 2.905 49.195 3.2 ;
      RECT 49.125 2.92 49.135 3.145 ;
      RECT 49.115 2.93 49.125 3.125 ;
      RECT 49.065 3.665 49.325 3.925 ;
      RECT 48.985 3.685 49.325 3.901 ;
      RECT 48.965 3.685 49.325 3.896 ;
      RECT 48.941 3.685 49.325 3.894 ;
      RECT 48.855 3.685 49.325 3.889 ;
      RECT 48.705 3.625 48.965 3.885 ;
      RECT 48.665 3.68 48.985 3.88 ;
      RECT 48.655 3.69 49.325 3.875 ;
      RECT 48.675 3.675 48.965 3.885 ;
      RECT 48.565 2.115 48.825 2.375 ;
      RECT 48.565 2.2 48.835 2.3 ;
      RECT 47.735 3.63 47.755 3.874 ;
      RECT 47.735 3.63 47.805 3.869 ;
      RECT 47.715 3.635 47.805 3.868 ;
      RECT 47.705 3.65 47.891 3.858 ;
      RECT 47.705 3.65 47.965 3.855 ;
      RECT 47.7 3.687 47.975 3.845 ;
      RECT 47.7 3.687 48.061 3.841 ;
      RECT 47.7 3.687 48.075 3.827 ;
      RECT 47.975 3.565 48.235 3.825 ;
      RECT 47.695 3.692 48.235 3.82 ;
      RECT 47.685 3.74 48.235 3.795 ;
      RECT 47.955 3.605 47.975 3.854 ;
      RECT 47.891 3.609 47.955 3.857 ;
      RECT 47.755 3.622 48.235 3.825 ;
      RECT 47.805 3.616 47.891 3.862 ;
      RECT 47.205 2.475 47.215 2.645 ;
      RECT 47.265 2.435 47.275 2.615 ;
      RECT 47.565 2.245 47.575 2.455 ;
      RECT 47.895 2.095 48.145 2.355 ;
      RECT 47.885 2.095 47.895 2.357 ;
      RECT 47.875 2.155 47.885 2.361 ;
      RECT 47.845 2.157 47.875 2.369 ;
      RECT 47.815 2.162 47.845 2.383 ;
      RECT 47.805 2.166 47.815 2.393 ;
      RECT 47.775 2.171 47.805 2.405 ;
      RECT 47.745 2.18 47.775 2.406 ;
      RECT 47.675 2.19 47.745 2.41 ;
      RECT 47.635 2.195 47.675 2.414 ;
      RECT 47.615 2.195 47.635 2.425 ;
      RECT 47.605 2.2 47.615 2.435 ;
      RECT 47.595 2.21 47.605 2.438 ;
      RECT 47.585 2.23 47.595 2.443 ;
      RECT 47.575 2.24 47.585 2.445 ;
      RECT 47.545 2.255 47.565 2.462 ;
      RECT 47.535 2.267 47.545 2.472 ;
      RECT 47.525 2.273 47.535 2.475 ;
      RECT 47.491 2.286 47.525 2.485 ;
      RECT 47.405 2.32 47.491 2.518 ;
      RECT 47.385 2.355 47.405 2.547 ;
      RECT 47.365 2.37 47.385 2.559 ;
      RECT 47.345 2.38 47.365 2.571 ;
      RECT 47.295 2.399 47.345 2.591 ;
      RECT 47.285 2.416 47.295 2.605 ;
      RECT 47.275 2.422 47.285 2.61 ;
      RECT 47.255 2.44 47.265 2.618 ;
      RECT 47.245 2.445 47.255 2.625 ;
      RECT 47.235 2.456 47.245 2.632 ;
      RECT 47.215 2.461 47.235 2.64 ;
      RECT 47.195 2.475 47.205 2.65 ;
      RECT 47.185 2.48 47.195 2.66 ;
      RECT 47.155 2.494 47.185 2.67 ;
      RECT 47.145 2.507 47.155 2.68 ;
      RECT 47.065 2.538 47.145 2.705 ;
      RECT 47.045 2.568 47.065 2.73 ;
      RECT 47.035 2.573 47.045 2.737 ;
      RECT 47.005 2.585 47.035 2.743 ;
      RECT 46.995 2.6 47.005 2.749 ;
      RECT 46.985 2.605 46.995 2.752 ;
      RECT 46.965 2.615 46.985 2.756 ;
      RECT 46.945 2.62 46.965 2.762 ;
      RECT 46.915 2.625 46.945 2.77 ;
      RECT 46.885 2.63 46.915 2.78 ;
      RECT 46.855 2.64 46.885 2.789 ;
      RECT 46.815 2.645 46.855 2.797 ;
      RECT 46.765 2.638 46.815 2.809 ;
      RECT 46.745 2.629 46.765 2.82 ;
      RECT 46.735 2.626 46.745 2.825 ;
      RECT 46.695 2.625 46.735 2.826 ;
      RECT 46.685 2.61 46.695 2.827 ;
      RECT 46.657 2.595 46.685 2.828 ;
      RECT 46.571 2.595 46.657 2.83 ;
      RECT 46.485 2.595 46.571 2.834 ;
      RECT 46.465 2.595 46.485 2.83 ;
      RECT 46.455 2.605 46.465 2.823 ;
      RECT 46.445 2.62 46.455 2.818 ;
      RECT 46.435 2.625 46.445 2.795 ;
      RECT 47.915 3.13 47.925 3.33 ;
      RECT 47.865 3.125 47.915 3.35 ;
      RECT 47.855 3.125 47.865 3.37 ;
      RECT 47.811 3.125 47.855 3.374 ;
      RECT 47.725 3.125 47.811 3.371 ;
      RECT 47.665 3.135 47.725 3.368 ;
      RECT 47.605 3.149 47.665 3.366 ;
      RECT 47.595 3.154 47.605 3.364 ;
      RECT 47.585 3.16 47.595 3.363 ;
      RECT 47.515 3.173 47.585 3.359 ;
      RECT 47.467 3.187 47.515 3.36 ;
      RECT 47.381 3.203 47.467 3.372 ;
      RECT 47.295 3.224 47.381 3.388 ;
      RECT 47.275 3.235 47.295 3.398 ;
      RECT 47.195 3.245 47.275 3.408 ;
      RECT 47.161 3.259 47.195 3.42 ;
      RECT 47.075 3.274 47.161 3.435 ;
      RECT 47.045 3.29 47.075 3.445 ;
      RECT 46.99 3.305 47.045 3.456 ;
      RECT 46.945 3.323 46.99 3.476 ;
      RECT 46.891 3.342 46.945 3.496 ;
      RECT 46.805 3.368 46.891 3.523 ;
      RECT 46.785 3.39 46.805 3.543 ;
      RECT 46.725 3.405 46.785 3.559 ;
      RECT 46.715 3.42 46.725 3.573 ;
      RECT 46.695 3.425 46.715 3.579 ;
      RECT 46.665 3.438 46.695 3.589 ;
      RECT 46.645 3.443 46.665 3.598 ;
      RECT 46.635 3.45 46.645 3.603 ;
      RECT 46.625 3.455 46.635 3.606 ;
      RECT 46.585 3.465 46.625 3.615 ;
      RECT 46.56 3.48 46.585 3.627 ;
      RECT 46.515 3.495 46.56 3.639 ;
      RECT 46.495 3.507 46.515 3.651 ;
      RECT 46.465 3.512 46.495 3.661 ;
      RECT 46.445 3.519 46.465 3.671 ;
      RECT 46.435 3.525 46.445 3.68 ;
      RECT 46.411 3.532 46.435 3.69 ;
      RECT 46.325 3.554 46.411 3.71 ;
      RECT 46.315 3.573 46.325 3.725 ;
      RECT 46.291 3.58 46.315 3.731 ;
      RECT 46.205 3.602 46.291 3.756 ;
      RECT 46.165 3.627 46.205 3.783 ;
      RECT 46.155 3.636 46.165 3.793 ;
      RECT 46.105 3.646 46.155 3.802 ;
      RECT 46.085 3.66 46.105 3.812 ;
      RECT 46.055 3.67 46.085 3.817 ;
      RECT 46.045 3.675 46.055 3.82 ;
      RECT 45.971 3.677 46.045 3.827 ;
      RECT 45.885 3.681 45.971 3.839 ;
      RECT 45.875 3.684 45.885 3.845 ;
      RECT 45.615 3.635 45.875 3.895 ;
      RECT 47.145 3.705 47.335 3.915 ;
      RECT 47.135 3.71 47.345 3.91 ;
      RECT 47.125 3.71 47.345 3.875 ;
      RECT 47.045 3.595 47.305 3.855 ;
      RECT 45.955 3.125 46.145 3.425 ;
      RECT 45.945 3.125 46.145 3.42 ;
      RECT 45.935 3.125 46.155 3.415 ;
      RECT 45.925 3.125 46.155 3.41 ;
      RECT 45.925 3.125 46.185 3.385 ;
      RECT 45.885 2.165 46.145 2.425 ;
      RECT 45.695 2.09 45.781 2.423 ;
      RECT 45.695 2.09 45.825 2.419 ;
      RECT 45.675 2.094 45.835 2.418 ;
      RECT 45.825 2.085 45.835 2.418 ;
      RECT 45.695 2.09 45.845 2.417 ;
      RECT 45.675 2.1 45.885 2.416 ;
      RECT 45.665 2.095 45.845 2.408 ;
      RECT 45.655 2.11 45.885 2.315 ;
      RECT 45.655 2.16 46.085 2.315 ;
      RECT 45.655 2.15 46.065 2.315 ;
      RECT 45.655 2.14 46.035 2.315 ;
      RECT 45.655 2.13 45.975 2.315 ;
      RECT 45.655 2.115 45.955 2.315 ;
      RECT 45.781 2.086 45.835 2.418 ;
      RECT 44.855 2.745 44.995 3.035 ;
      RECT 45.115 2.768 45.125 2.955 ;
      RECT 45.815 2.665 45.995 2.895 ;
      RECT 45.815 2.665 46.005 2.885 ;
      RECT 46.025 2.67 46.035 2.875 ;
      RECT 46.005 2.665 46.025 2.88 ;
      RECT 45.765 2.669 45.815 2.895 ;
      RECT 45.755 2.674 45.765 2.895 ;
      RECT 45.721 2.679 45.755 2.896 ;
      RECT 45.635 2.694 45.721 2.898 ;
      RECT 45.621 2.706 45.635 2.901 ;
      RECT 45.535 2.716 45.621 2.903 ;
      RECT 45.511 2.726 45.535 2.905 ;
      RECT 45.425 2.737 45.511 2.905 ;
      RECT 45.395 2.747 45.425 2.905 ;
      RECT 45.365 2.752 45.395 2.908 ;
      RECT 45.345 2.757 45.365 2.913 ;
      RECT 45.325 2.762 45.345 2.915 ;
      RECT 45.275 2.77 45.325 2.915 ;
      RECT 45.255 2.774 45.275 2.915 ;
      RECT 45.235 2.773 45.255 2.92 ;
      RECT 45.175 2.771 45.235 2.935 ;
      RECT 45.125 2.769 45.175 2.95 ;
      RECT 45.035 2.766 45.115 3.035 ;
      RECT 45.005 2.76 45.035 3.035 ;
      RECT 44.995 2.75 45.005 3.035 ;
      RECT 44.805 2.745 44.855 2.96 ;
      RECT 44.795 2.75 44.805 2.95 ;
      RECT 45.035 3.225 45.295 3.485 ;
      RECT 45.035 3.225 45.325 3.375 ;
      RECT 45.035 3.225 45.365 3.36 ;
      RECT 45.295 3.145 45.485 3.355 ;
      RECT 45.295 3.15 45.495 3.345 ;
      RECT 45.245 3.22 45.495 3.345 ;
      RECT 45.275 3.155 45.295 3.485 ;
      RECT 45.265 3.18 45.495 3.345 ;
      RECT 44.445 3.125 44.455 3.355 ;
      RECT 44.345 2.245 44.415 3.355 ;
      RECT 45.085 2.355 45.345 2.615 ;
      RECT 44.785 2.405 44.915 2.565 ;
      RECT 45.001 2.412 45.085 2.565 ;
      RECT 44.915 2.407 45.001 2.565 ;
      RECT 44.725 2.405 44.785 2.575 ;
      RECT 44.695 2.403 44.725 2.59 ;
      RECT 44.675 2.401 44.695 2.6 ;
      RECT 44.665 2.399 44.675 2.605 ;
      RECT 44.645 2.398 44.665 2.615 ;
      RECT 44.635 2.396 44.645 2.62 ;
      RECT 44.615 2.395 44.635 2.625 ;
      RECT 44.595 2.39 44.615 2.63 ;
      RECT 44.565 2.376 44.595 2.64 ;
      RECT 44.525 2.355 44.565 2.655 ;
      RECT 44.515 2.34 44.525 2.665 ;
      RECT 44.495 2.331 44.515 2.675 ;
      RECT 44.485 2.322 44.495 2.695 ;
      RECT 44.475 2.317 44.485 2.755 ;
      RECT 44.455 2.311 44.475 2.84 ;
      RECT 44.455 3.15 44.465 3.35 ;
      RECT 44.445 2.306 44.455 3.07 ;
      RECT 44.435 2.28 44.445 3.355 ;
      RECT 44.415 2.25 44.435 3.355 ;
      RECT 44.325 2.245 44.345 2.58 ;
      RECT 44.335 2.68 44.345 3.355 ;
      RECT 44.325 2.72 44.335 3.355 ;
      RECT 44.295 2.245 44.325 2.525 ;
      RECT 44.305 2.81 44.325 3.355 ;
      RECT 44.29 2.915 44.305 3.355 ;
      RECT 44.265 2.245 44.295 2.48 ;
      RECT 44.285 2.947 44.29 3.355 ;
      RECT 44.265 3.05 44.285 3.355 ;
      RECT 44.255 2.245 44.265 2.47 ;
      RECT 44.255 3.12 44.265 3.35 ;
      RECT 44.235 2.245 44.255 2.46 ;
      RECT 44.225 2.25 44.235 2.45 ;
      RECT 44.435 3.525 44.455 3.765 ;
      RECT 43.755 3.455 43.835 3.725 ;
      RECT 43.665 3.455 43.675 3.665 ;
      RECT 44.945 3.525 44.955 3.725 ;
      RECT 44.865 3.515 44.945 3.75 ;
      RECT 44.861 3.515 44.865 3.776 ;
      RECT 44.775 3.515 44.861 3.786 ;
      RECT 44.755 3.515 44.775 3.794 ;
      RECT 44.731 3.516 44.755 3.792 ;
      RECT 44.645 3.521 44.731 3.787 ;
      RECT 44.627 3.525 44.645 3.781 ;
      RECT 44.541 3.525 44.627 3.777 ;
      RECT 44.455 3.525 44.541 3.769 ;
      RECT 44.351 3.525 44.435 3.762 ;
      RECT 44.265 3.525 44.351 3.756 ;
      RECT 44.205 3.52 44.265 3.75 ;
      RECT 44.177 3.514 44.205 3.747 ;
      RECT 44.091 3.511 44.177 3.744 ;
      RECT 44.005 3.507 44.091 3.738 ;
      RECT 43.96 3.495 44.005 3.734 ;
      RECT 43.935 3.48 43.96 3.732 ;
      RECT 43.895 3.465 43.935 3.73 ;
      RECT 43.835 3.455 43.895 3.727 ;
      RECT 43.745 3.455 43.755 3.72 ;
      RECT 43.73 3.455 43.745 3.71 ;
      RECT 43.675 3.455 43.73 3.685 ;
      RECT 43.655 3.47 43.665 3.66 ;
      RECT 43.785 2.635 44.045 2.895 ;
      RECT 43.785 2.645 44.065 2.855 ;
      RECT 43.785 2.65 44.075 2.85 ;
      RECT 41.765 2.115 42.025 2.375 ;
      RECT 41.755 2.145 42.025 2.355 ;
      RECT 43.685 2.055 43.935 2.315 ;
      RECT 43.675 2.055 43.685 2.316 ;
      RECT 43.645 2.14 43.675 2.318 ;
      RECT 43.635 2.145 43.645 2.32 ;
      RECT 43.575 2.16 43.635 2.326 ;
      RECT 43.545 2.18 43.575 2.333 ;
      RECT 43.515 2.191 43.545 2.34 ;
      RECT 43.495 2.201 43.515 2.345 ;
      RECT 43.477 2.204 43.495 2.344 ;
      RECT 43.391 2.203 43.477 2.344 ;
      RECT 43.305 2.2 43.391 2.343 ;
      RECT 43.219 2.197 43.305 2.342 ;
      RECT 43.133 2.194 43.219 2.342 ;
      RECT 43.047 2.192 43.133 2.341 ;
      RECT 42.961 2.189 43.047 2.34 ;
      RECT 42.875 2.186 42.961 2.34 ;
      RECT 42.857 2.185 42.875 2.339 ;
      RECT 42.771 2.184 42.857 2.339 ;
      RECT 42.685 2.182 42.771 2.338 ;
      RECT 42.599 2.181 42.685 2.338 ;
      RECT 42.513 2.18 42.599 2.337 ;
      RECT 42.427 2.178 42.513 2.337 ;
      RECT 42.341 2.177 42.427 2.336 ;
      RECT 42.255 2.175 42.341 2.336 ;
      RECT 42.231 2.174 42.255 2.335 ;
      RECT 42.145 2.169 42.231 2.335 ;
      RECT 42.111 2.162 42.145 2.335 ;
      RECT 42.025 2.152 42.111 2.335 ;
      RECT 41.745 2.15 41.755 2.35 ;
      RECT 43.025 3.205 43.285 3.465 ;
      RECT 43.025 3.205 43.365 3.251 ;
      RECT 43.165 3.185 43.375 3.24 ;
      RECT 43.225 3.16 43.435 3.2 ;
      RECT 43.235 3.155 43.435 3.2 ;
      RECT 43.245 3.13 43.435 3.2 ;
      RECT 43.305 2.96 43.355 3.29 ;
      RECT 43.255 3.09 43.445 3.15 ;
      RECT 43.295 3.016 43.305 3.329 ;
      RECT 43.255 3.09 43.475 3.125 ;
      RECT 43.255 3.09 43.495 3.1 ;
      RECT 43.365 2.89 43.555 3.095 ;
      RECT 43.355 2.9 43.565 3.09 ;
      RECT 43.275 3.063 43.565 3.09 ;
      RECT 43.285 3.039 43.295 3.345 ;
      RECT 43.375 2.885 43.545 3.095 ;
      RECT 42.665 2.675 42.855 2.885 ;
      RECT 41.235 2.605 41.495 2.865 ;
      RECT 41.585 2.595 41.685 2.805 ;
      RECT 41.535 2.615 41.575 2.805 ;
      RECT 42.855 2.685 42.865 2.88 ;
      RECT 42.655 2.685 42.665 2.88 ;
      RECT 42.635 2.7 42.655 2.87 ;
      RECT 42.625 2.71 42.635 2.865 ;
      RECT 42.585 2.71 42.625 2.863 ;
      RECT 42.561 2.704 42.585 2.86 ;
      RECT 42.475 2.699 42.561 2.857 ;
      RECT 42.415 2.695 42.475 2.852 ;
      RECT 42.381 2.692 42.415 2.849 ;
      RECT 42.295 2.682 42.381 2.845 ;
      RECT 42.291 2.675 42.295 2.842 ;
      RECT 42.205 2.67 42.291 2.84 ;
      RECT 42.177 2.663 42.205 2.836 ;
      RECT 42.091 2.658 42.177 2.833 ;
      RECT 42.005 2.649 42.091 2.828 ;
      RECT 41.995 2.644 42.005 2.825 ;
      RECT 41.981 2.643 41.995 2.825 ;
      RECT 41.895 2.639 41.981 2.82 ;
      RECT 41.875 2.633 41.895 2.816 ;
      RECT 41.815 2.628 41.875 2.815 ;
      RECT 41.785 2.62 41.815 2.815 ;
      RECT 41.775 2.605 41.785 2.815 ;
      RECT 41.771 2.595 41.775 2.814 ;
      RECT 41.685 2.595 41.771 2.81 ;
      RECT 41.575 2.605 41.585 2.805 ;
      RECT 41.505 2.615 41.535 2.8 ;
      RECT 41.495 2.615 41.505 2.8 ;
      RECT 42.415 3.115 42.675 3.375 ;
      RECT 42.345 3.125 42.675 3.335 ;
      RECT 42.335 3.13 42.675 3.33 ;
      RECT 41.755 3.115 42.015 3.375 ;
      RECT 41.755 3.16 42.125 3.365 ;
      RECT 41.755 3.155 42.115 3.365 ;
      RECT 40.665 3.322 40.845 3.765 ;
      RECT 40.655 3.322 40.845 3.763 ;
      RECT 40.655 3.337 40.855 3.76 ;
      RECT 40.645 2.26 40.775 3.758 ;
      RECT 40.645 3.385 40.915 3.645 ;
      RECT 40.645 3.36 40.865 3.645 ;
      RECT 40.645 3.295 40.835 3.758 ;
      RECT 40.645 3.255 40.805 3.758 ;
      RECT 40.645 3.21 40.795 3.758 ;
      RECT 40.645 3.15 40.785 3.758 ;
      RECT 40.635 2.545 40.775 3.2 ;
      RECT 40.675 2.245 40.785 3.065 ;
      RECT 40.645 2.26 40.825 2.52 ;
      RECT 40.645 2.26 40.835 2.47 ;
      RECT 40.675 2.245 40.845 2.463 ;
      RECT 40.665 2.247 40.855 2.458 ;
      RECT 40.655 2.252 40.865 2.45 ;
      RECT 39.515 7.77 39.805 8 ;
      RECT 39.575 6.29 39.745 8 ;
      RECT 39.565 6.66 39.92 7.015 ;
      RECT 39.515 6.29 39.805 6.52 ;
      RECT 39.11 2.395 39.215 2.965 ;
      RECT 39.11 2.73 39.435 2.96 ;
      RECT 39.11 2.76 39.605 2.93 ;
      RECT 39.11 2.395 39.3 2.96 ;
      RECT 38.525 2.36 38.815 2.59 ;
      RECT 38.525 2.395 39.3 2.565 ;
      RECT 38.585 0.88 38.755 2.59 ;
      RECT 38.525 0.88 38.815 1.11 ;
      RECT 38.525 7.77 38.815 8 ;
      RECT 38.585 6.29 38.755 8 ;
      RECT 38.525 6.29 38.815 6.52 ;
      RECT 38.525 6.325 39.38 6.485 ;
      RECT 39.21 5.92 39.38 6.485 ;
      RECT 38.525 6.32 38.92 6.485 ;
      RECT 39.145 5.92 39.435 6.15 ;
      RECT 39.145 5.95 39.605 6.12 ;
      RECT 38.155 2.73 38.445 2.96 ;
      RECT 38.155 2.76 38.615 2.93 ;
      RECT 38.22 1.655 38.385 2.96 ;
      RECT 36.735 1.625 37.025 1.855 ;
      RECT 36.735 1.655 38.385 1.825 ;
      RECT 36.795 0.885 36.965 1.855 ;
      RECT 36.735 0.885 37.025 1.115 ;
      RECT 36.735 7.765 37.025 7.995 ;
      RECT 36.795 7.025 36.965 7.995 ;
      RECT 36.795 7.12 38.385 7.29 ;
      RECT 38.215 5.92 38.385 7.29 ;
      RECT 36.735 7.025 37.025 7.255 ;
      RECT 38.155 5.92 38.445 6.15 ;
      RECT 38.155 5.95 38.615 6.12 ;
      RECT 34.77 3.43 35.12 3.78 ;
      RECT 34.86 2.025 35.03 3.78 ;
      RECT 37.165 1.965 37.515 2.315 ;
      RECT 34.86 2.025 36.48 2.2 ;
      RECT 34.86 2.025 37.515 2.195 ;
      RECT 37.19 6.655 37.515 6.98 ;
      RECT 32.615 6.61 32.965 6.96 ;
      RECT 37.165 6.655 37.515 6.885 ;
      RECT 32.405 6.655 32.965 6.885 ;
      RECT 32.235 6.685 37.515 6.855 ;
      RECT 36.39 2.365 36.71 2.685 ;
      RECT 36.36 2.365 36.71 2.595 ;
      RECT 36.19 2.395 36.71 2.565 ;
      RECT 36.39 6.225 36.71 6.545 ;
      RECT 36.36 6.285 36.71 6.515 ;
      RECT 36.19 6.315 36.71 6.485 ;
      RECT 32.23 3.255 32.42 3.925 ;
      RECT 32.17 3.665 32.21 3.925 ;
      RECT 33.54 2.89 33.55 3.111 ;
      RECT 33.47 2.885 33.54 3.236 ;
      RECT 33.46 2.885 33.47 3.36 ;
      RECT 33.43 2.885 33.46 3.41 ;
      RECT 33.41 2.885 33.43 3.485 ;
      RECT 33.39 2.885 33.41 3.555 ;
      RECT 33.36 2.885 33.39 3.595 ;
      RECT 33.35 2.885 33.36 3.615 ;
      RECT 33.34 2.885 33.35 3.626 ;
      RECT 33.33 3.135 33.34 3.628 ;
      RECT 33.32 3.2 33.33 3.63 ;
      RECT 33.31 3.295 33.32 3.632 ;
      RECT 33.3 3.37 33.31 3.634 ;
      RECT 33.25 3.394 33.3 3.64 ;
      RECT 33.21 3.429 33.25 3.649 ;
      RECT 33.2 3.445 33.21 3.654 ;
      RECT 33.186 3.45 33.2 3.657 ;
      RECT 33.1 3.49 33.186 3.668 ;
      RECT 33.02 3.533 33.1 3.686 ;
      RECT 33 3.543 33.02 3.697 ;
      RECT 32.97 3.551 33 3.702 ;
      RECT 32.95 3.561 32.97 3.707 ;
      RECT 32.926 3.567 32.95 3.712 ;
      RECT 32.84 3.577 32.926 3.725 ;
      RECT 32.762 3.583 32.84 3.745 ;
      RECT 32.676 3.578 32.762 3.764 ;
      RECT 32.59 3.574 32.676 3.785 ;
      RECT 32.51 3.57 32.59 3.8 ;
      RECT 32.44 3.566 32.51 3.831 ;
      RECT 32.43 3.277 32.44 3.345 ;
      RECT 32.43 3.555 32.44 3.861 ;
      RECT 32.42 3.262 32.43 3.49 ;
      RECT 32.42 3.535 32.43 3.925 ;
      RECT 32.21 3.285 32.23 3.925 ;
      RECT 33.01 2.605 33.02 3.345 ;
      RECT 32.83 3.125 32.85 3.345 ;
      RECT 32.84 3.115 32.85 3.345 ;
      RECT 33.34 2.155 33.38 2.415 ;
      RECT 33.33 2.155 33.34 2.425 ;
      RECT 33.296 2.155 33.33 2.452 ;
      RECT 33.21 2.155 33.296 2.512 ;
      RECT 33.19 2.155 33.21 2.575 ;
      RECT 33.13 2.155 33.19 2.74 ;
      RECT 33.12 2.155 33.13 2.9 ;
      RECT 33.09 2.346 33.12 2.995 ;
      RECT 33.08 2.401 33.09 3.095 ;
      RECT 33.07 2.43 33.08 3.14 ;
      RECT 33.06 2.455 33.07 3.173 ;
      RECT 33.05 2.49 33.06 3.228 ;
      RECT 33.03 2.535 33.05 3.29 ;
      RECT 33.02 2.58 33.03 3.34 ;
      RECT 33 2.64 33.01 3.345 ;
      RECT 32.99 2.67 33 3.345 ;
      RECT 32.97 2.7 32.99 3.345 ;
      RECT 32.92 2.805 32.97 3.345 ;
      RECT 32.91 2.9 32.92 3.345 ;
      RECT 32.9 2.93 32.91 3.345 ;
      RECT 32.875 2.98 32.9 3.345 ;
      RECT 32.87 3.035 32.875 3.345 ;
      RECT 32.85 3.06 32.87 3.345 ;
      RECT 32.81 3.14 32.83 3.335 ;
      RECT 32.56 2.725 32.63 2.935 ;
      RECT 29.8 2.635 30.06 2.895 ;
      RECT 32.63 2.73 32.64 2.93 ;
      RECT 32.516 2.723 32.56 2.935 ;
      RECT 32.43 2.716 32.516 2.935 ;
      RECT 32.41 2.711 32.43 2.925 ;
      RECT 32.4 2.709 32.41 2.905 ;
      RECT 32.35 2.706 32.4 2.9 ;
      RECT 32.32 2.702 32.35 2.895 ;
      RECT 32.3 2.7 32.32 2.89 ;
      RECT 32.26 2.697 32.3 2.885 ;
      RECT 32.19 2.691 32.26 2.88 ;
      RECT 32.16 2.686 32.19 2.875 ;
      RECT 32.14 2.684 32.16 2.87 ;
      RECT 32.11 2.681 32.14 2.865 ;
      RECT 32.05 2.677 32.11 2.86 ;
      RECT 31.98 2.675 32.05 2.85 ;
      RECT 31.946 2.673 31.98 2.843 ;
      RECT 31.86 2.668 31.946 2.835 ;
      RECT 31.826 2.662 31.86 2.827 ;
      RECT 31.74 2.652 31.826 2.819 ;
      RECT 31.706 2.643 31.74 2.811 ;
      RECT 31.62 2.638 31.706 2.803 ;
      RECT 31.55 2.635 31.62 2.793 ;
      RECT 31.53 2.63 31.55 2.787 ;
      RECT 31.526 2.625 31.53 2.786 ;
      RECT 31.44 2.621 31.526 2.781 ;
      RECT 31.4 2.616 31.44 2.774 ;
      RECT 31.32 2.615 31.4 2.769 ;
      RECT 31.3 2.615 31.32 2.766 ;
      RECT 31.274 2.615 31.3 2.766 ;
      RECT 31.188 2.617 31.274 2.77 ;
      RECT 31.102 2.619 31.188 2.777 ;
      RECT 31.016 2.621 31.102 2.783 ;
      RECT 30.93 2.624 31.016 2.79 ;
      RECT 30.896 2.626 30.93 2.795 ;
      RECT 30.81 2.631 30.896 2.8 ;
      RECT 30.786 2.626 30.81 2.804 ;
      RECT 30.7 2.631 30.786 2.809 ;
      RECT 30.662 2.636 30.7 2.814 ;
      RECT 30.576 2.639 30.662 2.819 ;
      RECT 30.49 2.643 30.576 2.826 ;
      RECT 30.426 2.645 30.49 2.832 ;
      RECT 30.34 2.645 30.426 2.838 ;
      RECT 30.256 2.646 30.34 2.845 ;
      RECT 30.17 2.649 30.256 2.852 ;
      RECT 30.146 2.651 30.17 2.856 ;
      RECT 30.06 2.653 30.146 2.861 ;
      RECT 29.79 2.67 29.8 2.865 ;
      RECT 31.975 7.765 32.265 7.995 ;
      RECT 32.035 7.025 32.205 7.995 ;
      RECT 31.925 7.055 32.3 7.425 ;
      RECT 31.975 7.025 32.265 7.425 ;
      RECT 32.03 2.247 32.22 2.455 ;
      RECT 32.02 2.252 32.23 2.45 ;
      RECT 32.01 2.233 32.02 2.445 ;
      RECT 31.98 2.228 32.01 2.44 ;
      RECT 31.94 2.252 32.23 2.43 ;
      RECT 31.72 2.165 31.98 2.425 ;
      RECT 32.02 2.236 32.03 2.45 ;
      RECT 31.72 2.245 32.21 2.425 ;
      RECT 31.72 2.241 32.07 2.425 ;
      RECT 31.67 3.155 31.72 3.435 ;
      RECT 31.6 3.125 31.63 3.435 ;
      RECT 31.74 3.155 31.8 3.415 ;
      RECT 31.6 3.115 31.62 3.435 ;
      RECT 31.72 3.155 31.74 3.425 ;
      RECT 31.64 3.145 31.67 3.435 ;
      RECT 31.63 3.13 31.64 3.435 ;
      RECT 31.58 3.105 31.6 3.435 ;
      RECT 31.55 3.09 31.58 3.435 ;
      RECT 31.54 3.08 31.55 3.435 ;
      RECT 31.52 3.069 31.54 3.43 ;
      RECT 31.5 3.057 31.52 3.4 ;
      RECT 31.49 3.048 31.5 3.383 ;
      RECT 31.46 3.03 31.49 3.375 ;
      RECT 31.45 2.995 31.46 3.367 ;
      RECT 31.44 2.975 31.45 3.36 ;
      RECT 31.43 2.955 31.44 3.353 ;
      RECT 31.42 2.94 31.43 3.348 ;
      RECT 31.41 2.92 31.42 3.343 ;
      RECT 31.4 2.915 31.41 3.338 ;
      RECT 31.396 2.905 31.4 3.334 ;
      RECT 31.31 2.905 31.396 3.309 ;
      RECT 31.28 2.905 31.31 3.275 ;
      RECT 31.27 2.905 31.28 3.255 ;
      RECT 31.21 2.905 31.27 3.2 ;
      RECT 31.2 2.92 31.21 3.145 ;
      RECT 31.19 2.93 31.2 3.125 ;
      RECT 31.14 3.665 31.4 3.925 ;
      RECT 31.06 3.685 31.4 3.901 ;
      RECT 31.04 3.685 31.4 3.896 ;
      RECT 31.016 3.685 31.4 3.894 ;
      RECT 30.93 3.685 31.4 3.889 ;
      RECT 30.78 3.625 31.04 3.885 ;
      RECT 30.74 3.68 31.06 3.88 ;
      RECT 30.73 3.69 31.4 3.875 ;
      RECT 30.75 3.675 31.04 3.885 ;
      RECT 30.64 2.115 30.9 2.375 ;
      RECT 30.64 2.2 30.91 2.3 ;
      RECT 29.81 3.63 29.83 3.874 ;
      RECT 29.81 3.63 29.88 3.869 ;
      RECT 29.79 3.635 29.88 3.868 ;
      RECT 29.78 3.65 29.966 3.858 ;
      RECT 29.78 3.65 30.04 3.855 ;
      RECT 29.775 3.687 30.05 3.845 ;
      RECT 29.775 3.687 30.136 3.841 ;
      RECT 29.775 3.687 30.15 3.827 ;
      RECT 30.05 3.565 30.31 3.825 ;
      RECT 29.77 3.692 30.31 3.82 ;
      RECT 29.76 3.74 30.31 3.795 ;
      RECT 30.03 3.605 30.05 3.854 ;
      RECT 29.966 3.609 30.03 3.857 ;
      RECT 29.83 3.622 30.31 3.825 ;
      RECT 29.88 3.616 29.966 3.862 ;
      RECT 29.28 2.475 29.29 2.645 ;
      RECT 29.34 2.435 29.35 2.615 ;
      RECT 29.64 2.245 29.65 2.455 ;
      RECT 29.97 2.095 30.22 2.355 ;
      RECT 29.96 2.095 29.97 2.357 ;
      RECT 29.95 2.155 29.96 2.361 ;
      RECT 29.92 2.157 29.95 2.369 ;
      RECT 29.89 2.162 29.92 2.383 ;
      RECT 29.88 2.166 29.89 2.393 ;
      RECT 29.85 2.171 29.88 2.405 ;
      RECT 29.82 2.18 29.85 2.406 ;
      RECT 29.75 2.19 29.82 2.41 ;
      RECT 29.71 2.195 29.75 2.414 ;
      RECT 29.69 2.195 29.71 2.425 ;
      RECT 29.68 2.2 29.69 2.435 ;
      RECT 29.67 2.21 29.68 2.438 ;
      RECT 29.66 2.23 29.67 2.443 ;
      RECT 29.65 2.24 29.66 2.445 ;
      RECT 29.62 2.255 29.64 2.462 ;
      RECT 29.61 2.267 29.62 2.472 ;
      RECT 29.6 2.273 29.61 2.475 ;
      RECT 29.566 2.286 29.6 2.485 ;
      RECT 29.48 2.32 29.566 2.518 ;
      RECT 29.46 2.355 29.48 2.547 ;
      RECT 29.44 2.37 29.46 2.559 ;
      RECT 29.42 2.38 29.44 2.571 ;
      RECT 29.37 2.399 29.42 2.591 ;
      RECT 29.36 2.416 29.37 2.605 ;
      RECT 29.35 2.422 29.36 2.61 ;
      RECT 29.33 2.44 29.34 2.618 ;
      RECT 29.32 2.445 29.33 2.625 ;
      RECT 29.31 2.456 29.32 2.632 ;
      RECT 29.29 2.461 29.31 2.64 ;
      RECT 29.27 2.475 29.28 2.65 ;
      RECT 29.26 2.48 29.27 2.66 ;
      RECT 29.23 2.494 29.26 2.67 ;
      RECT 29.22 2.507 29.23 2.68 ;
      RECT 29.14 2.538 29.22 2.705 ;
      RECT 29.12 2.568 29.14 2.73 ;
      RECT 29.11 2.573 29.12 2.737 ;
      RECT 29.08 2.585 29.11 2.743 ;
      RECT 29.07 2.6 29.08 2.749 ;
      RECT 29.06 2.605 29.07 2.752 ;
      RECT 29.04 2.615 29.06 2.756 ;
      RECT 29.02 2.62 29.04 2.762 ;
      RECT 28.99 2.625 29.02 2.77 ;
      RECT 28.96 2.63 28.99 2.78 ;
      RECT 28.93 2.64 28.96 2.789 ;
      RECT 28.89 2.645 28.93 2.797 ;
      RECT 28.84 2.638 28.89 2.809 ;
      RECT 28.82 2.629 28.84 2.82 ;
      RECT 28.81 2.626 28.82 2.825 ;
      RECT 28.77 2.625 28.81 2.826 ;
      RECT 28.76 2.61 28.77 2.827 ;
      RECT 28.732 2.595 28.76 2.828 ;
      RECT 28.646 2.595 28.732 2.83 ;
      RECT 28.56 2.595 28.646 2.834 ;
      RECT 28.54 2.595 28.56 2.83 ;
      RECT 28.53 2.605 28.54 2.823 ;
      RECT 28.52 2.62 28.53 2.818 ;
      RECT 28.51 2.625 28.52 2.795 ;
      RECT 29.99 3.13 30 3.33 ;
      RECT 29.94 3.125 29.99 3.35 ;
      RECT 29.93 3.125 29.94 3.37 ;
      RECT 29.886 3.125 29.93 3.374 ;
      RECT 29.8 3.125 29.886 3.371 ;
      RECT 29.74 3.135 29.8 3.368 ;
      RECT 29.68 3.149 29.74 3.366 ;
      RECT 29.67 3.154 29.68 3.364 ;
      RECT 29.66 3.16 29.67 3.363 ;
      RECT 29.59 3.173 29.66 3.359 ;
      RECT 29.542 3.187 29.59 3.36 ;
      RECT 29.456 3.203 29.542 3.372 ;
      RECT 29.37 3.224 29.456 3.388 ;
      RECT 29.35 3.235 29.37 3.398 ;
      RECT 29.27 3.245 29.35 3.408 ;
      RECT 29.236 3.259 29.27 3.42 ;
      RECT 29.15 3.274 29.236 3.435 ;
      RECT 29.12 3.29 29.15 3.445 ;
      RECT 29.065 3.305 29.12 3.456 ;
      RECT 29.02 3.323 29.065 3.476 ;
      RECT 28.966 3.342 29.02 3.496 ;
      RECT 28.88 3.368 28.966 3.523 ;
      RECT 28.86 3.39 28.88 3.543 ;
      RECT 28.8 3.405 28.86 3.559 ;
      RECT 28.79 3.42 28.8 3.573 ;
      RECT 28.77 3.425 28.79 3.579 ;
      RECT 28.74 3.438 28.77 3.589 ;
      RECT 28.72 3.443 28.74 3.598 ;
      RECT 28.71 3.45 28.72 3.603 ;
      RECT 28.7 3.455 28.71 3.606 ;
      RECT 28.66 3.465 28.7 3.615 ;
      RECT 28.635 3.48 28.66 3.627 ;
      RECT 28.59 3.495 28.635 3.639 ;
      RECT 28.57 3.507 28.59 3.651 ;
      RECT 28.54 3.512 28.57 3.661 ;
      RECT 28.52 3.519 28.54 3.671 ;
      RECT 28.51 3.525 28.52 3.68 ;
      RECT 28.486 3.532 28.51 3.69 ;
      RECT 28.4 3.554 28.486 3.71 ;
      RECT 28.39 3.573 28.4 3.725 ;
      RECT 28.366 3.58 28.39 3.731 ;
      RECT 28.28 3.602 28.366 3.756 ;
      RECT 28.24 3.627 28.28 3.783 ;
      RECT 28.23 3.636 28.24 3.793 ;
      RECT 28.18 3.646 28.23 3.802 ;
      RECT 28.16 3.66 28.18 3.812 ;
      RECT 28.13 3.67 28.16 3.817 ;
      RECT 28.12 3.675 28.13 3.82 ;
      RECT 28.046 3.677 28.12 3.827 ;
      RECT 27.96 3.681 28.046 3.839 ;
      RECT 27.95 3.684 27.96 3.845 ;
      RECT 27.69 3.635 27.95 3.895 ;
      RECT 29.22 3.705 29.41 3.915 ;
      RECT 29.21 3.71 29.42 3.91 ;
      RECT 29.2 3.71 29.42 3.875 ;
      RECT 29.12 3.595 29.38 3.855 ;
      RECT 28.03 3.125 28.22 3.425 ;
      RECT 28.02 3.125 28.22 3.42 ;
      RECT 28.01 3.125 28.23 3.415 ;
      RECT 28 3.125 28.23 3.41 ;
      RECT 28 3.125 28.26 3.385 ;
      RECT 27.96 2.165 28.22 2.425 ;
      RECT 27.77 2.09 27.856 2.423 ;
      RECT 27.77 2.09 27.9 2.419 ;
      RECT 27.75 2.094 27.91 2.418 ;
      RECT 27.9 2.085 27.91 2.418 ;
      RECT 27.77 2.09 27.92 2.417 ;
      RECT 27.75 2.1 27.96 2.416 ;
      RECT 27.74 2.095 27.92 2.408 ;
      RECT 27.73 2.11 27.96 2.315 ;
      RECT 27.73 2.16 28.16 2.315 ;
      RECT 27.73 2.15 28.14 2.315 ;
      RECT 27.73 2.14 28.11 2.315 ;
      RECT 27.73 2.13 28.05 2.315 ;
      RECT 27.73 2.115 28.03 2.315 ;
      RECT 27.856 2.086 27.91 2.418 ;
      RECT 26.93 2.745 27.07 3.035 ;
      RECT 27.19 2.768 27.2 2.955 ;
      RECT 27.89 2.665 28.07 2.895 ;
      RECT 27.89 2.665 28.08 2.885 ;
      RECT 28.1 2.67 28.11 2.875 ;
      RECT 28.08 2.665 28.1 2.88 ;
      RECT 27.84 2.669 27.89 2.895 ;
      RECT 27.83 2.674 27.84 2.895 ;
      RECT 27.796 2.679 27.83 2.896 ;
      RECT 27.71 2.694 27.796 2.898 ;
      RECT 27.696 2.706 27.71 2.901 ;
      RECT 27.61 2.716 27.696 2.903 ;
      RECT 27.586 2.726 27.61 2.905 ;
      RECT 27.5 2.737 27.586 2.905 ;
      RECT 27.47 2.747 27.5 2.905 ;
      RECT 27.44 2.752 27.47 2.908 ;
      RECT 27.42 2.757 27.44 2.913 ;
      RECT 27.4 2.762 27.42 2.915 ;
      RECT 27.35 2.77 27.4 2.915 ;
      RECT 27.33 2.774 27.35 2.915 ;
      RECT 27.31 2.773 27.33 2.92 ;
      RECT 27.25 2.771 27.31 2.935 ;
      RECT 27.2 2.769 27.25 2.95 ;
      RECT 27.11 2.766 27.19 3.035 ;
      RECT 27.08 2.76 27.11 3.035 ;
      RECT 27.07 2.75 27.08 3.035 ;
      RECT 26.88 2.745 26.93 2.96 ;
      RECT 26.87 2.75 26.88 2.95 ;
      RECT 27.11 3.225 27.37 3.485 ;
      RECT 27.11 3.225 27.4 3.375 ;
      RECT 27.11 3.225 27.44 3.36 ;
      RECT 27.37 3.145 27.56 3.355 ;
      RECT 27.37 3.15 27.57 3.345 ;
      RECT 27.32 3.22 27.57 3.345 ;
      RECT 27.35 3.155 27.37 3.485 ;
      RECT 27.34 3.18 27.57 3.345 ;
      RECT 26.52 3.125 26.53 3.355 ;
      RECT 26.42 2.245 26.49 3.355 ;
      RECT 27.16 2.355 27.42 2.615 ;
      RECT 26.86 2.405 26.99 2.565 ;
      RECT 27.076 2.412 27.16 2.565 ;
      RECT 26.99 2.407 27.076 2.565 ;
      RECT 26.8 2.405 26.86 2.575 ;
      RECT 26.77 2.403 26.8 2.59 ;
      RECT 26.75 2.401 26.77 2.6 ;
      RECT 26.74 2.399 26.75 2.605 ;
      RECT 26.72 2.398 26.74 2.615 ;
      RECT 26.71 2.396 26.72 2.62 ;
      RECT 26.69 2.395 26.71 2.625 ;
      RECT 26.67 2.39 26.69 2.63 ;
      RECT 26.64 2.376 26.67 2.64 ;
      RECT 26.6 2.355 26.64 2.655 ;
      RECT 26.59 2.34 26.6 2.665 ;
      RECT 26.57 2.331 26.59 2.675 ;
      RECT 26.56 2.322 26.57 2.695 ;
      RECT 26.55 2.317 26.56 2.755 ;
      RECT 26.53 2.311 26.55 2.84 ;
      RECT 26.53 3.15 26.54 3.35 ;
      RECT 26.52 2.306 26.53 3.07 ;
      RECT 26.51 2.28 26.52 3.355 ;
      RECT 26.49 2.25 26.51 3.355 ;
      RECT 26.4 2.245 26.42 2.58 ;
      RECT 26.41 2.68 26.42 3.355 ;
      RECT 26.4 2.72 26.41 3.355 ;
      RECT 26.37 2.245 26.4 2.525 ;
      RECT 26.38 2.81 26.4 3.355 ;
      RECT 26.365 2.915 26.38 3.355 ;
      RECT 26.34 2.245 26.37 2.48 ;
      RECT 26.36 2.947 26.365 3.355 ;
      RECT 26.34 3.05 26.36 3.355 ;
      RECT 26.33 2.245 26.34 2.47 ;
      RECT 26.33 3.12 26.34 3.35 ;
      RECT 26.31 2.245 26.33 2.46 ;
      RECT 26.3 2.25 26.31 2.45 ;
      RECT 26.51 3.525 26.53 3.765 ;
      RECT 25.83 3.455 25.91 3.725 ;
      RECT 25.74 3.455 25.75 3.665 ;
      RECT 27.02 3.525 27.03 3.725 ;
      RECT 26.94 3.515 27.02 3.75 ;
      RECT 26.936 3.515 26.94 3.776 ;
      RECT 26.85 3.515 26.936 3.786 ;
      RECT 26.83 3.515 26.85 3.794 ;
      RECT 26.806 3.516 26.83 3.792 ;
      RECT 26.72 3.521 26.806 3.787 ;
      RECT 26.702 3.525 26.72 3.781 ;
      RECT 26.616 3.525 26.702 3.777 ;
      RECT 26.53 3.525 26.616 3.769 ;
      RECT 26.426 3.525 26.51 3.762 ;
      RECT 26.34 3.525 26.426 3.756 ;
      RECT 26.28 3.52 26.34 3.75 ;
      RECT 26.252 3.514 26.28 3.747 ;
      RECT 26.166 3.511 26.252 3.744 ;
      RECT 26.08 3.507 26.166 3.738 ;
      RECT 26.035 3.495 26.08 3.734 ;
      RECT 26.01 3.48 26.035 3.732 ;
      RECT 25.97 3.465 26.01 3.73 ;
      RECT 25.91 3.455 25.97 3.727 ;
      RECT 25.82 3.455 25.83 3.72 ;
      RECT 25.805 3.455 25.82 3.71 ;
      RECT 25.75 3.455 25.805 3.685 ;
      RECT 25.73 3.47 25.74 3.66 ;
      RECT 25.86 2.635 26.12 2.895 ;
      RECT 25.86 2.645 26.14 2.855 ;
      RECT 25.86 2.65 26.15 2.85 ;
      RECT 23.84 2.115 24.1 2.375 ;
      RECT 23.83 2.145 24.1 2.355 ;
      RECT 25.76 2.055 26.01 2.315 ;
      RECT 25.75 2.055 25.76 2.316 ;
      RECT 25.72 2.14 25.75 2.318 ;
      RECT 25.71 2.145 25.72 2.32 ;
      RECT 25.65 2.16 25.71 2.326 ;
      RECT 25.62 2.18 25.65 2.333 ;
      RECT 25.59 2.191 25.62 2.34 ;
      RECT 25.57 2.201 25.59 2.345 ;
      RECT 25.552 2.204 25.57 2.344 ;
      RECT 25.466 2.203 25.552 2.344 ;
      RECT 25.38 2.2 25.466 2.343 ;
      RECT 25.294 2.197 25.38 2.342 ;
      RECT 25.208 2.194 25.294 2.342 ;
      RECT 25.122 2.192 25.208 2.341 ;
      RECT 25.036 2.189 25.122 2.34 ;
      RECT 24.95 2.186 25.036 2.34 ;
      RECT 24.932 2.185 24.95 2.339 ;
      RECT 24.846 2.184 24.932 2.339 ;
      RECT 24.76 2.182 24.846 2.338 ;
      RECT 24.674 2.181 24.76 2.338 ;
      RECT 24.588 2.18 24.674 2.337 ;
      RECT 24.502 2.178 24.588 2.337 ;
      RECT 24.416 2.177 24.502 2.336 ;
      RECT 24.33 2.175 24.416 2.336 ;
      RECT 24.306 2.174 24.33 2.335 ;
      RECT 24.22 2.169 24.306 2.335 ;
      RECT 24.186 2.162 24.22 2.335 ;
      RECT 24.1 2.152 24.186 2.335 ;
      RECT 23.82 2.15 23.83 2.35 ;
      RECT 25.1 3.205 25.36 3.465 ;
      RECT 25.1 3.205 25.44 3.251 ;
      RECT 25.24 3.185 25.45 3.24 ;
      RECT 25.3 3.16 25.51 3.2 ;
      RECT 25.31 3.155 25.51 3.2 ;
      RECT 25.32 3.13 25.51 3.2 ;
      RECT 25.38 2.96 25.43 3.29 ;
      RECT 25.33 3.09 25.52 3.15 ;
      RECT 25.37 3.016 25.38 3.329 ;
      RECT 25.33 3.09 25.55 3.125 ;
      RECT 25.33 3.09 25.57 3.1 ;
      RECT 25.44 2.89 25.63 3.095 ;
      RECT 25.43 2.9 25.64 3.09 ;
      RECT 25.35 3.063 25.64 3.09 ;
      RECT 25.36 3.039 25.37 3.345 ;
      RECT 25.45 2.885 25.62 3.095 ;
      RECT 24.74 2.675 24.93 2.885 ;
      RECT 23.31 2.605 23.57 2.865 ;
      RECT 23.66 2.595 23.76 2.805 ;
      RECT 23.61 2.615 23.65 2.805 ;
      RECT 24.93 2.685 24.94 2.88 ;
      RECT 24.73 2.685 24.74 2.88 ;
      RECT 24.71 2.7 24.73 2.87 ;
      RECT 24.7 2.71 24.71 2.865 ;
      RECT 24.66 2.71 24.7 2.863 ;
      RECT 24.636 2.704 24.66 2.86 ;
      RECT 24.55 2.699 24.636 2.857 ;
      RECT 24.49 2.695 24.55 2.852 ;
      RECT 24.456 2.692 24.49 2.849 ;
      RECT 24.37 2.682 24.456 2.845 ;
      RECT 24.366 2.675 24.37 2.842 ;
      RECT 24.28 2.67 24.366 2.84 ;
      RECT 24.252 2.663 24.28 2.836 ;
      RECT 24.166 2.658 24.252 2.833 ;
      RECT 24.08 2.649 24.166 2.828 ;
      RECT 24.07 2.644 24.08 2.825 ;
      RECT 24.056 2.643 24.07 2.825 ;
      RECT 23.97 2.639 24.056 2.82 ;
      RECT 23.95 2.633 23.97 2.816 ;
      RECT 23.89 2.628 23.95 2.815 ;
      RECT 23.86 2.62 23.89 2.815 ;
      RECT 23.85 2.605 23.86 2.815 ;
      RECT 23.846 2.595 23.85 2.814 ;
      RECT 23.76 2.595 23.846 2.81 ;
      RECT 23.65 2.605 23.66 2.805 ;
      RECT 23.58 2.615 23.61 2.8 ;
      RECT 23.57 2.615 23.58 2.8 ;
      RECT 24.49 3.115 24.75 3.375 ;
      RECT 24.42 3.125 24.75 3.335 ;
      RECT 24.41 3.13 24.75 3.33 ;
      RECT 23.83 3.115 24.09 3.375 ;
      RECT 23.83 3.16 24.2 3.365 ;
      RECT 23.83 3.155 24.19 3.365 ;
      RECT 22.74 3.322 22.92 3.765 ;
      RECT 22.73 3.322 22.92 3.763 ;
      RECT 22.73 3.337 22.93 3.76 ;
      RECT 22.72 2.26 22.85 3.758 ;
      RECT 22.72 3.385 22.99 3.645 ;
      RECT 22.72 3.36 22.94 3.645 ;
      RECT 22.72 3.295 22.91 3.758 ;
      RECT 22.72 3.255 22.88 3.758 ;
      RECT 22.72 3.21 22.87 3.758 ;
      RECT 22.72 3.15 22.86 3.758 ;
      RECT 22.71 2.545 22.85 3.2 ;
      RECT 22.75 2.245 22.86 3.065 ;
      RECT 22.72 2.26 22.9 2.52 ;
      RECT 22.72 2.26 22.91 2.47 ;
      RECT 22.75 2.245 22.92 2.463 ;
      RECT 22.74 2.247 22.93 2.458 ;
      RECT 22.73 2.252 22.94 2.45 ;
      RECT 21.59 7.77 21.88 8 ;
      RECT 21.65 6.29 21.82 8 ;
      RECT 21.645 6.655 21.995 7.005 ;
      RECT 21.59 6.29 21.88 6.52 ;
      RECT 21.185 2.395 21.29 2.965 ;
      RECT 21.185 2.73 21.51 2.96 ;
      RECT 21.185 2.76 21.68 2.93 ;
      RECT 21.185 2.395 21.375 2.96 ;
      RECT 20.6 2.36 20.89 2.59 ;
      RECT 20.6 2.395 21.375 2.565 ;
      RECT 20.66 0.88 20.83 2.59 ;
      RECT 20.6 0.88 20.89 1.11 ;
      RECT 20.6 7.77 20.89 8 ;
      RECT 20.66 6.29 20.83 8 ;
      RECT 20.6 6.29 20.89 6.52 ;
      RECT 20.6 6.325 21.455 6.485 ;
      RECT 21.285 5.92 21.455 6.485 ;
      RECT 20.6 6.32 20.995 6.485 ;
      RECT 21.22 5.92 21.51 6.15 ;
      RECT 21.22 5.95 21.68 6.12 ;
      RECT 20.23 2.73 20.52 2.96 ;
      RECT 20.23 2.76 20.69 2.93 ;
      RECT 20.295 1.655 20.46 2.96 ;
      RECT 18.81 1.625 19.1 1.855 ;
      RECT 18.81 1.655 20.46 1.825 ;
      RECT 18.87 0.885 19.04 1.855 ;
      RECT 18.81 0.885 19.1 1.115 ;
      RECT 18.81 7.765 19.1 7.995 ;
      RECT 18.87 7.025 19.04 7.995 ;
      RECT 18.87 7.12 20.46 7.29 ;
      RECT 20.29 5.92 20.46 7.29 ;
      RECT 18.81 7.025 19.1 7.255 ;
      RECT 20.23 5.92 20.52 6.15 ;
      RECT 20.23 5.95 20.69 6.12 ;
      RECT 16.845 3.43 17.195 3.78 ;
      RECT 16.935 2.025 17.105 3.78 ;
      RECT 19.24 1.965 19.59 2.315 ;
      RECT 16.935 2.025 18.555 2.2 ;
      RECT 16.935 2.025 19.59 2.195 ;
      RECT 19.265 6.655 19.59 6.98 ;
      RECT 14.66 6.605 15.01 6.955 ;
      RECT 19.24 6.655 19.59 6.885 ;
      RECT 14.48 6.655 15.01 6.885 ;
      RECT 14.31 6.685 19.59 6.855 ;
      RECT 18.465 2.365 18.785 2.685 ;
      RECT 18.435 2.365 18.785 2.595 ;
      RECT 18.265 2.395 18.785 2.565 ;
      RECT 18.465 6.225 18.785 6.545 ;
      RECT 18.435 6.285 18.785 6.515 ;
      RECT 18.265 6.315 18.785 6.485 ;
      RECT 14.305 3.255 14.495 3.925 ;
      RECT 14.245 3.665 14.285 3.925 ;
      RECT 15.615 2.89 15.625 3.111 ;
      RECT 15.545 2.885 15.615 3.236 ;
      RECT 15.535 2.885 15.545 3.36 ;
      RECT 15.505 2.885 15.535 3.41 ;
      RECT 15.485 2.885 15.505 3.485 ;
      RECT 15.465 2.885 15.485 3.555 ;
      RECT 15.435 2.885 15.465 3.595 ;
      RECT 15.425 2.885 15.435 3.615 ;
      RECT 15.415 2.885 15.425 3.626 ;
      RECT 15.405 3.135 15.415 3.628 ;
      RECT 15.395 3.2 15.405 3.63 ;
      RECT 15.385 3.295 15.395 3.632 ;
      RECT 15.375 3.37 15.385 3.634 ;
      RECT 15.325 3.394 15.375 3.64 ;
      RECT 15.285 3.429 15.325 3.649 ;
      RECT 15.275 3.445 15.285 3.654 ;
      RECT 15.261 3.45 15.275 3.657 ;
      RECT 15.175 3.49 15.261 3.668 ;
      RECT 15.095 3.533 15.175 3.686 ;
      RECT 15.075 3.543 15.095 3.697 ;
      RECT 15.045 3.551 15.075 3.702 ;
      RECT 15.025 3.561 15.045 3.707 ;
      RECT 15.001 3.567 15.025 3.712 ;
      RECT 14.915 3.577 15.001 3.725 ;
      RECT 14.837 3.583 14.915 3.745 ;
      RECT 14.751 3.578 14.837 3.764 ;
      RECT 14.665 3.574 14.751 3.785 ;
      RECT 14.585 3.57 14.665 3.8 ;
      RECT 14.515 3.566 14.585 3.831 ;
      RECT 14.505 3.277 14.515 3.345 ;
      RECT 14.505 3.555 14.515 3.861 ;
      RECT 14.495 3.262 14.505 3.49 ;
      RECT 14.495 3.535 14.505 3.925 ;
      RECT 14.285 3.285 14.305 3.925 ;
      RECT 15.085 2.605 15.095 3.345 ;
      RECT 14.905 3.125 14.925 3.345 ;
      RECT 14.915 3.115 14.925 3.345 ;
      RECT 15.415 2.155 15.455 2.415 ;
      RECT 15.405 2.155 15.415 2.425 ;
      RECT 15.371 2.155 15.405 2.452 ;
      RECT 15.285 2.155 15.371 2.512 ;
      RECT 15.265 2.155 15.285 2.575 ;
      RECT 15.205 2.155 15.265 2.74 ;
      RECT 15.195 2.155 15.205 2.9 ;
      RECT 15.165 2.346 15.195 2.995 ;
      RECT 15.155 2.401 15.165 3.095 ;
      RECT 15.145 2.43 15.155 3.14 ;
      RECT 15.135 2.455 15.145 3.173 ;
      RECT 15.125 2.49 15.135 3.228 ;
      RECT 15.105 2.535 15.125 3.29 ;
      RECT 15.095 2.58 15.105 3.34 ;
      RECT 15.075 2.64 15.085 3.345 ;
      RECT 15.065 2.67 15.075 3.345 ;
      RECT 15.045 2.7 15.065 3.345 ;
      RECT 14.995 2.805 15.045 3.345 ;
      RECT 14.985 2.9 14.995 3.345 ;
      RECT 14.975 2.93 14.985 3.345 ;
      RECT 14.95 2.98 14.975 3.345 ;
      RECT 14.945 3.035 14.95 3.345 ;
      RECT 14.925 3.06 14.945 3.345 ;
      RECT 14.885 3.14 14.905 3.335 ;
      RECT 14.635 2.725 14.705 2.935 ;
      RECT 11.875 2.635 12.135 2.895 ;
      RECT 14.705 2.73 14.715 2.93 ;
      RECT 14.591 2.723 14.635 2.935 ;
      RECT 14.505 2.716 14.591 2.935 ;
      RECT 14.485 2.711 14.505 2.925 ;
      RECT 14.475 2.709 14.485 2.905 ;
      RECT 14.425 2.706 14.475 2.9 ;
      RECT 14.395 2.702 14.425 2.895 ;
      RECT 14.375 2.7 14.395 2.89 ;
      RECT 14.335 2.697 14.375 2.885 ;
      RECT 14.265 2.691 14.335 2.88 ;
      RECT 14.235 2.686 14.265 2.875 ;
      RECT 14.215 2.684 14.235 2.87 ;
      RECT 14.185 2.681 14.215 2.865 ;
      RECT 14.125 2.677 14.185 2.86 ;
      RECT 14.055 2.675 14.125 2.85 ;
      RECT 14.021 2.673 14.055 2.843 ;
      RECT 13.935 2.668 14.021 2.835 ;
      RECT 13.901 2.662 13.935 2.827 ;
      RECT 13.815 2.652 13.901 2.819 ;
      RECT 13.781 2.643 13.815 2.811 ;
      RECT 13.695 2.638 13.781 2.803 ;
      RECT 13.625 2.635 13.695 2.793 ;
      RECT 13.605 2.63 13.625 2.787 ;
      RECT 13.601 2.625 13.605 2.786 ;
      RECT 13.515 2.621 13.601 2.781 ;
      RECT 13.475 2.616 13.515 2.774 ;
      RECT 13.395 2.615 13.475 2.769 ;
      RECT 13.375 2.615 13.395 2.766 ;
      RECT 13.349 2.615 13.375 2.766 ;
      RECT 13.263 2.617 13.349 2.77 ;
      RECT 13.177 2.619 13.263 2.777 ;
      RECT 13.091 2.621 13.177 2.783 ;
      RECT 13.005 2.624 13.091 2.79 ;
      RECT 12.971 2.626 13.005 2.795 ;
      RECT 12.885 2.631 12.971 2.8 ;
      RECT 12.861 2.626 12.885 2.804 ;
      RECT 12.775 2.631 12.861 2.809 ;
      RECT 12.737 2.636 12.775 2.814 ;
      RECT 12.651 2.639 12.737 2.819 ;
      RECT 12.565 2.643 12.651 2.826 ;
      RECT 12.501 2.645 12.565 2.832 ;
      RECT 12.415 2.645 12.501 2.838 ;
      RECT 12.331 2.646 12.415 2.845 ;
      RECT 12.245 2.649 12.331 2.852 ;
      RECT 12.221 2.651 12.245 2.856 ;
      RECT 12.135 2.653 12.221 2.861 ;
      RECT 11.865 2.67 11.875 2.865 ;
      RECT 14.05 7.765 14.34 7.995 ;
      RECT 14.11 7.025 14.28 7.995 ;
      RECT 14 7.055 14.375 7.425 ;
      RECT 14.05 7.025 14.34 7.425 ;
      RECT 14.105 2.247 14.295 2.455 ;
      RECT 14.095 2.252 14.305 2.45 ;
      RECT 14.085 2.233 14.095 2.445 ;
      RECT 14.055 2.228 14.085 2.44 ;
      RECT 14.015 2.252 14.305 2.43 ;
      RECT 13.795 2.165 14.055 2.425 ;
      RECT 14.095 2.236 14.105 2.45 ;
      RECT 13.795 2.245 14.285 2.425 ;
      RECT 13.795 2.241 14.145 2.425 ;
      RECT 13.745 3.155 13.795 3.435 ;
      RECT 13.675 3.125 13.705 3.435 ;
      RECT 13.815 3.155 13.875 3.415 ;
      RECT 13.675 3.115 13.695 3.435 ;
      RECT 13.795 3.155 13.815 3.425 ;
      RECT 13.715 3.145 13.745 3.435 ;
      RECT 13.705 3.13 13.715 3.435 ;
      RECT 13.655 3.105 13.675 3.435 ;
      RECT 13.625 3.09 13.655 3.435 ;
      RECT 13.615 3.08 13.625 3.435 ;
      RECT 13.595 3.069 13.615 3.43 ;
      RECT 13.575 3.057 13.595 3.4 ;
      RECT 13.565 3.048 13.575 3.383 ;
      RECT 13.535 3.03 13.565 3.375 ;
      RECT 13.525 2.995 13.535 3.367 ;
      RECT 13.515 2.975 13.525 3.36 ;
      RECT 13.505 2.955 13.515 3.353 ;
      RECT 13.495 2.94 13.505 3.348 ;
      RECT 13.485 2.92 13.495 3.343 ;
      RECT 13.475 2.915 13.485 3.338 ;
      RECT 13.471 2.905 13.475 3.334 ;
      RECT 13.385 2.905 13.471 3.309 ;
      RECT 13.355 2.905 13.385 3.275 ;
      RECT 13.345 2.905 13.355 3.255 ;
      RECT 13.285 2.905 13.345 3.2 ;
      RECT 13.275 2.92 13.285 3.145 ;
      RECT 13.265 2.93 13.275 3.125 ;
      RECT 13.215 3.665 13.475 3.925 ;
      RECT 13.135 3.685 13.475 3.901 ;
      RECT 13.115 3.685 13.475 3.896 ;
      RECT 13.091 3.685 13.475 3.894 ;
      RECT 13.005 3.685 13.475 3.889 ;
      RECT 12.855 3.625 13.115 3.885 ;
      RECT 12.815 3.68 13.135 3.88 ;
      RECT 12.805 3.69 13.475 3.875 ;
      RECT 12.825 3.675 13.115 3.885 ;
      RECT 12.715 2.115 12.975 2.375 ;
      RECT 12.715 2.2 12.985 2.3 ;
      RECT 11.885 3.63 11.905 3.874 ;
      RECT 11.885 3.63 11.955 3.869 ;
      RECT 11.865 3.635 11.955 3.868 ;
      RECT 11.855 3.65 12.041 3.858 ;
      RECT 11.855 3.65 12.115 3.855 ;
      RECT 11.85 3.687 12.125 3.845 ;
      RECT 11.85 3.687 12.211 3.841 ;
      RECT 11.85 3.687 12.225 3.827 ;
      RECT 12.125 3.565 12.385 3.825 ;
      RECT 11.845 3.692 12.385 3.82 ;
      RECT 11.835 3.74 12.385 3.795 ;
      RECT 12.105 3.605 12.125 3.854 ;
      RECT 12.041 3.609 12.105 3.857 ;
      RECT 11.905 3.622 12.385 3.825 ;
      RECT 11.955 3.616 12.041 3.862 ;
      RECT 11.355 2.475 11.365 2.645 ;
      RECT 11.415 2.435 11.425 2.615 ;
      RECT 11.715 2.245 11.725 2.455 ;
      RECT 12.045 2.095 12.295 2.355 ;
      RECT 12.035 2.095 12.045 2.357 ;
      RECT 12.025 2.155 12.035 2.361 ;
      RECT 11.995 2.157 12.025 2.369 ;
      RECT 11.965 2.162 11.995 2.383 ;
      RECT 11.955 2.166 11.965 2.393 ;
      RECT 11.925 2.171 11.955 2.405 ;
      RECT 11.895 2.18 11.925 2.406 ;
      RECT 11.825 2.19 11.895 2.41 ;
      RECT 11.785 2.195 11.825 2.414 ;
      RECT 11.765 2.195 11.785 2.425 ;
      RECT 11.755 2.2 11.765 2.435 ;
      RECT 11.745 2.21 11.755 2.438 ;
      RECT 11.735 2.23 11.745 2.443 ;
      RECT 11.725 2.24 11.735 2.445 ;
      RECT 11.695 2.255 11.715 2.462 ;
      RECT 11.685 2.267 11.695 2.472 ;
      RECT 11.675 2.273 11.685 2.475 ;
      RECT 11.641 2.286 11.675 2.485 ;
      RECT 11.555 2.32 11.641 2.518 ;
      RECT 11.535 2.355 11.555 2.547 ;
      RECT 11.515 2.37 11.535 2.559 ;
      RECT 11.495 2.38 11.515 2.571 ;
      RECT 11.445 2.399 11.495 2.591 ;
      RECT 11.435 2.416 11.445 2.605 ;
      RECT 11.425 2.422 11.435 2.61 ;
      RECT 11.405 2.44 11.415 2.618 ;
      RECT 11.395 2.445 11.405 2.625 ;
      RECT 11.385 2.456 11.395 2.632 ;
      RECT 11.365 2.461 11.385 2.64 ;
      RECT 11.345 2.475 11.355 2.65 ;
      RECT 11.335 2.48 11.345 2.66 ;
      RECT 11.305 2.494 11.335 2.67 ;
      RECT 11.295 2.507 11.305 2.68 ;
      RECT 11.215 2.538 11.295 2.705 ;
      RECT 11.195 2.568 11.215 2.73 ;
      RECT 11.185 2.573 11.195 2.737 ;
      RECT 11.155 2.585 11.185 2.743 ;
      RECT 11.145 2.6 11.155 2.749 ;
      RECT 11.135 2.605 11.145 2.752 ;
      RECT 11.115 2.615 11.135 2.756 ;
      RECT 11.095 2.62 11.115 2.762 ;
      RECT 11.065 2.625 11.095 2.77 ;
      RECT 11.035 2.63 11.065 2.78 ;
      RECT 11.005 2.64 11.035 2.789 ;
      RECT 10.965 2.645 11.005 2.797 ;
      RECT 10.915 2.638 10.965 2.809 ;
      RECT 10.895 2.629 10.915 2.82 ;
      RECT 10.885 2.626 10.895 2.825 ;
      RECT 10.845 2.625 10.885 2.826 ;
      RECT 10.835 2.61 10.845 2.827 ;
      RECT 10.807 2.595 10.835 2.828 ;
      RECT 10.721 2.595 10.807 2.83 ;
      RECT 10.635 2.595 10.721 2.834 ;
      RECT 10.615 2.595 10.635 2.83 ;
      RECT 10.605 2.605 10.615 2.823 ;
      RECT 10.595 2.62 10.605 2.818 ;
      RECT 10.585 2.625 10.595 2.795 ;
      RECT 12.065 3.13 12.075 3.33 ;
      RECT 12.015 3.125 12.065 3.35 ;
      RECT 12.005 3.125 12.015 3.37 ;
      RECT 11.961 3.125 12.005 3.374 ;
      RECT 11.875 3.125 11.961 3.371 ;
      RECT 11.815 3.135 11.875 3.368 ;
      RECT 11.755 3.149 11.815 3.366 ;
      RECT 11.745 3.154 11.755 3.364 ;
      RECT 11.735 3.16 11.745 3.363 ;
      RECT 11.665 3.173 11.735 3.359 ;
      RECT 11.617 3.187 11.665 3.36 ;
      RECT 11.531 3.203 11.617 3.372 ;
      RECT 11.445 3.224 11.531 3.388 ;
      RECT 11.425 3.235 11.445 3.398 ;
      RECT 11.345 3.245 11.425 3.408 ;
      RECT 11.311 3.259 11.345 3.42 ;
      RECT 11.225 3.274 11.311 3.435 ;
      RECT 11.195 3.29 11.225 3.445 ;
      RECT 11.14 3.305 11.195 3.456 ;
      RECT 11.095 3.323 11.14 3.476 ;
      RECT 11.041 3.342 11.095 3.496 ;
      RECT 10.955 3.368 11.041 3.523 ;
      RECT 10.935 3.39 10.955 3.543 ;
      RECT 10.875 3.405 10.935 3.559 ;
      RECT 10.865 3.42 10.875 3.573 ;
      RECT 10.845 3.425 10.865 3.579 ;
      RECT 10.815 3.438 10.845 3.589 ;
      RECT 10.795 3.443 10.815 3.598 ;
      RECT 10.785 3.45 10.795 3.603 ;
      RECT 10.775 3.455 10.785 3.606 ;
      RECT 10.735 3.465 10.775 3.615 ;
      RECT 10.71 3.48 10.735 3.627 ;
      RECT 10.665 3.495 10.71 3.639 ;
      RECT 10.645 3.507 10.665 3.651 ;
      RECT 10.615 3.512 10.645 3.661 ;
      RECT 10.595 3.519 10.615 3.671 ;
      RECT 10.585 3.525 10.595 3.68 ;
      RECT 10.561 3.532 10.585 3.69 ;
      RECT 10.475 3.554 10.561 3.71 ;
      RECT 10.465 3.573 10.475 3.725 ;
      RECT 10.441 3.58 10.465 3.731 ;
      RECT 10.355 3.602 10.441 3.756 ;
      RECT 10.315 3.627 10.355 3.783 ;
      RECT 10.305 3.636 10.315 3.793 ;
      RECT 10.255 3.646 10.305 3.802 ;
      RECT 10.235 3.66 10.255 3.812 ;
      RECT 10.205 3.67 10.235 3.817 ;
      RECT 10.195 3.675 10.205 3.82 ;
      RECT 10.121 3.677 10.195 3.827 ;
      RECT 10.035 3.681 10.121 3.839 ;
      RECT 10.025 3.684 10.035 3.845 ;
      RECT 9.765 3.635 10.025 3.895 ;
      RECT 11.295 3.705 11.485 3.915 ;
      RECT 11.285 3.71 11.495 3.91 ;
      RECT 11.275 3.71 11.495 3.875 ;
      RECT 11.195 3.595 11.455 3.855 ;
      RECT 10.105 3.125 10.295 3.425 ;
      RECT 10.095 3.125 10.295 3.42 ;
      RECT 10.085 3.125 10.305 3.415 ;
      RECT 10.075 3.125 10.305 3.41 ;
      RECT 10.075 3.125 10.335 3.385 ;
      RECT 10.035 2.165 10.295 2.425 ;
      RECT 9.845 2.09 9.931 2.423 ;
      RECT 9.845 2.09 9.975 2.419 ;
      RECT 9.825 2.094 9.985 2.418 ;
      RECT 9.975 2.085 9.985 2.418 ;
      RECT 9.845 2.09 9.995 2.417 ;
      RECT 9.825 2.1 10.035 2.416 ;
      RECT 9.815 2.095 9.995 2.408 ;
      RECT 9.805 2.11 10.035 2.315 ;
      RECT 9.805 2.16 10.235 2.315 ;
      RECT 9.805 2.15 10.215 2.315 ;
      RECT 9.805 2.14 10.185 2.315 ;
      RECT 9.805 2.13 10.125 2.315 ;
      RECT 9.805 2.115 10.105 2.315 ;
      RECT 9.931 2.086 9.985 2.418 ;
      RECT 9.005 2.745 9.145 3.035 ;
      RECT 9.265 2.768 9.275 2.955 ;
      RECT 9.965 2.665 10.145 2.895 ;
      RECT 9.965 2.665 10.155 2.885 ;
      RECT 10.175 2.67 10.185 2.875 ;
      RECT 10.155 2.665 10.175 2.88 ;
      RECT 9.915 2.669 9.965 2.895 ;
      RECT 9.905 2.674 9.915 2.895 ;
      RECT 9.871 2.679 9.905 2.896 ;
      RECT 9.785 2.694 9.871 2.898 ;
      RECT 9.771 2.706 9.785 2.901 ;
      RECT 9.685 2.716 9.771 2.903 ;
      RECT 9.661 2.726 9.685 2.905 ;
      RECT 9.575 2.737 9.661 2.905 ;
      RECT 9.545 2.747 9.575 2.905 ;
      RECT 9.515 2.752 9.545 2.908 ;
      RECT 9.495 2.757 9.515 2.913 ;
      RECT 9.475 2.762 9.495 2.915 ;
      RECT 9.425 2.77 9.475 2.915 ;
      RECT 9.405 2.774 9.425 2.915 ;
      RECT 9.385 2.773 9.405 2.92 ;
      RECT 9.325 2.771 9.385 2.935 ;
      RECT 9.275 2.769 9.325 2.95 ;
      RECT 9.185 2.766 9.265 3.035 ;
      RECT 9.155 2.76 9.185 3.035 ;
      RECT 9.145 2.75 9.155 3.035 ;
      RECT 8.955 2.745 9.005 2.96 ;
      RECT 8.945 2.75 8.955 2.95 ;
      RECT 9.185 3.225 9.445 3.485 ;
      RECT 9.185 3.225 9.475 3.375 ;
      RECT 9.185 3.225 9.515 3.36 ;
      RECT 9.445 3.145 9.635 3.355 ;
      RECT 9.445 3.15 9.645 3.345 ;
      RECT 9.395 3.22 9.645 3.345 ;
      RECT 9.425 3.155 9.445 3.485 ;
      RECT 9.415 3.18 9.645 3.345 ;
      RECT 8.595 3.125 8.605 3.355 ;
      RECT 8.495 2.245 8.565 3.355 ;
      RECT 9.235 2.355 9.495 2.615 ;
      RECT 8.935 2.405 9.065 2.565 ;
      RECT 9.151 2.412 9.235 2.565 ;
      RECT 9.065 2.407 9.151 2.565 ;
      RECT 8.875 2.405 8.935 2.575 ;
      RECT 8.845 2.403 8.875 2.59 ;
      RECT 8.825 2.401 8.845 2.6 ;
      RECT 8.815 2.399 8.825 2.605 ;
      RECT 8.795 2.398 8.815 2.615 ;
      RECT 8.785 2.396 8.795 2.62 ;
      RECT 8.765 2.395 8.785 2.625 ;
      RECT 8.745 2.39 8.765 2.63 ;
      RECT 8.715 2.376 8.745 2.64 ;
      RECT 8.675 2.355 8.715 2.655 ;
      RECT 8.665 2.34 8.675 2.665 ;
      RECT 8.645 2.331 8.665 2.675 ;
      RECT 8.635 2.322 8.645 2.695 ;
      RECT 8.625 2.317 8.635 2.755 ;
      RECT 8.605 2.311 8.625 2.84 ;
      RECT 8.605 3.15 8.615 3.35 ;
      RECT 8.595 2.306 8.605 3.07 ;
      RECT 8.585 2.28 8.595 3.355 ;
      RECT 8.565 2.25 8.585 3.355 ;
      RECT 8.475 2.245 8.495 2.58 ;
      RECT 8.485 2.68 8.495 3.355 ;
      RECT 8.475 2.72 8.485 3.355 ;
      RECT 8.445 2.245 8.475 2.525 ;
      RECT 8.455 2.81 8.475 3.355 ;
      RECT 8.44 2.915 8.455 3.355 ;
      RECT 8.415 2.245 8.445 2.48 ;
      RECT 8.435 2.947 8.44 3.355 ;
      RECT 8.415 3.05 8.435 3.355 ;
      RECT 8.405 2.245 8.415 2.47 ;
      RECT 8.405 3.12 8.415 3.35 ;
      RECT 8.385 2.245 8.405 2.46 ;
      RECT 8.375 2.25 8.385 2.45 ;
      RECT 8.585 3.525 8.605 3.765 ;
      RECT 7.905 3.455 7.985 3.725 ;
      RECT 7.815 3.455 7.825 3.665 ;
      RECT 9.095 3.525 9.105 3.725 ;
      RECT 9.015 3.515 9.095 3.75 ;
      RECT 9.011 3.515 9.015 3.776 ;
      RECT 8.925 3.515 9.011 3.786 ;
      RECT 8.905 3.515 8.925 3.794 ;
      RECT 8.881 3.516 8.905 3.792 ;
      RECT 8.795 3.521 8.881 3.787 ;
      RECT 8.777 3.525 8.795 3.781 ;
      RECT 8.691 3.525 8.777 3.777 ;
      RECT 8.605 3.525 8.691 3.769 ;
      RECT 8.501 3.525 8.585 3.762 ;
      RECT 8.415 3.525 8.501 3.756 ;
      RECT 8.355 3.52 8.415 3.75 ;
      RECT 8.327 3.514 8.355 3.747 ;
      RECT 8.241 3.511 8.327 3.744 ;
      RECT 8.155 3.507 8.241 3.738 ;
      RECT 8.11 3.495 8.155 3.734 ;
      RECT 8.085 3.48 8.11 3.732 ;
      RECT 8.045 3.465 8.085 3.73 ;
      RECT 7.985 3.455 8.045 3.727 ;
      RECT 7.895 3.455 7.905 3.72 ;
      RECT 7.88 3.455 7.895 3.71 ;
      RECT 7.825 3.455 7.88 3.685 ;
      RECT 7.805 3.47 7.815 3.66 ;
      RECT 7.935 2.635 8.195 2.895 ;
      RECT 7.935 2.645 8.215 2.855 ;
      RECT 7.935 2.65 8.225 2.85 ;
      RECT 5.915 2.115 6.175 2.375 ;
      RECT 5.905 2.145 6.175 2.355 ;
      RECT 7.835 2.055 8.085 2.315 ;
      RECT 7.825 2.055 7.835 2.316 ;
      RECT 7.795 2.14 7.825 2.318 ;
      RECT 7.785 2.145 7.795 2.32 ;
      RECT 7.725 2.16 7.785 2.326 ;
      RECT 7.695 2.18 7.725 2.333 ;
      RECT 7.665 2.191 7.695 2.34 ;
      RECT 7.645 2.201 7.665 2.345 ;
      RECT 7.627 2.204 7.645 2.344 ;
      RECT 7.541 2.203 7.627 2.344 ;
      RECT 7.455 2.2 7.541 2.343 ;
      RECT 7.369 2.197 7.455 2.342 ;
      RECT 7.283 2.194 7.369 2.342 ;
      RECT 7.197 2.192 7.283 2.341 ;
      RECT 7.111 2.189 7.197 2.34 ;
      RECT 7.025 2.186 7.111 2.34 ;
      RECT 7.007 2.185 7.025 2.339 ;
      RECT 6.921 2.184 7.007 2.339 ;
      RECT 6.835 2.182 6.921 2.338 ;
      RECT 6.749 2.181 6.835 2.338 ;
      RECT 6.663 2.18 6.749 2.337 ;
      RECT 6.577 2.178 6.663 2.337 ;
      RECT 6.491 2.177 6.577 2.336 ;
      RECT 6.405 2.175 6.491 2.336 ;
      RECT 6.381 2.174 6.405 2.335 ;
      RECT 6.295 2.169 6.381 2.335 ;
      RECT 6.261 2.162 6.295 2.335 ;
      RECT 6.175 2.152 6.261 2.335 ;
      RECT 5.895 2.15 5.905 2.35 ;
      RECT 7.175 3.205 7.435 3.465 ;
      RECT 7.175 3.205 7.515 3.251 ;
      RECT 7.315 3.185 7.525 3.24 ;
      RECT 7.375 3.16 7.585 3.2 ;
      RECT 7.385 3.155 7.585 3.2 ;
      RECT 7.395 3.13 7.585 3.2 ;
      RECT 7.455 2.96 7.505 3.29 ;
      RECT 7.405 3.09 7.595 3.15 ;
      RECT 7.445 3.016 7.455 3.329 ;
      RECT 7.405 3.09 7.625 3.125 ;
      RECT 7.405 3.09 7.645 3.1 ;
      RECT 7.515 2.89 7.705 3.095 ;
      RECT 7.505 2.9 7.715 3.09 ;
      RECT 7.425 3.063 7.715 3.09 ;
      RECT 7.435 3.039 7.445 3.345 ;
      RECT 7.525 2.885 7.695 3.095 ;
      RECT 6.815 2.675 7.005 2.885 ;
      RECT 5.385 2.605 5.645 2.865 ;
      RECT 5.735 2.595 5.835 2.805 ;
      RECT 5.685 2.615 5.725 2.805 ;
      RECT 7.005 2.685 7.015 2.88 ;
      RECT 6.805 2.685 6.815 2.88 ;
      RECT 6.785 2.7 6.805 2.87 ;
      RECT 6.775 2.71 6.785 2.865 ;
      RECT 6.735 2.71 6.775 2.863 ;
      RECT 6.711 2.704 6.735 2.86 ;
      RECT 6.625 2.699 6.711 2.857 ;
      RECT 6.565 2.695 6.625 2.852 ;
      RECT 6.531 2.692 6.565 2.849 ;
      RECT 6.445 2.682 6.531 2.845 ;
      RECT 6.441 2.675 6.445 2.842 ;
      RECT 6.355 2.67 6.441 2.84 ;
      RECT 6.327 2.663 6.355 2.836 ;
      RECT 6.241 2.658 6.327 2.833 ;
      RECT 6.155 2.649 6.241 2.828 ;
      RECT 6.145 2.644 6.155 2.825 ;
      RECT 6.131 2.643 6.145 2.825 ;
      RECT 6.045 2.639 6.131 2.82 ;
      RECT 6.025 2.633 6.045 2.816 ;
      RECT 5.965 2.628 6.025 2.815 ;
      RECT 5.935 2.62 5.965 2.815 ;
      RECT 5.925 2.605 5.935 2.815 ;
      RECT 5.921 2.595 5.925 2.814 ;
      RECT 5.835 2.595 5.921 2.81 ;
      RECT 5.725 2.605 5.735 2.805 ;
      RECT 5.655 2.615 5.685 2.8 ;
      RECT 5.645 2.615 5.655 2.8 ;
      RECT 6.565 3.115 6.825 3.375 ;
      RECT 6.495 3.125 6.825 3.335 ;
      RECT 6.485 3.13 6.825 3.33 ;
      RECT 5.905 3.115 6.165 3.375 ;
      RECT 5.905 3.16 6.275 3.365 ;
      RECT 5.905 3.155 6.265 3.365 ;
      RECT 4.815 3.322 4.995 3.765 ;
      RECT 4.805 3.322 4.995 3.763 ;
      RECT 4.805 3.337 5.005 3.76 ;
      RECT 4.795 2.26 4.925 3.758 ;
      RECT 4.795 3.385 5.065 3.645 ;
      RECT 4.795 3.36 5.015 3.645 ;
      RECT 4.795 3.295 4.985 3.758 ;
      RECT 4.795 3.255 4.955 3.758 ;
      RECT 4.795 3.21 4.945 3.758 ;
      RECT 4.795 3.15 4.935 3.758 ;
      RECT 4.785 2.545 4.925 3.2 ;
      RECT 4.825 2.245 4.935 3.065 ;
      RECT 4.795 2.26 4.975 2.52 ;
      RECT 4.795 2.26 4.985 2.47 ;
      RECT 4.825 2.245 4.995 2.463 ;
      RECT 4.815 2.247 5.005 2.458 ;
      RECT 4.805 2.252 5.015 2.45 ;
      RECT 3.02 7.765 3.31 7.995 ;
      RECT 3.08 7.025 3.25 7.995 ;
      RECT 2.99 7.025 3.34 7.315 ;
      RECT 2.615 6.285 2.965 6.575 ;
      RECT 2.475 6.315 2.965 6.485 ;
      RECT 88.52 1.14 88.895 1.51 ;
      RECT 82.495 2.225 82.755 2.485 ;
      RECT 70.595 1.14 70.97 1.51 ;
      RECT 64.57 2.225 64.83 2.485 ;
      RECT 52.67 1.14 53.045 1.51 ;
      RECT 46.645 2.225 46.905 2.485 ;
      RECT 34.745 1.14 35.12 1.51 ;
      RECT 28.72 2.225 28.98 2.485 ;
      RECT 16.82 1.14 17.195 1.51 ;
      RECT 10.795 2.225 11.055 2.485 ;
    LAYER mcon ;
      RECT 93.35 6.32 93.52 6.49 ;
      RECT 93.355 6.315 93.525 6.485 ;
      RECT 75.425 6.32 75.595 6.49 ;
      RECT 75.43 6.315 75.6 6.485 ;
      RECT 57.5 6.32 57.67 6.49 ;
      RECT 57.505 6.315 57.675 6.485 ;
      RECT 39.575 6.32 39.745 6.49 ;
      RECT 39.58 6.315 39.75 6.485 ;
      RECT 21.65 6.32 21.82 6.49 ;
      RECT 21.655 6.315 21.825 6.485 ;
      RECT 93.35 7.8 93.52 7.97 ;
      RECT 93 0.1 93.17 0.27 ;
      RECT 93 8.61 93.17 8.78 ;
      RECT 92.98 2.76 93.15 2.93 ;
      RECT 92.98 5.95 93.15 6.12 ;
      RECT 92.36 0.91 92.53 1.08 ;
      RECT 92.36 2.39 92.53 2.56 ;
      RECT 92.36 6.32 92.53 6.49 ;
      RECT 92.36 7.8 92.53 7.97 ;
      RECT 92.01 0.1 92.18 0.27 ;
      RECT 92.01 8.61 92.18 8.78 ;
      RECT 91.99 2.76 92.16 2.93 ;
      RECT 91.99 5.95 92.16 6.12 ;
      RECT 91.31 0.105 91.48 0.275 ;
      RECT 91.31 8.605 91.48 8.775 ;
      RECT 91 2.025 91.17 2.195 ;
      RECT 91 6.685 91.17 6.855 ;
      RECT 90.63 0.105 90.8 0.275 ;
      RECT 90.63 8.605 90.8 8.775 ;
      RECT 90.57 0.915 90.74 1.085 ;
      RECT 90.57 1.655 90.74 1.825 ;
      RECT 90.57 7.055 90.74 7.225 ;
      RECT 90.57 7.795 90.74 7.965 ;
      RECT 90.195 2.395 90.365 2.565 ;
      RECT 90.195 6.315 90.365 6.485 ;
      RECT 89.95 0.105 90.12 0.275 ;
      RECT 89.95 8.605 90.12 8.775 ;
      RECT 89.27 0.105 89.44 0.275 ;
      RECT 89.27 8.605 89.44 8.775 ;
      RECT 87.985 1.565 88.155 1.735 ;
      RECT 87.525 1.565 87.695 1.735 ;
      RECT 87.135 2.905 87.305 3.075 ;
      RECT 87.065 1.565 87.235 1.735 ;
      RECT 86.925 2.245 87.095 2.415 ;
      RECT 86.605 1.565 86.775 1.735 ;
      RECT 86.605 3.155 86.775 3.325 ;
      RECT 86.55 8.605 86.72 8.775 ;
      RECT 86.24 6.685 86.41 6.855 ;
      RECT 86.225 2.745 86.395 2.915 ;
      RECT 86.145 1.565 86.315 1.735 ;
      RECT 86.005 3.315 86.175 3.485 ;
      RECT 85.985 3.715 86.155 3.885 ;
      RECT 85.87 8.605 86.04 8.775 ;
      RECT 85.815 2.265 85.985 2.435 ;
      RECT 85.81 7.055 85.98 7.225 ;
      RECT 85.81 7.795 85.98 7.965 ;
      RECT 85.685 1.565 85.855 1.735 ;
      RECT 85.435 6.315 85.605 6.485 ;
      RECT 85.315 3.245 85.485 3.415 ;
      RECT 85.225 1.565 85.395 1.735 ;
      RECT 85.19 8.605 85.36 8.775 ;
      RECT 84.995 2.935 85.165 3.105 ;
      RECT 84.925 3.715 85.095 3.885 ;
      RECT 84.765 1.565 84.935 1.735 ;
      RECT 84.525 3.695 84.695 3.865 ;
      RECT 84.51 8.605 84.68 8.775 ;
      RECT 84.485 2.185 84.655 2.355 ;
      RECT 84.305 1.565 84.475 1.735 ;
      RECT 83.845 1.565 84.015 1.735 ;
      RECT 83.585 2.685 83.755 2.855 ;
      RECT 83.585 3.145 83.755 3.315 ;
      RECT 83.585 3.655 83.755 3.825 ;
      RECT 83.475 2.215 83.645 2.385 ;
      RECT 83.385 1.565 83.555 1.735 ;
      RECT 83.005 3.725 83.175 3.895 ;
      RECT 82.925 1.565 83.095 1.735 ;
      RECT 82.525 2.255 82.695 2.425 ;
      RECT 82.465 1.565 82.635 1.735 ;
      RECT 82.315 2.635 82.485 2.805 ;
      RECT 82.005 1.565 82.175 1.735 ;
      RECT 81.815 3.235 81.985 3.405 ;
      RECT 81.695 2.685 81.865 2.855 ;
      RECT 81.545 1.565 81.715 1.735 ;
      RECT 81.525 2.135 81.695 2.305 ;
      RECT 81.155 3.165 81.325 3.335 ;
      RECT 81.085 1.565 81.255 1.735 ;
      RECT 80.665 2.765 80.835 2.935 ;
      RECT 80.625 1.565 80.795 1.735 ;
      RECT 80.615 3.535 80.785 3.705 ;
      RECT 80.165 1.565 80.335 1.735 ;
      RECT 80.125 3.165 80.295 3.335 ;
      RECT 80.095 2.265 80.265 2.435 ;
      RECT 79.735 2.665 79.905 2.835 ;
      RECT 79.705 1.565 79.875 1.735 ;
      RECT 79.525 3.475 79.695 3.645 ;
      RECT 79.245 1.565 79.415 1.735 ;
      RECT 79.225 2.905 79.395 3.075 ;
      RECT 78.785 1.565 78.955 1.735 ;
      RECT 78.525 2.695 78.695 2.865 ;
      RECT 78.325 1.565 78.495 1.735 ;
      RECT 78.205 3.145 78.375 3.315 ;
      RECT 77.865 1.565 78.035 1.735 ;
      RECT 77.785 3.175 77.955 3.345 ;
      RECT 77.615 2.165 77.785 2.335 ;
      RECT 77.445 2.615 77.615 2.785 ;
      RECT 77.405 1.565 77.575 1.735 ;
      RECT 76.945 1.565 77.115 1.735 ;
      RECT 76.525 2.265 76.695 2.435 ;
      RECT 76.515 3.585 76.685 3.755 ;
      RECT 76.485 1.565 76.655 1.735 ;
      RECT 75.425 7.8 75.595 7.97 ;
      RECT 75.075 0.1 75.245 0.27 ;
      RECT 75.075 8.61 75.245 8.78 ;
      RECT 75.055 2.76 75.225 2.93 ;
      RECT 75.055 5.95 75.225 6.12 ;
      RECT 74.435 0.91 74.605 1.08 ;
      RECT 74.435 2.39 74.605 2.56 ;
      RECT 74.435 6.32 74.605 6.49 ;
      RECT 74.435 7.8 74.605 7.97 ;
      RECT 74.085 0.1 74.255 0.27 ;
      RECT 74.085 8.61 74.255 8.78 ;
      RECT 74.065 2.76 74.235 2.93 ;
      RECT 74.065 5.95 74.235 6.12 ;
      RECT 73.385 0.105 73.555 0.275 ;
      RECT 73.385 8.605 73.555 8.775 ;
      RECT 73.075 2.025 73.245 2.195 ;
      RECT 73.075 6.685 73.245 6.855 ;
      RECT 72.705 0.105 72.875 0.275 ;
      RECT 72.705 8.605 72.875 8.775 ;
      RECT 72.645 0.915 72.815 1.085 ;
      RECT 72.645 1.655 72.815 1.825 ;
      RECT 72.645 7.055 72.815 7.225 ;
      RECT 72.645 7.795 72.815 7.965 ;
      RECT 72.27 2.395 72.44 2.565 ;
      RECT 72.27 6.315 72.44 6.485 ;
      RECT 72.025 0.105 72.195 0.275 ;
      RECT 72.025 8.605 72.195 8.775 ;
      RECT 71.345 0.105 71.515 0.275 ;
      RECT 71.345 8.605 71.515 8.775 ;
      RECT 70.06 1.565 70.23 1.735 ;
      RECT 69.6 1.565 69.77 1.735 ;
      RECT 69.21 2.905 69.38 3.075 ;
      RECT 69.14 1.565 69.31 1.735 ;
      RECT 69 2.245 69.17 2.415 ;
      RECT 68.68 1.565 68.85 1.735 ;
      RECT 68.68 3.155 68.85 3.325 ;
      RECT 68.625 8.605 68.795 8.775 ;
      RECT 68.315 6.685 68.485 6.855 ;
      RECT 68.3 2.745 68.47 2.915 ;
      RECT 68.22 1.565 68.39 1.735 ;
      RECT 68.08 3.315 68.25 3.485 ;
      RECT 68.06 3.715 68.23 3.885 ;
      RECT 67.945 8.605 68.115 8.775 ;
      RECT 67.89 2.265 68.06 2.435 ;
      RECT 67.885 7.055 68.055 7.225 ;
      RECT 67.885 7.795 68.055 7.965 ;
      RECT 67.76 1.565 67.93 1.735 ;
      RECT 67.51 6.315 67.68 6.485 ;
      RECT 67.39 3.245 67.56 3.415 ;
      RECT 67.3 1.565 67.47 1.735 ;
      RECT 67.265 8.605 67.435 8.775 ;
      RECT 67.07 2.935 67.24 3.105 ;
      RECT 67 3.715 67.17 3.885 ;
      RECT 66.84 1.565 67.01 1.735 ;
      RECT 66.6 3.695 66.77 3.865 ;
      RECT 66.585 8.605 66.755 8.775 ;
      RECT 66.56 2.185 66.73 2.355 ;
      RECT 66.38 1.565 66.55 1.735 ;
      RECT 65.92 1.565 66.09 1.735 ;
      RECT 65.66 2.685 65.83 2.855 ;
      RECT 65.66 3.145 65.83 3.315 ;
      RECT 65.66 3.655 65.83 3.825 ;
      RECT 65.55 2.215 65.72 2.385 ;
      RECT 65.46 1.565 65.63 1.735 ;
      RECT 65.08 3.725 65.25 3.895 ;
      RECT 65 1.565 65.17 1.735 ;
      RECT 64.6 2.255 64.77 2.425 ;
      RECT 64.54 1.565 64.71 1.735 ;
      RECT 64.39 2.635 64.56 2.805 ;
      RECT 64.08 1.565 64.25 1.735 ;
      RECT 63.89 3.235 64.06 3.405 ;
      RECT 63.77 2.685 63.94 2.855 ;
      RECT 63.62 1.565 63.79 1.735 ;
      RECT 63.6 2.135 63.77 2.305 ;
      RECT 63.23 3.165 63.4 3.335 ;
      RECT 63.16 1.565 63.33 1.735 ;
      RECT 62.74 2.765 62.91 2.935 ;
      RECT 62.7 1.565 62.87 1.735 ;
      RECT 62.69 3.535 62.86 3.705 ;
      RECT 62.24 1.565 62.41 1.735 ;
      RECT 62.2 3.165 62.37 3.335 ;
      RECT 62.17 2.265 62.34 2.435 ;
      RECT 61.81 2.665 61.98 2.835 ;
      RECT 61.78 1.565 61.95 1.735 ;
      RECT 61.6 3.475 61.77 3.645 ;
      RECT 61.32 1.565 61.49 1.735 ;
      RECT 61.3 2.905 61.47 3.075 ;
      RECT 60.86 1.565 61.03 1.735 ;
      RECT 60.6 2.695 60.77 2.865 ;
      RECT 60.4 1.565 60.57 1.735 ;
      RECT 60.28 3.145 60.45 3.315 ;
      RECT 59.94 1.565 60.11 1.735 ;
      RECT 59.86 3.175 60.03 3.345 ;
      RECT 59.69 2.165 59.86 2.335 ;
      RECT 59.52 2.615 59.69 2.785 ;
      RECT 59.48 1.565 59.65 1.735 ;
      RECT 59.02 1.565 59.19 1.735 ;
      RECT 58.6 2.265 58.77 2.435 ;
      RECT 58.59 3.585 58.76 3.755 ;
      RECT 58.56 1.565 58.73 1.735 ;
      RECT 57.5 7.8 57.67 7.97 ;
      RECT 57.15 0.1 57.32 0.27 ;
      RECT 57.15 8.61 57.32 8.78 ;
      RECT 57.13 2.76 57.3 2.93 ;
      RECT 57.13 5.95 57.3 6.12 ;
      RECT 56.51 0.91 56.68 1.08 ;
      RECT 56.51 2.39 56.68 2.56 ;
      RECT 56.51 6.32 56.68 6.49 ;
      RECT 56.51 7.8 56.68 7.97 ;
      RECT 56.16 0.1 56.33 0.27 ;
      RECT 56.16 8.61 56.33 8.78 ;
      RECT 56.14 2.76 56.31 2.93 ;
      RECT 56.14 5.95 56.31 6.12 ;
      RECT 55.46 0.105 55.63 0.275 ;
      RECT 55.46 8.605 55.63 8.775 ;
      RECT 55.15 2.025 55.32 2.195 ;
      RECT 55.15 6.685 55.32 6.855 ;
      RECT 54.78 0.105 54.95 0.275 ;
      RECT 54.78 8.605 54.95 8.775 ;
      RECT 54.72 0.915 54.89 1.085 ;
      RECT 54.72 1.655 54.89 1.825 ;
      RECT 54.72 7.055 54.89 7.225 ;
      RECT 54.72 7.795 54.89 7.965 ;
      RECT 54.345 2.395 54.515 2.565 ;
      RECT 54.345 6.315 54.515 6.485 ;
      RECT 54.1 0.105 54.27 0.275 ;
      RECT 54.1 8.605 54.27 8.775 ;
      RECT 53.42 0.105 53.59 0.275 ;
      RECT 53.42 8.605 53.59 8.775 ;
      RECT 52.135 1.565 52.305 1.735 ;
      RECT 51.675 1.565 51.845 1.735 ;
      RECT 51.285 2.905 51.455 3.075 ;
      RECT 51.215 1.565 51.385 1.735 ;
      RECT 51.075 2.245 51.245 2.415 ;
      RECT 50.755 1.565 50.925 1.735 ;
      RECT 50.755 3.155 50.925 3.325 ;
      RECT 50.7 8.605 50.87 8.775 ;
      RECT 50.39 6.685 50.56 6.855 ;
      RECT 50.375 2.745 50.545 2.915 ;
      RECT 50.295 1.565 50.465 1.735 ;
      RECT 50.155 3.315 50.325 3.485 ;
      RECT 50.135 3.715 50.305 3.885 ;
      RECT 50.02 8.605 50.19 8.775 ;
      RECT 49.965 2.265 50.135 2.435 ;
      RECT 49.96 7.055 50.13 7.225 ;
      RECT 49.96 7.795 50.13 7.965 ;
      RECT 49.835 1.565 50.005 1.735 ;
      RECT 49.585 6.315 49.755 6.485 ;
      RECT 49.465 3.245 49.635 3.415 ;
      RECT 49.375 1.565 49.545 1.735 ;
      RECT 49.34 8.605 49.51 8.775 ;
      RECT 49.145 2.935 49.315 3.105 ;
      RECT 49.075 3.715 49.245 3.885 ;
      RECT 48.915 1.565 49.085 1.735 ;
      RECT 48.675 3.695 48.845 3.865 ;
      RECT 48.66 8.605 48.83 8.775 ;
      RECT 48.635 2.185 48.805 2.355 ;
      RECT 48.455 1.565 48.625 1.735 ;
      RECT 47.995 1.565 48.165 1.735 ;
      RECT 47.735 2.685 47.905 2.855 ;
      RECT 47.735 3.145 47.905 3.315 ;
      RECT 47.735 3.655 47.905 3.825 ;
      RECT 47.625 2.215 47.795 2.385 ;
      RECT 47.535 1.565 47.705 1.735 ;
      RECT 47.155 3.725 47.325 3.895 ;
      RECT 47.075 1.565 47.245 1.735 ;
      RECT 46.675 2.255 46.845 2.425 ;
      RECT 46.615 1.565 46.785 1.735 ;
      RECT 46.465 2.635 46.635 2.805 ;
      RECT 46.155 1.565 46.325 1.735 ;
      RECT 45.965 3.235 46.135 3.405 ;
      RECT 45.845 2.685 46.015 2.855 ;
      RECT 45.695 1.565 45.865 1.735 ;
      RECT 45.675 2.135 45.845 2.305 ;
      RECT 45.305 3.165 45.475 3.335 ;
      RECT 45.235 1.565 45.405 1.735 ;
      RECT 44.815 2.765 44.985 2.935 ;
      RECT 44.775 1.565 44.945 1.735 ;
      RECT 44.765 3.535 44.935 3.705 ;
      RECT 44.315 1.565 44.485 1.735 ;
      RECT 44.275 3.165 44.445 3.335 ;
      RECT 44.245 2.265 44.415 2.435 ;
      RECT 43.885 2.665 44.055 2.835 ;
      RECT 43.855 1.565 44.025 1.735 ;
      RECT 43.675 3.475 43.845 3.645 ;
      RECT 43.395 1.565 43.565 1.735 ;
      RECT 43.375 2.905 43.545 3.075 ;
      RECT 42.935 1.565 43.105 1.735 ;
      RECT 42.675 2.695 42.845 2.865 ;
      RECT 42.475 1.565 42.645 1.735 ;
      RECT 42.355 3.145 42.525 3.315 ;
      RECT 42.015 1.565 42.185 1.735 ;
      RECT 41.935 3.175 42.105 3.345 ;
      RECT 41.765 2.165 41.935 2.335 ;
      RECT 41.595 2.615 41.765 2.785 ;
      RECT 41.555 1.565 41.725 1.735 ;
      RECT 41.095 1.565 41.265 1.735 ;
      RECT 40.675 2.265 40.845 2.435 ;
      RECT 40.665 3.585 40.835 3.755 ;
      RECT 40.635 1.565 40.805 1.735 ;
      RECT 39.575 7.8 39.745 7.97 ;
      RECT 39.225 0.1 39.395 0.27 ;
      RECT 39.225 8.61 39.395 8.78 ;
      RECT 39.205 2.76 39.375 2.93 ;
      RECT 39.205 5.95 39.375 6.12 ;
      RECT 38.585 0.91 38.755 1.08 ;
      RECT 38.585 2.39 38.755 2.56 ;
      RECT 38.585 6.32 38.755 6.49 ;
      RECT 38.585 7.8 38.755 7.97 ;
      RECT 38.235 0.1 38.405 0.27 ;
      RECT 38.235 8.61 38.405 8.78 ;
      RECT 38.215 2.76 38.385 2.93 ;
      RECT 38.215 5.95 38.385 6.12 ;
      RECT 37.535 0.105 37.705 0.275 ;
      RECT 37.535 8.605 37.705 8.775 ;
      RECT 37.225 2.025 37.395 2.195 ;
      RECT 37.225 6.685 37.395 6.855 ;
      RECT 36.855 0.105 37.025 0.275 ;
      RECT 36.855 8.605 37.025 8.775 ;
      RECT 36.795 0.915 36.965 1.085 ;
      RECT 36.795 1.655 36.965 1.825 ;
      RECT 36.795 7.055 36.965 7.225 ;
      RECT 36.795 7.795 36.965 7.965 ;
      RECT 36.42 2.395 36.59 2.565 ;
      RECT 36.42 6.315 36.59 6.485 ;
      RECT 36.175 0.105 36.345 0.275 ;
      RECT 36.175 8.605 36.345 8.775 ;
      RECT 35.495 0.105 35.665 0.275 ;
      RECT 35.495 8.605 35.665 8.775 ;
      RECT 34.21 1.565 34.38 1.735 ;
      RECT 33.75 1.565 33.92 1.735 ;
      RECT 33.36 2.905 33.53 3.075 ;
      RECT 33.29 1.565 33.46 1.735 ;
      RECT 33.15 2.245 33.32 2.415 ;
      RECT 32.83 1.565 33 1.735 ;
      RECT 32.83 3.155 33 3.325 ;
      RECT 32.775 8.605 32.945 8.775 ;
      RECT 32.465 6.685 32.635 6.855 ;
      RECT 32.45 2.745 32.62 2.915 ;
      RECT 32.37 1.565 32.54 1.735 ;
      RECT 32.23 3.315 32.4 3.485 ;
      RECT 32.21 3.715 32.38 3.885 ;
      RECT 32.095 8.605 32.265 8.775 ;
      RECT 32.04 2.265 32.21 2.435 ;
      RECT 32.035 7.055 32.205 7.225 ;
      RECT 32.035 7.795 32.205 7.965 ;
      RECT 31.91 1.565 32.08 1.735 ;
      RECT 31.66 6.315 31.83 6.485 ;
      RECT 31.54 3.245 31.71 3.415 ;
      RECT 31.45 1.565 31.62 1.735 ;
      RECT 31.415 8.605 31.585 8.775 ;
      RECT 31.22 2.935 31.39 3.105 ;
      RECT 31.15 3.715 31.32 3.885 ;
      RECT 30.99 1.565 31.16 1.735 ;
      RECT 30.75 3.695 30.92 3.865 ;
      RECT 30.735 8.605 30.905 8.775 ;
      RECT 30.71 2.185 30.88 2.355 ;
      RECT 30.53 1.565 30.7 1.735 ;
      RECT 30.07 1.565 30.24 1.735 ;
      RECT 29.81 2.685 29.98 2.855 ;
      RECT 29.81 3.145 29.98 3.315 ;
      RECT 29.81 3.655 29.98 3.825 ;
      RECT 29.7 2.215 29.87 2.385 ;
      RECT 29.61 1.565 29.78 1.735 ;
      RECT 29.23 3.725 29.4 3.895 ;
      RECT 29.15 1.565 29.32 1.735 ;
      RECT 28.75 2.255 28.92 2.425 ;
      RECT 28.69 1.565 28.86 1.735 ;
      RECT 28.54 2.635 28.71 2.805 ;
      RECT 28.23 1.565 28.4 1.735 ;
      RECT 28.04 3.235 28.21 3.405 ;
      RECT 27.92 2.685 28.09 2.855 ;
      RECT 27.77 1.565 27.94 1.735 ;
      RECT 27.75 2.135 27.92 2.305 ;
      RECT 27.38 3.165 27.55 3.335 ;
      RECT 27.31 1.565 27.48 1.735 ;
      RECT 26.89 2.765 27.06 2.935 ;
      RECT 26.85 1.565 27.02 1.735 ;
      RECT 26.84 3.535 27.01 3.705 ;
      RECT 26.39 1.565 26.56 1.735 ;
      RECT 26.35 3.165 26.52 3.335 ;
      RECT 26.32 2.265 26.49 2.435 ;
      RECT 25.96 2.665 26.13 2.835 ;
      RECT 25.93 1.565 26.1 1.735 ;
      RECT 25.75 3.475 25.92 3.645 ;
      RECT 25.47 1.565 25.64 1.735 ;
      RECT 25.45 2.905 25.62 3.075 ;
      RECT 25.01 1.565 25.18 1.735 ;
      RECT 24.75 2.695 24.92 2.865 ;
      RECT 24.55 1.565 24.72 1.735 ;
      RECT 24.43 3.145 24.6 3.315 ;
      RECT 24.09 1.565 24.26 1.735 ;
      RECT 24.01 3.175 24.18 3.345 ;
      RECT 23.84 2.165 24.01 2.335 ;
      RECT 23.67 2.615 23.84 2.785 ;
      RECT 23.63 1.565 23.8 1.735 ;
      RECT 23.17 1.565 23.34 1.735 ;
      RECT 22.75 2.265 22.92 2.435 ;
      RECT 22.74 3.585 22.91 3.755 ;
      RECT 22.71 1.565 22.88 1.735 ;
      RECT 21.65 7.8 21.82 7.97 ;
      RECT 21.3 0.1 21.47 0.27 ;
      RECT 21.3 8.61 21.47 8.78 ;
      RECT 21.28 2.76 21.45 2.93 ;
      RECT 21.28 5.95 21.45 6.12 ;
      RECT 20.66 0.91 20.83 1.08 ;
      RECT 20.66 2.39 20.83 2.56 ;
      RECT 20.66 6.32 20.83 6.49 ;
      RECT 20.66 7.8 20.83 7.97 ;
      RECT 20.31 0.1 20.48 0.27 ;
      RECT 20.31 8.61 20.48 8.78 ;
      RECT 20.29 2.76 20.46 2.93 ;
      RECT 20.29 5.95 20.46 6.12 ;
      RECT 19.61 0.105 19.78 0.275 ;
      RECT 19.61 8.605 19.78 8.775 ;
      RECT 19.3 2.025 19.47 2.195 ;
      RECT 19.3 6.685 19.47 6.855 ;
      RECT 18.93 0.105 19.1 0.275 ;
      RECT 18.93 8.605 19.1 8.775 ;
      RECT 18.87 0.915 19.04 1.085 ;
      RECT 18.87 1.655 19.04 1.825 ;
      RECT 18.87 7.055 19.04 7.225 ;
      RECT 18.87 7.795 19.04 7.965 ;
      RECT 18.495 2.395 18.665 2.565 ;
      RECT 18.495 6.315 18.665 6.485 ;
      RECT 18.25 0.105 18.42 0.275 ;
      RECT 18.25 8.605 18.42 8.775 ;
      RECT 17.57 0.105 17.74 0.275 ;
      RECT 17.57 8.605 17.74 8.775 ;
      RECT 16.285 1.565 16.455 1.735 ;
      RECT 15.825 1.565 15.995 1.735 ;
      RECT 15.435 2.905 15.605 3.075 ;
      RECT 15.365 1.565 15.535 1.735 ;
      RECT 15.225 2.245 15.395 2.415 ;
      RECT 14.905 1.565 15.075 1.735 ;
      RECT 14.905 3.155 15.075 3.325 ;
      RECT 14.85 8.605 15.02 8.775 ;
      RECT 14.54 6.685 14.71 6.855 ;
      RECT 14.525 2.745 14.695 2.915 ;
      RECT 14.445 1.565 14.615 1.735 ;
      RECT 14.305 3.315 14.475 3.485 ;
      RECT 14.285 3.715 14.455 3.885 ;
      RECT 14.17 8.605 14.34 8.775 ;
      RECT 14.115 2.265 14.285 2.435 ;
      RECT 14.11 7.055 14.28 7.225 ;
      RECT 14.11 7.795 14.28 7.965 ;
      RECT 13.985 1.565 14.155 1.735 ;
      RECT 13.735 6.315 13.905 6.485 ;
      RECT 13.615 3.245 13.785 3.415 ;
      RECT 13.525 1.565 13.695 1.735 ;
      RECT 13.49 8.605 13.66 8.775 ;
      RECT 13.295 2.935 13.465 3.105 ;
      RECT 13.225 3.715 13.395 3.885 ;
      RECT 13.065 1.565 13.235 1.735 ;
      RECT 12.825 3.695 12.995 3.865 ;
      RECT 12.81 8.605 12.98 8.775 ;
      RECT 12.785 2.185 12.955 2.355 ;
      RECT 12.605 1.565 12.775 1.735 ;
      RECT 12.145 1.565 12.315 1.735 ;
      RECT 11.885 2.685 12.055 2.855 ;
      RECT 11.885 3.145 12.055 3.315 ;
      RECT 11.885 3.655 12.055 3.825 ;
      RECT 11.775 2.215 11.945 2.385 ;
      RECT 11.685 1.565 11.855 1.735 ;
      RECT 11.305 3.725 11.475 3.895 ;
      RECT 11.225 1.565 11.395 1.735 ;
      RECT 10.825 2.255 10.995 2.425 ;
      RECT 10.765 1.565 10.935 1.735 ;
      RECT 10.615 2.635 10.785 2.805 ;
      RECT 10.305 1.565 10.475 1.735 ;
      RECT 10.115 3.235 10.285 3.405 ;
      RECT 9.995 2.685 10.165 2.855 ;
      RECT 9.845 1.565 10.015 1.735 ;
      RECT 9.825 2.135 9.995 2.305 ;
      RECT 9.455 3.165 9.625 3.335 ;
      RECT 9.385 1.565 9.555 1.735 ;
      RECT 8.965 2.765 9.135 2.935 ;
      RECT 8.925 1.565 9.095 1.735 ;
      RECT 8.915 3.535 9.085 3.705 ;
      RECT 8.465 1.565 8.635 1.735 ;
      RECT 8.425 3.165 8.595 3.335 ;
      RECT 8.395 2.265 8.565 2.435 ;
      RECT 8.035 2.665 8.205 2.835 ;
      RECT 8.005 1.565 8.175 1.735 ;
      RECT 7.825 3.475 7.995 3.645 ;
      RECT 7.545 1.565 7.715 1.735 ;
      RECT 7.525 2.905 7.695 3.075 ;
      RECT 7.085 1.565 7.255 1.735 ;
      RECT 6.825 2.695 6.995 2.865 ;
      RECT 6.625 1.565 6.795 1.735 ;
      RECT 6.505 3.145 6.675 3.315 ;
      RECT 6.165 1.565 6.335 1.735 ;
      RECT 6.085 3.175 6.255 3.345 ;
      RECT 5.915 2.165 6.085 2.335 ;
      RECT 5.745 2.615 5.915 2.785 ;
      RECT 5.705 1.565 5.875 1.735 ;
      RECT 5.245 1.565 5.415 1.735 ;
      RECT 4.825 2.265 4.995 2.435 ;
      RECT 4.815 3.585 4.985 3.755 ;
      RECT 4.785 1.565 4.955 1.735 ;
      RECT 3.82 8.605 3.99 8.775 ;
      RECT 3.14 8.605 3.31 8.775 ;
      RECT 3.08 7.055 3.25 7.225 ;
      RECT 3.08 7.795 3.25 7.965 ;
      RECT 2.705 6.315 2.875 6.485 ;
      RECT 2.46 8.605 2.63 8.775 ;
      RECT 1.78 8.605 1.95 8.775 ;
    LAYER li1 ;
      RECT 87.395 0 87.565 2.235 ;
      RECT 86.435 0 86.605 2.235 ;
      RECT 85.475 0 85.645 2.235 ;
      RECT 84.955 0 85.125 2.235 ;
      RECT 83.995 0 84.165 2.235 ;
      RECT 82.995 0 83.165 2.235 ;
      RECT 82.035 0 82.205 2.235 ;
      RECT 80.555 0 80.725 2.235 ;
      RECT 78.635 0 78.805 2.235 ;
      RECT 77.155 0 77.325 2.235 ;
      RECT 69.47 0 69.64 2.235 ;
      RECT 68.51 0 68.68 2.235 ;
      RECT 67.55 0 67.72 2.235 ;
      RECT 67.03 0 67.2 2.235 ;
      RECT 66.07 0 66.24 2.235 ;
      RECT 65.07 0 65.24 2.235 ;
      RECT 64.11 0 64.28 2.235 ;
      RECT 62.63 0 62.8 2.235 ;
      RECT 60.71 0 60.88 2.235 ;
      RECT 59.23 0 59.4 2.235 ;
      RECT 51.545 0 51.715 2.235 ;
      RECT 50.585 0 50.755 2.235 ;
      RECT 49.625 0 49.795 2.235 ;
      RECT 49.105 0 49.275 2.235 ;
      RECT 48.145 0 48.315 2.235 ;
      RECT 47.145 0 47.315 2.235 ;
      RECT 46.185 0 46.355 2.235 ;
      RECT 44.705 0 44.875 2.235 ;
      RECT 42.785 0 42.955 2.235 ;
      RECT 41.305 0 41.475 2.235 ;
      RECT 33.62 0 33.79 2.235 ;
      RECT 32.66 0 32.83 2.235 ;
      RECT 31.7 0 31.87 2.235 ;
      RECT 31.18 0 31.35 2.235 ;
      RECT 30.22 0 30.39 2.235 ;
      RECT 29.22 0 29.39 2.235 ;
      RECT 28.26 0 28.43 2.235 ;
      RECT 26.78 0 26.95 2.235 ;
      RECT 24.86 0 25.03 2.235 ;
      RECT 23.38 0 23.55 2.235 ;
      RECT 15.695 0 15.865 2.235 ;
      RECT 14.735 0 14.905 2.235 ;
      RECT 13.775 0 13.945 2.235 ;
      RECT 13.255 0 13.425 2.235 ;
      RECT 12.295 0 12.465 2.235 ;
      RECT 11.295 0 11.465 2.235 ;
      RECT 10.335 0 10.505 2.235 ;
      RECT 8.855 0 9.025 2.235 ;
      RECT 6.935 0 7.105 2.235 ;
      RECT 5.455 0 5.625 2.235 ;
      RECT 76.345 0 88.305 1.735 ;
      RECT 58.42 0 70.38 1.735 ;
      RECT 40.495 0 52.455 1.735 ;
      RECT 22.57 0 34.53 1.735 ;
      RECT 4.645 0 16.605 1.735 ;
      RECT 76.34 0 88.305 1.68 ;
      RECT 58.415 0 70.38 1.68 ;
      RECT 40.49 0 52.455 1.68 ;
      RECT 22.565 0 34.53 1.68 ;
      RECT 4.64 0 16.605 1.68 ;
      RECT 89.19 0 89.36 0.935 ;
      RECT 71.265 0 71.435 0.935 ;
      RECT 53.34 0 53.51 0.935 ;
      RECT 35.415 0 35.585 0.935 ;
      RECT 17.49 0 17.66 0.935 ;
      RECT 92.92 0 93.09 0.93 ;
      RECT 91.93 0 92.1 0.93 ;
      RECT 74.995 0 75.165 0.93 ;
      RECT 74.005 0 74.175 0.93 ;
      RECT 57.07 0 57.24 0.93 ;
      RECT 56.08 0 56.25 0.93 ;
      RECT 39.145 0 39.315 0.93 ;
      RECT 38.155 0 38.325 0.93 ;
      RECT 21.22 0 21.39 0.93 ;
      RECT 20.23 0 20.4 0.93 ;
      RECT 93.715 0 93.895 0.305 ;
      RECT 75.79 0 91.765 0.305 ;
      RECT 57.865 0 73.84 0.305 ;
      RECT 39.94 0 55.915 0.305 ;
      RECT 22.015 0 37.99 0.305 ;
      RECT 1.48 0 20.065 0.305 ;
      RECT 1.48 0 93.895 0.3 ;
      RECT 1.46 8.58 93.895 8.88 ;
      RECT 93.715 8.575 93.895 8.88 ;
      RECT 92.92 7.95 93.09 8.88 ;
      RECT 91.93 7.95 92.1 8.88 ;
      RECT 75.79 8.575 91.765 8.88 ;
      RECT 74.995 7.95 75.165 8.88 ;
      RECT 74.005 7.95 74.175 8.88 ;
      RECT 57.865 8.575 73.84 8.88 ;
      RECT 57.07 7.95 57.24 8.88 ;
      RECT 56.08 7.95 56.25 8.88 ;
      RECT 39.94 8.575 55.915 8.88 ;
      RECT 39.145 7.95 39.315 8.88 ;
      RECT 38.155 7.95 38.325 8.88 ;
      RECT 22.015 8.575 37.99 8.88 ;
      RECT 21.22 7.95 21.39 8.88 ;
      RECT 20.23 7.95 20.4 8.88 ;
      RECT 1.46 8.575 20.065 8.88 ;
      RECT 89.19 7.945 89.36 8.88 ;
      RECT 84.43 7.945 84.6 8.88 ;
      RECT 71.265 7.945 71.435 8.88 ;
      RECT 66.505 7.945 66.675 8.88 ;
      RECT 53.34 7.945 53.51 8.88 ;
      RECT 48.58 7.945 48.75 8.88 ;
      RECT 35.415 7.945 35.585 8.88 ;
      RECT 30.655 7.945 30.825 8.88 ;
      RECT 17.49 7.945 17.66 8.88 ;
      RECT 12.73 7.945 12.9 8.88 ;
      RECT 1.46 8.565 2.265 8.88 ;
      RECT 1.7 8.545 1.925 8.88 ;
      RECT 1.7 7.945 1.87 8.88 ;
      RECT 93.35 5.02 93.52 6.49 ;
      RECT 93.35 6.315 93.525 6.485 ;
      RECT 92.98 1.74 93.15 2.93 ;
      RECT 92.98 1.74 93.45 1.91 ;
      RECT 92.98 6.97 93.45 7.14 ;
      RECT 92.98 5.95 93.15 7.14 ;
      RECT 91.99 1.74 92.16 2.93 ;
      RECT 91.99 1.74 92.46 1.91 ;
      RECT 91.99 6.97 92.46 7.14 ;
      RECT 91.99 5.95 92.16 7.14 ;
      RECT 90.14 2.635 90.31 3.865 ;
      RECT 90.195 0.855 90.365 2.805 ;
      RECT 90.14 0.575 90.31 1.025 ;
      RECT 90.14 7.855 90.31 8.305 ;
      RECT 90.195 6.075 90.365 8.025 ;
      RECT 90.14 5.015 90.31 6.245 ;
      RECT 89.62 0.575 89.79 3.865 ;
      RECT 89.62 2.075 90.025 2.405 ;
      RECT 89.62 1.235 90.025 1.565 ;
      RECT 89.62 5.015 89.79 8.305 ;
      RECT 89.62 7.315 90.025 7.645 ;
      RECT 89.62 6.475 90.025 6.805 ;
      RECT 87.715 3.39 87.735 3.44 ;
      RECT 87.695 3.362 87.715 3.555 ;
      RECT 87.675 3.337 87.695 3.611 ;
      RECT 87.635 3.325 87.675 3.63 ;
      RECT 87.585 3.32 87.635 3.659 ;
      RECT 87.581 3.314 87.585 3.675 ;
      RECT 87.495 3.306 87.581 3.675 ;
      RECT 87.435 3.294 87.495 3.67 ;
      RECT 87.381 3.284 87.435 3.659 ;
      RECT 87.295 3.272 87.381 3.642 ;
      RECT 87.273 3.263 87.295 3.629 ;
      RECT 87.187 3.256 87.273 3.616 ;
      RECT 87.101 3.243 87.187 3.595 ;
      RECT 87.015 3.231 87.101 3.575 ;
      RECT 86.985 3.22 87.015 3.561 ;
      RECT 86.935 3.207 86.985 3.551 ;
      RECT 86.915 3.197 86.935 3.545 ;
      RECT 86.861 3.187 86.915 3.539 ;
      RECT 86.775 3.167 86.861 3.523 ;
      RECT 86.735 3.155 86.775 3.509 ;
      RECT 86.7 3.155 86.735 3.495 ;
      RECT 86.685 3.155 86.7 3.48 ;
      RECT 86.635 3.155 86.685 3.425 ;
      RECT 86.605 3.155 86.635 3.345 ;
      RECT 87.135 2.825 87.305 3.075 ;
      RECT 87.135 2.825 87.315 3.03 ;
      RECT 87.195 2.655 87.325 2.975 ;
      RECT 87.195 2.662 87.335 2.94 ;
      RECT 87.155 2.677 87.345 2.875 ;
      RECT 87.145 2.76 87.345 2.875 ;
      RECT 87.155 2.695 87.355 2.785 ;
      RECT 87.155 2.675 87.335 2.94 ;
      RECT 86.925 1.93 87.095 2.415 ;
      RECT 86.915 1.93 87.095 2.405 ;
      RECT 86.915 1.945 87.115 2.35 ;
      RECT 86.875 1.925 87.065 2.315 ;
      RECT 86.875 1.96 87.125 2.235 ;
      RECT 86.825 1.945 87.115 2.135 ;
      RECT 86.825 1.975 87.135 2.095 ;
      RECT 86.825 1.99 87.145 2.015 ;
      RECT 86.421 2.688 86.435 2.944 ;
      RECT 86.421 2.689 86.521 2.939 ;
      RECT 86.335 2.686 86.421 2.936 ;
      RECT 86.325 2.685 86.335 2.929 ;
      RECT 86.325 2.692 86.607 2.926 ;
      RECT 86.245 2.695 86.607 2.922 ;
      RECT 86.325 2.694 86.625 2.919 ;
      RECT 86.235 2.707 86.645 2.916 ;
      RECT 86.245 2.695 86.645 2.916 ;
      RECT 86.225 2.712 86.645 2.915 ;
      RECT 86.245 2.697 86.731 2.911 ;
      RECT 86.205 2.715 86.731 2.908 ;
      RECT 86.245 2.701 86.817 2.902 ;
      RECT 86.195 2.72 86.817 2.898 ;
      RECT 86.245 2.704 86.845 2.897 ;
      RECT 86.245 2.705 86.885 2.891 ;
      RECT 86.235 2.71 86.895 2.886 ;
      RECT 86.195 2.73 86.905 2.875 ;
      RECT 86.195 2.75 86.915 2.86 ;
      RECT 86.155 3.298 86.175 3.605 ;
      RECT 86.145 3.273 86.155 3.885 ;
      RECT 86.105 3.24 86.145 3.885 ;
      RECT 86.101 3.21 86.105 3.885 ;
      RECT 86.015 3.095 86.101 3.885 ;
      RECT 86.005 2.97 86.015 3.885 ;
      RECT 85.995 2.935 86.005 3.885 ;
      RECT 85.985 2.905 85.995 3.885 ;
      RECT 85.965 2.875 85.985 3.77 ;
      RECT 85.955 2.845 85.965 3.645 ;
      RECT 85.945 2.825 85.955 3.595 ;
      RECT 85.925 2.795 85.945 3.503 ;
      RECT 85.905 2.761 85.925 3.418 ;
      RECT 85.9 2.744 85.905 3.353 ;
      RECT 85.895 2.738 85.9 3.325 ;
      RECT 85.885 2.73 85.895 3.29 ;
      RECT 85.865 2.725 85.875 3.19 ;
      RECT 85.855 2.725 85.865 3.165 ;
      RECT 85.85 2.725 85.855 3.128 ;
      RECT 85.835 2.725 85.85 3.06 ;
      RECT 85.825 2.724 85.835 2.99 ;
      RECT 85.815 2.722 85.825 2.97 ;
      RECT 85.755 2.718 85.815 2.943 ;
      RECT 85.715 2.72 85.755 2.923 ;
      RECT 85.695 2.75 85.715 2.905 ;
      RECT 85.875 2.725 85.885 3.245 ;
      RECT 85.815 2.08 85.985 2.435 ;
      RECT 85.845 1.966 85.985 2.435 ;
      RECT 85.845 1.968 85.995 2.43 ;
      RECT 85.845 1.97 86.015 2.42 ;
      RECT 85.845 1.973 86.045 2.405 ;
      RECT 85.845 1.978 86.095 2.375 ;
      RECT 85.845 1.983 86.115 2.338 ;
      RECT 85.825 1.985 86.125 2.313 ;
      RECT 85.845 1.965 85.955 2.435 ;
      RECT 85.855 1.96 85.955 2.435 ;
      RECT 85.375 3.222 85.565 3.585 ;
      RECT 85.375 3.237 85.605 3.583 ;
      RECT 85.375 3.265 85.625 3.579 ;
      RECT 85.375 3.3 85.635 3.577 ;
      RECT 85.375 3.345 85.645 3.576 ;
      RECT 85.365 3.217 85.525 3.565 ;
      RECT 85.345 3.225 85.565 3.515 ;
      RECT 85.315 3.237 85.605 3.45 ;
      RECT 85.375 3.215 85.525 3.585 ;
      RECT 85.38 7.855 85.55 8.305 ;
      RECT 85.435 6.075 85.605 8.025 ;
      RECT 85.38 5.015 85.55 6.245 ;
      RECT 84.86 5.015 85.03 8.305 ;
      RECT 84.86 7.315 85.265 7.645 ;
      RECT 84.86 6.475 85.265 6.805 ;
      RECT 84.961 2.695 85.165 3.105 ;
      RECT 84.875 2.588 84.961 3.09 ;
      RECT 84.871 2.584 84.875 3.074 ;
      RECT 84.785 2.695 85.165 3.054 ;
      RECT 84.765 2.575 84.785 3.015 ;
      RECT 84.755 2.58 84.871 2.99 ;
      RECT 84.745 2.587 84.875 2.97 ;
      RECT 84.735 2.592 84.965 2.945 ;
      RECT 84.725 2.61 85.055 2.925 ;
      RECT 84.715 2.615 85.055 2.905 ;
      RECT 84.705 2.62 85.095 2.77 ;
      RECT 84.705 2.65 85.155 2.77 ;
      RECT 84.705 2.635 85.145 2.77 ;
      RECT 84.735 2.605 85.055 2.945 ;
      RECT 84.735 2.593 84.995 2.945 ;
      RECT 84.885 3.42 85.135 3.885 ;
      RECT 84.805 3.395 85.125 3.88 ;
      RECT 84.735 3.429 85.135 3.87 ;
      RECT 84.525 3.68 85.135 3.865 ;
      RECT 84.705 3.449 85.135 3.865 ;
      RECT 84.545 3.64 85.135 3.865 ;
      RECT 84.695 3.46 85.135 3.865 ;
      RECT 84.585 3.58 85.135 3.865 ;
      RECT 84.635 3.505 85.135 3.865 ;
      RECT 84.885 3.37 85.125 3.885 ;
      RECT 84.905 3.365 85.125 3.885 ;
      RECT 84.915 3.36 85.045 3.885 ;
      RECT 85.001 3.355 85.005 3.885 ;
      RECT 84.475 1.925 84.561 2.362 ;
      RECT 84.465 1.925 84.561 2.358 ;
      RECT 84.465 1.925 84.625 2.357 ;
      RECT 84.465 1.925 84.655 2.355 ;
      RECT 84.465 1.925 84.665 2.345 ;
      RECT 84.455 1.93 84.665 2.343 ;
      RECT 84.445 1.94 84.665 2.335 ;
      RECT 84.445 1.94 84.675 2.295 ;
      RECT 84.465 1.925 84.695 2.21 ;
      RECT 84.435 1.95 84.695 2.205 ;
      RECT 84.445 1.94 84.705 2.135 ;
      RECT 84.425 1.96 84.705 2.08 ;
      RECT 84.415 1.97 84.705 1.98 ;
      RECT 84.495 2.741 84.505 2.82 ;
      RECT 84.485 2.734 84.495 3.005 ;
      RECT 84.475 2.728 84.485 3.03 ;
      RECT 84.465 2.72 84.475 3.06 ;
      RECT 84.425 2.715 84.465 3.11 ;
      RECT 84.405 2.715 84.425 3.165 ;
      RECT 84.395 2.715 84.405 3.19 ;
      RECT 84.385 2.715 84.395 3.205 ;
      RECT 84.355 2.715 84.385 3.25 ;
      RECT 84.345 2.715 84.355 3.29 ;
      RECT 84.325 2.715 84.345 3.315 ;
      RECT 84.305 2.715 84.325 3.35 ;
      RECT 84.225 2.715 84.305 3.395 ;
      RECT 84.215 2.715 84.225 3.415 ;
      RECT 84.175 2.795 84.215 3.412 ;
      RECT 84.155 2.875 84.175 3.409 ;
      RECT 84.135 2.93 84.155 3.407 ;
      RECT 84.115 2.99 84.135 3.405 ;
      RECT 84.075 3.025 84.115 3.403 ;
      RECT 84.071 3.035 84.075 3.401 ;
      RECT 83.985 3.05 84.071 3.397 ;
      RECT 83.965 3.07 83.985 3.393 ;
      RECT 83.895 3.075 83.965 3.389 ;
      RECT 83.875 3.076 83.895 3.386 ;
      RECT 83.871 3.078 83.875 3.385 ;
      RECT 83.785 3.087 83.871 3.38 ;
      RECT 83.775 3.096 83.785 3.375 ;
      RECT 83.735 3.102 83.775 3.37 ;
      RECT 83.685 3.113 83.735 3.355 ;
      RECT 83.665 3.122 83.685 3.34 ;
      RECT 83.585 3.135 83.665 3.325 ;
      RECT 83.755 2.685 83.925 2.895 ;
      RECT 83.871 2.677 83.925 2.895 ;
      RECT 83.671 2.685 83.925 2.885 ;
      RECT 83.585 2.685 83.925 2.865 ;
      RECT 83.585 2.69 83.935 2.81 ;
      RECT 83.585 2.7 83.945 2.72 ;
      RECT 83.785 2.682 83.925 2.895 ;
      RECT 83.535 3.623 83.785 3.955 ;
      RECT 83.505 3.635 83.785 3.937 ;
      RECT 83.485 3.67 83.785 3.907 ;
      RECT 83.535 3.62 83.707 3.955 ;
      RECT 83.535 3.616 83.621 3.955 ;
      RECT 83.465 1.965 83.645 2.385 ;
      RECT 83.465 1.965 83.665 2.375 ;
      RECT 83.465 1.965 83.685 2.35 ;
      RECT 83.465 1.965 83.695 2.335 ;
      RECT 83.465 1.965 83.705 2.33 ;
      RECT 83.465 2.005 83.725 2.315 ;
      RECT 83.465 2.075 83.745 2.295 ;
      RECT 83.445 2.075 83.745 2.29 ;
      RECT 83.445 2.135 83.755 2.265 ;
      RECT 83.445 2.175 83.765 2.215 ;
      RECT 83.425 1.965 83.705 2.195 ;
      RECT 83.415 1.975 83.705 2.118 ;
      RECT 83.405 2.015 83.725 2.063 ;
      RECT 83.005 3.375 83.175 3.895 ;
      RECT 82.995 3.375 83.175 3.855 ;
      RECT 82.985 3.395 83.175 3.83 ;
      RECT 82.995 3.375 83.185 3.825 ;
      RECT 82.975 3.435 83.185 3.795 ;
      RECT 82.965 3.47 83.185 3.775 ;
      RECT 82.955 3.52 83.185 3.735 ;
      RECT 82.995 3.386 83.195 3.725 ;
      RECT 82.945 3.6 83.195 3.675 ;
      RECT 82.985 3.409 83.205 3.605 ;
      RECT 82.985 3.433 83.215 3.5 ;
      RECT 82.925 2.68 82.945 2.955 ;
      RECT 82.885 2.665 82.925 3 ;
      RECT 82.865 2.65 82.885 3.065 ;
      RECT 82.845 2.649 82.865 3.14 ;
      RECT 82.825 2.657 82.845 3.245 ;
      RECT 82.821 2.662 82.825 3.297 ;
      RECT 82.735 2.681 82.821 3.337 ;
      RECT 82.725 2.702 82.735 3.376 ;
      RECT 82.715 2.71 82.725 3.377 ;
      RECT 82.695 2.845 82.715 3.379 ;
      RECT 82.685 2.995 82.695 3.381 ;
      RECT 82.645 3.08 82.685 3.386 ;
      RECT 82.563 3.102 82.645 3.396 ;
      RECT 82.477 3.117 82.563 3.409 ;
      RECT 82.391 3.132 82.477 3.422 ;
      RECT 82.305 3.147 82.391 3.436 ;
      RECT 82.225 3.161 82.305 3.449 ;
      RECT 82.211 3.169 82.225 3.457 ;
      RECT 82.125 3.177 82.211 3.471 ;
      RECT 82.115 3.185 82.125 3.484 ;
      RECT 82.091 3.185 82.115 3.492 ;
      RECT 82.005 3.187 82.091 3.522 ;
      RECT 81.925 3.189 82.005 3.565 ;
      RECT 81.855 3.192 81.925 3.6 ;
      RECT 81.835 3.194 81.855 3.616 ;
      RECT 81.805 3.2 81.835 3.618 ;
      RECT 81.755 3.215 81.805 3.621 ;
      RECT 81.735 3.23 81.755 3.624 ;
      RECT 81.705 3.235 81.735 3.627 ;
      RECT 81.645 3.25 81.705 3.631 ;
      RECT 81.635 3.266 81.645 3.635 ;
      RECT 81.585 3.276 81.635 3.624 ;
      RECT 81.555 3.295 81.585 3.607 ;
      RECT 81.535 3.315 81.555 3.597 ;
      RECT 81.515 3.34 81.535 3.589 ;
      RECT 82.525 1.932 82.695 2.425 ;
      RECT 82.515 1.932 82.695 2.41 ;
      RECT 82.515 1.947 82.725 2.4 ;
      RECT 82.505 1.947 82.725 2.375 ;
      RECT 82.495 1.947 82.725 2.34 ;
      RECT 82.495 1.955 82.735 2.295 ;
      RECT 82.475 1.925 82.665 2.275 ;
      RECT 82.465 1.932 82.695 2.235 ;
      RECT 82.455 1.947 82.725 2.215 ;
      RECT 82.445 1.96 82.735 2.175 ;
      RECT 82.435 1.975 82.735 2.128 ;
      RECT 82.435 1.975 82.745 2.12 ;
      RECT 82.425 1.99 82.745 2.093 ;
      RECT 82.435 1.985 82.755 2.035 ;
      RECT 82.235 2.612 82.505 2.905 ;
      RECT 82.235 2.614 82.515 2.9 ;
      RECT 82.225 2.64 82.515 2.895 ;
      RECT 82.235 2.63 82.525 2.89 ;
      RECT 82.235 2.608 82.471 2.905 ;
      RECT 82.235 2.605 82.385 2.905 ;
      RECT 82.295 2.6 82.381 2.905 ;
      RECT 81.785 2.648 81.855 2.945 ;
      RECT 81.785 2.648 81.865 2.944 ;
      RECT 81.865 2.635 81.875 2.941 ;
      RECT 81.765 2.662 81.875 2.935 ;
      RECT 81.855 2.64 81.945 2.931 ;
      RECT 81.785 2.655 81.965 2.92 ;
      RECT 81.765 2.72 81.975 2.916 ;
      RECT 81.745 2.668 81.965 2.915 ;
      RECT 81.735 2.673 81.965 2.905 ;
      RECT 81.725 2.795 81.985 2.9 ;
      RECT 81.725 2.875 81.995 2.89 ;
      RECT 81.695 2.681 81.965 2.884 ;
      RECT 81.685 2.695 81.965 2.869 ;
      RECT 81.725 2.676 81.965 2.9 ;
      RECT 81.855 2.636 81.875 2.941 ;
      RECT 81.675 2.072 81.695 2.305 ;
      RECT 81.665 2.053 81.675 2.31 ;
      RECT 81.655 2.041 81.665 2.317 ;
      RECT 81.615 2.027 81.655 2.327 ;
      RECT 81.605 2.017 81.615 2.336 ;
      RECT 81.555 2.002 81.605 2.341 ;
      RECT 81.545 1.987 81.555 2.347 ;
      RECT 81.525 1.978 81.545 2.352 ;
      RECT 81.515 1.968 81.525 2.358 ;
      RECT 81.505 1.965 81.515 2.363 ;
      RECT 81.485 1.965 81.505 2.364 ;
      RECT 81.455 1.96 81.485 2.362 ;
      RECT 81.431 1.953 81.455 2.361 ;
      RECT 81.345 1.943 81.431 2.358 ;
      RECT 81.335 1.935 81.345 2.355 ;
      RECT 81.313 1.935 81.335 2.354 ;
      RECT 81.227 1.935 81.313 2.352 ;
      RECT 81.141 1.935 81.227 2.35 ;
      RECT 81.055 1.935 81.141 2.347 ;
      RECT 81.045 1.935 81.055 2.34 ;
      RECT 81.015 1.935 81.045 2.3 ;
      RECT 81.005 1.945 81.015 2.255 ;
      RECT 80.995 1.99 81.005 2.24 ;
      RECT 80.965 2.085 80.995 2.195 ;
      RECT 81.155 2.822 81.325 3.335 ;
      RECT 81.145 2.853 81.325 3.315 ;
      RECT 81.145 2.853 81.345 3.285 ;
      RECT 81.135 2.861 81.345 3.26 ;
      RECT 81.135 2.861 81.355 3.25 ;
      RECT 81.135 2.861 81.365 3.23 ;
      RECT 81.135 2.861 81.415 3.185 ;
      RECT 81.135 2.861 81.425 3.16 ;
      RECT 81.135 2.861 81.435 3.125 ;
      RECT 81.135 2.861 81.445 3.09 ;
      RECT 81.135 2.861 81.455 3.04 ;
      RECT 81.135 2.861 81.475 2.965 ;
      RECT 81.305 2.725 81.485 2.905 ;
      RECT 81.225 2.78 81.485 2.905 ;
      RECT 81.265 2.745 81.325 3.335 ;
      RECT 81.255 2.765 81.485 2.905 ;
      RECT 80.615 3.235 80.701 3.801 ;
      RECT 80.575 3.235 80.701 3.795 ;
      RECT 80.575 3.235 80.787 3.793 ;
      RECT 80.575 3.235 80.825 3.787 ;
      RECT 80.575 3.242 80.835 3.785 ;
      RECT 80.545 3.235 80.825 3.78 ;
      RECT 80.515 3.25 80.835 3.77 ;
      RECT 80.515 3.277 80.875 3.762 ;
      RECT 80.49 3.277 80.875 3.75 ;
      RECT 80.49 3.315 80.885 3.732 ;
      RECT 80.475 3.297 80.875 3.725 ;
      RECT 80.475 3.345 80.895 3.721 ;
      RECT 80.475 3.411 80.915 3.705 ;
      RECT 80.475 3.466 80.925 3.515 ;
      RECT 80.665 2.755 80.835 2.935 ;
      RECT 80.615 2.694 80.665 2.92 ;
      RECT 80.355 2.675 80.615 2.905 ;
      RECT 80.315 2.735 80.785 2.905 ;
      RECT 80.315 2.725 80.745 2.905 ;
      RECT 80.315 2.714 80.725 2.905 ;
      RECT 80.315 2.7 80.665 2.905 ;
      RECT 80.355 2.67 80.551 2.905 ;
      RECT 80.385 2.649 80.551 2.905 ;
      RECT 80.365 2.65 80.551 2.905 ;
      RECT 80.385 2.635 80.465 2.905 ;
      RECT 80.145 3.165 80.265 3.605 ;
      RECT 80.125 3.165 80.265 3.604 ;
      RECT 80.085 3.185 80.265 3.601 ;
      RECT 80.045 3.229 80.265 3.597 ;
      RECT 80.035 3.259 80.285 3.46 ;
      RECT 80.125 3.165 80.295 3.355 ;
      RECT 79.785 1.945 79.795 2.395 ;
      RECT 79.595 1.945 79.615 2.355 ;
      RECT 79.565 1.945 79.575 2.335 ;
      RECT 80.245 2.255 80.265 2.44 ;
      RECT 80.225 2.215 80.245 2.448 ;
      RECT 80.175 2.182 80.225 2.458 ;
      RECT 80.121 2.156 80.175 2.461 ;
      RECT 80.035 2.121 80.121 2.451 ;
      RECT 80.025 2.097 80.035 2.44 ;
      RECT 79.955 2.063 80.025 2.43 ;
      RECT 79.935 2.023 79.955 2.423 ;
      RECT 79.915 2.005 79.935 2.419 ;
      RECT 79.905 1.995 79.915 2.416 ;
      RECT 79.875 1.98 79.905 2.412 ;
      RECT 79.865 1.965 79.875 2.408 ;
      RECT 79.855 1.96 79.865 2.406 ;
      RECT 79.805 1.95 79.855 2.401 ;
      RECT 79.795 1.945 79.805 2.396 ;
      RECT 79.765 1.945 79.785 2.39 ;
      RECT 79.731 1.945 79.765 2.382 ;
      RECT 79.645 1.945 79.731 2.372 ;
      RECT 79.615 1.945 79.645 2.36 ;
      RECT 79.575 1.945 79.595 2.345 ;
      RECT 79.555 1.945 79.565 2.328 ;
      RECT 79.535 1.955 79.555 2.308 ;
      RECT 79.525 1.975 79.535 2.24 ;
      RECT 79.515 1.985 79.525 2 ;
      RECT 79.785 2.665 79.871 2.99 ;
      RECT 79.785 2.665 79.905 2.982 ;
      RECT 79.735 2.665 79.905 2.98 ;
      RECT 79.735 2.669 79.991 2.975 ;
      RECT 79.735 2.674 80.015 2.968 ;
      RECT 79.735 2.68 80.025 2.966 ;
      RECT 79.735 2.69 80.035 2.963 ;
      RECT 79.735 2.83 80.045 2.958 ;
      RECT 79.795 3.34 79.845 3.656 ;
      RECT 79.785 3.32 79.795 3.681 ;
      RECT 79.775 3.31 79.785 3.69 ;
      RECT 79.755 3.304 79.775 3.705 ;
      RECT 79.725 3.302 79.755 3.725 ;
      RECT 79.711 3.3 79.725 3.735 ;
      RECT 79.625 3.296 79.711 3.735 ;
      RECT 79.555 3.29 79.625 3.725 ;
      RECT 79.475 3.285 79.555 3.7 ;
      RECT 79.415 3.281 79.475 3.665 ;
      RECT 79.345 3.277 79.415 3.625 ;
      RECT 79.315 3.275 79.345 3.6 ;
      RECT 79.211 3.273 79.255 3.595 ;
      RECT 79.125 3.268 79.211 3.595 ;
      RECT 79.045 3.265 79.125 3.595 ;
      RECT 78.965 3.266 79.045 3.62 ;
      RECT 78.883 3.268 78.965 3.645 ;
      RECT 78.797 3.269 78.883 3.645 ;
      RECT 78.711 3.271 78.797 3.645 ;
      RECT 78.625 3.273 78.711 3.645 ;
      RECT 78.605 3.274 78.625 3.637 ;
      RECT 78.595 3.28 78.605 3.626 ;
      RECT 78.555 3.3 78.595 3.607 ;
      RECT 78.545 3.32 78.555 3.589 ;
      RECT 79.255 3.275 79.315 3.595 ;
      RECT 79.225 2.82 79.395 3.075 ;
      RECT 79.225 2.82 79.405 3.068 ;
      RECT 79.225 2.82 79.415 3.053 ;
      RECT 79.225 2.82 79.435 3.035 ;
      RECT 79.225 2.82 79.475 2.99 ;
      RECT 79.405 2.585 79.495 2.943 ;
      RECT 79.395 2.59 79.505 2.924 ;
      RECT 79.345 2.605 79.515 2.911 ;
      RECT 79.335 2.62 79.525 2.895 ;
      RECT 79.235 2.785 79.525 2.895 ;
      RECT 79.275 2.645 79.395 3.075 ;
      RECT 79.245 2.755 79.525 2.895 ;
      RECT 79.265 2.68 79.395 3.075 ;
      RECT 79.255 2.705 79.525 2.895 ;
      RECT 79.375 2.591 79.505 2.924 ;
      RECT 79.395 2.586 79.495 2.943 ;
      RECT 78.855 2.72 79.045 2.895 ;
      RECT 78.815 2.638 79.005 2.89 ;
      RECT 78.781 2.643 79.005 2.884 ;
      RECT 78.695 2.65 79.005 2.879 ;
      RECT 78.611 2.665 79.005 2.874 ;
      RECT 78.525 2.685 79.035 2.868 ;
      RECT 78.611 2.675 79.035 2.874 ;
      RECT 78.855 2.635 79.005 2.895 ;
      RECT 78.855 2.631 78.955 2.895 ;
      RECT 78.941 2.626 78.955 2.895 ;
      RECT 77.695 1.954 78.355 2.345 ;
      RECT 77.953 1.948 78.355 2.345 ;
      RECT 77.685 1.96 78.355 2.344 ;
      RECT 77.675 1.975 78.355 2.343 ;
      RECT 77.615 2.015 78.355 2.339 ;
      RECT 77.781 1.953 78.365 2.335 ;
      RECT 77.685 1.96 78.375 2.325 ;
      RECT 77.685 1.968 78.385 2.305 ;
      RECT 77.675 1.978 78.405 2.278 ;
      RECT 77.615 2.015 78.415 2.253 ;
      RECT 77.675 1.985 78.425 2.24 ;
      RECT 77.781 1.951 78.355 2.345 ;
      RECT 77.867 1.949 78.355 2.345 ;
      RECT 77.953 1.947 78.335 2.345 ;
      RECT 78.039 1.945 78.335 2.345 ;
      RECT 78.205 3.12 78.375 3.315 ;
      RECT 78.195 3.12 78.375 3.26 ;
      RECT 78.19 3.12 78.375 3.188 ;
      RECT 78.175 3.06 78.355 3.155 ;
      RECT 78.165 3.06 78.355 3.105 ;
      RECT 78.135 3.035 78.345 3.06 ;
      RECT 78.115 3.035 78.345 3.045 ;
      RECT 78.055 2.725 78.235 3.036 ;
      RECT 78.055 2.96 78.335 3.036 ;
      RECT 78.045 2.724 78.055 3.026 ;
      RECT 78.025 2.723 78.045 3.02 ;
      RECT 77.995 2.722 78.025 3 ;
      RECT 77.945 2.719 77.995 2.965 ;
      RECT 77.945 2.84 78.305 2.965 ;
      RECT 77.875 2.716 77.945 2.92 ;
      RECT 77.875 2.775 78.285 2.92 ;
      RECT 77.875 2.765 78.275 2.92 ;
      RECT 77.875 2.755 78.265 2.92 ;
      RECT 77.875 2.735 78.245 2.92 ;
      RECT 77.955 3.255 77.965 3.512 ;
      RECT 77.935 3.172 77.955 3.532 ;
      RECT 77.915 3.166 77.935 3.56 ;
      RECT 77.855 3.154 77.915 3.58 ;
      RECT 77.815 3.14 77.855 3.581 ;
      RECT 77.731 3.129 77.815 3.569 ;
      RECT 77.645 3.116 77.731 3.553 ;
      RECT 77.635 3.109 77.645 3.545 ;
      RECT 77.585 3.106 77.635 3.485 ;
      RECT 77.565 3.102 77.585 3.4 ;
      RECT 77.555 3.1 77.565 3.35 ;
      RECT 77.525 3.098 77.555 3.32 ;
      RECT 77.485 3.093 77.525 3.3 ;
      RECT 77.447 3.088 77.485 3.288 ;
      RECT 77.361 3.08 77.447 3.297 ;
      RECT 77.275 3.069 77.361 3.309 ;
      RECT 77.205 3.059 77.275 3.319 ;
      RECT 77.185 3.05 77.205 3.324 ;
      RECT 77.125 3.022 77.185 3.32 ;
      RECT 77.105 2.992 77.125 3.308 ;
      RECT 77.085 2.965 77.105 3.295 ;
      RECT 77.005 2.718 77.085 3.262 ;
      RECT 76.991 2.71 77.005 3.224 ;
      RECT 76.905 2.702 76.991 3.145 ;
      RECT 76.885 2.693 76.905 3.061 ;
      RECT 76.855 2.688 76.885 3.041 ;
      RECT 76.785 2.699 76.855 3.026 ;
      RECT 76.765 2.717 76.785 3 ;
      RECT 76.755 2.723 76.765 2.945 ;
      RECT 76.735 2.745 76.755 2.83 ;
      RECT 77.395 2.705 77.565 2.895 ;
      RECT 77.395 2.705 77.595 2.89 ;
      RECT 77.445 2.615 77.615 2.88 ;
      RECT 77.405 2.65 77.615 2.88 ;
      RECT 76.605 3.388 76.675 3.829 ;
      RECT 76.545 3.413 76.675 3.826 ;
      RECT 76.545 3.413 76.725 3.819 ;
      RECT 76.535 3.435 76.725 3.816 ;
      RECT 76.675 3.375 76.745 3.814 ;
      RECT 76.605 3.4 76.825 3.811 ;
      RECT 76.535 3.439 76.875 3.807 ;
      RECT 76.515 3.465 76.875 3.795 ;
      RECT 76.535 3.459 76.895 3.79 ;
      RECT 76.515 2.205 76.555 2.445 ;
      RECT 76.515 2.205 76.585 2.444 ;
      RECT 76.515 2.205 76.695 2.436 ;
      RECT 76.515 2.205 76.755 2.415 ;
      RECT 76.525 2.15 76.805 2.315 ;
      RECT 76.635 1.99 76.665 2.437 ;
      RECT 76.665 1.985 76.845 2.195 ;
      RECT 76.535 2.125 76.845 2.195 ;
      RECT 76.585 2.02 76.635 2.44 ;
      RECT 76.555 2.075 76.845 2.195 ;
      RECT 75.425 5.02 75.595 6.49 ;
      RECT 75.425 6.315 75.6 6.485 ;
      RECT 75.055 1.74 75.225 2.93 ;
      RECT 75.055 1.74 75.525 1.91 ;
      RECT 75.055 6.97 75.525 7.14 ;
      RECT 75.055 5.95 75.225 7.14 ;
      RECT 74.065 1.74 74.235 2.93 ;
      RECT 74.065 1.74 74.535 1.91 ;
      RECT 74.065 6.97 74.535 7.14 ;
      RECT 74.065 5.95 74.235 7.14 ;
      RECT 72.215 2.635 72.385 3.865 ;
      RECT 72.27 0.855 72.44 2.805 ;
      RECT 72.215 0.575 72.385 1.025 ;
      RECT 72.215 7.855 72.385 8.305 ;
      RECT 72.27 6.075 72.44 8.025 ;
      RECT 72.215 5.015 72.385 6.245 ;
      RECT 71.695 0.575 71.865 3.865 ;
      RECT 71.695 2.075 72.1 2.405 ;
      RECT 71.695 1.235 72.1 1.565 ;
      RECT 71.695 5.015 71.865 8.305 ;
      RECT 71.695 7.315 72.1 7.645 ;
      RECT 71.695 6.475 72.1 6.805 ;
      RECT 69.79 3.39 69.81 3.44 ;
      RECT 69.77 3.362 69.79 3.555 ;
      RECT 69.75 3.337 69.77 3.611 ;
      RECT 69.71 3.325 69.75 3.63 ;
      RECT 69.66 3.32 69.71 3.659 ;
      RECT 69.656 3.314 69.66 3.675 ;
      RECT 69.57 3.306 69.656 3.675 ;
      RECT 69.51 3.294 69.57 3.67 ;
      RECT 69.456 3.284 69.51 3.659 ;
      RECT 69.37 3.272 69.456 3.642 ;
      RECT 69.348 3.263 69.37 3.629 ;
      RECT 69.262 3.256 69.348 3.616 ;
      RECT 69.176 3.243 69.262 3.595 ;
      RECT 69.09 3.231 69.176 3.575 ;
      RECT 69.06 3.22 69.09 3.561 ;
      RECT 69.01 3.207 69.06 3.551 ;
      RECT 68.99 3.197 69.01 3.545 ;
      RECT 68.936 3.187 68.99 3.539 ;
      RECT 68.85 3.167 68.936 3.523 ;
      RECT 68.81 3.155 68.85 3.509 ;
      RECT 68.775 3.155 68.81 3.495 ;
      RECT 68.76 3.155 68.775 3.48 ;
      RECT 68.71 3.155 68.76 3.425 ;
      RECT 68.68 3.155 68.71 3.345 ;
      RECT 69.21 2.825 69.38 3.075 ;
      RECT 69.21 2.825 69.39 3.03 ;
      RECT 69.27 2.655 69.4 2.975 ;
      RECT 69.27 2.662 69.41 2.94 ;
      RECT 69.23 2.677 69.42 2.875 ;
      RECT 69.22 2.76 69.42 2.875 ;
      RECT 69.23 2.695 69.43 2.785 ;
      RECT 69.23 2.675 69.41 2.94 ;
      RECT 69 1.93 69.17 2.415 ;
      RECT 68.99 1.93 69.17 2.405 ;
      RECT 68.99 1.945 69.19 2.35 ;
      RECT 68.95 1.925 69.14 2.315 ;
      RECT 68.95 1.96 69.2 2.235 ;
      RECT 68.9 1.945 69.19 2.135 ;
      RECT 68.9 1.975 69.21 2.095 ;
      RECT 68.9 1.99 69.22 2.015 ;
      RECT 68.496 2.688 68.51 2.944 ;
      RECT 68.496 2.689 68.596 2.939 ;
      RECT 68.41 2.686 68.496 2.936 ;
      RECT 68.4 2.685 68.41 2.929 ;
      RECT 68.4 2.692 68.682 2.926 ;
      RECT 68.32 2.695 68.682 2.922 ;
      RECT 68.4 2.694 68.7 2.919 ;
      RECT 68.31 2.707 68.72 2.916 ;
      RECT 68.32 2.695 68.72 2.916 ;
      RECT 68.3 2.712 68.72 2.915 ;
      RECT 68.32 2.697 68.806 2.911 ;
      RECT 68.28 2.715 68.806 2.908 ;
      RECT 68.32 2.701 68.892 2.902 ;
      RECT 68.27 2.72 68.892 2.898 ;
      RECT 68.32 2.704 68.92 2.897 ;
      RECT 68.32 2.705 68.96 2.891 ;
      RECT 68.31 2.71 68.97 2.886 ;
      RECT 68.27 2.73 68.98 2.875 ;
      RECT 68.27 2.75 68.99 2.86 ;
      RECT 68.23 3.298 68.25 3.605 ;
      RECT 68.22 3.273 68.23 3.885 ;
      RECT 68.18 3.24 68.22 3.885 ;
      RECT 68.176 3.21 68.18 3.885 ;
      RECT 68.09 3.095 68.176 3.885 ;
      RECT 68.08 2.97 68.09 3.885 ;
      RECT 68.07 2.935 68.08 3.885 ;
      RECT 68.06 2.905 68.07 3.885 ;
      RECT 68.04 2.875 68.06 3.77 ;
      RECT 68.03 2.845 68.04 3.645 ;
      RECT 68.02 2.825 68.03 3.595 ;
      RECT 68 2.795 68.02 3.503 ;
      RECT 67.98 2.761 68 3.418 ;
      RECT 67.975 2.744 67.98 3.353 ;
      RECT 67.97 2.738 67.975 3.325 ;
      RECT 67.96 2.73 67.97 3.29 ;
      RECT 67.94 2.725 67.95 3.19 ;
      RECT 67.93 2.725 67.94 3.165 ;
      RECT 67.925 2.725 67.93 3.128 ;
      RECT 67.91 2.725 67.925 3.06 ;
      RECT 67.9 2.724 67.91 2.99 ;
      RECT 67.89 2.722 67.9 2.97 ;
      RECT 67.83 2.718 67.89 2.943 ;
      RECT 67.79 2.72 67.83 2.923 ;
      RECT 67.77 2.75 67.79 2.905 ;
      RECT 67.95 2.725 67.96 3.245 ;
      RECT 67.89 2.08 68.06 2.435 ;
      RECT 67.92 1.966 68.06 2.435 ;
      RECT 67.92 1.968 68.07 2.43 ;
      RECT 67.92 1.97 68.09 2.42 ;
      RECT 67.92 1.973 68.12 2.405 ;
      RECT 67.92 1.978 68.17 2.375 ;
      RECT 67.92 1.983 68.19 2.338 ;
      RECT 67.9 1.985 68.2 2.313 ;
      RECT 67.92 1.965 68.03 2.435 ;
      RECT 67.93 1.96 68.03 2.435 ;
      RECT 67.45 3.222 67.64 3.585 ;
      RECT 67.45 3.237 67.68 3.583 ;
      RECT 67.45 3.265 67.7 3.579 ;
      RECT 67.45 3.3 67.71 3.577 ;
      RECT 67.45 3.345 67.72 3.576 ;
      RECT 67.44 3.217 67.6 3.565 ;
      RECT 67.42 3.225 67.64 3.515 ;
      RECT 67.39 3.237 67.68 3.45 ;
      RECT 67.45 3.215 67.6 3.585 ;
      RECT 67.455 7.855 67.625 8.305 ;
      RECT 67.51 6.075 67.68 8.025 ;
      RECT 67.455 5.015 67.625 6.245 ;
      RECT 66.935 5.015 67.105 8.305 ;
      RECT 66.935 7.315 67.34 7.645 ;
      RECT 66.935 6.475 67.34 6.805 ;
      RECT 67.036 2.695 67.24 3.105 ;
      RECT 66.95 2.588 67.036 3.09 ;
      RECT 66.946 2.584 66.95 3.074 ;
      RECT 66.86 2.695 67.24 3.054 ;
      RECT 66.84 2.575 66.86 3.015 ;
      RECT 66.83 2.58 66.946 2.99 ;
      RECT 66.82 2.587 66.95 2.97 ;
      RECT 66.81 2.592 67.04 2.945 ;
      RECT 66.8 2.61 67.13 2.925 ;
      RECT 66.79 2.615 67.13 2.905 ;
      RECT 66.78 2.62 67.17 2.77 ;
      RECT 66.78 2.65 67.23 2.77 ;
      RECT 66.78 2.635 67.22 2.77 ;
      RECT 66.81 2.605 67.13 2.945 ;
      RECT 66.81 2.593 67.07 2.945 ;
      RECT 66.96 3.42 67.21 3.885 ;
      RECT 66.88 3.395 67.2 3.88 ;
      RECT 66.81 3.429 67.21 3.87 ;
      RECT 66.6 3.68 67.21 3.865 ;
      RECT 66.78 3.449 67.21 3.865 ;
      RECT 66.62 3.64 67.21 3.865 ;
      RECT 66.77 3.46 67.21 3.865 ;
      RECT 66.66 3.58 67.21 3.865 ;
      RECT 66.71 3.505 67.21 3.865 ;
      RECT 66.96 3.37 67.2 3.885 ;
      RECT 66.98 3.365 67.2 3.885 ;
      RECT 66.99 3.36 67.12 3.885 ;
      RECT 67.076 3.355 67.08 3.885 ;
      RECT 66.55 1.925 66.636 2.362 ;
      RECT 66.54 1.925 66.636 2.358 ;
      RECT 66.54 1.925 66.7 2.357 ;
      RECT 66.54 1.925 66.73 2.355 ;
      RECT 66.54 1.925 66.74 2.345 ;
      RECT 66.53 1.93 66.74 2.343 ;
      RECT 66.52 1.94 66.74 2.335 ;
      RECT 66.52 1.94 66.75 2.295 ;
      RECT 66.54 1.925 66.77 2.21 ;
      RECT 66.51 1.95 66.77 2.205 ;
      RECT 66.52 1.94 66.78 2.135 ;
      RECT 66.5 1.96 66.78 2.08 ;
      RECT 66.49 1.97 66.78 1.98 ;
      RECT 66.57 2.741 66.58 2.82 ;
      RECT 66.56 2.734 66.57 3.005 ;
      RECT 66.55 2.728 66.56 3.03 ;
      RECT 66.54 2.72 66.55 3.06 ;
      RECT 66.5 2.715 66.54 3.11 ;
      RECT 66.48 2.715 66.5 3.165 ;
      RECT 66.47 2.715 66.48 3.19 ;
      RECT 66.46 2.715 66.47 3.205 ;
      RECT 66.43 2.715 66.46 3.25 ;
      RECT 66.42 2.715 66.43 3.29 ;
      RECT 66.4 2.715 66.42 3.315 ;
      RECT 66.38 2.715 66.4 3.35 ;
      RECT 66.3 2.715 66.38 3.395 ;
      RECT 66.29 2.715 66.3 3.415 ;
      RECT 66.25 2.795 66.29 3.412 ;
      RECT 66.23 2.875 66.25 3.409 ;
      RECT 66.21 2.93 66.23 3.407 ;
      RECT 66.19 2.99 66.21 3.405 ;
      RECT 66.15 3.025 66.19 3.403 ;
      RECT 66.146 3.035 66.15 3.401 ;
      RECT 66.06 3.05 66.146 3.397 ;
      RECT 66.04 3.07 66.06 3.393 ;
      RECT 65.97 3.075 66.04 3.389 ;
      RECT 65.95 3.076 65.97 3.386 ;
      RECT 65.946 3.078 65.95 3.385 ;
      RECT 65.86 3.087 65.946 3.38 ;
      RECT 65.85 3.096 65.86 3.375 ;
      RECT 65.81 3.102 65.85 3.37 ;
      RECT 65.76 3.113 65.81 3.355 ;
      RECT 65.74 3.122 65.76 3.34 ;
      RECT 65.66 3.135 65.74 3.325 ;
      RECT 65.83 2.685 66 2.895 ;
      RECT 65.946 2.677 66 2.895 ;
      RECT 65.746 2.685 66 2.885 ;
      RECT 65.66 2.685 66 2.865 ;
      RECT 65.66 2.69 66.01 2.81 ;
      RECT 65.66 2.7 66.02 2.72 ;
      RECT 65.86 2.682 66 2.895 ;
      RECT 65.61 3.623 65.86 3.955 ;
      RECT 65.58 3.635 65.86 3.937 ;
      RECT 65.56 3.67 65.86 3.907 ;
      RECT 65.61 3.62 65.782 3.955 ;
      RECT 65.61 3.616 65.696 3.955 ;
      RECT 65.54 1.965 65.72 2.385 ;
      RECT 65.54 1.965 65.74 2.375 ;
      RECT 65.54 1.965 65.76 2.35 ;
      RECT 65.54 1.965 65.77 2.335 ;
      RECT 65.54 1.965 65.78 2.33 ;
      RECT 65.54 2.005 65.8 2.315 ;
      RECT 65.54 2.075 65.82 2.295 ;
      RECT 65.52 2.075 65.82 2.29 ;
      RECT 65.52 2.135 65.83 2.265 ;
      RECT 65.52 2.175 65.84 2.215 ;
      RECT 65.5 1.965 65.78 2.195 ;
      RECT 65.49 1.975 65.78 2.118 ;
      RECT 65.48 2.015 65.8 2.063 ;
      RECT 65.08 3.375 65.25 3.895 ;
      RECT 65.07 3.375 65.25 3.855 ;
      RECT 65.06 3.395 65.25 3.83 ;
      RECT 65.07 3.375 65.26 3.825 ;
      RECT 65.05 3.435 65.26 3.795 ;
      RECT 65.04 3.47 65.26 3.775 ;
      RECT 65.03 3.52 65.26 3.735 ;
      RECT 65.07 3.386 65.27 3.725 ;
      RECT 65.02 3.6 65.27 3.675 ;
      RECT 65.06 3.409 65.28 3.605 ;
      RECT 65.06 3.433 65.29 3.5 ;
      RECT 65 2.68 65.02 2.955 ;
      RECT 64.96 2.665 65 3 ;
      RECT 64.94 2.65 64.96 3.065 ;
      RECT 64.92 2.649 64.94 3.14 ;
      RECT 64.9 2.657 64.92 3.245 ;
      RECT 64.896 2.662 64.9 3.297 ;
      RECT 64.81 2.681 64.896 3.337 ;
      RECT 64.8 2.702 64.81 3.376 ;
      RECT 64.79 2.71 64.8 3.377 ;
      RECT 64.77 2.845 64.79 3.379 ;
      RECT 64.76 2.995 64.77 3.381 ;
      RECT 64.72 3.08 64.76 3.386 ;
      RECT 64.638 3.102 64.72 3.396 ;
      RECT 64.552 3.117 64.638 3.409 ;
      RECT 64.466 3.132 64.552 3.422 ;
      RECT 64.38 3.147 64.466 3.436 ;
      RECT 64.3 3.161 64.38 3.449 ;
      RECT 64.286 3.169 64.3 3.457 ;
      RECT 64.2 3.177 64.286 3.471 ;
      RECT 64.19 3.185 64.2 3.484 ;
      RECT 64.166 3.185 64.19 3.492 ;
      RECT 64.08 3.187 64.166 3.522 ;
      RECT 64 3.189 64.08 3.565 ;
      RECT 63.93 3.192 64 3.6 ;
      RECT 63.91 3.194 63.93 3.616 ;
      RECT 63.88 3.2 63.91 3.618 ;
      RECT 63.83 3.215 63.88 3.621 ;
      RECT 63.81 3.23 63.83 3.624 ;
      RECT 63.78 3.235 63.81 3.627 ;
      RECT 63.72 3.25 63.78 3.631 ;
      RECT 63.71 3.266 63.72 3.635 ;
      RECT 63.66 3.276 63.71 3.624 ;
      RECT 63.63 3.295 63.66 3.607 ;
      RECT 63.61 3.315 63.63 3.597 ;
      RECT 63.59 3.34 63.61 3.589 ;
      RECT 64.6 1.932 64.77 2.425 ;
      RECT 64.59 1.932 64.77 2.41 ;
      RECT 64.59 1.947 64.8 2.4 ;
      RECT 64.58 1.947 64.8 2.375 ;
      RECT 64.57 1.947 64.8 2.34 ;
      RECT 64.57 1.955 64.81 2.295 ;
      RECT 64.55 1.925 64.74 2.275 ;
      RECT 64.54 1.932 64.77 2.235 ;
      RECT 64.53 1.947 64.8 2.215 ;
      RECT 64.52 1.96 64.81 2.175 ;
      RECT 64.51 1.975 64.81 2.128 ;
      RECT 64.51 1.975 64.82 2.12 ;
      RECT 64.5 1.99 64.82 2.093 ;
      RECT 64.51 1.985 64.83 2.035 ;
      RECT 64.31 2.612 64.58 2.905 ;
      RECT 64.31 2.614 64.59 2.9 ;
      RECT 64.3 2.64 64.59 2.895 ;
      RECT 64.31 2.63 64.6 2.89 ;
      RECT 64.31 2.608 64.546 2.905 ;
      RECT 64.31 2.605 64.46 2.905 ;
      RECT 64.37 2.6 64.456 2.905 ;
      RECT 63.86 2.648 63.93 2.945 ;
      RECT 63.86 2.648 63.94 2.944 ;
      RECT 63.94 2.635 63.95 2.941 ;
      RECT 63.84 2.662 63.95 2.935 ;
      RECT 63.93 2.64 64.02 2.931 ;
      RECT 63.86 2.655 64.04 2.92 ;
      RECT 63.84 2.72 64.05 2.916 ;
      RECT 63.82 2.668 64.04 2.915 ;
      RECT 63.81 2.673 64.04 2.905 ;
      RECT 63.8 2.795 64.06 2.9 ;
      RECT 63.8 2.875 64.07 2.89 ;
      RECT 63.77 2.681 64.04 2.884 ;
      RECT 63.76 2.695 64.04 2.869 ;
      RECT 63.8 2.676 64.04 2.9 ;
      RECT 63.93 2.636 63.95 2.941 ;
      RECT 63.75 2.072 63.77 2.305 ;
      RECT 63.74 2.053 63.75 2.31 ;
      RECT 63.73 2.041 63.74 2.317 ;
      RECT 63.69 2.027 63.73 2.327 ;
      RECT 63.68 2.017 63.69 2.336 ;
      RECT 63.63 2.002 63.68 2.341 ;
      RECT 63.62 1.987 63.63 2.347 ;
      RECT 63.6 1.978 63.62 2.352 ;
      RECT 63.59 1.968 63.6 2.358 ;
      RECT 63.58 1.965 63.59 2.363 ;
      RECT 63.56 1.965 63.58 2.364 ;
      RECT 63.53 1.96 63.56 2.362 ;
      RECT 63.506 1.953 63.53 2.361 ;
      RECT 63.42 1.943 63.506 2.358 ;
      RECT 63.41 1.935 63.42 2.355 ;
      RECT 63.388 1.935 63.41 2.354 ;
      RECT 63.302 1.935 63.388 2.352 ;
      RECT 63.216 1.935 63.302 2.35 ;
      RECT 63.13 1.935 63.216 2.347 ;
      RECT 63.12 1.935 63.13 2.34 ;
      RECT 63.09 1.935 63.12 2.3 ;
      RECT 63.08 1.945 63.09 2.255 ;
      RECT 63.07 1.99 63.08 2.24 ;
      RECT 63.04 2.085 63.07 2.195 ;
      RECT 63.23 2.822 63.4 3.335 ;
      RECT 63.22 2.853 63.4 3.315 ;
      RECT 63.22 2.853 63.42 3.285 ;
      RECT 63.21 2.861 63.42 3.26 ;
      RECT 63.21 2.861 63.43 3.25 ;
      RECT 63.21 2.861 63.44 3.23 ;
      RECT 63.21 2.861 63.49 3.185 ;
      RECT 63.21 2.861 63.5 3.16 ;
      RECT 63.21 2.861 63.51 3.125 ;
      RECT 63.21 2.861 63.52 3.09 ;
      RECT 63.21 2.861 63.53 3.04 ;
      RECT 63.21 2.861 63.55 2.965 ;
      RECT 63.38 2.725 63.56 2.905 ;
      RECT 63.3 2.78 63.56 2.905 ;
      RECT 63.34 2.745 63.4 3.335 ;
      RECT 63.33 2.765 63.56 2.905 ;
      RECT 62.69 3.235 62.776 3.801 ;
      RECT 62.65 3.235 62.776 3.795 ;
      RECT 62.65 3.235 62.862 3.793 ;
      RECT 62.65 3.235 62.9 3.787 ;
      RECT 62.65 3.242 62.91 3.785 ;
      RECT 62.62 3.235 62.9 3.78 ;
      RECT 62.59 3.25 62.91 3.77 ;
      RECT 62.59 3.277 62.95 3.762 ;
      RECT 62.565 3.277 62.95 3.75 ;
      RECT 62.565 3.315 62.96 3.732 ;
      RECT 62.55 3.297 62.95 3.725 ;
      RECT 62.55 3.345 62.97 3.721 ;
      RECT 62.55 3.411 62.99 3.705 ;
      RECT 62.55 3.466 63 3.515 ;
      RECT 62.74 2.755 62.91 2.935 ;
      RECT 62.69 2.694 62.74 2.92 ;
      RECT 62.43 2.675 62.69 2.905 ;
      RECT 62.39 2.735 62.86 2.905 ;
      RECT 62.39 2.725 62.82 2.905 ;
      RECT 62.39 2.714 62.8 2.905 ;
      RECT 62.39 2.7 62.74 2.905 ;
      RECT 62.43 2.67 62.626 2.905 ;
      RECT 62.46 2.649 62.626 2.905 ;
      RECT 62.44 2.65 62.626 2.905 ;
      RECT 62.46 2.635 62.54 2.905 ;
      RECT 62.22 3.165 62.34 3.605 ;
      RECT 62.2 3.165 62.34 3.604 ;
      RECT 62.16 3.185 62.34 3.601 ;
      RECT 62.12 3.229 62.34 3.597 ;
      RECT 62.11 3.259 62.36 3.46 ;
      RECT 62.2 3.165 62.37 3.355 ;
      RECT 61.86 1.945 61.87 2.395 ;
      RECT 61.67 1.945 61.69 2.355 ;
      RECT 61.64 1.945 61.65 2.335 ;
      RECT 62.32 2.255 62.34 2.44 ;
      RECT 62.3 2.215 62.32 2.448 ;
      RECT 62.25 2.182 62.3 2.458 ;
      RECT 62.196 2.156 62.25 2.461 ;
      RECT 62.11 2.121 62.196 2.451 ;
      RECT 62.1 2.097 62.11 2.44 ;
      RECT 62.03 2.063 62.1 2.43 ;
      RECT 62.01 2.023 62.03 2.423 ;
      RECT 61.99 2.005 62.01 2.419 ;
      RECT 61.98 1.995 61.99 2.416 ;
      RECT 61.95 1.98 61.98 2.412 ;
      RECT 61.94 1.965 61.95 2.408 ;
      RECT 61.93 1.96 61.94 2.406 ;
      RECT 61.88 1.95 61.93 2.401 ;
      RECT 61.87 1.945 61.88 2.396 ;
      RECT 61.84 1.945 61.86 2.39 ;
      RECT 61.806 1.945 61.84 2.382 ;
      RECT 61.72 1.945 61.806 2.372 ;
      RECT 61.69 1.945 61.72 2.36 ;
      RECT 61.65 1.945 61.67 2.345 ;
      RECT 61.63 1.945 61.64 2.328 ;
      RECT 61.61 1.955 61.63 2.308 ;
      RECT 61.6 1.975 61.61 2.24 ;
      RECT 61.59 1.985 61.6 2 ;
      RECT 61.86 2.665 61.946 2.99 ;
      RECT 61.86 2.665 61.98 2.982 ;
      RECT 61.81 2.665 61.98 2.98 ;
      RECT 61.81 2.669 62.066 2.975 ;
      RECT 61.81 2.674 62.09 2.968 ;
      RECT 61.81 2.68 62.1 2.966 ;
      RECT 61.81 2.69 62.11 2.963 ;
      RECT 61.81 2.83 62.12 2.958 ;
      RECT 61.87 3.34 61.92 3.656 ;
      RECT 61.86 3.32 61.87 3.681 ;
      RECT 61.85 3.31 61.86 3.69 ;
      RECT 61.83 3.304 61.85 3.705 ;
      RECT 61.8 3.302 61.83 3.725 ;
      RECT 61.786 3.3 61.8 3.735 ;
      RECT 61.7 3.296 61.786 3.735 ;
      RECT 61.63 3.29 61.7 3.725 ;
      RECT 61.55 3.285 61.63 3.7 ;
      RECT 61.49 3.281 61.55 3.665 ;
      RECT 61.42 3.277 61.49 3.625 ;
      RECT 61.39 3.275 61.42 3.6 ;
      RECT 61.286 3.273 61.33 3.595 ;
      RECT 61.2 3.268 61.286 3.595 ;
      RECT 61.12 3.265 61.2 3.595 ;
      RECT 61.04 3.266 61.12 3.62 ;
      RECT 60.958 3.268 61.04 3.645 ;
      RECT 60.872 3.269 60.958 3.645 ;
      RECT 60.786 3.271 60.872 3.645 ;
      RECT 60.7 3.273 60.786 3.645 ;
      RECT 60.68 3.274 60.7 3.637 ;
      RECT 60.67 3.28 60.68 3.626 ;
      RECT 60.63 3.3 60.67 3.607 ;
      RECT 60.62 3.32 60.63 3.589 ;
      RECT 61.33 3.275 61.39 3.595 ;
      RECT 61.3 2.82 61.47 3.075 ;
      RECT 61.3 2.82 61.48 3.068 ;
      RECT 61.3 2.82 61.49 3.053 ;
      RECT 61.3 2.82 61.51 3.035 ;
      RECT 61.3 2.82 61.55 2.99 ;
      RECT 61.48 2.585 61.57 2.943 ;
      RECT 61.47 2.59 61.58 2.924 ;
      RECT 61.42 2.605 61.59 2.911 ;
      RECT 61.41 2.62 61.6 2.895 ;
      RECT 61.31 2.785 61.6 2.895 ;
      RECT 61.35 2.645 61.47 3.075 ;
      RECT 61.32 2.755 61.6 2.895 ;
      RECT 61.34 2.68 61.47 3.075 ;
      RECT 61.33 2.705 61.6 2.895 ;
      RECT 61.45 2.591 61.58 2.924 ;
      RECT 61.47 2.586 61.57 2.943 ;
      RECT 60.93 2.72 61.12 2.895 ;
      RECT 60.89 2.638 61.08 2.89 ;
      RECT 60.856 2.643 61.08 2.884 ;
      RECT 60.77 2.65 61.08 2.879 ;
      RECT 60.686 2.665 61.08 2.874 ;
      RECT 60.6 2.685 61.11 2.868 ;
      RECT 60.686 2.675 61.11 2.874 ;
      RECT 60.93 2.635 61.08 2.895 ;
      RECT 60.93 2.631 61.03 2.895 ;
      RECT 61.016 2.626 61.03 2.895 ;
      RECT 59.77 1.954 60.43 2.345 ;
      RECT 60.028 1.948 60.43 2.345 ;
      RECT 59.76 1.96 60.43 2.344 ;
      RECT 59.75 1.975 60.43 2.343 ;
      RECT 59.69 2.015 60.43 2.339 ;
      RECT 59.856 1.953 60.44 2.335 ;
      RECT 59.76 1.96 60.45 2.325 ;
      RECT 59.76 1.968 60.46 2.305 ;
      RECT 59.75 1.978 60.48 2.278 ;
      RECT 59.69 2.015 60.49 2.253 ;
      RECT 59.75 1.985 60.5 2.24 ;
      RECT 59.856 1.951 60.43 2.345 ;
      RECT 59.942 1.949 60.43 2.345 ;
      RECT 60.028 1.947 60.41 2.345 ;
      RECT 60.114 1.945 60.41 2.345 ;
      RECT 60.28 3.12 60.45 3.315 ;
      RECT 60.27 3.12 60.45 3.26 ;
      RECT 60.265 3.12 60.45 3.188 ;
      RECT 60.25 3.06 60.43 3.155 ;
      RECT 60.24 3.06 60.43 3.105 ;
      RECT 60.21 3.035 60.42 3.06 ;
      RECT 60.19 3.035 60.42 3.045 ;
      RECT 60.13 2.725 60.31 3.036 ;
      RECT 60.13 2.96 60.41 3.036 ;
      RECT 60.12 2.724 60.13 3.026 ;
      RECT 60.1 2.723 60.12 3.02 ;
      RECT 60.07 2.722 60.1 3 ;
      RECT 60.02 2.719 60.07 2.965 ;
      RECT 60.02 2.84 60.38 2.965 ;
      RECT 59.95 2.716 60.02 2.92 ;
      RECT 59.95 2.775 60.36 2.92 ;
      RECT 59.95 2.765 60.35 2.92 ;
      RECT 59.95 2.755 60.34 2.92 ;
      RECT 59.95 2.735 60.32 2.92 ;
      RECT 60.03 3.255 60.04 3.512 ;
      RECT 60.01 3.172 60.03 3.532 ;
      RECT 59.99 3.166 60.01 3.56 ;
      RECT 59.93 3.154 59.99 3.58 ;
      RECT 59.89 3.14 59.93 3.581 ;
      RECT 59.806 3.129 59.89 3.569 ;
      RECT 59.72 3.116 59.806 3.553 ;
      RECT 59.71 3.109 59.72 3.545 ;
      RECT 59.66 3.106 59.71 3.485 ;
      RECT 59.64 3.102 59.66 3.4 ;
      RECT 59.63 3.1 59.64 3.35 ;
      RECT 59.6 3.098 59.63 3.32 ;
      RECT 59.56 3.093 59.6 3.3 ;
      RECT 59.522 3.088 59.56 3.288 ;
      RECT 59.436 3.08 59.522 3.297 ;
      RECT 59.35 3.069 59.436 3.309 ;
      RECT 59.28 3.059 59.35 3.319 ;
      RECT 59.26 3.05 59.28 3.324 ;
      RECT 59.2 3.022 59.26 3.32 ;
      RECT 59.18 2.992 59.2 3.308 ;
      RECT 59.16 2.965 59.18 3.295 ;
      RECT 59.08 2.718 59.16 3.262 ;
      RECT 59.066 2.71 59.08 3.224 ;
      RECT 58.98 2.702 59.066 3.145 ;
      RECT 58.96 2.693 58.98 3.061 ;
      RECT 58.93 2.688 58.96 3.041 ;
      RECT 58.86 2.699 58.93 3.026 ;
      RECT 58.84 2.717 58.86 3 ;
      RECT 58.83 2.723 58.84 2.945 ;
      RECT 58.81 2.745 58.83 2.83 ;
      RECT 59.47 2.705 59.64 2.895 ;
      RECT 59.47 2.705 59.67 2.89 ;
      RECT 59.52 2.615 59.69 2.88 ;
      RECT 59.48 2.65 59.69 2.88 ;
      RECT 58.68 3.388 58.75 3.829 ;
      RECT 58.62 3.413 58.75 3.826 ;
      RECT 58.62 3.413 58.8 3.819 ;
      RECT 58.61 3.435 58.8 3.816 ;
      RECT 58.75 3.375 58.82 3.814 ;
      RECT 58.68 3.4 58.9 3.811 ;
      RECT 58.61 3.439 58.95 3.807 ;
      RECT 58.59 3.465 58.95 3.795 ;
      RECT 58.61 3.459 58.97 3.79 ;
      RECT 58.59 2.205 58.63 2.445 ;
      RECT 58.59 2.205 58.66 2.444 ;
      RECT 58.59 2.205 58.77 2.436 ;
      RECT 58.59 2.205 58.83 2.415 ;
      RECT 58.6 2.15 58.88 2.315 ;
      RECT 58.71 1.99 58.74 2.437 ;
      RECT 58.74 1.985 58.92 2.195 ;
      RECT 58.61 2.125 58.92 2.195 ;
      RECT 58.66 2.02 58.71 2.44 ;
      RECT 58.63 2.075 58.92 2.195 ;
      RECT 57.5 5.02 57.67 6.49 ;
      RECT 57.5 6.315 57.675 6.485 ;
      RECT 57.13 1.74 57.3 2.93 ;
      RECT 57.13 1.74 57.6 1.91 ;
      RECT 57.13 6.97 57.6 7.14 ;
      RECT 57.13 5.95 57.3 7.14 ;
      RECT 56.14 1.74 56.31 2.93 ;
      RECT 56.14 1.74 56.61 1.91 ;
      RECT 56.14 6.97 56.61 7.14 ;
      RECT 56.14 5.95 56.31 7.14 ;
      RECT 54.29 2.635 54.46 3.865 ;
      RECT 54.345 0.855 54.515 2.805 ;
      RECT 54.29 0.575 54.46 1.025 ;
      RECT 54.29 7.855 54.46 8.305 ;
      RECT 54.345 6.075 54.515 8.025 ;
      RECT 54.29 5.015 54.46 6.245 ;
      RECT 53.77 0.575 53.94 3.865 ;
      RECT 53.77 2.075 54.175 2.405 ;
      RECT 53.77 1.235 54.175 1.565 ;
      RECT 53.77 5.015 53.94 8.305 ;
      RECT 53.77 7.315 54.175 7.645 ;
      RECT 53.77 6.475 54.175 6.805 ;
      RECT 51.865 3.39 51.885 3.44 ;
      RECT 51.845 3.362 51.865 3.555 ;
      RECT 51.825 3.337 51.845 3.611 ;
      RECT 51.785 3.325 51.825 3.63 ;
      RECT 51.735 3.32 51.785 3.659 ;
      RECT 51.731 3.314 51.735 3.675 ;
      RECT 51.645 3.306 51.731 3.675 ;
      RECT 51.585 3.294 51.645 3.67 ;
      RECT 51.531 3.284 51.585 3.659 ;
      RECT 51.445 3.272 51.531 3.642 ;
      RECT 51.423 3.263 51.445 3.629 ;
      RECT 51.337 3.256 51.423 3.616 ;
      RECT 51.251 3.243 51.337 3.595 ;
      RECT 51.165 3.231 51.251 3.575 ;
      RECT 51.135 3.22 51.165 3.561 ;
      RECT 51.085 3.207 51.135 3.551 ;
      RECT 51.065 3.197 51.085 3.545 ;
      RECT 51.011 3.187 51.065 3.539 ;
      RECT 50.925 3.167 51.011 3.523 ;
      RECT 50.885 3.155 50.925 3.509 ;
      RECT 50.85 3.155 50.885 3.495 ;
      RECT 50.835 3.155 50.85 3.48 ;
      RECT 50.785 3.155 50.835 3.425 ;
      RECT 50.755 3.155 50.785 3.345 ;
      RECT 51.285 2.825 51.455 3.075 ;
      RECT 51.285 2.825 51.465 3.03 ;
      RECT 51.345 2.655 51.475 2.975 ;
      RECT 51.345 2.662 51.485 2.94 ;
      RECT 51.305 2.677 51.495 2.875 ;
      RECT 51.295 2.76 51.495 2.875 ;
      RECT 51.305 2.695 51.505 2.785 ;
      RECT 51.305 2.675 51.485 2.94 ;
      RECT 51.075 1.93 51.245 2.415 ;
      RECT 51.065 1.93 51.245 2.405 ;
      RECT 51.065 1.945 51.265 2.35 ;
      RECT 51.025 1.925 51.215 2.315 ;
      RECT 51.025 1.96 51.275 2.235 ;
      RECT 50.975 1.945 51.265 2.135 ;
      RECT 50.975 1.975 51.285 2.095 ;
      RECT 50.975 1.99 51.295 2.015 ;
      RECT 50.571 2.688 50.585 2.944 ;
      RECT 50.571 2.689 50.671 2.939 ;
      RECT 50.485 2.686 50.571 2.936 ;
      RECT 50.475 2.685 50.485 2.929 ;
      RECT 50.475 2.692 50.757 2.926 ;
      RECT 50.395 2.695 50.757 2.922 ;
      RECT 50.475 2.694 50.775 2.919 ;
      RECT 50.385 2.707 50.795 2.916 ;
      RECT 50.395 2.695 50.795 2.916 ;
      RECT 50.375 2.712 50.795 2.915 ;
      RECT 50.395 2.697 50.881 2.911 ;
      RECT 50.355 2.715 50.881 2.908 ;
      RECT 50.395 2.701 50.967 2.902 ;
      RECT 50.345 2.72 50.967 2.898 ;
      RECT 50.395 2.704 50.995 2.897 ;
      RECT 50.395 2.705 51.035 2.891 ;
      RECT 50.385 2.71 51.045 2.886 ;
      RECT 50.345 2.73 51.055 2.875 ;
      RECT 50.345 2.75 51.065 2.86 ;
      RECT 50.305 3.298 50.325 3.605 ;
      RECT 50.295 3.273 50.305 3.885 ;
      RECT 50.255 3.24 50.295 3.885 ;
      RECT 50.251 3.21 50.255 3.885 ;
      RECT 50.165 3.095 50.251 3.885 ;
      RECT 50.155 2.97 50.165 3.885 ;
      RECT 50.145 2.935 50.155 3.885 ;
      RECT 50.135 2.905 50.145 3.885 ;
      RECT 50.115 2.875 50.135 3.77 ;
      RECT 50.105 2.845 50.115 3.645 ;
      RECT 50.095 2.825 50.105 3.595 ;
      RECT 50.075 2.795 50.095 3.503 ;
      RECT 50.055 2.761 50.075 3.418 ;
      RECT 50.05 2.744 50.055 3.353 ;
      RECT 50.045 2.738 50.05 3.325 ;
      RECT 50.035 2.73 50.045 3.29 ;
      RECT 50.015 2.725 50.025 3.19 ;
      RECT 50.005 2.725 50.015 3.165 ;
      RECT 50 2.725 50.005 3.128 ;
      RECT 49.985 2.725 50 3.06 ;
      RECT 49.975 2.724 49.985 2.99 ;
      RECT 49.965 2.722 49.975 2.97 ;
      RECT 49.905 2.718 49.965 2.943 ;
      RECT 49.865 2.72 49.905 2.923 ;
      RECT 49.845 2.75 49.865 2.905 ;
      RECT 50.025 2.725 50.035 3.245 ;
      RECT 49.965 2.08 50.135 2.435 ;
      RECT 49.995 1.966 50.135 2.435 ;
      RECT 49.995 1.968 50.145 2.43 ;
      RECT 49.995 1.97 50.165 2.42 ;
      RECT 49.995 1.973 50.195 2.405 ;
      RECT 49.995 1.978 50.245 2.375 ;
      RECT 49.995 1.983 50.265 2.338 ;
      RECT 49.975 1.985 50.275 2.313 ;
      RECT 49.995 1.965 50.105 2.435 ;
      RECT 50.005 1.96 50.105 2.435 ;
      RECT 49.525 3.222 49.715 3.585 ;
      RECT 49.525 3.237 49.755 3.583 ;
      RECT 49.525 3.265 49.775 3.579 ;
      RECT 49.525 3.3 49.785 3.577 ;
      RECT 49.525 3.345 49.795 3.576 ;
      RECT 49.515 3.217 49.675 3.565 ;
      RECT 49.495 3.225 49.715 3.515 ;
      RECT 49.465 3.237 49.755 3.45 ;
      RECT 49.525 3.215 49.675 3.585 ;
      RECT 49.53 7.855 49.7 8.305 ;
      RECT 49.585 6.075 49.755 8.025 ;
      RECT 49.53 5.015 49.7 6.245 ;
      RECT 49.01 5.015 49.18 8.305 ;
      RECT 49.01 7.315 49.415 7.645 ;
      RECT 49.01 6.475 49.415 6.805 ;
      RECT 49.111 2.695 49.315 3.105 ;
      RECT 49.025 2.588 49.111 3.09 ;
      RECT 49.021 2.584 49.025 3.074 ;
      RECT 48.935 2.695 49.315 3.054 ;
      RECT 48.915 2.575 48.935 3.015 ;
      RECT 48.905 2.58 49.021 2.99 ;
      RECT 48.895 2.587 49.025 2.97 ;
      RECT 48.885 2.592 49.115 2.945 ;
      RECT 48.875 2.61 49.205 2.925 ;
      RECT 48.865 2.615 49.205 2.905 ;
      RECT 48.855 2.62 49.245 2.77 ;
      RECT 48.855 2.65 49.305 2.77 ;
      RECT 48.855 2.635 49.295 2.77 ;
      RECT 48.885 2.605 49.205 2.945 ;
      RECT 48.885 2.593 49.145 2.945 ;
      RECT 49.035 3.42 49.285 3.885 ;
      RECT 48.955 3.395 49.275 3.88 ;
      RECT 48.885 3.429 49.285 3.87 ;
      RECT 48.675 3.68 49.285 3.865 ;
      RECT 48.855 3.449 49.285 3.865 ;
      RECT 48.695 3.64 49.285 3.865 ;
      RECT 48.845 3.46 49.285 3.865 ;
      RECT 48.735 3.58 49.285 3.865 ;
      RECT 48.785 3.505 49.285 3.865 ;
      RECT 49.035 3.37 49.275 3.885 ;
      RECT 49.055 3.365 49.275 3.885 ;
      RECT 49.065 3.36 49.195 3.885 ;
      RECT 49.151 3.355 49.155 3.885 ;
      RECT 48.625 1.925 48.711 2.362 ;
      RECT 48.615 1.925 48.711 2.358 ;
      RECT 48.615 1.925 48.775 2.357 ;
      RECT 48.615 1.925 48.805 2.355 ;
      RECT 48.615 1.925 48.815 2.345 ;
      RECT 48.605 1.93 48.815 2.343 ;
      RECT 48.595 1.94 48.815 2.335 ;
      RECT 48.595 1.94 48.825 2.295 ;
      RECT 48.615 1.925 48.845 2.21 ;
      RECT 48.585 1.95 48.845 2.205 ;
      RECT 48.595 1.94 48.855 2.135 ;
      RECT 48.575 1.96 48.855 2.08 ;
      RECT 48.565 1.97 48.855 1.98 ;
      RECT 48.645 2.741 48.655 2.82 ;
      RECT 48.635 2.734 48.645 3.005 ;
      RECT 48.625 2.728 48.635 3.03 ;
      RECT 48.615 2.72 48.625 3.06 ;
      RECT 48.575 2.715 48.615 3.11 ;
      RECT 48.555 2.715 48.575 3.165 ;
      RECT 48.545 2.715 48.555 3.19 ;
      RECT 48.535 2.715 48.545 3.205 ;
      RECT 48.505 2.715 48.535 3.25 ;
      RECT 48.495 2.715 48.505 3.29 ;
      RECT 48.475 2.715 48.495 3.315 ;
      RECT 48.455 2.715 48.475 3.35 ;
      RECT 48.375 2.715 48.455 3.395 ;
      RECT 48.365 2.715 48.375 3.415 ;
      RECT 48.325 2.795 48.365 3.412 ;
      RECT 48.305 2.875 48.325 3.409 ;
      RECT 48.285 2.93 48.305 3.407 ;
      RECT 48.265 2.99 48.285 3.405 ;
      RECT 48.225 3.025 48.265 3.403 ;
      RECT 48.221 3.035 48.225 3.401 ;
      RECT 48.135 3.05 48.221 3.397 ;
      RECT 48.115 3.07 48.135 3.393 ;
      RECT 48.045 3.075 48.115 3.389 ;
      RECT 48.025 3.076 48.045 3.386 ;
      RECT 48.021 3.078 48.025 3.385 ;
      RECT 47.935 3.087 48.021 3.38 ;
      RECT 47.925 3.096 47.935 3.375 ;
      RECT 47.885 3.102 47.925 3.37 ;
      RECT 47.835 3.113 47.885 3.355 ;
      RECT 47.815 3.122 47.835 3.34 ;
      RECT 47.735 3.135 47.815 3.325 ;
      RECT 47.905 2.685 48.075 2.895 ;
      RECT 48.021 2.677 48.075 2.895 ;
      RECT 47.821 2.685 48.075 2.885 ;
      RECT 47.735 2.685 48.075 2.865 ;
      RECT 47.735 2.69 48.085 2.81 ;
      RECT 47.735 2.7 48.095 2.72 ;
      RECT 47.935 2.682 48.075 2.895 ;
      RECT 47.685 3.623 47.935 3.955 ;
      RECT 47.655 3.635 47.935 3.937 ;
      RECT 47.635 3.67 47.935 3.907 ;
      RECT 47.685 3.62 47.857 3.955 ;
      RECT 47.685 3.616 47.771 3.955 ;
      RECT 47.615 1.965 47.795 2.385 ;
      RECT 47.615 1.965 47.815 2.375 ;
      RECT 47.615 1.965 47.835 2.35 ;
      RECT 47.615 1.965 47.845 2.335 ;
      RECT 47.615 1.965 47.855 2.33 ;
      RECT 47.615 2.005 47.875 2.315 ;
      RECT 47.615 2.075 47.895 2.295 ;
      RECT 47.595 2.075 47.895 2.29 ;
      RECT 47.595 2.135 47.905 2.265 ;
      RECT 47.595 2.175 47.915 2.215 ;
      RECT 47.575 1.965 47.855 2.195 ;
      RECT 47.565 1.975 47.855 2.118 ;
      RECT 47.555 2.015 47.875 2.063 ;
      RECT 47.155 3.375 47.325 3.895 ;
      RECT 47.145 3.375 47.325 3.855 ;
      RECT 47.135 3.395 47.325 3.83 ;
      RECT 47.145 3.375 47.335 3.825 ;
      RECT 47.125 3.435 47.335 3.795 ;
      RECT 47.115 3.47 47.335 3.775 ;
      RECT 47.105 3.52 47.335 3.735 ;
      RECT 47.145 3.386 47.345 3.725 ;
      RECT 47.095 3.6 47.345 3.675 ;
      RECT 47.135 3.409 47.355 3.605 ;
      RECT 47.135 3.433 47.365 3.5 ;
      RECT 47.075 2.68 47.095 2.955 ;
      RECT 47.035 2.665 47.075 3 ;
      RECT 47.015 2.65 47.035 3.065 ;
      RECT 46.995 2.649 47.015 3.14 ;
      RECT 46.975 2.657 46.995 3.245 ;
      RECT 46.971 2.662 46.975 3.297 ;
      RECT 46.885 2.681 46.971 3.337 ;
      RECT 46.875 2.702 46.885 3.376 ;
      RECT 46.865 2.71 46.875 3.377 ;
      RECT 46.845 2.845 46.865 3.379 ;
      RECT 46.835 2.995 46.845 3.381 ;
      RECT 46.795 3.08 46.835 3.386 ;
      RECT 46.713 3.102 46.795 3.396 ;
      RECT 46.627 3.117 46.713 3.409 ;
      RECT 46.541 3.132 46.627 3.422 ;
      RECT 46.455 3.147 46.541 3.436 ;
      RECT 46.375 3.161 46.455 3.449 ;
      RECT 46.361 3.169 46.375 3.457 ;
      RECT 46.275 3.177 46.361 3.471 ;
      RECT 46.265 3.185 46.275 3.484 ;
      RECT 46.241 3.185 46.265 3.492 ;
      RECT 46.155 3.187 46.241 3.522 ;
      RECT 46.075 3.189 46.155 3.565 ;
      RECT 46.005 3.192 46.075 3.6 ;
      RECT 45.985 3.194 46.005 3.616 ;
      RECT 45.955 3.2 45.985 3.618 ;
      RECT 45.905 3.215 45.955 3.621 ;
      RECT 45.885 3.23 45.905 3.624 ;
      RECT 45.855 3.235 45.885 3.627 ;
      RECT 45.795 3.25 45.855 3.631 ;
      RECT 45.785 3.266 45.795 3.635 ;
      RECT 45.735 3.276 45.785 3.624 ;
      RECT 45.705 3.295 45.735 3.607 ;
      RECT 45.685 3.315 45.705 3.597 ;
      RECT 45.665 3.34 45.685 3.589 ;
      RECT 46.675 1.932 46.845 2.425 ;
      RECT 46.665 1.932 46.845 2.41 ;
      RECT 46.665 1.947 46.875 2.4 ;
      RECT 46.655 1.947 46.875 2.375 ;
      RECT 46.645 1.947 46.875 2.34 ;
      RECT 46.645 1.955 46.885 2.295 ;
      RECT 46.625 1.925 46.815 2.275 ;
      RECT 46.615 1.932 46.845 2.235 ;
      RECT 46.605 1.947 46.875 2.215 ;
      RECT 46.595 1.96 46.885 2.175 ;
      RECT 46.585 1.975 46.885 2.128 ;
      RECT 46.585 1.975 46.895 2.12 ;
      RECT 46.575 1.99 46.895 2.093 ;
      RECT 46.585 1.985 46.905 2.035 ;
      RECT 46.385 2.612 46.655 2.905 ;
      RECT 46.385 2.614 46.665 2.9 ;
      RECT 46.375 2.64 46.665 2.895 ;
      RECT 46.385 2.63 46.675 2.89 ;
      RECT 46.385 2.608 46.621 2.905 ;
      RECT 46.385 2.605 46.535 2.905 ;
      RECT 46.445 2.6 46.531 2.905 ;
      RECT 45.935 2.648 46.005 2.945 ;
      RECT 45.935 2.648 46.015 2.944 ;
      RECT 46.015 2.635 46.025 2.941 ;
      RECT 45.915 2.662 46.025 2.935 ;
      RECT 46.005 2.64 46.095 2.931 ;
      RECT 45.935 2.655 46.115 2.92 ;
      RECT 45.915 2.72 46.125 2.916 ;
      RECT 45.895 2.668 46.115 2.915 ;
      RECT 45.885 2.673 46.115 2.905 ;
      RECT 45.875 2.795 46.135 2.9 ;
      RECT 45.875 2.875 46.145 2.89 ;
      RECT 45.845 2.681 46.115 2.884 ;
      RECT 45.835 2.695 46.115 2.869 ;
      RECT 45.875 2.676 46.115 2.9 ;
      RECT 46.005 2.636 46.025 2.941 ;
      RECT 45.825 2.072 45.845 2.305 ;
      RECT 45.815 2.053 45.825 2.31 ;
      RECT 45.805 2.041 45.815 2.317 ;
      RECT 45.765 2.027 45.805 2.327 ;
      RECT 45.755 2.017 45.765 2.336 ;
      RECT 45.705 2.002 45.755 2.341 ;
      RECT 45.695 1.987 45.705 2.347 ;
      RECT 45.675 1.978 45.695 2.352 ;
      RECT 45.665 1.968 45.675 2.358 ;
      RECT 45.655 1.965 45.665 2.363 ;
      RECT 45.635 1.965 45.655 2.364 ;
      RECT 45.605 1.96 45.635 2.362 ;
      RECT 45.581 1.953 45.605 2.361 ;
      RECT 45.495 1.943 45.581 2.358 ;
      RECT 45.485 1.935 45.495 2.355 ;
      RECT 45.463 1.935 45.485 2.354 ;
      RECT 45.377 1.935 45.463 2.352 ;
      RECT 45.291 1.935 45.377 2.35 ;
      RECT 45.205 1.935 45.291 2.347 ;
      RECT 45.195 1.935 45.205 2.34 ;
      RECT 45.165 1.935 45.195 2.3 ;
      RECT 45.155 1.945 45.165 2.255 ;
      RECT 45.145 1.99 45.155 2.24 ;
      RECT 45.115 2.085 45.145 2.195 ;
      RECT 45.305 2.822 45.475 3.335 ;
      RECT 45.295 2.853 45.475 3.315 ;
      RECT 45.295 2.853 45.495 3.285 ;
      RECT 45.285 2.861 45.495 3.26 ;
      RECT 45.285 2.861 45.505 3.25 ;
      RECT 45.285 2.861 45.515 3.23 ;
      RECT 45.285 2.861 45.565 3.185 ;
      RECT 45.285 2.861 45.575 3.16 ;
      RECT 45.285 2.861 45.585 3.125 ;
      RECT 45.285 2.861 45.595 3.09 ;
      RECT 45.285 2.861 45.605 3.04 ;
      RECT 45.285 2.861 45.625 2.965 ;
      RECT 45.455 2.725 45.635 2.905 ;
      RECT 45.375 2.78 45.635 2.905 ;
      RECT 45.415 2.745 45.475 3.335 ;
      RECT 45.405 2.765 45.635 2.905 ;
      RECT 44.765 3.235 44.851 3.801 ;
      RECT 44.725 3.235 44.851 3.795 ;
      RECT 44.725 3.235 44.937 3.793 ;
      RECT 44.725 3.235 44.975 3.787 ;
      RECT 44.725 3.242 44.985 3.785 ;
      RECT 44.695 3.235 44.975 3.78 ;
      RECT 44.665 3.25 44.985 3.77 ;
      RECT 44.665 3.277 45.025 3.762 ;
      RECT 44.64 3.277 45.025 3.75 ;
      RECT 44.64 3.315 45.035 3.732 ;
      RECT 44.625 3.297 45.025 3.725 ;
      RECT 44.625 3.345 45.045 3.721 ;
      RECT 44.625 3.411 45.065 3.705 ;
      RECT 44.625 3.466 45.075 3.515 ;
      RECT 44.815 2.755 44.985 2.935 ;
      RECT 44.765 2.694 44.815 2.92 ;
      RECT 44.505 2.675 44.765 2.905 ;
      RECT 44.465 2.735 44.935 2.905 ;
      RECT 44.465 2.725 44.895 2.905 ;
      RECT 44.465 2.714 44.875 2.905 ;
      RECT 44.465 2.7 44.815 2.905 ;
      RECT 44.505 2.67 44.701 2.905 ;
      RECT 44.535 2.649 44.701 2.905 ;
      RECT 44.515 2.65 44.701 2.905 ;
      RECT 44.535 2.635 44.615 2.905 ;
      RECT 44.295 3.165 44.415 3.605 ;
      RECT 44.275 3.165 44.415 3.604 ;
      RECT 44.235 3.185 44.415 3.601 ;
      RECT 44.195 3.229 44.415 3.597 ;
      RECT 44.185 3.259 44.435 3.46 ;
      RECT 44.275 3.165 44.445 3.355 ;
      RECT 43.935 1.945 43.945 2.395 ;
      RECT 43.745 1.945 43.765 2.355 ;
      RECT 43.715 1.945 43.725 2.335 ;
      RECT 44.395 2.255 44.415 2.44 ;
      RECT 44.375 2.215 44.395 2.448 ;
      RECT 44.325 2.182 44.375 2.458 ;
      RECT 44.271 2.156 44.325 2.461 ;
      RECT 44.185 2.121 44.271 2.451 ;
      RECT 44.175 2.097 44.185 2.44 ;
      RECT 44.105 2.063 44.175 2.43 ;
      RECT 44.085 2.023 44.105 2.423 ;
      RECT 44.065 2.005 44.085 2.419 ;
      RECT 44.055 1.995 44.065 2.416 ;
      RECT 44.025 1.98 44.055 2.412 ;
      RECT 44.015 1.965 44.025 2.408 ;
      RECT 44.005 1.96 44.015 2.406 ;
      RECT 43.955 1.95 44.005 2.401 ;
      RECT 43.945 1.945 43.955 2.396 ;
      RECT 43.915 1.945 43.935 2.39 ;
      RECT 43.881 1.945 43.915 2.382 ;
      RECT 43.795 1.945 43.881 2.372 ;
      RECT 43.765 1.945 43.795 2.36 ;
      RECT 43.725 1.945 43.745 2.345 ;
      RECT 43.705 1.945 43.715 2.328 ;
      RECT 43.685 1.955 43.705 2.308 ;
      RECT 43.675 1.975 43.685 2.24 ;
      RECT 43.665 1.985 43.675 2 ;
      RECT 43.935 2.665 44.021 2.99 ;
      RECT 43.935 2.665 44.055 2.982 ;
      RECT 43.885 2.665 44.055 2.98 ;
      RECT 43.885 2.669 44.141 2.975 ;
      RECT 43.885 2.674 44.165 2.968 ;
      RECT 43.885 2.68 44.175 2.966 ;
      RECT 43.885 2.69 44.185 2.963 ;
      RECT 43.885 2.83 44.195 2.958 ;
      RECT 43.945 3.34 43.995 3.656 ;
      RECT 43.935 3.32 43.945 3.681 ;
      RECT 43.925 3.31 43.935 3.69 ;
      RECT 43.905 3.304 43.925 3.705 ;
      RECT 43.875 3.302 43.905 3.725 ;
      RECT 43.861 3.3 43.875 3.735 ;
      RECT 43.775 3.296 43.861 3.735 ;
      RECT 43.705 3.29 43.775 3.725 ;
      RECT 43.625 3.285 43.705 3.7 ;
      RECT 43.565 3.281 43.625 3.665 ;
      RECT 43.495 3.277 43.565 3.625 ;
      RECT 43.465 3.275 43.495 3.6 ;
      RECT 43.361 3.273 43.405 3.595 ;
      RECT 43.275 3.268 43.361 3.595 ;
      RECT 43.195 3.265 43.275 3.595 ;
      RECT 43.115 3.266 43.195 3.62 ;
      RECT 43.033 3.268 43.115 3.645 ;
      RECT 42.947 3.269 43.033 3.645 ;
      RECT 42.861 3.271 42.947 3.645 ;
      RECT 42.775 3.273 42.861 3.645 ;
      RECT 42.755 3.274 42.775 3.637 ;
      RECT 42.745 3.28 42.755 3.626 ;
      RECT 42.705 3.3 42.745 3.607 ;
      RECT 42.695 3.32 42.705 3.589 ;
      RECT 43.405 3.275 43.465 3.595 ;
      RECT 43.375 2.82 43.545 3.075 ;
      RECT 43.375 2.82 43.555 3.068 ;
      RECT 43.375 2.82 43.565 3.053 ;
      RECT 43.375 2.82 43.585 3.035 ;
      RECT 43.375 2.82 43.625 2.99 ;
      RECT 43.555 2.585 43.645 2.943 ;
      RECT 43.545 2.59 43.655 2.924 ;
      RECT 43.495 2.605 43.665 2.911 ;
      RECT 43.485 2.62 43.675 2.895 ;
      RECT 43.385 2.785 43.675 2.895 ;
      RECT 43.425 2.645 43.545 3.075 ;
      RECT 43.395 2.755 43.675 2.895 ;
      RECT 43.415 2.68 43.545 3.075 ;
      RECT 43.405 2.705 43.675 2.895 ;
      RECT 43.525 2.591 43.655 2.924 ;
      RECT 43.545 2.586 43.645 2.943 ;
      RECT 43.005 2.72 43.195 2.895 ;
      RECT 42.965 2.638 43.155 2.89 ;
      RECT 42.931 2.643 43.155 2.884 ;
      RECT 42.845 2.65 43.155 2.879 ;
      RECT 42.761 2.665 43.155 2.874 ;
      RECT 42.675 2.685 43.185 2.868 ;
      RECT 42.761 2.675 43.185 2.874 ;
      RECT 43.005 2.635 43.155 2.895 ;
      RECT 43.005 2.631 43.105 2.895 ;
      RECT 43.091 2.626 43.105 2.895 ;
      RECT 41.845 1.954 42.505 2.345 ;
      RECT 42.103 1.948 42.505 2.345 ;
      RECT 41.835 1.96 42.505 2.344 ;
      RECT 41.825 1.975 42.505 2.343 ;
      RECT 41.765 2.015 42.505 2.339 ;
      RECT 41.931 1.953 42.515 2.335 ;
      RECT 41.835 1.96 42.525 2.325 ;
      RECT 41.835 1.968 42.535 2.305 ;
      RECT 41.825 1.978 42.555 2.278 ;
      RECT 41.765 2.015 42.565 2.253 ;
      RECT 41.825 1.985 42.575 2.24 ;
      RECT 41.931 1.951 42.505 2.345 ;
      RECT 42.017 1.949 42.505 2.345 ;
      RECT 42.103 1.947 42.485 2.345 ;
      RECT 42.189 1.945 42.485 2.345 ;
      RECT 42.355 3.12 42.525 3.315 ;
      RECT 42.345 3.12 42.525 3.26 ;
      RECT 42.34 3.12 42.525 3.188 ;
      RECT 42.325 3.06 42.505 3.155 ;
      RECT 42.315 3.06 42.505 3.105 ;
      RECT 42.285 3.035 42.495 3.06 ;
      RECT 42.265 3.035 42.495 3.045 ;
      RECT 42.205 2.725 42.385 3.036 ;
      RECT 42.205 2.96 42.485 3.036 ;
      RECT 42.195 2.724 42.205 3.026 ;
      RECT 42.175 2.723 42.195 3.02 ;
      RECT 42.145 2.722 42.175 3 ;
      RECT 42.095 2.719 42.145 2.965 ;
      RECT 42.095 2.84 42.455 2.965 ;
      RECT 42.025 2.716 42.095 2.92 ;
      RECT 42.025 2.775 42.435 2.92 ;
      RECT 42.025 2.765 42.425 2.92 ;
      RECT 42.025 2.755 42.415 2.92 ;
      RECT 42.025 2.735 42.395 2.92 ;
      RECT 42.105 3.255 42.115 3.512 ;
      RECT 42.085 3.172 42.105 3.532 ;
      RECT 42.065 3.166 42.085 3.56 ;
      RECT 42.005 3.154 42.065 3.58 ;
      RECT 41.965 3.14 42.005 3.581 ;
      RECT 41.881 3.129 41.965 3.569 ;
      RECT 41.795 3.116 41.881 3.553 ;
      RECT 41.785 3.109 41.795 3.545 ;
      RECT 41.735 3.106 41.785 3.485 ;
      RECT 41.715 3.102 41.735 3.4 ;
      RECT 41.705 3.1 41.715 3.35 ;
      RECT 41.675 3.098 41.705 3.32 ;
      RECT 41.635 3.093 41.675 3.3 ;
      RECT 41.597 3.088 41.635 3.288 ;
      RECT 41.511 3.08 41.597 3.297 ;
      RECT 41.425 3.069 41.511 3.309 ;
      RECT 41.355 3.059 41.425 3.319 ;
      RECT 41.335 3.05 41.355 3.324 ;
      RECT 41.275 3.022 41.335 3.32 ;
      RECT 41.255 2.992 41.275 3.308 ;
      RECT 41.235 2.965 41.255 3.295 ;
      RECT 41.155 2.718 41.235 3.262 ;
      RECT 41.141 2.71 41.155 3.224 ;
      RECT 41.055 2.702 41.141 3.145 ;
      RECT 41.035 2.693 41.055 3.061 ;
      RECT 41.005 2.688 41.035 3.041 ;
      RECT 40.935 2.699 41.005 3.026 ;
      RECT 40.915 2.717 40.935 3 ;
      RECT 40.905 2.723 40.915 2.945 ;
      RECT 40.885 2.745 40.905 2.83 ;
      RECT 41.545 2.705 41.715 2.895 ;
      RECT 41.545 2.705 41.745 2.89 ;
      RECT 41.595 2.615 41.765 2.88 ;
      RECT 41.555 2.65 41.765 2.88 ;
      RECT 40.755 3.388 40.825 3.829 ;
      RECT 40.695 3.413 40.825 3.826 ;
      RECT 40.695 3.413 40.875 3.819 ;
      RECT 40.685 3.435 40.875 3.816 ;
      RECT 40.825 3.375 40.895 3.814 ;
      RECT 40.755 3.4 40.975 3.811 ;
      RECT 40.685 3.439 41.025 3.807 ;
      RECT 40.665 3.465 41.025 3.795 ;
      RECT 40.685 3.459 41.045 3.79 ;
      RECT 40.665 2.205 40.705 2.445 ;
      RECT 40.665 2.205 40.735 2.444 ;
      RECT 40.665 2.205 40.845 2.436 ;
      RECT 40.665 2.205 40.905 2.415 ;
      RECT 40.675 2.15 40.955 2.315 ;
      RECT 40.785 1.99 40.815 2.437 ;
      RECT 40.815 1.985 40.995 2.195 ;
      RECT 40.685 2.125 40.995 2.195 ;
      RECT 40.735 2.02 40.785 2.44 ;
      RECT 40.705 2.075 40.995 2.195 ;
      RECT 39.575 5.02 39.745 6.49 ;
      RECT 39.575 6.315 39.75 6.485 ;
      RECT 39.205 1.74 39.375 2.93 ;
      RECT 39.205 1.74 39.675 1.91 ;
      RECT 39.205 6.97 39.675 7.14 ;
      RECT 39.205 5.95 39.375 7.14 ;
      RECT 38.215 1.74 38.385 2.93 ;
      RECT 38.215 1.74 38.685 1.91 ;
      RECT 38.215 6.97 38.685 7.14 ;
      RECT 38.215 5.95 38.385 7.14 ;
      RECT 36.365 2.635 36.535 3.865 ;
      RECT 36.42 0.855 36.59 2.805 ;
      RECT 36.365 0.575 36.535 1.025 ;
      RECT 36.365 7.855 36.535 8.305 ;
      RECT 36.42 6.075 36.59 8.025 ;
      RECT 36.365 5.015 36.535 6.245 ;
      RECT 35.845 0.575 36.015 3.865 ;
      RECT 35.845 2.075 36.25 2.405 ;
      RECT 35.845 1.235 36.25 1.565 ;
      RECT 35.845 5.015 36.015 8.305 ;
      RECT 35.845 7.315 36.25 7.645 ;
      RECT 35.845 6.475 36.25 6.805 ;
      RECT 33.94 3.39 33.96 3.44 ;
      RECT 33.92 3.362 33.94 3.555 ;
      RECT 33.9 3.337 33.92 3.611 ;
      RECT 33.86 3.325 33.9 3.63 ;
      RECT 33.81 3.32 33.86 3.659 ;
      RECT 33.806 3.314 33.81 3.675 ;
      RECT 33.72 3.306 33.806 3.675 ;
      RECT 33.66 3.294 33.72 3.67 ;
      RECT 33.606 3.284 33.66 3.659 ;
      RECT 33.52 3.272 33.606 3.642 ;
      RECT 33.498 3.263 33.52 3.629 ;
      RECT 33.412 3.256 33.498 3.616 ;
      RECT 33.326 3.243 33.412 3.595 ;
      RECT 33.24 3.231 33.326 3.575 ;
      RECT 33.21 3.22 33.24 3.561 ;
      RECT 33.16 3.207 33.21 3.551 ;
      RECT 33.14 3.197 33.16 3.545 ;
      RECT 33.086 3.187 33.14 3.539 ;
      RECT 33 3.167 33.086 3.523 ;
      RECT 32.96 3.155 33 3.509 ;
      RECT 32.925 3.155 32.96 3.495 ;
      RECT 32.91 3.155 32.925 3.48 ;
      RECT 32.86 3.155 32.91 3.425 ;
      RECT 32.83 3.155 32.86 3.345 ;
      RECT 33.36 2.825 33.53 3.075 ;
      RECT 33.36 2.825 33.54 3.03 ;
      RECT 33.42 2.655 33.55 2.975 ;
      RECT 33.42 2.662 33.56 2.94 ;
      RECT 33.38 2.677 33.57 2.875 ;
      RECT 33.37 2.76 33.57 2.875 ;
      RECT 33.38 2.695 33.58 2.785 ;
      RECT 33.38 2.675 33.56 2.94 ;
      RECT 33.15 1.93 33.32 2.415 ;
      RECT 33.14 1.93 33.32 2.405 ;
      RECT 33.14 1.945 33.34 2.35 ;
      RECT 33.1 1.925 33.29 2.315 ;
      RECT 33.1 1.96 33.35 2.235 ;
      RECT 33.05 1.945 33.34 2.135 ;
      RECT 33.05 1.975 33.36 2.095 ;
      RECT 33.05 1.99 33.37 2.015 ;
      RECT 32.646 2.688 32.66 2.944 ;
      RECT 32.646 2.689 32.746 2.939 ;
      RECT 32.56 2.686 32.646 2.936 ;
      RECT 32.55 2.685 32.56 2.929 ;
      RECT 32.55 2.692 32.832 2.926 ;
      RECT 32.47 2.695 32.832 2.922 ;
      RECT 32.55 2.694 32.85 2.919 ;
      RECT 32.46 2.707 32.87 2.916 ;
      RECT 32.47 2.695 32.87 2.916 ;
      RECT 32.45 2.712 32.87 2.915 ;
      RECT 32.47 2.697 32.956 2.911 ;
      RECT 32.43 2.715 32.956 2.908 ;
      RECT 32.47 2.701 33.042 2.902 ;
      RECT 32.42 2.72 33.042 2.898 ;
      RECT 32.47 2.704 33.07 2.897 ;
      RECT 32.47 2.705 33.11 2.891 ;
      RECT 32.46 2.71 33.12 2.886 ;
      RECT 32.42 2.73 33.13 2.875 ;
      RECT 32.42 2.75 33.14 2.86 ;
      RECT 32.38 3.298 32.4 3.605 ;
      RECT 32.37 3.273 32.38 3.885 ;
      RECT 32.33 3.24 32.37 3.885 ;
      RECT 32.326 3.21 32.33 3.885 ;
      RECT 32.24 3.095 32.326 3.885 ;
      RECT 32.23 2.97 32.24 3.885 ;
      RECT 32.22 2.935 32.23 3.885 ;
      RECT 32.21 2.905 32.22 3.885 ;
      RECT 32.19 2.875 32.21 3.77 ;
      RECT 32.18 2.845 32.19 3.645 ;
      RECT 32.17 2.825 32.18 3.595 ;
      RECT 32.15 2.795 32.17 3.503 ;
      RECT 32.13 2.761 32.15 3.418 ;
      RECT 32.125 2.744 32.13 3.353 ;
      RECT 32.12 2.738 32.125 3.325 ;
      RECT 32.11 2.73 32.12 3.29 ;
      RECT 32.09 2.725 32.1 3.19 ;
      RECT 32.08 2.725 32.09 3.165 ;
      RECT 32.075 2.725 32.08 3.128 ;
      RECT 32.06 2.725 32.075 3.06 ;
      RECT 32.05 2.724 32.06 2.99 ;
      RECT 32.04 2.722 32.05 2.97 ;
      RECT 31.98 2.718 32.04 2.943 ;
      RECT 31.94 2.72 31.98 2.923 ;
      RECT 31.92 2.75 31.94 2.905 ;
      RECT 32.1 2.725 32.11 3.245 ;
      RECT 32.04 2.08 32.21 2.435 ;
      RECT 32.07 1.966 32.21 2.435 ;
      RECT 32.07 1.968 32.22 2.43 ;
      RECT 32.07 1.97 32.24 2.42 ;
      RECT 32.07 1.973 32.27 2.405 ;
      RECT 32.07 1.978 32.32 2.375 ;
      RECT 32.07 1.983 32.34 2.338 ;
      RECT 32.05 1.985 32.35 2.313 ;
      RECT 32.07 1.965 32.18 2.435 ;
      RECT 32.08 1.96 32.18 2.435 ;
      RECT 31.6 3.222 31.79 3.585 ;
      RECT 31.6 3.237 31.83 3.583 ;
      RECT 31.6 3.265 31.85 3.579 ;
      RECT 31.6 3.3 31.86 3.577 ;
      RECT 31.6 3.345 31.87 3.576 ;
      RECT 31.59 3.217 31.75 3.565 ;
      RECT 31.57 3.225 31.79 3.515 ;
      RECT 31.54 3.237 31.83 3.45 ;
      RECT 31.6 3.215 31.75 3.585 ;
      RECT 31.605 7.855 31.775 8.305 ;
      RECT 31.66 6.075 31.83 8.025 ;
      RECT 31.605 5.015 31.775 6.245 ;
      RECT 31.085 5.015 31.255 8.305 ;
      RECT 31.085 7.315 31.49 7.645 ;
      RECT 31.085 6.475 31.49 6.805 ;
      RECT 31.186 2.695 31.39 3.105 ;
      RECT 31.1 2.588 31.186 3.09 ;
      RECT 31.096 2.584 31.1 3.074 ;
      RECT 31.01 2.695 31.39 3.054 ;
      RECT 30.99 2.575 31.01 3.015 ;
      RECT 30.98 2.58 31.096 2.99 ;
      RECT 30.97 2.587 31.1 2.97 ;
      RECT 30.96 2.592 31.19 2.945 ;
      RECT 30.95 2.61 31.28 2.925 ;
      RECT 30.94 2.615 31.28 2.905 ;
      RECT 30.93 2.62 31.32 2.77 ;
      RECT 30.93 2.65 31.38 2.77 ;
      RECT 30.93 2.635 31.37 2.77 ;
      RECT 30.96 2.605 31.28 2.945 ;
      RECT 30.96 2.593 31.22 2.945 ;
      RECT 31.11 3.42 31.36 3.885 ;
      RECT 31.03 3.395 31.35 3.88 ;
      RECT 30.96 3.429 31.36 3.87 ;
      RECT 30.75 3.68 31.36 3.865 ;
      RECT 30.93 3.449 31.36 3.865 ;
      RECT 30.77 3.64 31.36 3.865 ;
      RECT 30.92 3.46 31.36 3.865 ;
      RECT 30.81 3.58 31.36 3.865 ;
      RECT 30.86 3.505 31.36 3.865 ;
      RECT 31.11 3.37 31.35 3.885 ;
      RECT 31.13 3.365 31.35 3.885 ;
      RECT 31.14 3.36 31.27 3.885 ;
      RECT 31.226 3.355 31.23 3.885 ;
      RECT 30.7 1.925 30.786 2.362 ;
      RECT 30.69 1.925 30.786 2.358 ;
      RECT 30.69 1.925 30.85 2.357 ;
      RECT 30.69 1.925 30.88 2.355 ;
      RECT 30.69 1.925 30.89 2.345 ;
      RECT 30.68 1.93 30.89 2.343 ;
      RECT 30.67 1.94 30.89 2.335 ;
      RECT 30.67 1.94 30.9 2.295 ;
      RECT 30.69 1.925 30.92 2.21 ;
      RECT 30.66 1.95 30.92 2.205 ;
      RECT 30.67 1.94 30.93 2.135 ;
      RECT 30.65 1.96 30.93 2.08 ;
      RECT 30.64 1.97 30.93 1.98 ;
      RECT 30.72 2.741 30.73 2.82 ;
      RECT 30.71 2.734 30.72 3.005 ;
      RECT 30.7 2.728 30.71 3.03 ;
      RECT 30.69 2.72 30.7 3.06 ;
      RECT 30.65 2.715 30.69 3.11 ;
      RECT 30.63 2.715 30.65 3.165 ;
      RECT 30.62 2.715 30.63 3.19 ;
      RECT 30.61 2.715 30.62 3.205 ;
      RECT 30.58 2.715 30.61 3.25 ;
      RECT 30.57 2.715 30.58 3.29 ;
      RECT 30.55 2.715 30.57 3.315 ;
      RECT 30.53 2.715 30.55 3.35 ;
      RECT 30.45 2.715 30.53 3.395 ;
      RECT 30.44 2.715 30.45 3.415 ;
      RECT 30.4 2.795 30.44 3.412 ;
      RECT 30.38 2.875 30.4 3.409 ;
      RECT 30.36 2.93 30.38 3.407 ;
      RECT 30.34 2.99 30.36 3.405 ;
      RECT 30.3 3.025 30.34 3.403 ;
      RECT 30.296 3.035 30.3 3.401 ;
      RECT 30.21 3.05 30.296 3.397 ;
      RECT 30.19 3.07 30.21 3.393 ;
      RECT 30.12 3.075 30.19 3.389 ;
      RECT 30.1 3.076 30.12 3.386 ;
      RECT 30.096 3.078 30.1 3.385 ;
      RECT 30.01 3.087 30.096 3.38 ;
      RECT 30 3.096 30.01 3.375 ;
      RECT 29.96 3.102 30 3.37 ;
      RECT 29.91 3.113 29.96 3.355 ;
      RECT 29.89 3.122 29.91 3.34 ;
      RECT 29.81 3.135 29.89 3.325 ;
      RECT 29.98 2.685 30.15 2.895 ;
      RECT 30.096 2.677 30.15 2.895 ;
      RECT 29.896 2.685 30.15 2.885 ;
      RECT 29.81 2.685 30.15 2.865 ;
      RECT 29.81 2.69 30.16 2.81 ;
      RECT 29.81 2.7 30.17 2.72 ;
      RECT 30.01 2.682 30.15 2.895 ;
      RECT 29.76 3.623 30.01 3.955 ;
      RECT 29.73 3.635 30.01 3.937 ;
      RECT 29.71 3.67 30.01 3.907 ;
      RECT 29.76 3.62 29.932 3.955 ;
      RECT 29.76 3.616 29.846 3.955 ;
      RECT 29.69 1.965 29.87 2.385 ;
      RECT 29.69 1.965 29.89 2.375 ;
      RECT 29.69 1.965 29.91 2.35 ;
      RECT 29.69 1.965 29.92 2.335 ;
      RECT 29.69 1.965 29.93 2.33 ;
      RECT 29.69 2.005 29.95 2.315 ;
      RECT 29.69 2.075 29.97 2.295 ;
      RECT 29.67 2.075 29.97 2.29 ;
      RECT 29.67 2.135 29.98 2.265 ;
      RECT 29.67 2.175 29.99 2.215 ;
      RECT 29.65 1.965 29.93 2.195 ;
      RECT 29.64 1.975 29.93 2.118 ;
      RECT 29.63 2.015 29.95 2.063 ;
      RECT 29.23 3.375 29.4 3.895 ;
      RECT 29.22 3.375 29.4 3.855 ;
      RECT 29.21 3.395 29.4 3.83 ;
      RECT 29.22 3.375 29.41 3.825 ;
      RECT 29.2 3.435 29.41 3.795 ;
      RECT 29.19 3.47 29.41 3.775 ;
      RECT 29.18 3.52 29.41 3.735 ;
      RECT 29.22 3.386 29.42 3.725 ;
      RECT 29.17 3.6 29.42 3.675 ;
      RECT 29.21 3.409 29.43 3.605 ;
      RECT 29.21 3.433 29.44 3.5 ;
      RECT 29.15 2.68 29.17 2.955 ;
      RECT 29.11 2.665 29.15 3 ;
      RECT 29.09 2.65 29.11 3.065 ;
      RECT 29.07 2.649 29.09 3.14 ;
      RECT 29.05 2.657 29.07 3.245 ;
      RECT 29.046 2.662 29.05 3.297 ;
      RECT 28.96 2.681 29.046 3.337 ;
      RECT 28.95 2.702 28.96 3.376 ;
      RECT 28.94 2.71 28.95 3.377 ;
      RECT 28.92 2.845 28.94 3.379 ;
      RECT 28.91 2.995 28.92 3.381 ;
      RECT 28.87 3.08 28.91 3.386 ;
      RECT 28.788 3.102 28.87 3.396 ;
      RECT 28.702 3.117 28.788 3.409 ;
      RECT 28.616 3.132 28.702 3.422 ;
      RECT 28.53 3.147 28.616 3.436 ;
      RECT 28.45 3.161 28.53 3.449 ;
      RECT 28.436 3.169 28.45 3.457 ;
      RECT 28.35 3.177 28.436 3.471 ;
      RECT 28.34 3.185 28.35 3.484 ;
      RECT 28.316 3.185 28.34 3.492 ;
      RECT 28.23 3.187 28.316 3.522 ;
      RECT 28.15 3.189 28.23 3.565 ;
      RECT 28.08 3.192 28.15 3.6 ;
      RECT 28.06 3.194 28.08 3.616 ;
      RECT 28.03 3.2 28.06 3.618 ;
      RECT 27.98 3.215 28.03 3.621 ;
      RECT 27.96 3.23 27.98 3.624 ;
      RECT 27.93 3.235 27.96 3.627 ;
      RECT 27.87 3.25 27.93 3.631 ;
      RECT 27.86 3.266 27.87 3.635 ;
      RECT 27.81 3.276 27.86 3.624 ;
      RECT 27.78 3.295 27.81 3.607 ;
      RECT 27.76 3.315 27.78 3.597 ;
      RECT 27.74 3.34 27.76 3.589 ;
      RECT 28.75 1.932 28.92 2.425 ;
      RECT 28.74 1.932 28.92 2.41 ;
      RECT 28.74 1.947 28.95 2.4 ;
      RECT 28.73 1.947 28.95 2.375 ;
      RECT 28.72 1.947 28.95 2.34 ;
      RECT 28.72 1.955 28.96 2.295 ;
      RECT 28.7 1.925 28.89 2.275 ;
      RECT 28.69 1.932 28.92 2.235 ;
      RECT 28.68 1.947 28.95 2.215 ;
      RECT 28.67 1.96 28.96 2.175 ;
      RECT 28.66 1.975 28.96 2.128 ;
      RECT 28.66 1.975 28.97 2.12 ;
      RECT 28.65 1.99 28.97 2.093 ;
      RECT 28.66 1.985 28.98 2.035 ;
      RECT 28.46 2.612 28.73 2.905 ;
      RECT 28.46 2.614 28.74 2.9 ;
      RECT 28.45 2.64 28.74 2.895 ;
      RECT 28.46 2.63 28.75 2.89 ;
      RECT 28.46 2.608 28.696 2.905 ;
      RECT 28.46 2.605 28.61 2.905 ;
      RECT 28.52 2.6 28.606 2.905 ;
      RECT 28.01 2.648 28.08 2.945 ;
      RECT 28.01 2.648 28.09 2.944 ;
      RECT 28.09 2.635 28.1 2.941 ;
      RECT 27.99 2.662 28.1 2.935 ;
      RECT 28.08 2.64 28.17 2.931 ;
      RECT 28.01 2.655 28.19 2.92 ;
      RECT 27.99 2.72 28.2 2.916 ;
      RECT 27.97 2.668 28.19 2.915 ;
      RECT 27.96 2.673 28.19 2.905 ;
      RECT 27.95 2.795 28.21 2.9 ;
      RECT 27.95 2.875 28.22 2.89 ;
      RECT 27.92 2.681 28.19 2.884 ;
      RECT 27.91 2.695 28.19 2.869 ;
      RECT 27.95 2.676 28.19 2.9 ;
      RECT 28.08 2.636 28.1 2.941 ;
      RECT 27.9 2.072 27.92 2.305 ;
      RECT 27.89 2.053 27.9 2.31 ;
      RECT 27.88 2.041 27.89 2.317 ;
      RECT 27.84 2.027 27.88 2.327 ;
      RECT 27.83 2.017 27.84 2.336 ;
      RECT 27.78 2.002 27.83 2.341 ;
      RECT 27.77 1.987 27.78 2.347 ;
      RECT 27.75 1.978 27.77 2.352 ;
      RECT 27.74 1.968 27.75 2.358 ;
      RECT 27.73 1.965 27.74 2.363 ;
      RECT 27.71 1.965 27.73 2.364 ;
      RECT 27.68 1.96 27.71 2.362 ;
      RECT 27.656 1.953 27.68 2.361 ;
      RECT 27.57 1.943 27.656 2.358 ;
      RECT 27.56 1.935 27.57 2.355 ;
      RECT 27.538 1.935 27.56 2.354 ;
      RECT 27.452 1.935 27.538 2.352 ;
      RECT 27.366 1.935 27.452 2.35 ;
      RECT 27.28 1.935 27.366 2.347 ;
      RECT 27.27 1.935 27.28 2.34 ;
      RECT 27.24 1.935 27.27 2.3 ;
      RECT 27.23 1.945 27.24 2.255 ;
      RECT 27.22 1.99 27.23 2.24 ;
      RECT 27.19 2.085 27.22 2.195 ;
      RECT 27.38 2.822 27.55 3.335 ;
      RECT 27.37 2.853 27.55 3.315 ;
      RECT 27.37 2.853 27.57 3.285 ;
      RECT 27.36 2.861 27.57 3.26 ;
      RECT 27.36 2.861 27.58 3.25 ;
      RECT 27.36 2.861 27.59 3.23 ;
      RECT 27.36 2.861 27.64 3.185 ;
      RECT 27.36 2.861 27.65 3.16 ;
      RECT 27.36 2.861 27.66 3.125 ;
      RECT 27.36 2.861 27.67 3.09 ;
      RECT 27.36 2.861 27.68 3.04 ;
      RECT 27.36 2.861 27.7 2.965 ;
      RECT 27.53 2.725 27.71 2.905 ;
      RECT 27.45 2.78 27.71 2.905 ;
      RECT 27.49 2.745 27.55 3.335 ;
      RECT 27.48 2.765 27.71 2.905 ;
      RECT 26.84 3.235 26.926 3.801 ;
      RECT 26.8 3.235 26.926 3.795 ;
      RECT 26.8 3.235 27.012 3.793 ;
      RECT 26.8 3.235 27.05 3.787 ;
      RECT 26.8 3.242 27.06 3.785 ;
      RECT 26.77 3.235 27.05 3.78 ;
      RECT 26.74 3.25 27.06 3.77 ;
      RECT 26.74 3.277 27.1 3.762 ;
      RECT 26.715 3.277 27.1 3.75 ;
      RECT 26.715 3.315 27.11 3.732 ;
      RECT 26.7 3.297 27.1 3.725 ;
      RECT 26.7 3.345 27.12 3.721 ;
      RECT 26.7 3.411 27.14 3.705 ;
      RECT 26.7 3.466 27.15 3.515 ;
      RECT 26.89 2.755 27.06 2.935 ;
      RECT 26.84 2.694 26.89 2.92 ;
      RECT 26.58 2.675 26.84 2.905 ;
      RECT 26.54 2.735 27.01 2.905 ;
      RECT 26.54 2.725 26.97 2.905 ;
      RECT 26.54 2.714 26.95 2.905 ;
      RECT 26.54 2.7 26.89 2.905 ;
      RECT 26.58 2.67 26.776 2.905 ;
      RECT 26.61 2.649 26.776 2.905 ;
      RECT 26.59 2.65 26.776 2.905 ;
      RECT 26.61 2.635 26.69 2.905 ;
      RECT 26.37 3.165 26.49 3.605 ;
      RECT 26.35 3.165 26.49 3.604 ;
      RECT 26.31 3.185 26.49 3.601 ;
      RECT 26.27 3.229 26.49 3.597 ;
      RECT 26.26 3.259 26.51 3.46 ;
      RECT 26.35 3.165 26.52 3.355 ;
      RECT 26.01 1.945 26.02 2.395 ;
      RECT 25.82 1.945 25.84 2.355 ;
      RECT 25.79 1.945 25.8 2.335 ;
      RECT 26.47 2.255 26.49 2.44 ;
      RECT 26.45 2.215 26.47 2.448 ;
      RECT 26.4 2.182 26.45 2.458 ;
      RECT 26.346 2.156 26.4 2.461 ;
      RECT 26.26 2.121 26.346 2.451 ;
      RECT 26.25 2.097 26.26 2.44 ;
      RECT 26.18 2.063 26.25 2.43 ;
      RECT 26.16 2.023 26.18 2.423 ;
      RECT 26.14 2.005 26.16 2.419 ;
      RECT 26.13 1.995 26.14 2.416 ;
      RECT 26.1 1.98 26.13 2.412 ;
      RECT 26.09 1.965 26.1 2.408 ;
      RECT 26.08 1.96 26.09 2.406 ;
      RECT 26.03 1.95 26.08 2.401 ;
      RECT 26.02 1.945 26.03 2.396 ;
      RECT 25.99 1.945 26.01 2.39 ;
      RECT 25.956 1.945 25.99 2.382 ;
      RECT 25.87 1.945 25.956 2.372 ;
      RECT 25.84 1.945 25.87 2.36 ;
      RECT 25.8 1.945 25.82 2.345 ;
      RECT 25.78 1.945 25.79 2.328 ;
      RECT 25.76 1.955 25.78 2.308 ;
      RECT 25.75 1.975 25.76 2.24 ;
      RECT 25.74 1.985 25.75 2 ;
      RECT 26.01 2.665 26.096 2.99 ;
      RECT 26.01 2.665 26.13 2.982 ;
      RECT 25.96 2.665 26.13 2.98 ;
      RECT 25.96 2.669 26.216 2.975 ;
      RECT 25.96 2.674 26.24 2.968 ;
      RECT 25.96 2.68 26.25 2.966 ;
      RECT 25.96 2.69 26.26 2.963 ;
      RECT 25.96 2.83 26.27 2.958 ;
      RECT 26.02 3.34 26.07 3.656 ;
      RECT 26.01 3.32 26.02 3.681 ;
      RECT 26 3.31 26.01 3.69 ;
      RECT 25.98 3.304 26 3.705 ;
      RECT 25.95 3.302 25.98 3.725 ;
      RECT 25.936 3.3 25.95 3.735 ;
      RECT 25.85 3.296 25.936 3.735 ;
      RECT 25.78 3.29 25.85 3.725 ;
      RECT 25.7 3.285 25.78 3.7 ;
      RECT 25.64 3.281 25.7 3.665 ;
      RECT 25.57 3.277 25.64 3.625 ;
      RECT 25.54 3.275 25.57 3.6 ;
      RECT 25.436 3.273 25.48 3.595 ;
      RECT 25.35 3.268 25.436 3.595 ;
      RECT 25.27 3.265 25.35 3.595 ;
      RECT 25.19 3.266 25.27 3.62 ;
      RECT 25.108 3.268 25.19 3.645 ;
      RECT 25.022 3.269 25.108 3.645 ;
      RECT 24.936 3.271 25.022 3.645 ;
      RECT 24.85 3.273 24.936 3.645 ;
      RECT 24.83 3.274 24.85 3.637 ;
      RECT 24.82 3.28 24.83 3.626 ;
      RECT 24.78 3.3 24.82 3.607 ;
      RECT 24.77 3.32 24.78 3.589 ;
      RECT 25.48 3.275 25.54 3.595 ;
      RECT 25.45 2.82 25.62 3.075 ;
      RECT 25.45 2.82 25.63 3.068 ;
      RECT 25.45 2.82 25.64 3.053 ;
      RECT 25.45 2.82 25.66 3.035 ;
      RECT 25.45 2.82 25.7 2.99 ;
      RECT 25.63 2.585 25.72 2.943 ;
      RECT 25.62 2.59 25.73 2.924 ;
      RECT 25.57 2.605 25.74 2.911 ;
      RECT 25.56 2.62 25.75 2.895 ;
      RECT 25.46 2.785 25.75 2.895 ;
      RECT 25.5 2.645 25.62 3.075 ;
      RECT 25.47 2.755 25.75 2.895 ;
      RECT 25.49 2.68 25.62 3.075 ;
      RECT 25.48 2.705 25.75 2.895 ;
      RECT 25.6 2.591 25.73 2.924 ;
      RECT 25.62 2.586 25.72 2.943 ;
      RECT 25.08 2.72 25.27 2.895 ;
      RECT 25.04 2.638 25.23 2.89 ;
      RECT 25.006 2.643 25.23 2.884 ;
      RECT 24.92 2.65 25.23 2.879 ;
      RECT 24.836 2.665 25.23 2.874 ;
      RECT 24.75 2.685 25.26 2.868 ;
      RECT 24.836 2.675 25.26 2.874 ;
      RECT 25.08 2.635 25.23 2.895 ;
      RECT 25.08 2.631 25.18 2.895 ;
      RECT 25.166 2.626 25.18 2.895 ;
      RECT 23.92 1.954 24.58 2.345 ;
      RECT 24.178 1.948 24.58 2.345 ;
      RECT 23.91 1.96 24.58 2.344 ;
      RECT 23.9 1.975 24.58 2.343 ;
      RECT 23.84 2.015 24.58 2.339 ;
      RECT 24.006 1.953 24.59 2.335 ;
      RECT 23.91 1.96 24.6 2.325 ;
      RECT 23.91 1.968 24.61 2.305 ;
      RECT 23.9 1.978 24.63 2.278 ;
      RECT 23.84 2.015 24.64 2.253 ;
      RECT 23.9 1.985 24.65 2.24 ;
      RECT 24.006 1.951 24.58 2.345 ;
      RECT 24.092 1.949 24.58 2.345 ;
      RECT 24.178 1.947 24.56 2.345 ;
      RECT 24.264 1.945 24.56 2.345 ;
      RECT 24.43 3.12 24.6 3.315 ;
      RECT 24.42 3.12 24.6 3.26 ;
      RECT 24.415 3.12 24.6 3.188 ;
      RECT 24.4 3.06 24.58 3.155 ;
      RECT 24.39 3.06 24.58 3.105 ;
      RECT 24.36 3.035 24.57 3.06 ;
      RECT 24.34 3.035 24.57 3.045 ;
      RECT 24.28 2.725 24.46 3.036 ;
      RECT 24.28 2.96 24.56 3.036 ;
      RECT 24.27 2.724 24.28 3.026 ;
      RECT 24.25 2.723 24.27 3.02 ;
      RECT 24.22 2.722 24.25 3 ;
      RECT 24.17 2.719 24.22 2.965 ;
      RECT 24.17 2.84 24.53 2.965 ;
      RECT 24.1 2.716 24.17 2.92 ;
      RECT 24.1 2.775 24.51 2.92 ;
      RECT 24.1 2.765 24.5 2.92 ;
      RECT 24.1 2.755 24.49 2.92 ;
      RECT 24.1 2.735 24.47 2.92 ;
      RECT 24.18 3.255 24.19 3.512 ;
      RECT 24.16 3.172 24.18 3.532 ;
      RECT 24.14 3.166 24.16 3.56 ;
      RECT 24.08 3.154 24.14 3.58 ;
      RECT 24.04 3.14 24.08 3.581 ;
      RECT 23.956 3.129 24.04 3.569 ;
      RECT 23.87 3.116 23.956 3.553 ;
      RECT 23.86 3.109 23.87 3.545 ;
      RECT 23.81 3.106 23.86 3.485 ;
      RECT 23.79 3.102 23.81 3.4 ;
      RECT 23.78 3.1 23.79 3.35 ;
      RECT 23.75 3.098 23.78 3.32 ;
      RECT 23.71 3.093 23.75 3.3 ;
      RECT 23.672 3.088 23.71 3.288 ;
      RECT 23.586 3.08 23.672 3.297 ;
      RECT 23.5 3.069 23.586 3.309 ;
      RECT 23.43 3.059 23.5 3.319 ;
      RECT 23.41 3.05 23.43 3.324 ;
      RECT 23.35 3.022 23.41 3.32 ;
      RECT 23.33 2.992 23.35 3.308 ;
      RECT 23.31 2.965 23.33 3.295 ;
      RECT 23.23 2.718 23.31 3.262 ;
      RECT 23.216 2.71 23.23 3.224 ;
      RECT 23.13 2.702 23.216 3.145 ;
      RECT 23.11 2.693 23.13 3.061 ;
      RECT 23.08 2.688 23.11 3.041 ;
      RECT 23.01 2.699 23.08 3.026 ;
      RECT 22.99 2.717 23.01 3 ;
      RECT 22.98 2.723 22.99 2.945 ;
      RECT 22.96 2.745 22.98 2.83 ;
      RECT 23.62 2.705 23.79 2.895 ;
      RECT 23.62 2.705 23.82 2.89 ;
      RECT 23.67 2.615 23.84 2.88 ;
      RECT 23.63 2.65 23.84 2.88 ;
      RECT 22.83 3.388 22.9 3.829 ;
      RECT 22.77 3.413 22.9 3.826 ;
      RECT 22.77 3.413 22.95 3.819 ;
      RECT 22.76 3.435 22.95 3.816 ;
      RECT 22.9 3.375 22.97 3.814 ;
      RECT 22.83 3.4 23.05 3.811 ;
      RECT 22.76 3.439 23.1 3.807 ;
      RECT 22.74 3.465 23.1 3.795 ;
      RECT 22.76 3.459 23.12 3.79 ;
      RECT 22.74 2.205 22.78 2.445 ;
      RECT 22.74 2.205 22.81 2.444 ;
      RECT 22.74 2.205 22.92 2.436 ;
      RECT 22.74 2.205 22.98 2.415 ;
      RECT 22.75 2.15 23.03 2.315 ;
      RECT 22.86 1.99 22.89 2.437 ;
      RECT 22.89 1.985 23.07 2.195 ;
      RECT 22.76 2.125 23.07 2.195 ;
      RECT 22.81 2.02 22.86 2.44 ;
      RECT 22.78 2.075 23.07 2.195 ;
      RECT 21.65 5.02 21.82 6.49 ;
      RECT 21.65 6.315 21.825 6.485 ;
      RECT 21.28 1.74 21.45 2.93 ;
      RECT 21.28 1.74 21.75 1.91 ;
      RECT 21.28 6.97 21.75 7.14 ;
      RECT 21.28 5.95 21.45 7.14 ;
      RECT 20.29 1.74 20.46 2.93 ;
      RECT 20.29 1.74 20.76 1.91 ;
      RECT 20.29 6.97 20.76 7.14 ;
      RECT 20.29 5.95 20.46 7.14 ;
      RECT 18.44 2.635 18.61 3.865 ;
      RECT 18.495 0.855 18.665 2.805 ;
      RECT 18.44 0.575 18.61 1.025 ;
      RECT 18.44 7.855 18.61 8.305 ;
      RECT 18.495 6.075 18.665 8.025 ;
      RECT 18.44 5.015 18.61 6.245 ;
      RECT 17.92 0.575 18.09 3.865 ;
      RECT 17.92 2.075 18.325 2.405 ;
      RECT 17.92 1.235 18.325 1.565 ;
      RECT 17.92 5.015 18.09 8.305 ;
      RECT 17.92 7.315 18.325 7.645 ;
      RECT 17.92 6.475 18.325 6.805 ;
      RECT 16.015 3.39 16.035 3.44 ;
      RECT 15.995 3.362 16.015 3.555 ;
      RECT 15.975 3.337 15.995 3.611 ;
      RECT 15.935 3.325 15.975 3.63 ;
      RECT 15.885 3.32 15.935 3.659 ;
      RECT 15.881 3.314 15.885 3.675 ;
      RECT 15.795 3.306 15.881 3.675 ;
      RECT 15.735 3.294 15.795 3.67 ;
      RECT 15.681 3.284 15.735 3.659 ;
      RECT 15.595 3.272 15.681 3.642 ;
      RECT 15.573 3.263 15.595 3.629 ;
      RECT 15.487 3.256 15.573 3.616 ;
      RECT 15.401 3.243 15.487 3.595 ;
      RECT 15.315 3.231 15.401 3.575 ;
      RECT 15.285 3.22 15.315 3.561 ;
      RECT 15.235 3.207 15.285 3.551 ;
      RECT 15.215 3.197 15.235 3.545 ;
      RECT 15.161 3.187 15.215 3.539 ;
      RECT 15.075 3.167 15.161 3.523 ;
      RECT 15.035 3.155 15.075 3.509 ;
      RECT 15 3.155 15.035 3.495 ;
      RECT 14.985 3.155 15 3.48 ;
      RECT 14.935 3.155 14.985 3.425 ;
      RECT 14.905 3.155 14.935 3.345 ;
      RECT 15.435 2.825 15.605 3.075 ;
      RECT 15.435 2.825 15.615 3.03 ;
      RECT 15.495 2.655 15.625 2.975 ;
      RECT 15.495 2.662 15.635 2.94 ;
      RECT 15.455 2.677 15.645 2.875 ;
      RECT 15.445 2.76 15.645 2.875 ;
      RECT 15.455 2.695 15.655 2.785 ;
      RECT 15.455 2.675 15.635 2.94 ;
      RECT 15.225 1.93 15.395 2.415 ;
      RECT 15.215 1.93 15.395 2.405 ;
      RECT 15.215 1.945 15.415 2.35 ;
      RECT 15.175 1.925 15.365 2.315 ;
      RECT 15.175 1.96 15.425 2.235 ;
      RECT 15.125 1.945 15.415 2.135 ;
      RECT 15.125 1.975 15.435 2.095 ;
      RECT 15.125 1.99 15.445 2.015 ;
      RECT 14.721 2.688 14.735 2.944 ;
      RECT 14.721 2.689 14.821 2.939 ;
      RECT 14.635 2.686 14.721 2.936 ;
      RECT 14.625 2.685 14.635 2.929 ;
      RECT 14.625 2.692 14.907 2.926 ;
      RECT 14.545 2.695 14.907 2.922 ;
      RECT 14.625 2.694 14.925 2.919 ;
      RECT 14.535 2.707 14.945 2.916 ;
      RECT 14.545 2.695 14.945 2.916 ;
      RECT 14.525 2.712 14.945 2.915 ;
      RECT 14.545 2.697 15.031 2.911 ;
      RECT 14.505 2.715 15.031 2.908 ;
      RECT 14.545 2.701 15.117 2.902 ;
      RECT 14.495 2.72 15.117 2.898 ;
      RECT 14.545 2.704 15.145 2.897 ;
      RECT 14.545 2.705 15.185 2.891 ;
      RECT 14.535 2.71 15.195 2.886 ;
      RECT 14.495 2.73 15.205 2.875 ;
      RECT 14.495 2.75 15.215 2.86 ;
      RECT 14.455 3.298 14.475 3.605 ;
      RECT 14.445 3.273 14.455 3.885 ;
      RECT 14.405 3.24 14.445 3.885 ;
      RECT 14.401 3.21 14.405 3.885 ;
      RECT 14.315 3.095 14.401 3.885 ;
      RECT 14.305 2.97 14.315 3.885 ;
      RECT 14.295 2.935 14.305 3.885 ;
      RECT 14.285 2.905 14.295 3.885 ;
      RECT 14.265 2.875 14.285 3.77 ;
      RECT 14.255 2.845 14.265 3.645 ;
      RECT 14.245 2.825 14.255 3.595 ;
      RECT 14.225 2.795 14.245 3.503 ;
      RECT 14.205 2.761 14.225 3.418 ;
      RECT 14.2 2.744 14.205 3.353 ;
      RECT 14.195 2.738 14.2 3.325 ;
      RECT 14.185 2.73 14.195 3.29 ;
      RECT 14.165 2.725 14.175 3.19 ;
      RECT 14.155 2.725 14.165 3.165 ;
      RECT 14.15 2.725 14.155 3.128 ;
      RECT 14.135 2.725 14.15 3.06 ;
      RECT 14.125 2.724 14.135 2.99 ;
      RECT 14.115 2.722 14.125 2.97 ;
      RECT 14.055 2.718 14.115 2.943 ;
      RECT 14.015 2.72 14.055 2.923 ;
      RECT 13.995 2.75 14.015 2.905 ;
      RECT 14.175 2.725 14.185 3.245 ;
      RECT 14.115 2.08 14.285 2.435 ;
      RECT 14.145 1.966 14.285 2.435 ;
      RECT 14.145 1.968 14.295 2.43 ;
      RECT 14.145 1.97 14.315 2.42 ;
      RECT 14.145 1.973 14.345 2.405 ;
      RECT 14.145 1.978 14.395 2.375 ;
      RECT 14.145 1.983 14.415 2.338 ;
      RECT 14.125 1.985 14.425 2.313 ;
      RECT 14.145 1.965 14.255 2.435 ;
      RECT 14.155 1.96 14.255 2.435 ;
      RECT 13.675 3.222 13.865 3.585 ;
      RECT 13.675 3.237 13.905 3.583 ;
      RECT 13.675 3.265 13.925 3.579 ;
      RECT 13.675 3.3 13.935 3.577 ;
      RECT 13.675 3.345 13.945 3.576 ;
      RECT 13.665 3.217 13.825 3.565 ;
      RECT 13.645 3.225 13.865 3.515 ;
      RECT 13.615 3.237 13.905 3.45 ;
      RECT 13.675 3.215 13.825 3.585 ;
      RECT 13.68 7.855 13.85 8.305 ;
      RECT 13.735 6.075 13.905 8.025 ;
      RECT 13.68 5.015 13.85 6.245 ;
      RECT 13.16 5.015 13.33 8.305 ;
      RECT 13.16 7.315 13.565 7.645 ;
      RECT 13.16 6.475 13.565 6.805 ;
      RECT 13.261 2.695 13.465 3.105 ;
      RECT 13.175 2.588 13.261 3.09 ;
      RECT 13.171 2.584 13.175 3.074 ;
      RECT 13.085 2.695 13.465 3.054 ;
      RECT 13.065 2.575 13.085 3.015 ;
      RECT 13.055 2.58 13.171 2.99 ;
      RECT 13.045 2.587 13.175 2.97 ;
      RECT 13.035 2.592 13.265 2.945 ;
      RECT 13.025 2.61 13.355 2.925 ;
      RECT 13.015 2.615 13.355 2.905 ;
      RECT 13.005 2.62 13.395 2.77 ;
      RECT 13.005 2.65 13.455 2.77 ;
      RECT 13.005 2.635 13.445 2.77 ;
      RECT 13.035 2.605 13.355 2.945 ;
      RECT 13.035 2.593 13.295 2.945 ;
      RECT 13.185 3.42 13.435 3.885 ;
      RECT 13.105 3.395 13.425 3.88 ;
      RECT 13.035 3.429 13.435 3.87 ;
      RECT 12.825 3.68 13.435 3.865 ;
      RECT 13.005 3.449 13.435 3.865 ;
      RECT 12.845 3.64 13.435 3.865 ;
      RECT 12.995 3.46 13.435 3.865 ;
      RECT 12.885 3.58 13.435 3.865 ;
      RECT 12.935 3.505 13.435 3.865 ;
      RECT 13.185 3.37 13.425 3.885 ;
      RECT 13.205 3.365 13.425 3.885 ;
      RECT 13.215 3.36 13.345 3.885 ;
      RECT 13.301 3.355 13.305 3.885 ;
      RECT 12.775 1.925 12.861 2.362 ;
      RECT 12.765 1.925 12.861 2.358 ;
      RECT 12.765 1.925 12.925 2.357 ;
      RECT 12.765 1.925 12.955 2.355 ;
      RECT 12.765 1.925 12.965 2.345 ;
      RECT 12.755 1.93 12.965 2.343 ;
      RECT 12.745 1.94 12.965 2.335 ;
      RECT 12.745 1.94 12.975 2.295 ;
      RECT 12.765 1.925 12.995 2.21 ;
      RECT 12.735 1.95 12.995 2.205 ;
      RECT 12.745 1.94 13.005 2.135 ;
      RECT 12.725 1.96 13.005 2.08 ;
      RECT 12.715 1.97 13.005 1.98 ;
      RECT 12.795 2.741 12.805 2.82 ;
      RECT 12.785 2.734 12.795 3.005 ;
      RECT 12.775 2.728 12.785 3.03 ;
      RECT 12.765 2.72 12.775 3.06 ;
      RECT 12.725 2.715 12.765 3.11 ;
      RECT 12.705 2.715 12.725 3.165 ;
      RECT 12.695 2.715 12.705 3.19 ;
      RECT 12.685 2.715 12.695 3.205 ;
      RECT 12.655 2.715 12.685 3.25 ;
      RECT 12.645 2.715 12.655 3.29 ;
      RECT 12.625 2.715 12.645 3.315 ;
      RECT 12.605 2.715 12.625 3.35 ;
      RECT 12.525 2.715 12.605 3.395 ;
      RECT 12.515 2.715 12.525 3.415 ;
      RECT 12.475 2.795 12.515 3.412 ;
      RECT 12.455 2.875 12.475 3.409 ;
      RECT 12.435 2.93 12.455 3.407 ;
      RECT 12.415 2.99 12.435 3.405 ;
      RECT 12.375 3.025 12.415 3.403 ;
      RECT 12.371 3.035 12.375 3.401 ;
      RECT 12.285 3.05 12.371 3.397 ;
      RECT 12.265 3.07 12.285 3.393 ;
      RECT 12.195 3.075 12.265 3.389 ;
      RECT 12.175 3.076 12.195 3.386 ;
      RECT 12.171 3.078 12.175 3.385 ;
      RECT 12.085 3.087 12.171 3.38 ;
      RECT 12.075 3.096 12.085 3.375 ;
      RECT 12.035 3.102 12.075 3.37 ;
      RECT 11.985 3.113 12.035 3.355 ;
      RECT 11.965 3.122 11.985 3.34 ;
      RECT 11.885 3.135 11.965 3.325 ;
      RECT 12.055 2.685 12.225 2.895 ;
      RECT 12.171 2.677 12.225 2.895 ;
      RECT 11.971 2.685 12.225 2.885 ;
      RECT 11.885 2.685 12.225 2.865 ;
      RECT 11.885 2.69 12.235 2.81 ;
      RECT 11.885 2.7 12.245 2.72 ;
      RECT 12.085 2.682 12.225 2.895 ;
      RECT 11.835 3.623 12.085 3.955 ;
      RECT 11.805 3.635 12.085 3.937 ;
      RECT 11.785 3.67 12.085 3.907 ;
      RECT 11.835 3.62 12.007 3.955 ;
      RECT 11.835 3.616 11.921 3.955 ;
      RECT 11.765 1.965 11.945 2.385 ;
      RECT 11.765 1.965 11.965 2.375 ;
      RECT 11.765 1.965 11.985 2.35 ;
      RECT 11.765 1.965 11.995 2.335 ;
      RECT 11.765 1.965 12.005 2.33 ;
      RECT 11.765 2.005 12.025 2.315 ;
      RECT 11.765 2.075 12.045 2.295 ;
      RECT 11.745 2.075 12.045 2.29 ;
      RECT 11.745 2.135 12.055 2.265 ;
      RECT 11.745 2.175 12.065 2.215 ;
      RECT 11.725 1.965 12.005 2.195 ;
      RECT 11.715 1.975 12.005 2.118 ;
      RECT 11.705 2.015 12.025 2.063 ;
      RECT 11.305 3.375 11.475 3.895 ;
      RECT 11.295 3.375 11.475 3.855 ;
      RECT 11.285 3.395 11.475 3.83 ;
      RECT 11.295 3.375 11.485 3.825 ;
      RECT 11.275 3.435 11.485 3.795 ;
      RECT 11.265 3.47 11.485 3.775 ;
      RECT 11.255 3.52 11.485 3.735 ;
      RECT 11.295 3.386 11.495 3.725 ;
      RECT 11.245 3.6 11.495 3.675 ;
      RECT 11.285 3.409 11.505 3.605 ;
      RECT 11.285 3.433 11.515 3.5 ;
      RECT 11.225 2.68 11.245 2.955 ;
      RECT 11.185 2.665 11.225 3 ;
      RECT 11.165 2.65 11.185 3.065 ;
      RECT 11.145 2.649 11.165 3.14 ;
      RECT 11.125 2.657 11.145 3.245 ;
      RECT 11.121 2.662 11.125 3.297 ;
      RECT 11.035 2.681 11.121 3.337 ;
      RECT 11.025 2.702 11.035 3.376 ;
      RECT 11.015 2.71 11.025 3.377 ;
      RECT 10.995 2.845 11.015 3.379 ;
      RECT 10.985 2.995 10.995 3.381 ;
      RECT 10.945 3.08 10.985 3.386 ;
      RECT 10.863 3.102 10.945 3.396 ;
      RECT 10.777 3.117 10.863 3.409 ;
      RECT 10.691 3.132 10.777 3.422 ;
      RECT 10.605 3.147 10.691 3.436 ;
      RECT 10.525 3.161 10.605 3.449 ;
      RECT 10.511 3.169 10.525 3.457 ;
      RECT 10.425 3.177 10.511 3.471 ;
      RECT 10.415 3.185 10.425 3.484 ;
      RECT 10.391 3.185 10.415 3.492 ;
      RECT 10.305 3.187 10.391 3.522 ;
      RECT 10.225 3.189 10.305 3.565 ;
      RECT 10.155 3.192 10.225 3.6 ;
      RECT 10.135 3.194 10.155 3.616 ;
      RECT 10.105 3.2 10.135 3.618 ;
      RECT 10.055 3.215 10.105 3.621 ;
      RECT 10.035 3.23 10.055 3.624 ;
      RECT 10.005 3.235 10.035 3.627 ;
      RECT 9.945 3.25 10.005 3.631 ;
      RECT 9.935 3.266 9.945 3.635 ;
      RECT 9.885 3.276 9.935 3.624 ;
      RECT 9.855 3.295 9.885 3.607 ;
      RECT 9.835 3.315 9.855 3.597 ;
      RECT 9.815 3.34 9.835 3.589 ;
      RECT 10.825 1.932 10.995 2.425 ;
      RECT 10.815 1.932 10.995 2.41 ;
      RECT 10.815 1.947 11.025 2.4 ;
      RECT 10.805 1.947 11.025 2.375 ;
      RECT 10.795 1.947 11.025 2.34 ;
      RECT 10.795 1.955 11.035 2.295 ;
      RECT 10.775 1.925 10.965 2.275 ;
      RECT 10.765 1.932 10.995 2.235 ;
      RECT 10.755 1.947 11.025 2.215 ;
      RECT 10.745 1.96 11.035 2.175 ;
      RECT 10.735 1.975 11.035 2.128 ;
      RECT 10.735 1.975 11.045 2.12 ;
      RECT 10.725 1.99 11.045 2.093 ;
      RECT 10.735 1.985 11.055 2.035 ;
      RECT 10.535 2.612 10.805 2.905 ;
      RECT 10.535 2.614 10.815 2.9 ;
      RECT 10.525 2.64 10.815 2.895 ;
      RECT 10.535 2.63 10.825 2.89 ;
      RECT 10.535 2.608 10.771 2.905 ;
      RECT 10.535 2.605 10.685 2.905 ;
      RECT 10.595 2.6 10.681 2.905 ;
      RECT 10.085 2.648 10.155 2.945 ;
      RECT 10.085 2.648 10.165 2.944 ;
      RECT 10.165 2.635 10.175 2.941 ;
      RECT 10.065 2.662 10.175 2.935 ;
      RECT 10.155 2.64 10.245 2.931 ;
      RECT 10.085 2.655 10.265 2.92 ;
      RECT 10.065 2.72 10.275 2.916 ;
      RECT 10.045 2.668 10.265 2.915 ;
      RECT 10.035 2.673 10.265 2.905 ;
      RECT 10.025 2.795 10.285 2.9 ;
      RECT 10.025 2.875 10.295 2.89 ;
      RECT 9.995 2.681 10.265 2.884 ;
      RECT 9.985 2.695 10.265 2.869 ;
      RECT 10.025 2.676 10.265 2.9 ;
      RECT 10.155 2.636 10.175 2.941 ;
      RECT 9.975 2.072 9.995 2.305 ;
      RECT 9.965 2.053 9.975 2.31 ;
      RECT 9.955 2.041 9.965 2.317 ;
      RECT 9.915 2.027 9.955 2.327 ;
      RECT 9.905 2.017 9.915 2.336 ;
      RECT 9.855 2.002 9.905 2.341 ;
      RECT 9.845 1.987 9.855 2.347 ;
      RECT 9.825 1.978 9.845 2.352 ;
      RECT 9.815 1.968 9.825 2.358 ;
      RECT 9.805 1.965 9.815 2.363 ;
      RECT 9.785 1.965 9.805 2.364 ;
      RECT 9.755 1.96 9.785 2.362 ;
      RECT 9.731 1.953 9.755 2.361 ;
      RECT 9.645 1.943 9.731 2.358 ;
      RECT 9.635 1.935 9.645 2.355 ;
      RECT 9.613 1.935 9.635 2.354 ;
      RECT 9.527 1.935 9.613 2.352 ;
      RECT 9.441 1.935 9.527 2.35 ;
      RECT 9.355 1.935 9.441 2.347 ;
      RECT 9.345 1.935 9.355 2.34 ;
      RECT 9.315 1.935 9.345 2.3 ;
      RECT 9.305 1.945 9.315 2.255 ;
      RECT 9.295 1.99 9.305 2.24 ;
      RECT 9.265 2.085 9.295 2.195 ;
      RECT 9.455 2.822 9.625 3.335 ;
      RECT 9.445 2.853 9.625 3.315 ;
      RECT 9.445 2.853 9.645 3.285 ;
      RECT 9.435 2.861 9.645 3.26 ;
      RECT 9.435 2.861 9.655 3.25 ;
      RECT 9.435 2.861 9.665 3.23 ;
      RECT 9.435 2.861 9.715 3.185 ;
      RECT 9.435 2.861 9.725 3.16 ;
      RECT 9.435 2.861 9.735 3.125 ;
      RECT 9.435 2.861 9.745 3.09 ;
      RECT 9.435 2.861 9.755 3.04 ;
      RECT 9.435 2.861 9.775 2.965 ;
      RECT 9.605 2.725 9.785 2.905 ;
      RECT 9.525 2.78 9.785 2.905 ;
      RECT 9.565 2.745 9.625 3.335 ;
      RECT 9.555 2.765 9.785 2.905 ;
      RECT 8.915 3.235 9.001 3.801 ;
      RECT 8.875 3.235 9.001 3.795 ;
      RECT 8.875 3.235 9.087 3.793 ;
      RECT 8.875 3.235 9.125 3.787 ;
      RECT 8.875 3.242 9.135 3.785 ;
      RECT 8.845 3.235 9.125 3.78 ;
      RECT 8.815 3.25 9.135 3.77 ;
      RECT 8.815 3.277 9.175 3.762 ;
      RECT 8.79 3.277 9.175 3.75 ;
      RECT 8.79 3.315 9.185 3.732 ;
      RECT 8.775 3.297 9.175 3.725 ;
      RECT 8.775 3.345 9.195 3.721 ;
      RECT 8.775 3.411 9.215 3.705 ;
      RECT 8.775 3.466 9.225 3.515 ;
      RECT 8.965 2.755 9.135 2.935 ;
      RECT 8.915 2.694 8.965 2.92 ;
      RECT 8.655 2.675 8.915 2.905 ;
      RECT 8.615 2.735 9.085 2.905 ;
      RECT 8.615 2.725 9.045 2.905 ;
      RECT 8.615 2.714 9.025 2.905 ;
      RECT 8.615 2.7 8.965 2.905 ;
      RECT 8.655 2.67 8.851 2.905 ;
      RECT 8.685 2.649 8.851 2.905 ;
      RECT 8.665 2.65 8.851 2.905 ;
      RECT 8.685 2.635 8.765 2.905 ;
      RECT 8.445 3.165 8.565 3.605 ;
      RECT 8.425 3.165 8.565 3.604 ;
      RECT 8.385 3.185 8.565 3.601 ;
      RECT 8.345 3.229 8.565 3.597 ;
      RECT 8.335 3.259 8.585 3.46 ;
      RECT 8.425 3.165 8.595 3.355 ;
      RECT 8.085 1.945 8.095 2.395 ;
      RECT 7.895 1.945 7.915 2.355 ;
      RECT 7.865 1.945 7.875 2.335 ;
      RECT 8.545 2.255 8.565 2.44 ;
      RECT 8.525 2.215 8.545 2.448 ;
      RECT 8.475 2.182 8.525 2.458 ;
      RECT 8.421 2.156 8.475 2.461 ;
      RECT 8.335 2.121 8.421 2.451 ;
      RECT 8.325 2.097 8.335 2.44 ;
      RECT 8.255 2.063 8.325 2.43 ;
      RECT 8.235 2.023 8.255 2.423 ;
      RECT 8.215 2.005 8.235 2.419 ;
      RECT 8.205 1.995 8.215 2.416 ;
      RECT 8.175 1.98 8.205 2.412 ;
      RECT 8.165 1.965 8.175 2.408 ;
      RECT 8.155 1.96 8.165 2.406 ;
      RECT 8.105 1.95 8.155 2.401 ;
      RECT 8.095 1.945 8.105 2.396 ;
      RECT 8.065 1.945 8.085 2.39 ;
      RECT 8.031 1.945 8.065 2.382 ;
      RECT 7.945 1.945 8.031 2.372 ;
      RECT 7.915 1.945 7.945 2.36 ;
      RECT 7.875 1.945 7.895 2.345 ;
      RECT 7.855 1.945 7.865 2.328 ;
      RECT 7.835 1.955 7.855 2.308 ;
      RECT 7.825 1.975 7.835 2.24 ;
      RECT 7.815 1.985 7.825 2 ;
      RECT 8.085 2.665 8.171 2.99 ;
      RECT 8.085 2.665 8.205 2.982 ;
      RECT 8.035 2.665 8.205 2.98 ;
      RECT 8.035 2.669 8.291 2.975 ;
      RECT 8.035 2.674 8.315 2.968 ;
      RECT 8.035 2.68 8.325 2.966 ;
      RECT 8.035 2.69 8.335 2.963 ;
      RECT 8.035 2.83 8.345 2.958 ;
      RECT 8.095 3.34 8.145 3.656 ;
      RECT 8.085 3.32 8.095 3.681 ;
      RECT 8.075 3.31 8.085 3.69 ;
      RECT 8.055 3.304 8.075 3.705 ;
      RECT 8.025 3.302 8.055 3.725 ;
      RECT 8.011 3.3 8.025 3.735 ;
      RECT 7.925 3.296 8.011 3.735 ;
      RECT 7.855 3.29 7.925 3.725 ;
      RECT 7.775 3.285 7.855 3.7 ;
      RECT 7.715 3.281 7.775 3.665 ;
      RECT 7.645 3.277 7.715 3.625 ;
      RECT 7.615 3.275 7.645 3.6 ;
      RECT 7.511 3.273 7.555 3.595 ;
      RECT 7.425 3.268 7.511 3.595 ;
      RECT 7.345 3.265 7.425 3.595 ;
      RECT 7.265 3.266 7.345 3.62 ;
      RECT 7.183 3.268 7.265 3.645 ;
      RECT 7.097 3.269 7.183 3.645 ;
      RECT 7.011 3.271 7.097 3.645 ;
      RECT 6.925 3.273 7.011 3.645 ;
      RECT 6.905 3.274 6.925 3.637 ;
      RECT 6.895 3.28 6.905 3.626 ;
      RECT 6.855 3.3 6.895 3.607 ;
      RECT 6.845 3.32 6.855 3.589 ;
      RECT 7.555 3.275 7.615 3.595 ;
      RECT 7.525 2.82 7.695 3.075 ;
      RECT 7.525 2.82 7.705 3.068 ;
      RECT 7.525 2.82 7.715 3.053 ;
      RECT 7.525 2.82 7.735 3.035 ;
      RECT 7.525 2.82 7.775 2.99 ;
      RECT 7.705 2.585 7.795 2.943 ;
      RECT 7.695 2.59 7.805 2.924 ;
      RECT 7.645 2.605 7.815 2.911 ;
      RECT 7.635 2.62 7.825 2.895 ;
      RECT 7.535 2.785 7.825 2.895 ;
      RECT 7.575 2.645 7.695 3.075 ;
      RECT 7.545 2.755 7.825 2.895 ;
      RECT 7.565 2.68 7.695 3.075 ;
      RECT 7.555 2.705 7.825 2.895 ;
      RECT 7.675 2.591 7.805 2.924 ;
      RECT 7.695 2.586 7.795 2.943 ;
      RECT 7.155 2.72 7.345 2.895 ;
      RECT 7.115 2.638 7.305 2.89 ;
      RECT 7.081 2.643 7.305 2.884 ;
      RECT 6.995 2.65 7.305 2.879 ;
      RECT 6.911 2.665 7.305 2.874 ;
      RECT 6.825 2.685 7.335 2.868 ;
      RECT 6.911 2.675 7.335 2.874 ;
      RECT 7.155 2.635 7.305 2.895 ;
      RECT 7.155 2.631 7.255 2.895 ;
      RECT 7.241 2.626 7.255 2.895 ;
      RECT 5.995 1.954 6.655 2.345 ;
      RECT 6.253 1.948 6.655 2.345 ;
      RECT 5.985 1.96 6.655 2.344 ;
      RECT 5.975 1.975 6.655 2.343 ;
      RECT 5.915 2.015 6.655 2.339 ;
      RECT 6.081 1.953 6.665 2.335 ;
      RECT 5.985 1.96 6.675 2.325 ;
      RECT 5.985 1.968 6.685 2.305 ;
      RECT 5.975 1.978 6.705 2.278 ;
      RECT 5.915 2.015 6.715 2.253 ;
      RECT 5.975 1.985 6.725 2.24 ;
      RECT 6.081 1.951 6.655 2.345 ;
      RECT 6.167 1.949 6.655 2.345 ;
      RECT 6.253 1.947 6.635 2.345 ;
      RECT 6.339 1.945 6.635 2.345 ;
      RECT 6.505 3.12 6.675 3.315 ;
      RECT 6.495 3.12 6.675 3.26 ;
      RECT 6.49 3.12 6.675 3.188 ;
      RECT 6.475 3.06 6.655 3.155 ;
      RECT 6.465 3.06 6.655 3.105 ;
      RECT 6.435 3.035 6.645 3.06 ;
      RECT 6.415 3.035 6.645 3.045 ;
      RECT 6.355 2.725 6.535 3.036 ;
      RECT 6.355 2.96 6.635 3.036 ;
      RECT 6.345 2.724 6.355 3.026 ;
      RECT 6.325 2.723 6.345 3.02 ;
      RECT 6.295 2.722 6.325 3 ;
      RECT 6.245 2.719 6.295 2.965 ;
      RECT 6.245 2.84 6.605 2.965 ;
      RECT 6.175 2.716 6.245 2.92 ;
      RECT 6.175 2.775 6.585 2.92 ;
      RECT 6.175 2.765 6.575 2.92 ;
      RECT 6.175 2.755 6.565 2.92 ;
      RECT 6.175 2.735 6.545 2.92 ;
      RECT 6.255 3.255 6.265 3.512 ;
      RECT 6.235 3.172 6.255 3.532 ;
      RECT 6.215 3.166 6.235 3.56 ;
      RECT 6.155 3.154 6.215 3.58 ;
      RECT 6.115 3.14 6.155 3.581 ;
      RECT 6.031 3.129 6.115 3.569 ;
      RECT 5.945 3.116 6.031 3.553 ;
      RECT 5.935 3.109 5.945 3.545 ;
      RECT 5.885 3.106 5.935 3.485 ;
      RECT 5.865 3.102 5.885 3.4 ;
      RECT 5.855 3.1 5.865 3.35 ;
      RECT 5.825 3.098 5.855 3.32 ;
      RECT 5.785 3.093 5.825 3.3 ;
      RECT 5.747 3.088 5.785 3.288 ;
      RECT 5.661 3.08 5.747 3.297 ;
      RECT 5.575 3.069 5.661 3.309 ;
      RECT 5.505 3.059 5.575 3.319 ;
      RECT 5.485 3.05 5.505 3.324 ;
      RECT 5.425 3.022 5.485 3.32 ;
      RECT 5.405 2.992 5.425 3.308 ;
      RECT 5.385 2.965 5.405 3.295 ;
      RECT 5.305 2.718 5.385 3.262 ;
      RECT 5.291 2.71 5.305 3.224 ;
      RECT 5.205 2.702 5.291 3.145 ;
      RECT 5.185 2.693 5.205 3.061 ;
      RECT 5.155 2.688 5.185 3.041 ;
      RECT 5.085 2.699 5.155 3.026 ;
      RECT 5.065 2.717 5.085 3 ;
      RECT 5.055 2.723 5.065 2.945 ;
      RECT 5.035 2.745 5.055 2.83 ;
      RECT 5.695 2.705 5.865 2.895 ;
      RECT 5.695 2.705 5.895 2.89 ;
      RECT 5.745 2.615 5.915 2.88 ;
      RECT 5.705 2.65 5.915 2.88 ;
      RECT 4.905 3.388 4.975 3.829 ;
      RECT 4.845 3.413 4.975 3.826 ;
      RECT 4.845 3.413 5.025 3.819 ;
      RECT 4.835 3.435 5.025 3.816 ;
      RECT 4.975 3.375 5.045 3.814 ;
      RECT 4.905 3.4 5.125 3.811 ;
      RECT 4.835 3.439 5.175 3.807 ;
      RECT 4.815 3.465 5.175 3.795 ;
      RECT 4.835 3.459 5.195 3.79 ;
      RECT 4.815 2.205 4.855 2.445 ;
      RECT 4.815 2.205 4.885 2.444 ;
      RECT 4.815 2.205 4.995 2.436 ;
      RECT 4.815 2.205 5.055 2.415 ;
      RECT 4.825 2.15 5.105 2.315 ;
      RECT 4.935 1.99 4.965 2.437 ;
      RECT 4.965 1.985 5.145 2.195 ;
      RECT 4.835 2.125 5.145 2.195 ;
      RECT 4.885 2.02 4.935 2.44 ;
      RECT 4.855 2.075 5.145 2.195 ;
      RECT 2.65 7.855 2.82 8.305 ;
      RECT 2.705 6.075 2.875 8.025 ;
      RECT 2.65 5.015 2.82 6.245 ;
      RECT 2.13 5.015 2.3 8.305 ;
      RECT 2.13 7.315 2.535 7.645 ;
      RECT 2.13 6.475 2.535 6.805 ;
      RECT 93.35 7.8 93.52 8.31 ;
      RECT 92.36 0.57 92.53 1.08 ;
      RECT 92.36 2.39 92.53 3.86 ;
      RECT 92.36 5.02 92.53 6.49 ;
      RECT 92.36 7.8 92.53 8.31 ;
      RECT 91 0.575 91.17 3.865 ;
      RECT 91 5.015 91.17 8.305 ;
      RECT 90.57 0.575 90.74 1.085 ;
      RECT 90.57 1.655 90.74 3.865 ;
      RECT 90.57 5.015 90.74 7.225 ;
      RECT 90.57 7.795 90.74 8.305 ;
      RECT 86.24 5.015 86.41 8.305 ;
      RECT 85.81 5.015 85.98 7.225 ;
      RECT 85.81 7.795 85.98 8.305 ;
      RECT 75.425 7.8 75.595 8.31 ;
      RECT 74.435 0.57 74.605 1.08 ;
      RECT 74.435 2.39 74.605 3.86 ;
      RECT 74.435 5.02 74.605 6.49 ;
      RECT 74.435 7.8 74.605 8.31 ;
      RECT 73.075 0.575 73.245 3.865 ;
      RECT 73.075 5.015 73.245 8.305 ;
      RECT 72.645 0.575 72.815 1.085 ;
      RECT 72.645 1.655 72.815 3.865 ;
      RECT 72.645 5.015 72.815 7.225 ;
      RECT 72.645 7.795 72.815 8.305 ;
      RECT 68.315 5.015 68.485 8.305 ;
      RECT 67.885 5.015 68.055 7.225 ;
      RECT 67.885 7.795 68.055 8.305 ;
      RECT 57.5 7.8 57.67 8.31 ;
      RECT 56.51 0.57 56.68 1.08 ;
      RECT 56.51 2.39 56.68 3.86 ;
      RECT 56.51 5.02 56.68 6.49 ;
      RECT 56.51 7.8 56.68 8.31 ;
      RECT 55.15 0.575 55.32 3.865 ;
      RECT 55.15 5.015 55.32 8.305 ;
      RECT 54.72 0.575 54.89 1.085 ;
      RECT 54.72 1.655 54.89 3.865 ;
      RECT 54.72 5.015 54.89 7.225 ;
      RECT 54.72 7.795 54.89 8.305 ;
      RECT 50.39 5.015 50.56 8.305 ;
      RECT 49.96 5.015 50.13 7.225 ;
      RECT 49.96 7.795 50.13 8.305 ;
      RECT 39.575 7.8 39.745 8.31 ;
      RECT 38.585 0.57 38.755 1.08 ;
      RECT 38.585 2.39 38.755 3.86 ;
      RECT 38.585 5.02 38.755 6.49 ;
      RECT 38.585 7.8 38.755 8.31 ;
      RECT 37.225 0.575 37.395 3.865 ;
      RECT 37.225 5.015 37.395 8.305 ;
      RECT 36.795 0.575 36.965 1.085 ;
      RECT 36.795 1.655 36.965 3.865 ;
      RECT 36.795 5.015 36.965 7.225 ;
      RECT 36.795 7.795 36.965 8.305 ;
      RECT 32.465 5.015 32.635 8.305 ;
      RECT 32.035 5.015 32.205 7.225 ;
      RECT 32.035 7.795 32.205 8.305 ;
      RECT 21.65 7.8 21.82 8.31 ;
      RECT 20.66 0.57 20.83 1.08 ;
      RECT 20.66 2.39 20.83 3.86 ;
      RECT 20.66 5.02 20.83 6.49 ;
      RECT 20.66 7.8 20.83 8.31 ;
      RECT 19.3 0.575 19.47 3.865 ;
      RECT 19.3 5.015 19.47 8.305 ;
      RECT 18.87 0.575 19.04 1.085 ;
      RECT 18.87 1.655 19.04 3.865 ;
      RECT 18.87 5.015 19.04 7.225 ;
      RECT 18.87 7.795 19.04 8.305 ;
      RECT 14.54 5.015 14.71 8.305 ;
      RECT 14.11 5.015 14.28 7.225 ;
      RECT 14.11 7.795 14.28 8.305 ;
      RECT 3.08 5.015 3.25 7.225 ;
      RECT 3.08 7.795 3.25 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8_b0r2 ;
  SIZE 92.575 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 20.335 0.915 20.505 1.085 ;
        RECT 20.33 0.91 20.5 1.08 ;
        RECT 20.33 2.39 20.5 2.56 ;
      LAYER li1 ;
        RECT 20.335 0.915 20.505 1.085 ;
        RECT 20.33 0.57 20.5 1.08 ;
        RECT 20.33 2.39 20.5 3.86 ;
      LAYER met1 ;
        RECT 20.27 2.36 20.56 2.59 ;
        RECT 20.27 0.88 20.56 1.11 ;
        RECT 20.33 0.88 20.5 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 38.26 0.915 38.43 1.085 ;
        RECT 38.255 0.91 38.425 1.08 ;
        RECT 38.255 2.39 38.425 2.56 ;
      LAYER li1 ;
        RECT 38.26 0.915 38.43 1.085 ;
        RECT 38.255 0.57 38.425 1.08 ;
        RECT 38.255 2.39 38.425 3.86 ;
      LAYER met1 ;
        RECT 38.195 2.36 38.485 2.59 ;
        RECT 38.195 0.88 38.485 1.11 ;
        RECT 38.255 0.88 38.425 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 56.185 0.915 56.355 1.085 ;
        RECT 56.18 0.91 56.35 1.08 ;
        RECT 56.18 2.39 56.35 2.56 ;
      LAYER li1 ;
        RECT 56.185 0.915 56.355 1.085 ;
        RECT 56.18 0.57 56.35 1.08 ;
        RECT 56.18 2.39 56.35 3.86 ;
      LAYER met1 ;
        RECT 56.12 2.36 56.41 2.59 ;
        RECT 56.12 0.88 56.41 1.11 ;
        RECT 56.18 0.88 56.35 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 74.11 0.915 74.28 1.085 ;
        RECT 74.105 0.91 74.275 1.08 ;
        RECT 74.105 2.39 74.275 2.56 ;
      LAYER li1 ;
        RECT 74.11 0.915 74.28 1.085 ;
        RECT 74.105 0.57 74.275 1.08 ;
        RECT 74.105 2.39 74.275 3.86 ;
      LAYER met1 ;
        RECT 74.045 2.36 74.335 2.59 ;
        RECT 74.045 0.88 74.335 1.11 ;
        RECT 74.105 0.88 74.275 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 92.035 0.915 92.205 1.085 ;
        RECT 92.03 0.91 92.2 1.08 ;
        RECT 92.03 2.39 92.2 2.56 ;
      LAYER li1 ;
        RECT 92.035 0.915 92.205 1.085 ;
        RECT 92.03 0.57 92.2 1.08 ;
        RECT 92.03 2.39 92.2 3.86 ;
      LAYER met1 ;
        RECT 91.97 2.36 92.26 2.59 ;
        RECT 91.97 0.88 92.26 1.11 ;
        RECT 92.03 0.88 92.2 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 16.18 1.66 16.35 2.935 ;
        RECT 16.18 5.945 16.35 7.22 ;
        RECT 11.42 5.945 11.59 7.22 ;
      LAYER met2 ;
        RECT 16.1 2.705 16.45 3.055 ;
        RECT 16.09 5.84 16.44 6.19 ;
        RECT 16.165 2.705 16.34 6.19 ;
      LAYER met1 ;
        RECT 16.1 2.765 16.58 2.935 ;
        RECT 16.1 2.705 16.45 3.055 ;
        RECT 11.36 5.945 16.58 6.115 ;
        RECT 16.09 5.84 16.44 6.19 ;
        RECT 11.36 5.915 11.65 6.145 ;
      LAYER mcon ;
        RECT 11.42 5.945 11.59 6.115 ;
        RECT 16.18 5.945 16.35 6.115 ;
        RECT 16.18 2.765 16.35 2.935 ;
      LAYER via1 ;
        RECT 16.19 5.94 16.34 6.09 ;
        RECT 16.2 2.805 16.35 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 34.105 1.66 34.275 2.935 ;
        RECT 34.105 5.945 34.275 7.22 ;
        RECT 29.345 5.945 29.515 7.22 ;
      LAYER met2 ;
        RECT 34.025 2.705 34.375 3.055 ;
        RECT 34.015 5.84 34.365 6.19 ;
        RECT 34.09 2.705 34.265 6.19 ;
      LAYER met1 ;
        RECT 34.025 2.765 34.505 2.935 ;
        RECT 34.025 2.705 34.375 3.055 ;
        RECT 29.285 5.945 34.505 6.115 ;
        RECT 34.015 5.84 34.365 6.19 ;
        RECT 29.285 5.915 29.575 6.145 ;
      LAYER mcon ;
        RECT 29.345 5.945 29.515 6.115 ;
        RECT 34.105 5.945 34.275 6.115 ;
        RECT 34.105 2.765 34.275 2.935 ;
      LAYER via1 ;
        RECT 34.115 5.94 34.265 6.09 ;
        RECT 34.125 2.805 34.275 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 52.03 1.66 52.2 2.935 ;
        RECT 52.03 5.945 52.2 7.22 ;
        RECT 47.27 5.945 47.44 7.22 ;
      LAYER met2 ;
        RECT 51.95 2.705 52.3 3.055 ;
        RECT 51.94 5.84 52.29 6.19 ;
        RECT 52.015 2.705 52.19 6.19 ;
      LAYER met1 ;
        RECT 51.95 2.765 52.43 2.935 ;
        RECT 51.95 2.705 52.3 3.055 ;
        RECT 47.21 5.945 52.43 6.115 ;
        RECT 51.94 5.84 52.29 6.19 ;
        RECT 47.21 5.915 47.5 6.145 ;
      LAYER mcon ;
        RECT 47.27 5.945 47.44 6.115 ;
        RECT 52.03 5.945 52.2 6.115 ;
        RECT 52.03 2.765 52.2 2.935 ;
      LAYER via1 ;
        RECT 52.04 5.94 52.19 6.09 ;
        RECT 52.05 2.805 52.2 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 69.955 1.66 70.125 2.935 ;
        RECT 69.955 5.945 70.125 7.22 ;
        RECT 65.195 5.945 65.365 7.22 ;
      LAYER met2 ;
        RECT 69.875 2.705 70.225 3.055 ;
        RECT 69.865 5.84 70.215 6.19 ;
        RECT 69.94 2.705 70.115 6.19 ;
      LAYER met1 ;
        RECT 69.875 2.765 70.355 2.935 ;
        RECT 69.875 2.705 70.225 3.055 ;
        RECT 65.135 5.945 70.355 6.115 ;
        RECT 69.865 5.84 70.215 6.19 ;
        RECT 65.135 5.915 65.425 6.145 ;
      LAYER mcon ;
        RECT 65.195 5.945 65.365 6.115 ;
        RECT 69.955 5.945 70.125 6.115 ;
        RECT 69.955 2.765 70.125 2.935 ;
      LAYER via1 ;
        RECT 69.965 5.94 70.115 6.09 ;
        RECT 69.975 2.805 70.125 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 87.88 1.66 88.05 2.935 ;
        RECT 87.88 5.945 88.05 7.22 ;
        RECT 83.12 5.945 83.29 7.22 ;
      LAYER met2 ;
        RECT 87.8 2.705 88.15 3.055 ;
        RECT 87.79 5.84 88.14 6.19 ;
        RECT 87.865 2.705 88.04 6.19 ;
      LAYER met1 ;
        RECT 87.8 2.765 88.28 2.935 ;
        RECT 87.8 2.705 88.15 3.055 ;
        RECT 83.06 5.945 88.28 6.115 ;
        RECT 87.79 5.84 88.14 6.19 ;
        RECT 83.06 5.915 83.35 6.145 ;
      LAYER mcon ;
        RECT 83.12 5.945 83.29 6.115 ;
        RECT 87.88 5.945 88.05 6.115 ;
        RECT 87.88 2.765 88.05 2.935 ;
      LAYER via1 ;
        RECT 87.89 5.94 88.04 6.09 ;
        RECT 87.9 2.805 88.05 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.39 5.945 0.56 7.22 ;
      LAYER met1 ;
        RECT 0.33 5.945 0.79 6.115 ;
        RECT 0.33 5.915 0.62 6.145 ;
      LAYER mcon ;
        RECT 0.39 5.945 0.56 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.385 4.33 2.19 4.71 ;
      LAYER li1 ;
        RECT 0 4.44 92.575 4.745 ;
        RECT 86.615 4.135 92.575 4.745 ;
        RECT 90.44 4.13 92.42 4.75 ;
        RECT 91.6 3.4 91.77 5.48 ;
        RECT 90.61 3.4 90.78 5.48 ;
        RECT 87.87 3.405 88.04 5.475 ;
        RECT 1.85 4.285 92.575 4.745 ;
        RECT 85.115 3.785 85.285 4.745 ;
        RECT 83.11 4.285 83.28 5.475 ;
        RECT 82.675 3.785 82.845 4.745 ;
        RECT 80.715 3.785 80.885 4.745 ;
        RECT 79.755 3.785 79.925 4.745 ;
        RECT 77.795 3.785 77.965 4.745 ;
        RECT 76.795 3.785 76.965 4.745 ;
        RECT 75.835 3.785 76.005 4.745 ;
        RECT 68.69 4.135 74.65 4.745 ;
        RECT 72.515 4.13 74.495 4.75 ;
        RECT 73.675 3.4 73.845 5.48 ;
        RECT 72.685 3.4 72.855 5.48 ;
        RECT 69.945 3.405 70.115 5.475 ;
        RECT 67.19 3.785 67.36 4.745 ;
        RECT 65.185 4.285 65.355 5.475 ;
        RECT 64.75 3.785 64.92 4.745 ;
        RECT 62.79 3.785 62.96 4.745 ;
        RECT 61.83 3.785 62 4.745 ;
        RECT 59.87 3.785 60.04 4.745 ;
        RECT 58.87 3.785 59.04 4.745 ;
        RECT 57.91 3.785 58.08 4.745 ;
        RECT 50.765 4.135 56.725 4.745 ;
        RECT 54.59 4.13 56.57 4.75 ;
        RECT 55.75 3.4 55.92 5.48 ;
        RECT 54.76 3.4 54.93 5.48 ;
        RECT 52.02 3.405 52.19 5.475 ;
        RECT 49.265 3.785 49.435 4.745 ;
        RECT 47.26 4.285 47.43 5.475 ;
        RECT 46.825 3.785 46.995 4.745 ;
        RECT 44.865 3.785 45.035 4.745 ;
        RECT 43.905 3.785 44.075 4.745 ;
        RECT 41.945 3.785 42.115 4.745 ;
        RECT 40.945 3.785 41.115 4.745 ;
        RECT 39.985 3.785 40.155 4.745 ;
        RECT 32.84 4.135 38.8 4.745 ;
        RECT 36.665 4.13 38.645 4.75 ;
        RECT 37.825 3.4 37.995 5.48 ;
        RECT 36.835 3.4 37.005 5.48 ;
        RECT 34.095 3.405 34.265 5.475 ;
        RECT 31.34 3.785 31.51 4.745 ;
        RECT 29.335 4.285 29.505 5.475 ;
        RECT 28.9 3.785 29.07 4.745 ;
        RECT 26.94 3.785 27.11 4.745 ;
        RECT 25.98 3.785 26.15 4.745 ;
        RECT 24.02 3.785 24.19 4.745 ;
        RECT 23.02 3.785 23.19 4.745 ;
        RECT 22.06 3.785 22.23 4.745 ;
        RECT 14.915 4.135 20.875 4.745 ;
        RECT 18.74 4.13 20.72 4.75 ;
        RECT 19.9 3.4 20.07 5.48 ;
        RECT 18.91 3.4 19.08 5.48 ;
        RECT 16.17 3.405 16.34 5.475 ;
        RECT 13.415 3.785 13.585 4.745 ;
        RECT 11.41 4.285 11.58 5.475 ;
        RECT 10.975 3.785 11.145 4.745 ;
        RECT 9.015 3.785 9.185 4.745 ;
        RECT 8.055 3.785 8.225 4.745 ;
        RECT 6.095 3.785 6.265 4.745 ;
        RECT 5.095 3.785 5.265 4.745 ;
        RECT 4.135 3.785 4.305 4.745 ;
        RECT 2.19 4.285 2.36 8.305 ;
        RECT 0 4.285 92.575 4.405 ;
        RECT 0 4.285 1.68 4.745 ;
        RECT 0.38 4.285 0.55 5.475 ;
      LAYER met2 ;
        RECT 1.575 4.33 1.955 4.71 ;
      LAYER met1 ;
        RECT 0 4.285 92.575 4.745 ;
        RECT 75.025 4.135 92.575 4.745 ;
        RECT 90.44 4.13 92.42 4.75 ;
        RECT 75.025 4.125 86.985 4.745 ;
        RECT 57.1 4.135 74.65 4.745 ;
        RECT 72.515 4.13 74.495 4.75 ;
        RECT 57.1 4.125 69.06 4.745 ;
        RECT 39.175 4.135 56.725 4.745 ;
        RECT 54.59 4.13 56.57 4.75 ;
        RECT 39.175 4.125 51.135 4.745 ;
        RECT 21.25 4.135 38.8 4.745 ;
        RECT 36.665 4.13 38.645 4.75 ;
        RECT 21.25 4.125 33.21 4.745 ;
        RECT 3.325 4.135 20.875 4.745 ;
        RECT 18.74 4.13 20.72 4.75 ;
        RECT 3.325 4.125 15.285 4.745 ;
        RECT 2.13 6.655 2.42 6.885 ;
        RECT 1.96 6.685 2.42 6.855 ;
      LAYER via2 ;
        RECT 1.665 4.42 1.865 4.62 ;
      LAYER mcon ;
        RECT 2.19 6.685 2.36 6.855 ;
        RECT 2.5 4.545 2.67 4.715 ;
        RECT 3.465 4.285 3.635 4.455 ;
        RECT 3.925 4.285 4.095 4.455 ;
        RECT 4.385 4.285 4.555 4.455 ;
        RECT 4.845 4.285 5.015 4.455 ;
        RECT 5.305 4.285 5.475 4.455 ;
        RECT 5.765 4.285 5.935 4.455 ;
        RECT 6.225 4.285 6.395 4.455 ;
        RECT 6.685 4.285 6.855 4.455 ;
        RECT 7.145 4.285 7.315 4.455 ;
        RECT 7.605 4.285 7.775 4.455 ;
        RECT 8.065 4.285 8.235 4.455 ;
        RECT 8.525 4.285 8.695 4.455 ;
        RECT 8.985 4.285 9.155 4.455 ;
        RECT 9.445 4.285 9.615 4.455 ;
        RECT 9.905 4.285 10.075 4.455 ;
        RECT 10.365 4.285 10.535 4.455 ;
        RECT 10.825 4.285 10.995 4.455 ;
        RECT 11.285 4.285 11.455 4.455 ;
        RECT 11.745 4.285 11.915 4.455 ;
        RECT 12.205 4.285 12.375 4.455 ;
        RECT 12.665 4.285 12.835 4.455 ;
        RECT 13.125 4.285 13.295 4.455 ;
        RECT 13.53 4.545 13.7 4.715 ;
        RECT 13.585 4.285 13.755 4.455 ;
        RECT 14.045 4.285 14.215 4.455 ;
        RECT 14.505 4.285 14.675 4.455 ;
        RECT 14.965 4.285 15.135 4.455 ;
        RECT 18.29 4.545 18.46 4.715 ;
        RECT 18.29 4.165 18.46 4.335 ;
        RECT 18.99 4.55 19.16 4.72 ;
        RECT 18.99 4.16 19.16 4.33 ;
        RECT 19.98 4.55 20.15 4.72 ;
        RECT 19.98 4.16 20.15 4.33 ;
        RECT 21.39 4.285 21.56 4.455 ;
        RECT 21.85 4.285 22.02 4.455 ;
        RECT 22.31 4.285 22.48 4.455 ;
        RECT 22.77 4.285 22.94 4.455 ;
        RECT 23.23 4.285 23.4 4.455 ;
        RECT 23.69 4.285 23.86 4.455 ;
        RECT 24.15 4.285 24.32 4.455 ;
        RECT 24.61 4.285 24.78 4.455 ;
        RECT 25.07 4.285 25.24 4.455 ;
        RECT 25.53 4.285 25.7 4.455 ;
        RECT 25.99 4.285 26.16 4.455 ;
        RECT 26.45 4.285 26.62 4.455 ;
        RECT 26.91 4.285 27.08 4.455 ;
        RECT 27.37 4.285 27.54 4.455 ;
        RECT 27.83 4.285 28 4.455 ;
        RECT 28.29 4.285 28.46 4.455 ;
        RECT 28.75 4.285 28.92 4.455 ;
        RECT 29.21 4.285 29.38 4.455 ;
        RECT 29.67 4.285 29.84 4.455 ;
        RECT 30.13 4.285 30.3 4.455 ;
        RECT 30.59 4.285 30.76 4.455 ;
        RECT 31.05 4.285 31.22 4.455 ;
        RECT 31.455 4.545 31.625 4.715 ;
        RECT 31.51 4.285 31.68 4.455 ;
        RECT 31.97 4.285 32.14 4.455 ;
        RECT 32.43 4.285 32.6 4.455 ;
        RECT 32.89 4.285 33.06 4.455 ;
        RECT 36.215 4.545 36.385 4.715 ;
        RECT 36.215 4.165 36.385 4.335 ;
        RECT 36.915 4.55 37.085 4.72 ;
        RECT 36.915 4.16 37.085 4.33 ;
        RECT 37.905 4.55 38.075 4.72 ;
        RECT 37.905 4.16 38.075 4.33 ;
        RECT 39.315 4.285 39.485 4.455 ;
        RECT 39.775 4.285 39.945 4.455 ;
        RECT 40.235 4.285 40.405 4.455 ;
        RECT 40.695 4.285 40.865 4.455 ;
        RECT 41.155 4.285 41.325 4.455 ;
        RECT 41.615 4.285 41.785 4.455 ;
        RECT 42.075 4.285 42.245 4.455 ;
        RECT 42.535 4.285 42.705 4.455 ;
        RECT 42.995 4.285 43.165 4.455 ;
        RECT 43.455 4.285 43.625 4.455 ;
        RECT 43.915 4.285 44.085 4.455 ;
        RECT 44.375 4.285 44.545 4.455 ;
        RECT 44.835 4.285 45.005 4.455 ;
        RECT 45.295 4.285 45.465 4.455 ;
        RECT 45.755 4.285 45.925 4.455 ;
        RECT 46.215 4.285 46.385 4.455 ;
        RECT 46.675 4.285 46.845 4.455 ;
        RECT 47.135 4.285 47.305 4.455 ;
        RECT 47.595 4.285 47.765 4.455 ;
        RECT 48.055 4.285 48.225 4.455 ;
        RECT 48.515 4.285 48.685 4.455 ;
        RECT 48.975 4.285 49.145 4.455 ;
        RECT 49.38 4.545 49.55 4.715 ;
        RECT 49.435 4.285 49.605 4.455 ;
        RECT 49.895 4.285 50.065 4.455 ;
        RECT 50.355 4.285 50.525 4.455 ;
        RECT 50.815 4.285 50.985 4.455 ;
        RECT 54.14 4.545 54.31 4.715 ;
        RECT 54.14 4.165 54.31 4.335 ;
        RECT 54.84 4.55 55.01 4.72 ;
        RECT 54.84 4.16 55.01 4.33 ;
        RECT 55.83 4.55 56 4.72 ;
        RECT 55.83 4.16 56 4.33 ;
        RECT 57.24 4.285 57.41 4.455 ;
        RECT 57.7 4.285 57.87 4.455 ;
        RECT 58.16 4.285 58.33 4.455 ;
        RECT 58.62 4.285 58.79 4.455 ;
        RECT 59.08 4.285 59.25 4.455 ;
        RECT 59.54 4.285 59.71 4.455 ;
        RECT 60 4.285 60.17 4.455 ;
        RECT 60.46 4.285 60.63 4.455 ;
        RECT 60.92 4.285 61.09 4.455 ;
        RECT 61.38 4.285 61.55 4.455 ;
        RECT 61.84 4.285 62.01 4.455 ;
        RECT 62.3 4.285 62.47 4.455 ;
        RECT 62.76 4.285 62.93 4.455 ;
        RECT 63.22 4.285 63.39 4.455 ;
        RECT 63.68 4.285 63.85 4.455 ;
        RECT 64.14 4.285 64.31 4.455 ;
        RECT 64.6 4.285 64.77 4.455 ;
        RECT 65.06 4.285 65.23 4.455 ;
        RECT 65.52 4.285 65.69 4.455 ;
        RECT 65.98 4.285 66.15 4.455 ;
        RECT 66.44 4.285 66.61 4.455 ;
        RECT 66.9 4.285 67.07 4.455 ;
        RECT 67.305 4.545 67.475 4.715 ;
        RECT 67.36 4.285 67.53 4.455 ;
        RECT 67.82 4.285 67.99 4.455 ;
        RECT 68.28 4.285 68.45 4.455 ;
        RECT 68.74 4.285 68.91 4.455 ;
        RECT 72.065 4.545 72.235 4.715 ;
        RECT 72.065 4.165 72.235 4.335 ;
        RECT 72.765 4.55 72.935 4.72 ;
        RECT 72.765 4.16 72.935 4.33 ;
        RECT 73.755 4.55 73.925 4.72 ;
        RECT 73.755 4.16 73.925 4.33 ;
        RECT 75.165 4.285 75.335 4.455 ;
        RECT 75.625 4.285 75.795 4.455 ;
        RECT 76.085 4.285 76.255 4.455 ;
        RECT 76.545 4.285 76.715 4.455 ;
        RECT 77.005 4.285 77.175 4.455 ;
        RECT 77.465 4.285 77.635 4.455 ;
        RECT 77.925 4.285 78.095 4.455 ;
        RECT 78.385 4.285 78.555 4.455 ;
        RECT 78.845 4.285 79.015 4.455 ;
        RECT 79.305 4.285 79.475 4.455 ;
        RECT 79.765 4.285 79.935 4.455 ;
        RECT 80.225 4.285 80.395 4.455 ;
        RECT 80.685 4.285 80.855 4.455 ;
        RECT 81.145 4.285 81.315 4.455 ;
        RECT 81.605 4.285 81.775 4.455 ;
        RECT 82.065 4.285 82.235 4.455 ;
        RECT 82.525 4.285 82.695 4.455 ;
        RECT 82.985 4.285 83.155 4.455 ;
        RECT 83.445 4.285 83.615 4.455 ;
        RECT 83.905 4.285 84.075 4.455 ;
        RECT 84.365 4.285 84.535 4.455 ;
        RECT 84.825 4.285 84.995 4.455 ;
        RECT 85.23 4.545 85.4 4.715 ;
        RECT 85.285 4.285 85.455 4.455 ;
        RECT 85.745 4.285 85.915 4.455 ;
        RECT 86.205 4.285 86.375 4.455 ;
        RECT 86.665 4.285 86.835 4.455 ;
        RECT 89.99 4.545 90.16 4.715 ;
        RECT 89.99 4.165 90.16 4.335 ;
        RECT 90.69 4.55 90.86 4.72 ;
        RECT 90.69 4.16 90.86 4.33 ;
        RECT 91.68 4.55 91.85 4.72 ;
        RECT 91.68 4.16 91.85 4.33 ;
      LAYER via1 ;
        RECT 1.69 4.445 1.84 4.595 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 84.415 4.925 84.725 7.425 ;
      RECT 84.415 4.925 87.51 5.235 ;
      RECT 87.2 1.125 87.51 5.235 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 84.325 3.685 84.885 4.015 ;
      RECT 84.325 2.015 84.625 4.015 ;
      RECT 80.395 3.125 80.945 3.455 ;
      RECT 80.645 2.015 80.945 3.455 ;
      RECT 81.445 1.885 81.595 2.535 ;
      RECT 80.645 2.015 84.625 2.315 ;
      RECT 79.165 0.96 79.465 3.91 ;
      RECT 79.155 2.565 79.885 2.895 ;
      RECT 79.12 0.96 79.495 1.33 ;
      RECT 77.715 3.125 78.445 3.455 ;
      RECT 77.73 0.96 78.03 3.455 ;
      RECT 75.605 2.565 76.335 2.895 ;
      RECT 75.76 0.93 76.06 2.895 ;
      RECT 77.685 0.96 78.06 1.33 ;
      RECT 75.715 0.93 76.09 1.3 ;
      RECT 75.715 0.97 78.06 1.27 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 66.49 4.925 66.8 7.425 ;
      RECT 66.49 4.925 69.585 5.235 ;
      RECT 69.275 1.125 69.585 5.235 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 66.4 3.685 66.96 4.015 ;
      RECT 66.4 2.015 66.7 4.015 ;
      RECT 62.47 3.125 63.02 3.455 ;
      RECT 62.72 2.015 63.02 3.455 ;
      RECT 63.52 1.885 63.67 2.535 ;
      RECT 62.72 2.015 66.7 2.315 ;
      RECT 61.24 0.96 61.54 3.91 ;
      RECT 61.23 2.565 61.96 2.895 ;
      RECT 61.195 0.96 61.57 1.33 ;
      RECT 59.79 3.125 60.52 3.455 ;
      RECT 59.805 0.96 60.105 3.455 ;
      RECT 57.68 2.565 58.41 2.895 ;
      RECT 57.835 0.93 58.135 2.895 ;
      RECT 59.76 0.96 60.135 1.33 ;
      RECT 57.79 0.93 58.165 1.3 ;
      RECT 57.79 0.97 60.135 1.27 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 48.565 4.925 48.875 7.425 ;
      RECT 48.565 4.925 51.66 5.235 ;
      RECT 51.35 1.125 51.66 5.235 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 48.475 3.685 49.035 4.015 ;
      RECT 48.475 2.015 48.775 4.015 ;
      RECT 44.545 3.125 45.095 3.455 ;
      RECT 44.795 2.015 45.095 3.455 ;
      RECT 45.595 1.885 45.745 2.535 ;
      RECT 44.795 2.015 48.775 2.315 ;
      RECT 43.315 0.96 43.615 3.91 ;
      RECT 43.305 2.565 44.035 2.895 ;
      RECT 43.27 0.96 43.645 1.33 ;
      RECT 41.865 3.125 42.595 3.455 ;
      RECT 41.88 0.96 42.18 3.455 ;
      RECT 39.755 2.565 40.485 2.895 ;
      RECT 39.91 0.93 40.21 2.895 ;
      RECT 41.835 0.96 42.21 1.33 ;
      RECT 39.865 0.93 40.24 1.3 ;
      RECT 39.865 0.97 42.21 1.27 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 30.64 4.925 30.95 7.425 ;
      RECT 30.64 4.925 33.735 5.235 ;
      RECT 33.425 1.125 33.735 5.235 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 30.55 3.685 31.11 4.015 ;
      RECT 30.55 2.015 30.85 4.015 ;
      RECT 26.62 3.125 27.17 3.455 ;
      RECT 26.87 2.015 27.17 3.455 ;
      RECT 27.67 1.885 27.82 2.535 ;
      RECT 26.87 2.015 30.85 2.315 ;
      RECT 25.39 0.96 25.69 3.91 ;
      RECT 25.38 2.565 26.11 2.895 ;
      RECT 25.345 0.96 25.72 1.33 ;
      RECT 23.94 3.125 24.67 3.455 ;
      RECT 23.955 0.96 24.255 3.455 ;
      RECT 21.83 2.565 22.56 2.895 ;
      RECT 21.985 0.93 22.285 2.895 ;
      RECT 23.91 0.96 24.285 1.33 ;
      RECT 21.94 0.93 22.315 1.3 ;
      RECT 21.94 0.97 24.285 1.27 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 12.715 4.925 13.025 7.425 ;
      RECT 12.715 4.925 15.81 5.235 ;
      RECT 15.5 1.125 15.81 5.235 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 12.625 3.685 13.185 4.015 ;
      RECT 12.625 2.015 12.925 4.015 ;
      RECT 8.695 3.125 9.245 3.455 ;
      RECT 8.945 2.015 9.245 3.455 ;
      RECT 9.745 1.885 9.895 2.535 ;
      RECT 8.945 2.015 12.925 2.315 ;
      RECT 7.465 0.96 7.765 3.91 ;
      RECT 7.455 2.565 8.185 2.895 ;
      RECT 7.42 0.96 7.795 1.33 ;
      RECT 6.015 3.125 6.745 3.455 ;
      RECT 6.03 0.96 6.33 3.455 ;
      RECT 3.905 2.565 4.635 2.895 ;
      RECT 4.06 0.93 4.36 2.895 ;
      RECT 5.985 0.96 6.36 1.33 ;
      RECT 4.015 0.93 4.39 1.3 ;
      RECT 4.015 0.97 6.36 1.27 ;
      RECT 85.515 2.005 86.245 2.335 ;
      RECT 83.295 3.685 84.025 4.015 ;
      RECT 81.595 3.685 82.325 4.015 ;
      RECT 76.635 2.565 77.365 2.895 ;
      RECT 75.275 3.685 76.005 4.015 ;
      RECT 67.59 2.005 68.32 2.335 ;
      RECT 65.37 3.685 66.1 4.015 ;
      RECT 63.67 3.685 64.4 4.015 ;
      RECT 58.71 2.565 59.44 2.895 ;
      RECT 57.35 3.685 58.08 4.015 ;
      RECT 49.665 2.005 50.395 2.335 ;
      RECT 47.445 3.685 48.175 4.015 ;
      RECT 45.745 3.685 46.475 4.015 ;
      RECT 40.785 2.565 41.515 2.895 ;
      RECT 39.425 3.685 40.155 4.015 ;
      RECT 31.74 2.005 32.47 2.335 ;
      RECT 29.52 3.685 30.25 4.015 ;
      RECT 27.82 3.685 28.55 4.015 ;
      RECT 22.86 2.565 23.59 2.895 ;
      RECT 21.5 3.685 22.23 4.015 ;
      RECT 13.815 2.005 14.545 2.335 ;
      RECT 11.595 3.685 12.325 4.015 ;
      RECT 9.895 3.685 10.625 4.015 ;
      RECT 4.935 2.565 5.665 2.895 ;
      RECT 3.575 3.685 4.305 4.015 ;
      RECT 0.025 8.5 0.83 8.88 ;
    LAYER via2 ;
      RECT 77.04 2.63 77.24 2.83 ;
      RECT 77.035 2.625 77.235 2.825 ;
      RECT 59.115 2.63 59.315 2.83 ;
      RECT 59.11 2.625 59.31 2.825 ;
      RECT 41.19 2.63 41.39 2.83 ;
      RECT 41.185 2.625 41.385 2.825 ;
      RECT 23.265 2.63 23.465 2.83 ;
      RECT 23.26 2.625 23.46 2.825 ;
      RECT 5.34 2.63 5.54 2.83 ;
      RECT 5.335 2.625 5.535 2.825 ;
      RECT 87.29 1.225 87.49 1.425 ;
      RECT 85.575 2.065 85.775 2.265 ;
      RECT 84.615 3.745 84.815 3.945 ;
      RECT 84.47 7.14 84.67 7.34 ;
      RECT 83.615 3.745 83.815 3.945 ;
      RECT 81.655 3.745 81.855 3.945 ;
      RECT 80.455 3.185 80.655 3.385 ;
      RECT 79.215 2.625 79.415 2.825 ;
      RECT 79.21 1.045 79.41 1.245 ;
      RECT 77.775 1.04 77.975 1.24 ;
      RECT 77.775 3.185 77.975 3.385 ;
      RECT 75.815 2.625 76.015 2.825 ;
      RECT 75.805 1.015 76.005 1.215 ;
      RECT 75.335 3.745 75.535 3.945 ;
      RECT 69.365 1.225 69.565 1.425 ;
      RECT 67.65 2.065 67.85 2.265 ;
      RECT 66.69 3.745 66.89 3.945 ;
      RECT 66.545 7.14 66.745 7.34 ;
      RECT 65.69 3.745 65.89 3.945 ;
      RECT 63.73 3.745 63.93 3.945 ;
      RECT 62.53 3.185 62.73 3.385 ;
      RECT 61.29 2.625 61.49 2.825 ;
      RECT 61.285 1.045 61.485 1.245 ;
      RECT 59.85 1.04 60.05 1.24 ;
      RECT 59.85 3.185 60.05 3.385 ;
      RECT 57.89 2.625 58.09 2.825 ;
      RECT 57.88 1.015 58.08 1.215 ;
      RECT 57.41 3.745 57.61 3.945 ;
      RECT 51.44 1.225 51.64 1.425 ;
      RECT 49.725 2.065 49.925 2.265 ;
      RECT 48.765 3.745 48.965 3.945 ;
      RECT 48.62 7.14 48.82 7.34 ;
      RECT 47.765 3.745 47.965 3.945 ;
      RECT 45.805 3.745 46.005 3.945 ;
      RECT 44.605 3.185 44.805 3.385 ;
      RECT 43.365 2.625 43.565 2.825 ;
      RECT 43.36 1.045 43.56 1.245 ;
      RECT 41.925 1.04 42.125 1.24 ;
      RECT 41.925 3.185 42.125 3.385 ;
      RECT 39.965 2.625 40.165 2.825 ;
      RECT 39.955 1.015 40.155 1.215 ;
      RECT 39.485 3.745 39.685 3.945 ;
      RECT 33.515 1.225 33.715 1.425 ;
      RECT 31.8 2.065 32 2.265 ;
      RECT 30.84 3.745 31.04 3.945 ;
      RECT 30.695 7.14 30.895 7.34 ;
      RECT 29.84 3.745 30.04 3.945 ;
      RECT 27.88 3.745 28.08 3.945 ;
      RECT 26.68 3.185 26.88 3.385 ;
      RECT 25.44 2.625 25.64 2.825 ;
      RECT 25.435 1.045 25.635 1.245 ;
      RECT 24 1.04 24.2 1.24 ;
      RECT 24 3.185 24.2 3.385 ;
      RECT 22.04 2.625 22.24 2.825 ;
      RECT 22.03 1.015 22.23 1.215 ;
      RECT 21.56 3.745 21.76 3.945 ;
      RECT 15.59 1.225 15.79 1.425 ;
      RECT 13.875 2.065 14.075 2.265 ;
      RECT 12.915 3.745 13.115 3.945 ;
      RECT 12.77 7.14 12.97 7.34 ;
      RECT 11.915 3.745 12.115 3.945 ;
      RECT 9.955 3.745 10.155 3.945 ;
      RECT 8.755 3.185 8.955 3.385 ;
      RECT 7.515 2.625 7.715 2.825 ;
      RECT 7.51 1.045 7.71 1.245 ;
      RECT 6.075 1.04 6.275 1.24 ;
      RECT 6.075 3.185 6.275 3.385 ;
      RECT 4.115 2.625 4.315 2.825 ;
      RECT 4.105 1.015 4.305 1.215 ;
      RECT 3.635 3.745 3.835 3.945 ;
      RECT 0.305 8.59 0.505 8.79 ;
    LAYER met2 ;
      RECT 1.385 8.4 92.2 8.57 ;
      RECT 92.03 7.275 92.2 8.57 ;
      RECT 1.385 6.255 1.555 8.57 ;
      RECT 92 7.275 92.35 7.625 ;
      RECT 1.325 6.255 1.615 6.605 ;
      RECT 88.845 6.225 89.165 6.545 ;
      RECT 88.875 5.695 89.045 6.545 ;
      RECT 88.875 5.695 89.05 6.045 ;
      RECT 88.875 5.695 89.85 5.87 ;
      RECT 89.675 1.965 89.85 5.87 ;
      RECT 89.62 1.965 89.97 2.315 ;
      RECT 89.645 6.655 89.97 6.98 ;
      RECT 88.53 6.745 89.97 6.915 ;
      RECT 88.53 2.395 88.69 6.915 ;
      RECT 88.845 2.365 89.165 2.685 ;
      RECT 88.53 2.395 89.165 2.565 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 79.12 0.96 79.495 1.33 ;
      RECT 77.685 0.96 78.06 1.33 ;
      RECT 77.685 1.08 87.505 1.25 ;
      RECT 81.805 4.36 87.485 4.53 ;
      RECT 87.315 3.425 87.485 4.53 ;
      RECT 81.615 3.595 81.635 4.53 ;
      RECT 81.865 3.705 81.895 3.985 ;
      RECT 81.575 3.595 81.635 3.855 ;
      RECT 87.225 3.43 87.575 3.78 ;
      RECT 81.405 2.225 81.435 2.485 ;
      RECT 81.175 2.225 81.235 2.485 ;
      RECT 81.855 3.685 81.865 3.985 ;
      RECT 81.835 3.605 81.855 3.985 ;
      RECT 81.825 3.545 81.835 3.985 ;
      RECT 81.805 3.495 81.825 3.985 ;
      RECT 81.775 3.395 81.805 4.53 ;
      RECT 81.765 3.305 81.775 4.53 ;
      RECT 81.725 3.245 81.765 4.53 ;
      RECT 81.721 3.214 81.725 4.53 ;
      RECT 81.635 3.205 81.721 4.53 ;
      RECT 81.625 3.196 81.635 3.55 ;
      RECT 81.595 3.175 81.625 3.517 ;
      RECT 81.585 3.125 81.595 3.493 ;
      RECT 81.575 3.09 81.585 3.481 ;
      RECT 81.535 3.015 81.575 3.45 ;
      RECT 81.515 2.925 81.535 3.415 ;
      RECT 81.505 2.866 81.515 3.4 ;
      RECT 81.455 2.756 81.505 3.36 ;
      RECT 81.445 2.65 81.455 3.315 ;
      RECT 81.415 2.579 81.445 3.235 ;
      RECT 81.405 2.511 81.415 3.16 ;
      RECT 81.395 2.225 81.405 3.125 ;
      RECT 81.365 2.225 81.395 3.055 ;
      RECT 81.355 2.225 81.365 2.95 ;
      RECT 81.345 2.225 81.355 2.915 ;
      RECT 81.275 2.225 81.345 2.775 ;
      RECT 81.245 2.225 81.275 2.575 ;
      RECT 81.235 2.225 81.245 2.5 ;
      RECT 85.575 2.155 85.835 2.415 ;
      RECT 85.565 2.155 85.835 2.365 ;
      RECT 85.535 2.025 85.815 2.305 ;
      RECT 74.055 6.655 74.405 7.005 ;
      RECT 85.3 6.61 85.65 6.96 ;
      RECT 74.055 6.685 85.65 6.885 ;
      RECT 84.575 3.705 84.855 3.985 ;
      RECT 84.615 3.665 84.885 3.925 ;
      RECT 84.605 3.7 84.885 3.925 ;
      RECT 84.615 3.66 84.825 3.985 ;
      RECT 84.615 3.655 84.815 3.985 ;
      RECT 84.655 3.645 84.815 3.985 ;
      RECT 84.625 3.65 84.815 3.985 ;
      RECT 84.665 3.64 84.755 3.985 ;
      RECT 84.685 3.635 84.755 3.985 ;
      RECT 83.995 3.155 84.255 3.415 ;
      RECT 84.045 3.065 84.235 3.415 ;
      RECT 84.075 2.85 84.235 3.415 ;
      RECT 84.165 2.455 84.235 3.415 ;
      RECT 84.185 2.165 84.321 2.893 ;
      RECT 84.125 2.66 84.321 2.893 ;
      RECT 84.145 2.54 84.235 3.415 ;
      RECT 84.185 2.165 84.345 2.558 ;
      RECT 84.185 2.165 84.355 2.455 ;
      RECT 84.175 2.165 84.435 2.425 ;
      RECT 83.575 3.705 83.855 3.985 ;
      RECT 83.595 3.665 83.855 3.985 ;
      RECT 83.235 3.625 83.345 3.885 ;
      RECT 83.095 2.115 83.185 2.375 ;
      RECT 83.625 3.17 83.635 3.3 ;
      RECT 83.615 3.135 83.625 3.454 ;
      RECT 83.535 3.067 83.615 3.534 ;
      RECT 83.565 3.71 83.575 3.93 ;
      RECT 83.545 3.705 83.565 3.919 ;
      RECT 83.515 3.7 83.545 3.904 ;
      RECT 83.525 3.002 83.535 3.61 ;
      RECT 83.505 2.946 83.525 3.625 ;
      RECT 83.495 3.685 83.515 3.89 ;
      RECT 83.495 2.874 83.505 3.645 ;
      RECT 83.465 2.777 83.495 3.885 ;
      RECT 83.445 2.66 83.465 3.885 ;
      RECT 83.415 2.54 83.445 3.885 ;
      RECT 83.405 2.455 83.415 3.885 ;
      RECT 83.395 2.4 83.405 3.885 ;
      RECT 83.385 2.355 83.395 3.104 ;
      RECT 83.375 3.315 83.395 3.885 ;
      RECT 83.375 2.285 83.385 3.061 ;
      RECT 83.355 2.235 83.375 2.996 ;
      RECT 83.365 3.395 83.375 3.885 ;
      RECT 83.345 3.495 83.365 3.885 ;
      RECT 83.295 2.115 83.355 2.824 ;
      RECT 83.285 2.115 83.295 2.66 ;
      RECT 83.275 2.115 83.285 2.61 ;
      RECT 83.225 2.115 83.275 2.54 ;
      RECT 83.205 2.115 83.225 2.455 ;
      RECT 83.185 2.115 83.205 2.41 ;
      RECT 82.505 3.565 82.555 3.825 ;
      RECT 82.415 2.095 82.555 2.355 ;
      RECT 82.915 2.72 82.925 2.808 ;
      RECT 82.905 2.655 82.915 2.854 ;
      RECT 82.895 2.605 82.905 2.9 ;
      RECT 82.845 2.552 82.895 3.039 ;
      RECT 82.835 2.501 82.845 3.23 ;
      RECT 82.795 2.459 82.835 3.335 ;
      RECT 82.775 2.405 82.795 3.472 ;
      RECT 82.765 2.38 82.775 2.688 ;
      RECT 82.765 2.77 82.775 3.542 ;
      RECT 82.755 2.366 82.765 2.673 ;
      RECT 82.755 2.825 82.765 3.825 ;
      RECT 82.735 2.341 82.755 2.655 ;
      RECT 82.715 3 82.755 3.825 ;
      RECT 82.725 2.315 82.735 2.635 ;
      RECT 82.695 2.28 82.725 2.589 ;
      RECT 82.705 3.125 82.715 3.825 ;
      RECT 82.695 3.205 82.705 3.825 ;
      RECT 82.685 2.245 82.695 2.554 ;
      RECT 82.645 3.275 82.695 3.825 ;
      RECT 82.675 2.225 82.685 2.53 ;
      RECT 82.645 2.095 82.675 2.495 ;
      RECT 82.635 2.095 82.645 2.46 ;
      RECT 82.615 3.375 82.645 3.825 ;
      RECT 82.615 2.095 82.635 2.435 ;
      RECT 82.605 2.095 82.615 2.41 ;
      RECT 82.565 3.475 82.615 3.825 ;
      RECT 82.585 2.095 82.605 2.38 ;
      RECT 82.555 2.095 82.585 2.365 ;
      RECT 82.555 3.55 82.565 3.825 ;
      RECT 82.475 2.635 82.515 2.895 ;
      RECT 78.205 2.055 78.465 2.315 ;
      RECT 78.205 2.085 78.485 2.295 ;
      RECT 80.415 1.905 80.595 2.055 ;
      RECT 82.465 2.63 82.475 2.895 ;
      RECT 82.445 2.62 82.465 2.895 ;
      RECT 82.427 2.613 82.445 2.895 ;
      RECT 82.341 2.602 82.427 2.895 ;
      RECT 82.255 2.585 82.341 2.895 ;
      RECT 82.205 2.572 82.255 2.82 ;
      RECT 82.171 2.564 82.205 2.795 ;
      RECT 82.085 2.553 82.171 2.76 ;
      RECT 82.045 2.53 82.085 2.723 ;
      RECT 82.035 2.495 82.045 2.708 ;
      RECT 82.025 2.455 82.035 2.703 ;
      RECT 82.015 2.435 82.025 2.698 ;
      RECT 82 2.395 82.015 2.693 ;
      RECT 81.985 2.347 82 2.689 ;
      RECT 81.975 2.306 81.985 2.686 ;
      RECT 81.965 2.268 81.975 2.675 ;
      RECT 81.945 2.212 81.965 2.655 ;
      RECT 81.925 2.16 81.945 2.591 ;
      RECT 81.905 2.11 81.925 2.543 ;
      RECT 81.895 2.08 81.905 2.507 ;
      RECT 81.89 2.062 81.895 2.493 ;
      RECT 81.875 2.053 81.89 2.475 ;
      RECT 81.845 2.034 81.875 2.415 ;
      RECT 81.835 2.017 81.845 2.37 ;
      RECT 81.825 2.009 81.835 2.34 ;
      RECT 81.795 1.997 81.825 2.29 ;
      RECT 81.775 1.985 81.795 2.225 ;
      RECT 81.765 1.977 81.775 2.185 ;
      RECT 81.745 1.974 81.765 2.175 ;
      RECT 81.73 1.972 81.745 2.17 ;
      RECT 81.71 1.971 81.73 2.16 ;
      RECT 81.695 1.97 81.71 2.15 ;
      RECT 81.675 1.969 81.695 2.145 ;
      RECT 81.673 1.969 81.675 2.145 ;
      RECT 81.587 1.966 81.673 2.142 ;
      RECT 81.501 1.961 81.587 2.135 ;
      RECT 81.415 1.956 81.501 2.129 ;
      RECT 81.365 1.953 81.415 2.12 ;
      RECT 81.321 1.951 81.365 2.114 ;
      RECT 81.235 1.947 81.321 2.109 ;
      RECT 81.231 1.945 81.235 2.105 ;
      RECT 81.145 1.942 81.231 2.1 ;
      RECT 81.091 1.938 81.145 2.093 ;
      RECT 81.005 1.935 81.091 2.088 ;
      RECT 80.981 1.932 81.005 2.084 ;
      RECT 80.895 1.93 80.981 2.079 ;
      RECT 80.835 1.926 80.895 2.073 ;
      RECT 80.827 1.924 80.835 2.07 ;
      RECT 80.741 1.92 80.827 2.066 ;
      RECT 80.655 1.913 80.741 2.059 ;
      RECT 80.595 1.907 80.655 2.055 ;
      RECT 80.395 1.905 80.415 2.058 ;
      RECT 80.345 1.915 80.395 2.068 ;
      RECT 80.315 1.925 80.345 2.08 ;
      RECT 80.291 1.927 80.315 2.086 ;
      RECT 80.205 1.93 80.291 2.091 ;
      RECT 80.135 1.935 80.205 2.1 ;
      RECT 80.121 1.937 80.135 2.106 ;
      RECT 80.035 1.941 80.121 2.111 ;
      RECT 79.995 1.945 80.035 2.12 ;
      RECT 79.981 1.947 79.995 2.126 ;
      RECT 79.895 1.951 79.981 2.131 ;
      RECT 79.811 1.957 79.895 2.138 ;
      RECT 79.725 1.963 79.811 2.143 ;
      RECT 79.701 1.967 79.725 2.146 ;
      RECT 79.615 1.971 79.701 2.151 ;
      RECT 79.565 1.976 79.615 2.16 ;
      RECT 79.485 1.981 79.565 2.17 ;
      RECT 79.405 1.987 79.485 2.185 ;
      RECT 79.385 1.991 79.405 2.195 ;
      RECT 79.315 1.994 79.385 2.205 ;
      RECT 79.265 1.999 79.315 2.22 ;
      RECT 79.235 2.002 79.265 2.24 ;
      RECT 79.225 2.004 79.235 2.256 ;
      RECT 79.165 2.016 79.225 2.266 ;
      RECT 79.145 2.031 79.165 2.275 ;
      RECT 79.135 2.05 79.145 2.275 ;
      RECT 79.125 2.07 79.135 2.275 ;
      RECT 79.105 2.08 79.125 2.275 ;
      RECT 79.055 2.09 79.105 2.275 ;
      RECT 79.025 2.096 79.055 2.275 ;
      RECT 78.955 2.101 79.025 2.277 ;
      RECT 78.875 2.102 78.955 2.282 ;
      RECT 78.871 2.1 78.875 2.285 ;
      RECT 78.785 2.097 78.871 2.286 ;
      RECT 78.743 2.094 78.785 2.288 ;
      RECT 78.657 2.092 78.743 2.289 ;
      RECT 78.571 2.089 78.657 2.292 ;
      RECT 78.485 2.086 78.571 2.294 ;
      RECT 80.415 3.145 80.695 3.425 ;
      RECT 80.445 3.125 80.715 3.385 ;
      RECT 80.445 3.075 80.675 3.425 ;
      RECT 80.515 3.065 80.675 3.425 ;
      RECT 80.515 2.775 80.665 3.425 ;
      RECT 80.505 2.455 80.655 2.825 ;
      RECT 80.495 2.455 80.655 2.695 ;
      RECT 80.475 2.165 80.645 2.5 ;
      RECT 80.455 2.165 80.645 2.45 ;
      RECT 80.415 2.165 80.675 2.425 ;
      RECT 80.325 3.635 80.405 3.895 ;
      RECT 79.615 2.355 79.735 2.615 ;
      RECT 80.3 3.615 80.325 3.895 ;
      RECT 80.285 3.577 80.3 3.895 ;
      RECT 80.245 3.52 80.285 3.895 ;
      RECT 80.215 3.43 80.245 3.895 ;
      RECT 80.175 3.33 80.215 3.895 ;
      RECT 80.145 3.23 80.175 3.895 ;
      RECT 80.14 3.177 80.145 3.718 ;
      RECT 80.125 3.147 80.14 3.684 ;
      RECT 80.115 3.108 80.125 3.649 ;
      RECT 80.105 3.075 80.115 3.605 ;
      RECT 80.095 3.042 80.105 3.57 ;
      RECT 80.065 2.976 80.095 3.505 ;
      RECT 80.055 2.911 80.065 3.43 ;
      RECT 80.045 2.881 80.055 3.4 ;
      RECT 80.005 2.811 80.045 3.33 ;
      RECT 79.995 2.746 80.005 3.245 ;
      RECT 79.985 2.728 79.995 3.23 ;
      RECT 79.975 2.711 79.985 3.195 ;
      RECT 79.965 2.694 79.975 3.165 ;
      RECT 79.955 2.677 79.965 3.135 ;
      RECT 79.935 2.652 79.955 3.075 ;
      RECT 79.925 2.626 79.935 3.02 ;
      RECT 79.905 2.601 79.925 2.98 ;
      RECT 79.895 2.57 79.905 2.945 ;
      RECT 79.885 2.557 79.895 2.9 ;
      RECT 79.875 2.542 79.885 2.875 ;
      RECT 79.865 2.355 79.875 2.835 ;
      RECT 79.855 2.355 79.865 2.805 ;
      RECT 79.85 2.355 79.855 2.788 ;
      RECT 79.845 2.355 79.85 2.77 ;
      RECT 79.775 2.355 79.845 2.71 ;
      RECT 79.735 2.355 79.775 2.645 ;
      RECT 79.565 3.225 79.825 3.485 ;
      RECT 77.735 3.145 77.815 3.465 ;
      RECT 77.555 3.205 77.705 3.465 ;
      RECT 77.735 3.145 77.845 3.425 ;
      RECT 79.555 3.317 79.565 3.48 ;
      RECT 79.525 3.327 79.555 3.488 ;
      RECT 79.505 3.335 79.525 3.493 ;
      RECT 79.437 3.343 79.505 3.503 ;
      RECT 79.351 3.363 79.437 3.52 ;
      RECT 79.265 3.384 79.351 3.539 ;
      RECT 79.255 3.4 79.265 3.55 ;
      RECT 79.215 3.41 79.255 3.556 ;
      RECT 79.195 3.415 79.215 3.563 ;
      RECT 79.157 3.416 79.195 3.566 ;
      RECT 79.071 3.419 79.157 3.567 ;
      RECT 78.985 3.423 79.071 3.568 ;
      RECT 78.931 3.425 78.985 3.57 ;
      RECT 78.845 3.425 78.931 3.572 ;
      RECT 78.805 3.42 78.845 3.574 ;
      RECT 78.795 3.414 78.805 3.575 ;
      RECT 78.755 3.409 78.795 3.571 ;
      RECT 78.745 3.4 78.755 3.567 ;
      RECT 78.713 3.391 78.745 3.564 ;
      RECT 78.627 3.379 78.713 3.554 ;
      RECT 78.541 3.362 78.627 3.539 ;
      RECT 78.455 3.344 78.541 3.525 ;
      RECT 78.435 3.335 78.455 3.516 ;
      RECT 78.365 3.325 78.435 3.509 ;
      RECT 78.315 3.31 78.365 3.499 ;
      RECT 78.255 3.3 78.315 3.49 ;
      RECT 78.215 3.29 78.255 3.485 ;
      RECT 78.165 3.28 78.215 3.479 ;
      RECT 78.125 3.268 78.165 3.469 ;
      RECT 78.105 3.258 78.125 3.465 ;
      RECT 78.085 3.248 78.105 3.465 ;
      RECT 78.075 3.238 78.085 3.464 ;
      RECT 78.055 3.23 78.075 3.46 ;
      RECT 78.015 3.205 78.055 3.454 ;
      RECT 77.995 3.145 78.015 3.447 ;
      RECT 77.971 3.145 77.995 3.444 ;
      RECT 77.885 3.145 77.971 3.439 ;
      RECT 77.845 3.145 77.885 3.43 ;
      RECT 77.705 3.195 77.735 3.465 ;
      RECT 79.385 2.775 79.645 3.035 ;
      RECT 79.345 2.775 79.645 2.915 ;
      RECT 79.315 2.775 79.645 2.9 ;
      RECT 79.255 2.775 79.645 2.88 ;
      RECT 79.175 2.585 79.455 2.865 ;
      RECT 79.175 2.77 79.525 2.865 ;
      RECT 79.175 2.71 79.515 2.865 ;
      RECT 79.175 2.66 79.465 2.865 ;
      RECT 76.945 3.115 77.205 3.375 ;
      RECT 77.09 1.205 77.205 3.375 ;
      RECT 77.005 2.585 77.205 3.375 ;
      RECT 78.315 2.635 78.575 2.895 ;
      RECT 77 2.585 77.205 2.87 ;
      RECT 76.995 2.585 77.205 2.865 ;
      RECT 78.295 2.645 78.575 2.825 ;
      RECT 77.885 2.615 78.025 2.765 ;
      RECT 77.26 1.205 77.34 1.55 ;
      RECT 76.995 1.205 77.205 1.55 ;
      RECT 78.285 2.644 78.295 2.825 ;
      RECT 78.281 2.644 78.285 2.825 ;
      RECT 78.195 2.639 78.281 2.814 ;
      RECT 78.121 2.63 78.195 2.794 ;
      RECT 78.035 2.621 78.121 2.775 ;
      RECT 78.025 2.615 78.035 2.765 ;
      RECT 77.845 2.615 77.885 2.768 ;
      RECT 77.759 2.615 77.845 2.776 ;
      RECT 77.673 2.615 77.759 2.787 ;
      RECT 77.587 2.615 77.673 2.798 ;
      RECT 77.501 2.615 77.587 2.809 ;
      RECT 77.415 2.615 77.501 2.82 ;
      RECT 77.385 2.615 77.415 2.86 ;
      RECT 77.355 2.615 77.385 2.91 ;
      RECT 77.28 2.615 77.355 2.93 ;
      RECT 77.275 2.59 77.28 2.935 ;
      RECT 77.26 2.585 77.275 2.943 ;
      RECT 77.255 1.205 77.26 2.953 ;
      RECT 77.225 1.205 77.255 2.995 ;
      RECT 77.205 1.205 77.225 3.075 ;
      RECT 76.335 2.965 76.355 3.404 ;
      RECT 76.335 2.965 76.441 3.401 ;
      RECT 76.325 3.08 76.441 3.4 ;
      RECT 76.355 2.115 76.485 3.397 ;
      RECT 76.335 2.985 76.495 3.395 ;
      RECT 76.335 3.07 76.505 3.39 ;
      RECT 76.305 3.115 76.505 3.385 ;
      RECT 76.305 3.115 76.515 3.38 ;
      RECT 76.285 3.115 76.545 3.375 ;
      RECT 76.355 2.115 76.515 2.765 ;
      RECT 76.345 2.115 76.515 2.74 ;
      RECT 76.345 2.115 76.535 2.505 ;
      RECT 76.295 2.115 76.555 2.375 ;
      RECT 75.765 2.605 76.055 2.865 ;
      RECT 75.775 2.585 76.055 2.865 ;
      RECT 75.725 2.665 76.055 2.86 ;
      RECT 75.795 2.578 75.965 2.865 ;
      RECT 75.795 2.565 75.921 2.865 ;
      RECT 75.835 2.558 75.921 2.865 ;
      RECT 75.295 3.705 75.575 3.985 ;
      RECT 75.255 3.67 75.555 3.78 ;
      RECT 75.245 3.62 75.535 3.675 ;
      RECT 75.185 3.385 75.445 3.645 ;
      RECT 75.185 3.525 75.525 3.645 ;
      RECT 75.185 3.475 75.505 3.645 ;
      RECT 75.185 3.43 75.495 3.645 ;
      RECT 75.185 3.415 75.465 3.645 ;
      RECT 70.92 6.225 71.24 6.545 ;
      RECT 70.95 5.695 71.12 6.545 ;
      RECT 70.95 5.695 71.125 6.045 ;
      RECT 70.95 5.695 71.925 5.87 ;
      RECT 71.75 1.965 71.925 5.87 ;
      RECT 71.695 1.965 72.045 2.315 ;
      RECT 71.72 6.655 72.045 6.98 ;
      RECT 70.605 6.745 72.045 6.915 ;
      RECT 70.605 2.395 70.765 6.915 ;
      RECT 70.92 2.365 71.24 2.685 ;
      RECT 70.605 2.395 71.24 2.565 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 61.195 0.96 61.57 1.33 ;
      RECT 59.76 0.96 60.135 1.33 ;
      RECT 59.76 1.08 69.58 1.25 ;
      RECT 63.88 4.36 69.56 4.53 ;
      RECT 69.39 3.425 69.56 4.53 ;
      RECT 63.69 3.595 63.71 4.53 ;
      RECT 63.94 3.705 63.97 3.985 ;
      RECT 63.65 3.595 63.71 3.855 ;
      RECT 69.3 3.43 69.65 3.78 ;
      RECT 63.48 2.225 63.51 2.485 ;
      RECT 63.25 2.225 63.31 2.485 ;
      RECT 63.93 3.685 63.94 3.985 ;
      RECT 63.91 3.605 63.93 3.985 ;
      RECT 63.9 3.545 63.91 3.985 ;
      RECT 63.88 3.495 63.9 3.985 ;
      RECT 63.85 3.395 63.88 4.53 ;
      RECT 63.84 3.305 63.85 4.53 ;
      RECT 63.8 3.245 63.84 4.53 ;
      RECT 63.796 3.214 63.8 4.53 ;
      RECT 63.71 3.205 63.796 4.53 ;
      RECT 63.7 3.196 63.71 3.55 ;
      RECT 63.67 3.175 63.7 3.517 ;
      RECT 63.66 3.125 63.67 3.493 ;
      RECT 63.65 3.09 63.66 3.481 ;
      RECT 63.61 3.015 63.65 3.45 ;
      RECT 63.59 2.925 63.61 3.415 ;
      RECT 63.58 2.866 63.59 3.4 ;
      RECT 63.53 2.756 63.58 3.36 ;
      RECT 63.52 2.65 63.53 3.315 ;
      RECT 63.49 2.579 63.52 3.235 ;
      RECT 63.48 2.511 63.49 3.16 ;
      RECT 63.47 2.225 63.48 3.125 ;
      RECT 63.44 2.225 63.47 3.055 ;
      RECT 63.43 2.225 63.44 2.95 ;
      RECT 63.42 2.225 63.43 2.915 ;
      RECT 63.35 2.225 63.42 2.775 ;
      RECT 63.32 2.225 63.35 2.575 ;
      RECT 63.31 2.225 63.32 2.5 ;
      RECT 67.65 2.155 67.91 2.415 ;
      RECT 67.64 2.155 67.91 2.365 ;
      RECT 67.61 2.025 67.89 2.305 ;
      RECT 56.13 6.655 56.48 7.005 ;
      RECT 67.095 6.61 67.445 6.96 ;
      RECT 56.13 6.685 67.445 6.885 ;
      RECT 66.65 3.705 66.93 3.985 ;
      RECT 66.69 3.665 66.96 3.925 ;
      RECT 66.68 3.7 66.96 3.925 ;
      RECT 66.69 3.66 66.9 3.985 ;
      RECT 66.69 3.655 66.89 3.985 ;
      RECT 66.73 3.645 66.89 3.985 ;
      RECT 66.7 3.65 66.89 3.985 ;
      RECT 66.74 3.64 66.83 3.985 ;
      RECT 66.76 3.635 66.83 3.985 ;
      RECT 66.07 3.155 66.33 3.415 ;
      RECT 66.12 3.065 66.31 3.415 ;
      RECT 66.15 2.85 66.31 3.415 ;
      RECT 66.24 2.455 66.31 3.415 ;
      RECT 66.26 2.165 66.396 2.893 ;
      RECT 66.2 2.66 66.396 2.893 ;
      RECT 66.22 2.54 66.31 3.415 ;
      RECT 66.26 2.165 66.42 2.558 ;
      RECT 66.26 2.165 66.43 2.455 ;
      RECT 66.25 2.165 66.51 2.425 ;
      RECT 65.65 3.705 65.93 3.985 ;
      RECT 65.67 3.665 65.93 3.985 ;
      RECT 65.31 3.625 65.42 3.885 ;
      RECT 65.17 2.115 65.26 2.375 ;
      RECT 65.7 3.17 65.71 3.3 ;
      RECT 65.69 3.135 65.7 3.454 ;
      RECT 65.61 3.067 65.69 3.534 ;
      RECT 65.64 3.71 65.65 3.93 ;
      RECT 65.62 3.705 65.64 3.919 ;
      RECT 65.59 3.7 65.62 3.904 ;
      RECT 65.6 3.002 65.61 3.61 ;
      RECT 65.58 2.946 65.6 3.625 ;
      RECT 65.57 3.685 65.59 3.89 ;
      RECT 65.57 2.874 65.58 3.645 ;
      RECT 65.54 2.777 65.57 3.885 ;
      RECT 65.52 2.66 65.54 3.885 ;
      RECT 65.49 2.54 65.52 3.885 ;
      RECT 65.48 2.455 65.49 3.885 ;
      RECT 65.47 2.4 65.48 3.885 ;
      RECT 65.46 2.355 65.47 3.104 ;
      RECT 65.45 3.315 65.47 3.885 ;
      RECT 65.45 2.285 65.46 3.061 ;
      RECT 65.43 2.235 65.45 2.996 ;
      RECT 65.44 3.395 65.45 3.885 ;
      RECT 65.42 3.495 65.44 3.885 ;
      RECT 65.37 2.115 65.43 2.824 ;
      RECT 65.36 2.115 65.37 2.66 ;
      RECT 65.35 2.115 65.36 2.61 ;
      RECT 65.3 2.115 65.35 2.54 ;
      RECT 65.28 2.115 65.3 2.455 ;
      RECT 65.26 2.115 65.28 2.41 ;
      RECT 64.58 3.565 64.63 3.825 ;
      RECT 64.49 2.095 64.63 2.355 ;
      RECT 64.99 2.72 65 2.808 ;
      RECT 64.98 2.655 64.99 2.854 ;
      RECT 64.97 2.605 64.98 2.9 ;
      RECT 64.92 2.552 64.97 3.039 ;
      RECT 64.91 2.501 64.92 3.23 ;
      RECT 64.87 2.459 64.91 3.335 ;
      RECT 64.85 2.405 64.87 3.472 ;
      RECT 64.84 2.38 64.85 2.688 ;
      RECT 64.84 2.77 64.85 3.542 ;
      RECT 64.83 2.366 64.84 2.673 ;
      RECT 64.83 2.825 64.84 3.825 ;
      RECT 64.81 2.341 64.83 2.655 ;
      RECT 64.79 3 64.83 3.825 ;
      RECT 64.8 2.315 64.81 2.635 ;
      RECT 64.77 2.28 64.8 2.589 ;
      RECT 64.78 3.125 64.79 3.825 ;
      RECT 64.77 3.205 64.78 3.825 ;
      RECT 64.76 2.245 64.77 2.554 ;
      RECT 64.72 3.275 64.77 3.825 ;
      RECT 64.75 2.225 64.76 2.53 ;
      RECT 64.72 2.095 64.75 2.495 ;
      RECT 64.71 2.095 64.72 2.46 ;
      RECT 64.69 3.375 64.72 3.825 ;
      RECT 64.69 2.095 64.71 2.435 ;
      RECT 64.68 2.095 64.69 2.41 ;
      RECT 64.64 3.475 64.69 3.825 ;
      RECT 64.66 2.095 64.68 2.38 ;
      RECT 64.63 2.095 64.66 2.365 ;
      RECT 64.63 3.55 64.64 3.825 ;
      RECT 64.55 2.635 64.59 2.895 ;
      RECT 60.28 2.055 60.54 2.315 ;
      RECT 60.28 2.085 60.56 2.295 ;
      RECT 62.49 1.905 62.67 2.055 ;
      RECT 64.54 2.63 64.55 2.895 ;
      RECT 64.52 2.62 64.54 2.895 ;
      RECT 64.502 2.613 64.52 2.895 ;
      RECT 64.416 2.602 64.502 2.895 ;
      RECT 64.33 2.585 64.416 2.895 ;
      RECT 64.28 2.572 64.33 2.82 ;
      RECT 64.246 2.564 64.28 2.795 ;
      RECT 64.16 2.553 64.246 2.76 ;
      RECT 64.12 2.53 64.16 2.723 ;
      RECT 64.11 2.495 64.12 2.708 ;
      RECT 64.1 2.455 64.11 2.703 ;
      RECT 64.09 2.435 64.1 2.698 ;
      RECT 64.075 2.395 64.09 2.693 ;
      RECT 64.06 2.347 64.075 2.689 ;
      RECT 64.05 2.306 64.06 2.686 ;
      RECT 64.04 2.268 64.05 2.675 ;
      RECT 64.02 2.212 64.04 2.655 ;
      RECT 64 2.16 64.02 2.591 ;
      RECT 63.98 2.11 64 2.543 ;
      RECT 63.97 2.08 63.98 2.507 ;
      RECT 63.965 2.062 63.97 2.493 ;
      RECT 63.95 2.053 63.965 2.475 ;
      RECT 63.92 2.034 63.95 2.415 ;
      RECT 63.91 2.017 63.92 2.37 ;
      RECT 63.9 2.009 63.91 2.34 ;
      RECT 63.87 1.997 63.9 2.29 ;
      RECT 63.85 1.985 63.87 2.225 ;
      RECT 63.84 1.977 63.85 2.185 ;
      RECT 63.82 1.974 63.84 2.175 ;
      RECT 63.805 1.972 63.82 2.17 ;
      RECT 63.785 1.971 63.805 2.16 ;
      RECT 63.77 1.97 63.785 2.15 ;
      RECT 63.75 1.969 63.77 2.145 ;
      RECT 63.748 1.969 63.75 2.145 ;
      RECT 63.662 1.966 63.748 2.142 ;
      RECT 63.576 1.961 63.662 2.135 ;
      RECT 63.49 1.956 63.576 2.129 ;
      RECT 63.44 1.953 63.49 2.12 ;
      RECT 63.396 1.951 63.44 2.114 ;
      RECT 63.31 1.947 63.396 2.109 ;
      RECT 63.306 1.945 63.31 2.105 ;
      RECT 63.22 1.942 63.306 2.1 ;
      RECT 63.166 1.938 63.22 2.093 ;
      RECT 63.08 1.935 63.166 2.088 ;
      RECT 63.056 1.932 63.08 2.084 ;
      RECT 62.97 1.93 63.056 2.079 ;
      RECT 62.91 1.926 62.97 2.073 ;
      RECT 62.902 1.924 62.91 2.07 ;
      RECT 62.816 1.92 62.902 2.066 ;
      RECT 62.73 1.913 62.816 2.059 ;
      RECT 62.67 1.907 62.73 2.055 ;
      RECT 62.47 1.905 62.49 2.058 ;
      RECT 62.42 1.915 62.47 2.068 ;
      RECT 62.39 1.925 62.42 2.08 ;
      RECT 62.366 1.927 62.39 2.086 ;
      RECT 62.28 1.93 62.366 2.091 ;
      RECT 62.21 1.935 62.28 2.1 ;
      RECT 62.196 1.937 62.21 2.106 ;
      RECT 62.11 1.941 62.196 2.111 ;
      RECT 62.07 1.945 62.11 2.12 ;
      RECT 62.056 1.947 62.07 2.126 ;
      RECT 61.97 1.951 62.056 2.131 ;
      RECT 61.886 1.957 61.97 2.138 ;
      RECT 61.8 1.963 61.886 2.143 ;
      RECT 61.776 1.967 61.8 2.146 ;
      RECT 61.69 1.971 61.776 2.151 ;
      RECT 61.64 1.976 61.69 2.16 ;
      RECT 61.56 1.981 61.64 2.17 ;
      RECT 61.48 1.987 61.56 2.185 ;
      RECT 61.46 1.991 61.48 2.195 ;
      RECT 61.39 1.994 61.46 2.205 ;
      RECT 61.34 1.999 61.39 2.22 ;
      RECT 61.31 2.002 61.34 2.24 ;
      RECT 61.3 2.004 61.31 2.256 ;
      RECT 61.24 2.016 61.3 2.266 ;
      RECT 61.22 2.031 61.24 2.275 ;
      RECT 61.21 2.05 61.22 2.275 ;
      RECT 61.2 2.07 61.21 2.275 ;
      RECT 61.18 2.08 61.2 2.275 ;
      RECT 61.13 2.09 61.18 2.275 ;
      RECT 61.1 2.096 61.13 2.275 ;
      RECT 61.03 2.101 61.1 2.277 ;
      RECT 60.95 2.102 61.03 2.282 ;
      RECT 60.946 2.1 60.95 2.285 ;
      RECT 60.86 2.097 60.946 2.286 ;
      RECT 60.818 2.094 60.86 2.288 ;
      RECT 60.732 2.092 60.818 2.289 ;
      RECT 60.646 2.089 60.732 2.292 ;
      RECT 60.56 2.086 60.646 2.294 ;
      RECT 62.49 3.145 62.77 3.425 ;
      RECT 62.52 3.125 62.79 3.385 ;
      RECT 62.52 3.075 62.75 3.425 ;
      RECT 62.59 3.065 62.75 3.425 ;
      RECT 62.59 2.775 62.74 3.425 ;
      RECT 62.58 2.455 62.73 2.825 ;
      RECT 62.57 2.455 62.73 2.695 ;
      RECT 62.55 2.165 62.72 2.5 ;
      RECT 62.53 2.165 62.72 2.45 ;
      RECT 62.49 2.165 62.75 2.425 ;
      RECT 62.4 3.635 62.48 3.895 ;
      RECT 61.69 2.355 61.81 2.615 ;
      RECT 62.375 3.615 62.4 3.895 ;
      RECT 62.36 3.577 62.375 3.895 ;
      RECT 62.32 3.52 62.36 3.895 ;
      RECT 62.29 3.43 62.32 3.895 ;
      RECT 62.25 3.33 62.29 3.895 ;
      RECT 62.22 3.23 62.25 3.895 ;
      RECT 62.215 3.177 62.22 3.718 ;
      RECT 62.2 3.147 62.215 3.684 ;
      RECT 62.19 3.108 62.2 3.649 ;
      RECT 62.18 3.075 62.19 3.605 ;
      RECT 62.17 3.042 62.18 3.57 ;
      RECT 62.14 2.976 62.17 3.505 ;
      RECT 62.13 2.911 62.14 3.43 ;
      RECT 62.12 2.881 62.13 3.4 ;
      RECT 62.08 2.811 62.12 3.33 ;
      RECT 62.07 2.746 62.08 3.245 ;
      RECT 62.06 2.728 62.07 3.23 ;
      RECT 62.05 2.711 62.06 3.195 ;
      RECT 62.04 2.694 62.05 3.165 ;
      RECT 62.03 2.677 62.04 3.135 ;
      RECT 62.01 2.652 62.03 3.075 ;
      RECT 62 2.626 62.01 3.02 ;
      RECT 61.98 2.601 62 2.98 ;
      RECT 61.97 2.57 61.98 2.945 ;
      RECT 61.96 2.557 61.97 2.9 ;
      RECT 61.95 2.542 61.96 2.875 ;
      RECT 61.94 2.355 61.95 2.835 ;
      RECT 61.93 2.355 61.94 2.805 ;
      RECT 61.925 2.355 61.93 2.788 ;
      RECT 61.92 2.355 61.925 2.77 ;
      RECT 61.85 2.355 61.92 2.71 ;
      RECT 61.81 2.355 61.85 2.645 ;
      RECT 61.64 3.225 61.9 3.485 ;
      RECT 59.81 3.145 59.89 3.465 ;
      RECT 59.63 3.205 59.78 3.465 ;
      RECT 59.81 3.145 59.92 3.425 ;
      RECT 61.63 3.317 61.64 3.48 ;
      RECT 61.6 3.327 61.63 3.488 ;
      RECT 61.58 3.335 61.6 3.493 ;
      RECT 61.512 3.343 61.58 3.503 ;
      RECT 61.426 3.363 61.512 3.52 ;
      RECT 61.34 3.384 61.426 3.539 ;
      RECT 61.33 3.4 61.34 3.55 ;
      RECT 61.29 3.41 61.33 3.556 ;
      RECT 61.27 3.415 61.29 3.563 ;
      RECT 61.232 3.416 61.27 3.566 ;
      RECT 61.146 3.419 61.232 3.567 ;
      RECT 61.06 3.423 61.146 3.568 ;
      RECT 61.006 3.425 61.06 3.57 ;
      RECT 60.92 3.425 61.006 3.572 ;
      RECT 60.88 3.42 60.92 3.574 ;
      RECT 60.87 3.414 60.88 3.575 ;
      RECT 60.83 3.409 60.87 3.571 ;
      RECT 60.82 3.4 60.83 3.567 ;
      RECT 60.788 3.391 60.82 3.564 ;
      RECT 60.702 3.379 60.788 3.554 ;
      RECT 60.616 3.362 60.702 3.539 ;
      RECT 60.53 3.344 60.616 3.525 ;
      RECT 60.51 3.335 60.53 3.516 ;
      RECT 60.44 3.325 60.51 3.509 ;
      RECT 60.39 3.31 60.44 3.499 ;
      RECT 60.33 3.3 60.39 3.49 ;
      RECT 60.29 3.29 60.33 3.485 ;
      RECT 60.24 3.28 60.29 3.479 ;
      RECT 60.2 3.268 60.24 3.469 ;
      RECT 60.18 3.258 60.2 3.465 ;
      RECT 60.16 3.248 60.18 3.465 ;
      RECT 60.15 3.238 60.16 3.464 ;
      RECT 60.13 3.23 60.15 3.46 ;
      RECT 60.09 3.205 60.13 3.454 ;
      RECT 60.07 3.145 60.09 3.447 ;
      RECT 60.046 3.145 60.07 3.444 ;
      RECT 59.96 3.145 60.046 3.439 ;
      RECT 59.92 3.145 59.96 3.43 ;
      RECT 59.78 3.195 59.81 3.465 ;
      RECT 61.46 2.775 61.72 3.035 ;
      RECT 61.42 2.775 61.72 2.915 ;
      RECT 61.39 2.775 61.72 2.9 ;
      RECT 61.33 2.775 61.72 2.88 ;
      RECT 61.25 2.585 61.53 2.865 ;
      RECT 61.25 2.77 61.6 2.865 ;
      RECT 61.25 2.71 61.59 2.865 ;
      RECT 61.25 2.66 61.54 2.865 ;
      RECT 59.02 3.115 59.28 3.375 ;
      RECT 59.165 1.205 59.28 3.375 ;
      RECT 59.08 2.585 59.28 3.375 ;
      RECT 60.39 2.635 60.65 2.895 ;
      RECT 59.075 2.585 59.28 2.87 ;
      RECT 59.07 2.585 59.28 2.865 ;
      RECT 60.37 2.645 60.65 2.825 ;
      RECT 59.96 2.615 60.1 2.765 ;
      RECT 59.335 1.205 59.415 1.55 ;
      RECT 59.07 1.205 59.28 1.55 ;
      RECT 60.36 2.644 60.37 2.825 ;
      RECT 60.356 2.644 60.36 2.825 ;
      RECT 60.27 2.639 60.356 2.814 ;
      RECT 60.196 2.63 60.27 2.794 ;
      RECT 60.11 2.621 60.196 2.775 ;
      RECT 60.1 2.615 60.11 2.765 ;
      RECT 59.92 2.615 59.96 2.768 ;
      RECT 59.834 2.615 59.92 2.776 ;
      RECT 59.748 2.615 59.834 2.787 ;
      RECT 59.662 2.615 59.748 2.798 ;
      RECT 59.576 2.615 59.662 2.809 ;
      RECT 59.49 2.615 59.576 2.82 ;
      RECT 59.46 2.615 59.49 2.86 ;
      RECT 59.43 2.615 59.46 2.91 ;
      RECT 59.355 2.615 59.43 2.93 ;
      RECT 59.35 2.59 59.355 2.935 ;
      RECT 59.335 2.585 59.35 2.943 ;
      RECT 59.33 1.205 59.335 2.953 ;
      RECT 59.3 1.205 59.33 2.995 ;
      RECT 59.28 1.205 59.3 3.075 ;
      RECT 58.41 2.965 58.43 3.404 ;
      RECT 58.41 2.965 58.516 3.401 ;
      RECT 58.4 3.08 58.516 3.4 ;
      RECT 58.43 2.115 58.56 3.397 ;
      RECT 58.41 2.985 58.57 3.395 ;
      RECT 58.41 3.07 58.58 3.39 ;
      RECT 58.38 3.115 58.58 3.385 ;
      RECT 58.38 3.115 58.59 3.38 ;
      RECT 58.36 3.115 58.62 3.375 ;
      RECT 58.43 2.115 58.59 2.765 ;
      RECT 58.42 2.115 58.59 2.74 ;
      RECT 58.42 2.115 58.61 2.505 ;
      RECT 58.37 2.115 58.63 2.375 ;
      RECT 57.84 2.605 58.13 2.865 ;
      RECT 57.85 2.585 58.13 2.865 ;
      RECT 57.8 2.665 58.13 2.86 ;
      RECT 57.87 2.578 58.04 2.865 ;
      RECT 57.87 2.565 57.996 2.865 ;
      RECT 57.91 2.558 57.996 2.865 ;
      RECT 57.37 3.705 57.65 3.985 ;
      RECT 57.33 3.67 57.63 3.78 ;
      RECT 57.32 3.62 57.61 3.675 ;
      RECT 57.26 3.385 57.52 3.645 ;
      RECT 57.26 3.525 57.6 3.645 ;
      RECT 57.26 3.475 57.58 3.645 ;
      RECT 57.26 3.43 57.57 3.645 ;
      RECT 57.26 3.415 57.54 3.645 ;
      RECT 52.995 6.225 53.315 6.545 ;
      RECT 53.025 5.695 53.195 6.545 ;
      RECT 53.025 5.695 53.2 6.045 ;
      RECT 53.025 5.695 54 5.87 ;
      RECT 53.825 1.965 54 5.87 ;
      RECT 53.77 1.965 54.12 2.315 ;
      RECT 53.795 6.655 54.12 6.98 ;
      RECT 52.68 6.745 54.12 6.915 ;
      RECT 52.68 2.395 52.84 6.915 ;
      RECT 52.995 2.365 53.315 2.685 ;
      RECT 52.68 2.395 53.315 2.565 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 43.27 0.96 43.645 1.33 ;
      RECT 41.835 0.96 42.21 1.33 ;
      RECT 41.835 1.08 51.655 1.25 ;
      RECT 45.955 4.36 51.635 4.53 ;
      RECT 51.465 3.425 51.635 4.53 ;
      RECT 45.765 3.595 45.785 4.53 ;
      RECT 46.015 3.705 46.045 3.985 ;
      RECT 45.725 3.595 45.785 3.855 ;
      RECT 51.375 3.43 51.725 3.78 ;
      RECT 45.555 2.225 45.585 2.485 ;
      RECT 45.325 2.225 45.385 2.485 ;
      RECT 46.005 3.685 46.015 3.985 ;
      RECT 45.985 3.605 46.005 3.985 ;
      RECT 45.975 3.545 45.985 3.985 ;
      RECT 45.955 3.495 45.975 3.985 ;
      RECT 45.925 3.395 45.955 4.53 ;
      RECT 45.915 3.305 45.925 4.53 ;
      RECT 45.875 3.245 45.915 4.53 ;
      RECT 45.871 3.214 45.875 4.53 ;
      RECT 45.785 3.205 45.871 4.53 ;
      RECT 45.775 3.196 45.785 3.55 ;
      RECT 45.745 3.175 45.775 3.517 ;
      RECT 45.735 3.125 45.745 3.493 ;
      RECT 45.725 3.09 45.735 3.481 ;
      RECT 45.685 3.015 45.725 3.45 ;
      RECT 45.665 2.925 45.685 3.415 ;
      RECT 45.655 2.866 45.665 3.4 ;
      RECT 45.605 2.756 45.655 3.36 ;
      RECT 45.595 2.65 45.605 3.315 ;
      RECT 45.565 2.579 45.595 3.235 ;
      RECT 45.555 2.511 45.565 3.16 ;
      RECT 45.545 2.225 45.555 3.125 ;
      RECT 45.515 2.225 45.545 3.055 ;
      RECT 45.505 2.225 45.515 2.95 ;
      RECT 45.495 2.225 45.505 2.915 ;
      RECT 45.425 2.225 45.495 2.775 ;
      RECT 45.395 2.225 45.425 2.575 ;
      RECT 45.385 2.225 45.395 2.5 ;
      RECT 49.725 2.155 49.985 2.415 ;
      RECT 49.715 2.155 49.985 2.365 ;
      RECT 49.685 2.025 49.965 2.305 ;
      RECT 38.25 6.66 38.6 7.01 ;
      RECT 49.225 6.615 49.575 6.965 ;
      RECT 38.25 6.69 49.575 6.89 ;
      RECT 48.725 3.705 49.005 3.985 ;
      RECT 48.765 3.665 49.035 3.925 ;
      RECT 48.755 3.7 49.035 3.925 ;
      RECT 48.765 3.66 48.975 3.985 ;
      RECT 48.765 3.655 48.965 3.985 ;
      RECT 48.805 3.645 48.965 3.985 ;
      RECT 48.775 3.65 48.965 3.985 ;
      RECT 48.815 3.64 48.905 3.985 ;
      RECT 48.835 3.635 48.905 3.985 ;
      RECT 48.145 3.155 48.405 3.415 ;
      RECT 48.195 3.065 48.385 3.415 ;
      RECT 48.225 2.85 48.385 3.415 ;
      RECT 48.315 2.455 48.385 3.415 ;
      RECT 48.335 2.165 48.471 2.893 ;
      RECT 48.275 2.66 48.471 2.893 ;
      RECT 48.295 2.54 48.385 3.415 ;
      RECT 48.335 2.165 48.495 2.558 ;
      RECT 48.335 2.165 48.505 2.455 ;
      RECT 48.325 2.165 48.585 2.425 ;
      RECT 47.725 3.705 48.005 3.985 ;
      RECT 47.745 3.665 48.005 3.985 ;
      RECT 47.385 3.625 47.495 3.885 ;
      RECT 47.245 2.115 47.335 2.375 ;
      RECT 47.775 3.17 47.785 3.3 ;
      RECT 47.765 3.135 47.775 3.454 ;
      RECT 47.685 3.067 47.765 3.534 ;
      RECT 47.715 3.71 47.725 3.93 ;
      RECT 47.695 3.705 47.715 3.919 ;
      RECT 47.665 3.7 47.695 3.904 ;
      RECT 47.675 3.002 47.685 3.61 ;
      RECT 47.655 2.946 47.675 3.625 ;
      RECT 47.645 3.685 47.665 3.89 ;
      RECT 47.645 2.874 47.655 3.645 ;
      RECT 47.615 2.777 47.645 3.885 ;
      RECT 47.595 2.66 47.615 3.885 ;
      RECT 47.565 2.54 47.595 3.885 ;
      RECT 47.555 2.455 47.565 3.885 ;
      RECT 47.545 2.4 47.555 3.885 ;
      RECT 47.535 2.355 47.545 3.104 ;
      RECT 47.525 3.315 47.545 3.885 ;
      RECT 47.525 2.285 47.535 3.061 ;
      RECT 47.505 2.235 47.525 2.996 ;
      RECT 47.515 3.395 47.525 3.885 ;
      RECT 47.495 3.495 47.515 3.885 ;
      RECT 47.445 2.115 47.505 2.824 ;
      RECT 47.435 2.115 47.445 2.66 ;
      RECT 47.425 2.115 47.435 2.61 ;
      RECT 47.375 2.115 47.425 2.54 ;
      RECT 47.355 2.115 47.375 2.455 ;
      RECT 47.335 2.115 47.355 2.41 ;
      RECT 46.655 3.565 46.705 3.825 ;
      RECT 46.565 2.095 46.705 2.355 ;
      RECT 47.065 2.72 47.075 2.808 ;
      RECT 47.055 2.655 47.065 2.854 ;
      RECT 47.045 2.605 47.055 2.9 ;
      RECT 46.995 2.552 47.045 3.039 ;
      RECT 46.985 2.501 46.995 3.23 ;
      RECT 46.945 2.459 46.985 3.335 ;
      RECT 46.925 2.405 46.945 3.472 ;
      RECT 46.915 2.38 46.925 2.688 ;
      RECT 46.915 2.77 46.925 3.542 ;
      RECT 46.905 2.366 46.915 2.673 ;
      RECT 46.905 2.825 46.915 3.825 ;
      RECT 46.885 2.341 46.905 2.655 ;
      RECT 46.865 3 46.905 3.825 ;
      RECT 46.875 2.315 46.885 2.635 ;
      RECT 46.845 2.28 46.875 2.589 ;
      RECT 46.855 3.125 46.865 3.825 ;
      RECT 46.845 3.205 46.855 3.825 ;
      RECT 46.835 2.245 46.845 2.554 ;
      RECT 46.795 3.275 46.845 3.825 ;
      RECT 46.825 2.225 46.835 2.53 ;
      RECT 46.795 2.095 46.825 2.495 ;
      RECT 46.785 2.095 46.795 2.46 ;
      RECT 46.765 3.375 46.795 3.825 ;
      RECT 46.765 2.095 46.785 2.435 ;
      RECT 46.755 2.095 46.765 2.41 ;
      RECT 46.715 3.475 46.765 3.825 ;
      RECT 46.735 2.095 46.755 2.38 ;
      RECT 46.705 2.095 46.735 2.365 ;
      RECT 46.705 3.55 46.715 3.825 ;
      RECT 46.625 2.635 46.665 2.895 ;
      RECT 42.355 2.055 42.615 2.315 ;
      RECT 42.355 2.085 42.635 2.295 ;
      RECT 44.565 1.905 44.745 2.055 ;
      RECT 46.615 2.63 46.625 2.895 ;
      RECT 46.595 2.62 46.615 2.895 ;
      RECT 46.577 2.613 46.595 2.895 ;
      RECT 46.491 2.602 46.577 2.895 ;
      RECT 46.405 2.585 46.491 2.895 ;
      RECT 46.355 2.572 46.405 2.82 ;
      RECT 46.321 2.564 46.355 2.795 ;
      RECT 46.235 2.553 46.321 2.76 ;
      RECT 46.195 2.53 46.235 2.723 ;
      RECT 46.185 2.495 46.195 2.708 ;
      RECT 46.175 2.455 46.185 2.703 ;
      RECT 46.165 2.435 46.175 2.698 ;
      RECT 46.15 2.395 46.165 2.693 ;
      RECT 46.135 2.347 46.15 2.689 ;
      RECT 46.125 2.306 46.135 2.686 ;
      RECT 46.115 2.268 46.125 2.675 ;
      RECT 46.095 2.212 46.115 2.655 ;
      RECT 46.075 2.16 46.095 2.591 ;
      RECT 46.055 2.11 46.075 2.543 ;
      RECT 46.045 2.08 46.055 2.507 ;
      RECT 46.04 2.062 46.045 2.493 ;
      RECT 46.025 2.053 46.04 2.475 ;
      RECT 45.995 2.034 46.025 2.415 ;
      RECT 45.985 2.017 45.995 2.37 ;
      RECT 45.975 2.009 45.985 2.34 ;
      RECT 45.945 1.997 45.975 2.29 ;
      RECT 45.925 1.985 45.945 2.225 ;
      RECT 45.915 1.977 45.925 2.185 ;
      RECT 45.895 1.974 45.915 2.175 ;
      RECT 45.88 1.972 45.895 2.17 ;
      RECT 45.86 1.971 45.88 2.16 ;
      RECT 45.845 1.97 45.86 2.15 ;
      RECT 45.825 1.969 45.845 2.145 ;
      RECT 45.823 1.969 45.825 2.145 ;
      RECT 45.737 1.966 45.823 2.142 ;
      RECT 45.651 1.961 45.737 2.135 ;
      RECT 45.565 1.956 45.651 2.129 ;
      RECT 45.515 1.953 45.565 2.12 ;
      RECT 45.471 1.951 45.515 2.114 ;
      RECT 45.385 1.947 45.471 2.109 ;
      RECT 45.381 1.945 45.385 2.105 ;
      RECT 45.295 1.942 45.381 2.1 ;
      RECT 45.241 1.938 45.295 2.093 ;
      RECT 45.155 1.935 45.241 2.088 ;
      RECT 45.131 1.932 45.155 2.084 ;
      RECT 45.045 1.93 45.131 2.079 ;
      RECT 44.985 1.926 45.045 2.073 ;
      RECT 44.977 1.924 44.985 2.07 ;
      RECT 44.891 1.92 44.977 2.066 ;
      RECT 44.805 1.913 44.891 2.059 ;
      RECT 44.745 1.907 44.805 2.055 ;
      RECT 44.545 1.905 44.565 2.058 ;
      RECT 44.495 1.915 44.545 2.068 ;
      RECT 44.465 1.925 44.495 2.08 ;
      RECT 44.441 1.927 44.465 2.086 ;
      RECT 44.355 1.93 44.441 2.091 ;
      RECT 44.285 1.935 44.355 2.1 ;
      RECT 44.271 1.937 44.285 2.106 ;
      RECT 44.185 1.941 44.271 2.111 ;
      RECT 44.145 1.945 44.185 2.12 ;
      RECT 44.131 1.947 44.145 2.126 ;
      RECT 44.045 1.951 44.131 2.131 ;
      RECT 43.961 1.957 44.045 2.138 ;
      RECT 43.875 1.963 43.961 2.143 ;
      RECT 43.851 1.967 43.875 2.146 ;
      RECT 43.765 1.971 43.851 2.151 ;
      RECT 43.715 1.976 43.765 2.16 ;
      RECT 43.635 1.981 43.715 2.17 ;
      RECT 43.555 1.987 43.635 2.185 ;
      RECT 43.535 1.991 43.555 2.195 ;
      RECT 43.465 1.994 43.535 2.205 ;
      RECT 43.415 1.999 43.465 2.22 ;
      RECT 43.385 2.002 43.415 2.24 ;
      RECT 43.375 2.004 43.385 2.256 ;
      RECT 43.315 2.016 43.375 2.266 ;
      RECT 43.295 2.031 43.315 2.275 ;
      RECT 43.285 2.05 43.295 2.275 ;
      RECT 43.275 2.07 43.285 2.275 ;
      RECT 43.255 2.08 43.275 2.275 ;
      RECT 43.205 2.09 43.255 2.275 ;
      RECT 43.175 2.096 43.205 2.275 ;
      RECT 43.105 2.101 43.175 2.277 ;
      RECT 43.025 2.102 43.105 2.282 ;
      RECT 43.021 2.1 43.025 2.285 ;
      RECT 42.935 2.097 43.021 2.286 ;
      RECT 42.893 2.094 42.935 2.288 ;
      RECT 42.807 2.092 42.893 2.289 ;
      RECT 42.721 2.089 42.807 2.292 ;
      RECT 42.635 2.086 42.721 2.294 ;
      RECT 44.565 3.145 44.845 3.425 ;
      RECT 44.595 3.125 44.865 3.385 ;
      RECT 44.595 3.075 44.825 3.425 ;
      RECT 44.665 3.065 44.825 3.425 ;
      RECT 44.665 2.775 44.815 3.425 ;
      RECT 44.655 2.455 44.805 2.825 ;
      RECT 44.645 2.455 44.805 2.695 ;
      RECT 44.625 2.165 44.795 2.5 ;
      RECT 44.605 2.165 44.795 2.45 ;
      RECT 44.565 2.165 44.825 2.425 ;
      RECT 44.475 3.635 44.555 3.895 ;
      RECT 43.765 2.355 43.885 2.615 ;
      RECT 44.45 3.615 44.475 3.895 ;
      RECT 44.435 3.577 44.45 3.895 ;
      RECT 44.395 3.52 44.435 3.895 ;
      RECT 44.365 3.43 44.395 3.895 ;
      RECT 44.325 3.33 44.365 3.895 ;
      RECT 44.295 3.23 44.325 3.895 ;
      RECT 44.29 3.177 44.295 3.718 ;
      RECT 44.275 3.147 44.29 3.684 ;
      RECT 44.265 3.108 44.275 3.649 ;
      RECT 44.255 3.075 44.265 3.605 ;
      RECT 44.245 3.042 44.255 3.57 ;
      RECT 44.215 2.976 44.245 3.505 ;
      RECT 44.205 2.911 44.215 3.43 ;
      RECT 44.195 2.881 44.205 3.4 ;
      RECT 44.155 2.811 44.195 3.33 ;
      RECT 44.145 2.746 44.155 3.245 ;
      RECT 44.135 2.728 44.145 3.23 ;
      RECT 44.125 2.711 44.135 3.195 ;
      RECT 44.115 2.694 44.125 3.165 ;
      RECT 44.105 2.677 44.115 3.135 ;
      RECT 44.085 2.652 44.105 3.075 ;
      RECT 44.075 2.626 44.085 3.02 ;
      RECT 44.055 2.601 44.075 2.98 ;
      RECT 44.045 2.57 44.055 2.945 ;
      RECT 44.035 2.557 44.045 2.9 ;
      RECT 44.025 2.542 44.035 2.875 ;
      RECT 44.015 2.355 44.025 2.835 ;
      RECT 44.005 2.355 44.015 2.805 ;
      RECT 44 2.355 44.005 2.788 ;
      RECT 43.995 2.355 44 2.77 ;
      RECT 43.925 2.355 43.995 2.71 ;
      RECT 43.885 2.355 43.925 2.645 ;
      RECT 43.715 3.225 43.975 3.485 ;
      RECT 41.885 3.145 41.965 3.465 ;
      RECT 41.705 3.205 41.855 3.465 ;
      RECT 41.885 3.145 41.995 3.425 ;
      RECT 43.705 3.317 43.715 3.48 ;
      RECT 43.675 3.327 43.705 3.488 ;
      RECT 43.655 3.335 43.675 3.493 ;
      RECT 43.587 3.343 43.655 3.503 ;
      RECT 43.501 3.363 43.587 3.52 ;
      RECT 43.415 3.384 43.501 3.539 ;
      RECT 43.405 3.4 43.415 3.55 ;
      RECT 43.365 3.41 43.405 3.556 ;
      RECT 43.345 3.415 43.365 3.563 ;
      RECT 43.307 3.416 43.345 3.566 ;
      RECT 43.221 3.419 43.307 3.567 ;
      RECT 43.135 3.423 43.221 3.568 ;
      RECT 43.081 3.425 43.135 3.57 ;
      RECT 42.995 3.425 43.081 3.572 ;
      RECT 42.955 3.42 42.995 3.574 ;
      RECT 42.945 3.414 42.955 3.575 ;
      RECT 42.905 3.409 42.945 3.571 ;
      RECT 42.895 3.4 42.905 3.567 ;
      RECT 42.863 3.391 42.895 3.564 ;
      RECT 42.777 3.379 42.863 3.554 ;
      RECT 42.691 3.362 42.777 3.539 ;
      RECT 42.605 3.344 42.691 3.525 ;
      RECT 42.585 3.335 42.605 3.516 ;
      RECT 42.515 3.325 42.585 3.509 ;
      RECT 42.465 3.31 42.515 3.499 ;
      RECT 42.405 3.3 42.465 3.49 ;
      RECT 42.365 3.29 42.405 3.485 ;
      RECT 42.315 3.28 42.365 3.479 ;
      RECT 42.275 3.268 42.315 3.469 ;
      RECT 42.255 3.258 42.275 3.465 ;
      RECT 42.235 3.248 42.255 3.465 ;
      RECT 42.225 3.238 42.235 3.464 ;
      RECT 42.205 3.23 42.225 3.46 ;
      RECT 42.165 3.205 42.205 3.454 ;
      RECT 42.145 3.145 42.165 3.447 ;
      RECT 42.121 3.145 42.145 3.444 ;
      RECT 42.035 3.145 42.121 3.439 ;
      RECT 41.995 3.145 42.035 3.43 ;
      RECT 41.855 3.195 41.885 3.465 ;
      RECT 43.535 2.775 43.795 3.035 ;
      RECT 43.495 2.775 43.795 2.915 ;
      RECT 43.465 2.775 43.795 2.9 ;
      RECT 43.405 2.775 43.795 2.88 ;
      RECT 43.325 2.585 43.605 2.865 ;
      RECT 43.325 2.77 43.675 2.865 ;
      RECT 43.325 2.71 43.665 2.865 ;
      RECT 43.325 2.66 43.615 2.865 ;
      RECT 41.095 3.115 41.355 3.375 ;
      RECT 41.24 1.205 41.355 3.375 ;
      RECT 41.155 2.585 41.355 3.375 ;
      RECT 42.465 2.635 42.725 2.895 ;
      RECT 41.15 2.585 41.355 2.87 ;
      RECT 41.145 2.585 41.355 2.865 ;
      RECT 42.445 2.645 42.725 2.825 ;
      RECT 42.035 2.615 42.175 2.765 ;
      RECT 41.41 1.205 41.49 1.55 ;
      RECT 41.145 1.205 41.355 1.55 ;
      RECT 42.435 2.644 42.445 2.825 ;
      RECT 42.431 2.644 42.435 2.825 ;
      RECT 42.345 2.639 42.431 2.814 ;
      RECT 42.271 2.63 42.345 2.794 ;
      RECT 42.185 2.621 42.271 2.775 ;
      RECT 42.175 2.615 42.185 2.765 ;
      RECT 41.995 2.615 42.035 2.768 ;
      RECT 41.909 2.615 41.995 2.776 ;
      RECT 41.823 2.615 41.909 2.787 ;
      RECT 41.737 2.615 41.823 2.798 ;
      RECT 41.651 2.615 41.737 2.809 ;
      RECT 41.565 2.615 41.651 2.82 ;
      RECT 41.535 2.615 41.565 2.86 ;
      RECT 41.505 2.615 41.535 2.91 ;
      RECT 41.43 2.615 41.505 2.93 ;
      RECT 41.425 2.59 41.43 2.935 ;
      RECT 41.41 2.585 41.425 2.943 ;
      RECT 41.405 1.205 41.41 2.953 ;
      RECT 41.375 1.205 41.405 2.995 ;
      RECT 41.355 1.205 41.375 3.075 ;
      RECT 40.485 2.965 40.505 3.404 ;
      RECT 40.485 2.965 40.591 3.401 ;
      RECT 40.475 3.08 40.591 3.4 ;
      RECT 40.505 2.115 40.635 3.397 ;
      RECT 40.485 2.985 40.645 3.395 ;
      RECT 40.485 3.07 40.655 3.39 ;
      RECT 40.455 3.115 40.655 3.385 ;
      RECT 40.455 3.115 40.665 3.38 ;
      RECT 40.435 3.115 40.695 3.375 ;
      RECT 40.505 2.115 40.665 2.765 ;
      RECT 40.495 2.115 40.665 2.74 ;
      RECT 40.495 2.115 40.685 2.505 ;
      RECT 40.445 2.115 40.705 2.375 ;
      RECT 39.915 2.605 40.205 2.865 ;
      RECT 39.925 2.585 40.205 2.865 ;
      RECT 39.875 2.665 40.205 2.86 ;
      RECT 39.945 2.578 40.115 2.865 ;
      RECT 39.945 2.565 40.071 2.865 ;
      RECT 39.985 2.558 40.071 2.865 ;
      RECT 39.445 3.705 39.725 3.985 ;
      RECT 39.405 3.67 39.705 3.78 ;
      RECT 39.395 3.62 39.685 3.675 ;
      RECT 39.335 3.385 39.595 3.645 ;
      RECT 39.335 3.525 39.675 3.645 ;
      RECT 39.335 3.475 39.655 3.645 ;
      RECT 39.335 3.43 39.645 3.645 ;
      RECT 39.335 3.415 39.615 3.645 ;
      RECT 35.07 6.225 35.39 6.545 ;
      RECT 35.1 5.695 35.27 6.545 ;
      RECT 35.1 5.695 35.275 6.045 ;
      RECT 35.1 5.695 36.075 5.87 ;
      RECT 35.9 1.965 36.075 5.87 ;
      RECT 35.845 1.965 36.195 2.315 ;
      RECT 35.87 6.655 36.195 6.98 ;
      RECT 34.755 6.745 36.195 6.915 ;
      RECT 34.755 2.395 34.915 6.915 ;
      RECT 35.07 2.365 35.39 2.685 ;
      RECT 34.755 2.395 35.39 2.565 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 25.345 0.96 25.72 1.33 ;
      RECT 23.91 0.96 24.285 1.33 ;
      RECT 23.91 1.08 33.73 1.25 ;
      RECT 28.03 4.36 33.71 4.53 ;
      RECT 33.54 3.425 33.71 4.53 ;
      RECT 27.84 3.595 27.86 4.53 ;
      RECT 28.09 3.705 28.12 3.985 ;
      RECT 27.8 3.595 27.86 3.855 ;
      RECT 33.45 3.43 33.8 3.78 ;
      RECT 27.63 2.225 27.66 2.485 ;
      RECT 27.4 2.225 27.46 2.485 ;
      RECT 28.08 3.685 28.09 3.985 ;
      RECT 28.06 3.605 28.08 3.985 ;
      RECT 28.05 3.545 28.06 3.985 ;
      RECT 28.03 3.495 28.05 3.985 ;
      RECT 28 3.395 28.03 4.53 ;
      RECT 27.99 3.305 28 4.53 ;
      RECT 27.95 3.245 27.99 4.53 ;
      RECT 27.946 3.214 27.95 4.53 ;
      RECT 27.86 3.205 27.946 4.53 ;
      RECT 27.85 3.196 27.86 3.55 ;
      RECT 27.82 3.175 27.85 3.517 ;
      RECT 27.81 3.125 27.82 3.493 ;
      RECT 27.8 3.09 27.81 3.481 ;
      RECT 27.76 3.015 27.8 3.45 ;
      RECT 27.74 2.925 27.76 3.415 ;
      RECT 27.73 2.866 27.74 3.4 ;
      RECT 27.68 2.756 27.73 3.36 ;
      RECT 27.67 2.65 27.68 3.315 ;
      RECT 27.64 2.579 27.67 3.235 ;
      RECT 27.63 2.511 27.64 3.16 ;
      RECT 27.62 2.225 27.63 3.125 ;
      RECT 27.59 2.225 27.62 3.055 ;
      RECT 27.58 2.225 27.59 2.95 ;
      RECT 27.57 2.225 27.58 2.915 ;
      RECT 27.5 2.225 27.57 2.775 ;
      RECT 27.47 2.225 27.5 2.575 ;
      RECT 27.46 2.225 27.47 2.5 ;
      RECT 31.8 2.155 32.06 2.415 ;
      RECT 31.79 2.155 32.06 2.365 ;
      RECT 31.76 2.025 32.04 2.305 ;
      RECT 20.325 6.655 20.675 7.005 ;
      RECT 31.295 6.61 31.645 6.96 ;
      RECT 20.325 6.685 31.645 6.885 ;
      RECT 30.8 3.705 31.08 3.985 ;
      RECT 30.84 3.665 31.11 3.925 ;
      RECT 30.83 3.7 31.11 3.925 ;
      RECT 30.84 3.66 31.05 3.985 ;
      RECT 30.84 3.655 31.04 3.985 ;
      RECT 30.88 3.645 31.04 3.985 ;
      RECT 30.85 3.65 31.04 3.985 ;
      RECT 30.89 3.64 30.98 3.985 ;
      RECT 30.91 3.635 30.98 3.985 ;
      RECT 30.22 3.155 30.48 3.415 ;
      RECT 30.27 3.065 30.46 3.415 ;
      RECT 30.3 2.85 30.46 3.415 ;
      RECT 30.39 2.455 30.46 3.415 ;
      RECT 30.41 2.165 30.546 2.893 ;
      RECT 30.35 2.66 30.546 2.893 ;
      RECT 30.37 2.54 30.46 3.415 ;
      RECT 30.41 2.165 30.57 2.558 ;
      RECT 30.41 2.165 30.58 2.455 ;
      RECT 30.4 2.165 30.66 2.425 ;
      RECT 29.8 3.705 30.08 3.985 ;
      RECT 29.82 3.665 30.08 3.985 ;
      RECT 29.46 3.625 29.57 3.885 ;
      RECT 29.32 2.115 29.41 2.375 ;
      RECT 29.85 3.17 29.86 3.3 ;
      RECT 29.84 3.135 29.85 3.454 ;
      RECT 29.76 3.067 29.84 3.534 ;
      RECT 29.79 3.71 29.8 3.93 ;
      RECT 29.77 3.705 29.79 3.919 ;
      RECT 29.74 3.7 29.77 3.904 ;
      RECT 29.75 3.002 29.76 3.61 ;
      RECT 29.73 2.946 29.75 3.625 ;
      RECT 29.72 3.685 29.74 3.89 ;
      RECT 29.72 2.874 29.73 3.645 ;
      RECT 29.69 2.777 29.72 3.885 ;
      RECT 29.67 2.66 29.69 3.885 ;
      RECT 29.64 2.54 29.67 3.885 ;
      RECT 29.63 2.455 29.64 3.885 ;
      RECT 29.62 2.4 29.63 3.885 ;
      RECT 29.61 2.355 29.62 3.104 ;
      RECT 29.6 3.315 29.62 3.885 ;
      RECT 29.6 2.285 29.61 3.061 ;
      RECT 29.58 2.235 29.6 2.996 ;
      RECT 29.59 3.395 29.6 3.885 ;
      RECT 29.57 3.495 29.59 3.885 ;
      RECT 29.52 2.115 29.58 2.824 ;
      RECT 29.51 2.115 29.52 2.66 ;
      RECT 29.5 2.115 29.51 2.61 ;
      RECT 29.45 2.115 29.5 2.54 ;
      RECT 29.43 2.115 29.45 2.455 ;
      RECT 29.41 2.115 29.43 2.41 ;
      RECT 28.73 3.565 28.78 3.825 ;
      RECT 28.64 2.095 28.78 2.355 ;
      RECT 29.14 2.72 29.15 2.808 ;
      RECT 29.13 2.655 29.14 2.854 ;
      RECT 29.12 2.605 29.13 2.9 ;
      RECT 29.07 2.552 29.12 3.039 ;
      RECT 29.06 2.501 29.07 3.23 ;
      RECT 29.02 2.459 29.06 3.335 ;
      RECT 29 2.405 29.02 3.472 ;
      RECT 28.99 2.38 29 2.688 ;
      RECT 28.99 2.77 29 3.542 ;
      RECT 28.98 2.366 28.99 2.673 ;
      RECT 28.98 2.825 28.99 3.825 ;
      RECT 28.96 2.341 28.98 2.655 ;
      RECT 28.94 3 28.98 3.825 ;
      RECT 28.95 2.315 28.96 2.635 ;
      RECT 28.92 2.28 28.95 2.589 ;
      RECT 28.93 3.125 28.94 3.825 ;
      RECT 28.92 3.205 28.93 3.825 ;
      RECT 28.91 2.245 28.92 2.554 ;
      RECT 28.87 3.275 28.92 3.825 ;
      RECT 28.9 2.225 28.91 2.53 ;
      RECT 28.87 2.095 28.9 2.495 ;
      RECT 28.86 2.095 28.87 2.46 ;
      RECT 28.84 3.375 28.87 3.825 ;
      RECT 28.84 2.095 28.86 2.435 ;
      RECT 28.83 2.095 28.84 2.41 ;
      RECT 28.79 3.475 28.84 3.825 ;
      RECT 28.81 2.095 28.83 2.38 ;
      RECT 28.78 2.095 28.81 2.365 ;
      RECT 28.78 3.55 28.79 3.825 ;
      RECT 28.7 2.635 28.74 2.895 ;
      RECT 24.43 2.055 24.69 2.315 ;
      RECT 24.43 2.085 24.71 2.295 ;
      RECT 26.64 1.905 26.82 2.055 ;
      RECT 28.69 2.63 28.7 2.895 ;
      RECT 28.67 2.62 28.69 2.895 ;
      RECT 28.652 2.613 28.67 2.895 ;
      RECT 28.566 2.602 28.652 2.895 ;
      RECT 28.48 2.585 28.566 2.895 ;
      RECT 28.43 2.572 28.48 2.82 ;
      RECT 28.396 2.564 28.43 2.795 ;
      RECT 28.31 2.553 28.396 2.76 ;
      RECT 28.27 2.53 28.31 2.723 ;
      RECT 28.26 2.495 28.27 2.708 ;
      RECT 28.25 2.455 28.26 2.703 ;
      RECT 28.24 2.435 28.25 2.698 ;
      RECT 28.225 2.395 28.24 2.693 ;
      RECT 28.21 2.347 28.225 2.689 ;
      RECT 28.2 2.306 28.21 2.686 ;
      RECT 28.19 2.268 28.2 2.675 ;
      RECT 28.17 2.212 28.19 2.655 ;
      RECT 28.15 2.16 28.17 2.591 ;
      RECT 28.13 2.11 28.15 2.543 ;
      RECT 28.12 2.08 28.13 2.507 ;
      RECT 28.115 2.062 28.12 2.493 ;
      RECT 28.1 2.053 28.115 2.475 ;
      RECT 28.07 2.034 28.1 2.415 ;
      RECT 28.06 2.017 28.07 2.37 ;
      RECT 28.05 2.009 28.06 2.34 ;
      RECT 28.02 1.997 28.05 2.29 ;
      RECT 28 1.985 28.02 2.225 ;
      RECT 27.99 1.977 28 2.185 ;
      RECT 27.97 1.974 27.99 2.175 ;
      RECT 27.955 1.972 27.97 2.17 ;
      RECT 27.935 1.971 27.955 2.16 ;
      RECT 27.92 1.97 27.935 2.15 ;
      RECT 27.9 1.969 27.92 2.145 ;
      RECT 27.898 1.969 27.9 2.145 ;
      RECT 27.812 1.966 27.898 2.142 ;
      RECT 27.726 1.961 27.812 2.135 ;
      RECT 27.64 1.956 27.726 2.129 ;
      RECT 27.59 1.953 27.64 2.12 ;
      RECT 27.546 1.951 27.59 2.114 ;
      RECT 27.46 1.947 27.546 2.109 ;
      RECT 27.456 1.945 27.46 2.105 ;
      RECT 27.37 1.942 27.456 2.1 ;
      RECT 27.316 1.938 27.37 2.093 ;
      RECT 27.23 1.935 27.316 2.088 ;
      RECT 27.206 1.932 27.23 2.084 ;
      RECT 27.12 1.93 27.206 2.079 ;
      RECT 27.06 1.926 27.12 2.073 ;
      RECT 27.052 1.924 27.06 2.07 ;
      RECT 26.966 1.92 27.052 2.066 ;
      RECT 26.88 1.913 26.966 2.059 ;
      RECT 26.82 1.907 26.88 2.055 ;
      RECT 26.62 1.905 26.64 2.058 ;
      RECT 26.57 1.915 26.62 2.068 ;
      RECT 26.54 1.925 26.57 2.08 ;
      RECT 26.516 1.927 26.54 2.086 ;
      RECT 26.43 1.93 26.516 2.091 ;
      RECT 26.36 1.935 26.43 2.1 ;
      RECT 26.346 1.937 26.36 2.106 ;
      RECT 26.26 1.941 26.346 2.111 ;
      RECT 26.22 1.945 26.26 2.12 ;
      RECT 26.206 1.947 26.22 2.126 ;
      RECT 26.12 1.951 26.206 2.131 ;
      RECT 26.036 1.957 26.12 2.138 ;
      RECT 25.95 1.963 26.036 2.143 ;
      RECT 25.926 1.967 25.95 2.146 ;
      RECT 25.84 1.971 25.926 2.151 ;
      RECT 25.79 1.976 25.84 2.16 ;
      RECT 25.71 1.981 25.79 2.17 ;
      RECT 25.63 1.987 25.71 2.185 ;
      RECT 25.61 1.991 25.63 2.195 ;
      RECT 25.54 1.994 25.61 2.205 ;
      RECT 25.49 1.999 25.54 2.22 ;
      RECT 25.46 2.002 25.49 2.24 ;
      RECT 25.45 2.004 25.46 2.256 ;
      RECT 25.39 2.016 25.45 2.266 ;
      RECT 25.37 2.031 25.39 2.275 ;
      RECT 25.36 2.05 25.37 2.275 ;
      RECT 25.35 2.07 25.36 2.275 ;
      RECT 25.33 2.08 25.35 2.275 ;
      RECT 25.28 2.09 25.33 2.275 ;
      RECT 25.25 2.096 25.28 2.275 ;
      RECT 25.18 2.101 25.25 2.277 ;
      RECT 25.1 2.102 25.18 2.282 ;
      RECT 25.096 2.1 25.1 2.285 ;
      RECT 25.01 2.097 25.096 2.286 ;
      RECT 24.968 2.094 25.01 2.288 ;
      RECT 24.882 2.092 24.968 2.289 ;
      RECT 24.796 2.089 24.882 2.292 ;
      RECT 24.71 2.086 24.796 2.294 ;
      RECT 26.64 3.145 26.92 3.425 ;
      RECT 26.67 3.125 26.94 3.385 ;
      RECT 26.67 3.075 26.9 3.425 ;
      RECT 26.74 3.065 26.9 3.425 ;
      RECT 26.74 2.775 26.89 3.425 ;
      RECT 26.73 2.455 26.88 2.825 ;
      RECT 26.72 2.455 26.88 2.695 ;
      RECT 26.7 2.165 26.87 2.5 ;
      RECT 26.68 2.165 26.87 2.45 ;
      RECT 26.64 2.165 26.9 2.425 ;
      RECT 26.55 3.635 26.63 3.895 ;
      RECT 25.84 2.355 25.96 2.615 ;
      RECT 26.525 3.615 26.55 3.895 ;
      RECT 26.51 3.577 26.525 3.895 ;
      RECT 26.47 3.52 26.51 3.895 ;
      RECT 26.44 3.43 26.47 3.895 ;
      RECT 26.4 3.33 26.44 3.895 ;
      RECT 26.37 3.23 26.4 3.895 ;
      RECT 26.365 3.177 26.37 3.718 ;
      RECT 26.35 3.147 26.365 3.684 ;
      RECT 26.34 3.108 26.35 3.649 ;
      RECT 26.33 3.075 26.34 3.605 ;
      RECT 26.32 3.042 26.33 3.57 ;
      RECT 26.29 2.976 26.32 3.505 ;
      RECT 26.28 2.911 26.29 3.43 ;
      RECT 26.27 2.881 26.28 3.4 ;
      RECT 26.23 2.811 26.27 3.33 ;
      RECT 26.22 2.746 26.23 3.245 ;
      RECT 26.21 2.728 26.22 3.23 ;
      RECT 26.2 2.711 26.21 3.195 ;
      RECT 26.19 2.694 26.2 3.165 ;
      RECT 26.18 2.677 26.19 3.135 ;
      RECT 26.16 2.652 26.18 3.075 ;
      RECT 26.15 2.626 26.16 3.02 ;
      RECT 26.13 2.601 26.15 2.98 ;
      RECT 26.12 2.57 26.13 2.945 ;
      RECT 26.11 2.557 26.12 2.9 ;
      RECT 26.1 2.542 26.11 2.875 ;
      RECT 26.09 2.355 26.1 2.835 ;
      RECT 26.08 2.355 26.09 2.805 ;
      RECT 26.075 2.355 26.08 2.788 ;
      RECT 26.07 2.355 26.075 2.77 ;
      RECT 26 2.355 26.07 2.71 ;
      RECT 25.96 2.355 26 2.645 ;
      RECT 25.79 3.225 26.05 3.485 ;
      RECT 23.96 3.145 24.04 3.465 ;
      RECT 23.78 3.205 23.93 3.465 ;
      RECT 23.96 3.145 24.07 3.425 ;
      RECT 25.78 3.317 25.79 3.48 ;
      RECT 25.75 3.327 25.78 3.488 ;
      RECT 25.73 3.335 25.75 3.493 ;
      RECT 25.662 3.343 25.73 3.503 ;
      RECT 25.576 3.363 25.662 3.52 ;
      RECT 25.49 3.384 25.576 3.539 ;
      RECT 25.48 3.4 25.49 3.55 ;
      RECT 25.44 3.41 25.48 3.556 ;
      RECT 25.42 3.415 25.44 3.563 ;
      RECT 25.382 3.416 25.42 3.566 ;
      RECT 25.296 3.419 25.382 3.567 ;
      RECT 25.21 3.423 25.296 3.568 ;
      RECT 25.156 3.425 25.21 3.57 ;
      RECT 25.07 3.425 25.156 3.572 ;
      RECT 25.03 3.42 25.07 3.574 ;
      RECT 25.02 3.414 25.03 3.575 ;
      RECT 24.98 3.409 25.02 3.571 ;
      RECT 24.97 3.4 24.98 3.567 ;
      RECT 24.938 3.391 24.97 3.564 ;
      RECT 24.852 3.379 24.938 3.554 ;
      RECT 24.766 3.362 24.852 3.539 ;
      RECT 24.68 3.344 24.766 3.525 ;
      RECT 24.66 3.335 24.68 3.516 ;
      RECT 24.59 3.325 24.66 3.509 ;
      RECT 24.54 3.31 24.59 3.499 ;
      RECT 24.48 3.3 24.54 3.49 ;
      RECT 24.44 3.29 24.48 3.485 ;
      RECT 24.39 3.28 24.44 3.479 ;
      RECT 24.35 3.268 24.39 3.469 ;
      RECT 24.33 3.258 24.35 3.465 ;
      RECT 24.31 3.248 24.33 3.465 ;
      RECT 24.3 3.238 24.31 3.464 ;
      RECT 24.28 3.23 24.3 3.46 ;
      RECT 24.24 3.205 24.28 3.454 ;
      RECT 24.22 3.145 24.24 3.447 ;
      RECT 24.196 3.145 24.22 3.444 ;
      RECT 24.11 3.145 24.196 3.439 ;
      RECT 24.07 3.145 24.11 3.43 ;
      RECT 23.93 3.195 23.96 3.465 ;
      RECT 25.61 2.775 25.87 3.035 ;
      RECT 25.57 2.775 25.87 2.915 ;
      RECT 25.54 2.775 25.87 2.9 ;
      RECT 25.48 2.775 25.87 2.88 ;
      RECT 25.4 2.585 25.68 2.865 ;
      RECT 25.4 2.77 25.75 2.865 ;
      RECT 25.4 2.71 25.74 2.865 ;
      RECT 25.4 2.66 25.69 2.865 ;
      RECT 23.17 3.115 23.43 3.375 ;
      RECT 23.315 1.205 23.43 3.375 ;
      RECT 23.23 2.585 23.43 3.375 ;
      RECT 24.54 2.635 24.8 2.895 ;
      RECT 23.225 2.585 23.43 2.87 ;
      RECT 23.22 2.585 23.43 2.865 ;
      RECT 24.52 2.645 24.8 2.825 ;
      RECT 24.11 2.615 24.25 2.765 ;
      RECT 23.485 1.205 23.565 1.55 ;
      RECT 23.22 1.205 23.43 1.55 ;
      RECT 24.51 2.644 24.52 2.825 ;
      RECT 24.506 2.644 24.51 2.825 ;
      RECT 24.42 2.639 24.506 2.814 ;
      RECT 24.346 2.63 24.42 2.794 ;
      RECT 24.26 2.621 24.346 2.775 ;
      RECT 24.25 2.615 24.26 2.765 ;
      RECT 24.07 2.615 24.11 2.768 ;
      RECT 23.984 2.615 24.07 2.776 ;
      RECT 23.898 2.615 23.984 2.787 ;
      RECT 23.812 2.615 23.898 2.798 ;
      RECT 23.726 2.615 23.812 2.809 ;
      RECT 23.64 2.615 23.726 2.82 ;
      RECT 23.61 2.615 23.64 2.86 ;
      RECT 23.58 2.615 23.61 2.91 ;
      RECT 23.505 2.615 23.58 2.93 ;
      RECT 23.5 2.59 23.505 2.935 ;
      RECT 23.485 2.585 23.5 2.943 ;
      RECT 23.48 1.205 23.485 2.953 ;
      RECT 23.45 1.205 23.48 2.995 ;
      RECT 23.43 1.205 23.45 3.075 ;
      RECT 22.56 2.965 22.58 3.404 ;
      RECT 22.56 2.965 22.666 3.401 ;
      RECT 22.55 3.08 22.666 3.4 ;
      RECT 22.58 2.115 22.71 3.397 ;
      RECT 22.56 2.985 22.72 3.395 ;
      RECT 22.56 3.07 22.73 3.39 ;
      RECT 22.53 3.115 22.73 3.385 ;
      RECT 22.53 3.115 22.74 3.38 ;
      RECT 22.51 3.115 22.77 3.375 ;
      RECT 22.58 2.115 22.74 2.765 ;
      RECT 22.57 2.115 22.74 2.74 ;
      RECT 22.57 2.115 22.76 2.505 ;
      RECT 22.52 2.115 22.78 2.375 ;
      RECT 21.99 2.605 22.28 2.865 ;
      RECT 22 2.585 22.28 2.865 ;
      RECT 21.95 2.665 22.28 2.86 ;
      RECT 22.02 2.578 22.19 2.865 ;
      RECT 22.02 2.565 22.146 2.865 ;
      RECT 22.06 2.558 22.146 2.865 ;
      RECT 21.52 3.705 21.8 3.985 ;
      RECT 21.48 3.67 21.78 3.78 ;
      RECT 21.47 3.62 21.76 3.675 ;
      RECT 21.41 3.385 21.67 3.645 ;
      RECT 21.41 3.525 21.75 3.645 ;
      RECT 21.41 3.475 21.73 3.645 ;
      RECT 21.41 3.43 21.72 3.645 ;
      RECT 21.41 3.415 21.69 3.645 ;
      RECT 17.145 6.225 17.465 6.545 ;
      RECT 17.175 5.695 17.345 6.545 ;
      RECT 17.175 5.695 17.35 6.045 ;
      RECT 17.175 5.695 18.15 5.87 ;
      RECT 17.975 1.965 18.15 5.87 ;
      RECT 17.92 1.965 18.27 2.315 ;
      RECT 17.945 6.655 18.27 6.98 ;
      RECT 16.83 6.745 18.27 6.915 ;
      RECT 16.83 2.395 16.99 6.915 ;
      RECT 17.145 2.365 17.465 2.685 ;
      RECT 16.83 2.395 17.465 2.565 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 7.42 0.96 7.795 1.33 ;
      RECT 5.985 0.96 6.36 1.33 ;
      RECT 5.985 1.08 15.805 1.25 ;
      RECT 10.105 4.36 15.785 4.53 ;
      RECT 15.615 3.425 15.785 4.53 ;
      RECT 9.915 3.595 9.935 4.53 ;
      RECT 10.165 3.705 10.195 3.985 ;
      RECT 9.875 3.595 9.935 3.855 ;
      RECT 15.525 3.43 15.875 3.78 ;
      RECT 9.705 2.225 9.735 2.485 ;
      RECT 9.475 2.225 9.535 2.485 ;
      RECT 10.155 3.685 10.165 3.985 ;
      RECT 10.135 3.605 10.155 3.985 ;
      RECT 10.125 3.545 10.135 3.985 ;
      RECT 10.105 3.495 10.125 3.985 ;
      RECT 10.075 3.395 10.105 4.53 ;
      RECT 10.065 3.305 10.075 4.53 ;
      RECT 10.025 3.245 10.065 4.53 ;
      RECT 10.021 3.214 10.025 4.53 ;
      RECT 9.935 3.205 10.021 4.53 ;
      RECT 9.925 3.196 9.935 3.55 ;
      RECT 9.895 3.175 9.925 3.517 ;
      RECT 9.885 3.125 9.895 3.493 ;
      RECT 9.875 3.09 9.885 3.481 ;
      RECT 9.835 3.015 9.875 3.45 ;
      RECT 9.815 2.925 9.835 3.415 ;
      RECT 9.805 2.866 9.815 3.4 ;
      RECT 9.755 2.756 9.805 3.36 ;
      RECT 9.745 2.65 9.755 3.315 ;
      RECT 9.715 2.579 9.745 3.235 ;
      RECT 9.705 2.511 9.715 3.16 ;
      RECT 9.695 2.225 9.705 3.125 ;
      RECT 9.665 2.225 9.695 3.055 ;
      RECT 9.655 2.225 9.665 2.95 ;
      RECT 9.645 2.225 9.655 2.915 ;
      RECT 9.575 2.225 9.645 2.775 ;
      RECT 9.545 2.225 9.575 2.575 ;
      RECT 9.535 2.225 9.545 2.5 ;
      RECT 13.875 2.155 14.135 2.415 ;
      RECT 13.865 2.155 14.135 2.365 ;
      RECT 13.835 2.025 14.115 2.305 ;
      RECT 1.7 6.995 1.99 7.345 ;
      RECT 1.7 7.055 3.01 7.225 ;
      RECT 2.84 6.685 3.01 7.225 ;
      RECT 13.34 6.605 13.69 6.955 ;
      RECT 2.84 6.685 13.69 6.855 ;
      RECT 12.875 3.705 13.155 3.985 ;
      RECT 12.915 3.665 13.185 3.925 ;
      RECT 12.905 3.7 13.185 3.925 ;
      RECT 12.915 3.66 13.125 3.985 ;
      RECT 12.915 3.655 13.115 3.985 ;
      RECT 12.955 3.645 13.115 3.985 ;
      RECT 12.925 3.65 13.115 3.985 ;
      RECT 12.965 3.64 13.055 3.985 ;
      RECT 12.985 3.635 13.055 3.985 ;
      RECT 12.295 3.155 12.555 3.415 ;
      RECT 12.345 3.065 12.535 3.415 ;
      RECT 12.375 2.85 12.535 3.415 ;
      RECT 12.465 2.455 12.535 3.415 ;
      RECT 12.485 2.165 12.621 2.893 ;
      RECT 12.425 2.66 12.621 2.893 ;
      RECT 12.445 2.54 12.535 3.415 ;
      RECT 12.485 2.165 12.645 2.558 ;
      RECT 12.485 2.165 12.655 2.455 ;
      RECT 12.475 2.165 12.735 2.425 ;
      RECT 11.875 3.705 12.155 3.985 ;
      RECT 11.895 3.665 12.155 3.985 ;
      RECT 11.535 3.625 11.645 3.885 ;
      RECT 11.395 2.115 11.485 2.375 ;
      RECT 11.925 3.17 11.935 3.3 ;
      RECT 11.915 3.135 11.925 3.454 ;
      RECT 11.835 3.067 11.915 3.534 ;
      RECT 11.865 3.71 11.875 3.93 ;
      RECT 11.845 3.705 11.865 3.919 ;
      RECT 11.815 3.7 11.845 3.904 ;
      RECT 11.825 3.002 11.835 3.61 ;
      RECT 11.805 2.946 11.825 3.625 ;
      RECT 11.795 3.685 11.815 3.89 ;
      RECT 11.795 2.874 11.805 3.645 ;
      RECT 11.765 2.777 11.795 3.885 ;
      RECT 11.745 2.66 11.765 3.885 ;
      RECT 11.715 2.54 11.745 3.885 ;
      RECT 11.705 2.455 11.715 3.885 ;
      RECT 11.695 2.4 11.705 3.885 ;
      RECT 11.685 2.355 11.695 3.104 ;
      RECT 11.675 3.315 11.695 3.885 ;
      RECT 11.675 2.285 11.685 3.061 ;
      RECT 11.655 2.235 11.675 2.996 ;
      RECT 11.665 3.395 11.675 3.885 ;
      RECT 11.645 3.495 11.665 3.885 ;
      RECT 11.595 2.115 11.655 2.824 ;
      RECT 11.585 2.115 11.595 2.66 ;
      RECT 11.575 2.115 11.585 2.61 ;
      RECT 11.525 2.115 11.575 2.54 ;
      RECT 11.505 2.115 11.525 2.455 ;
      RECT 11.485 2.115 11.505 2.41 ;
      RECT 10.805 3.565 10.855 3.825 ;
      RECT 10.715 2.095 10.855 2.355 ;
      RECT 11.215 2.72 11.225 2.808 ;
      RECT 11.205 2.655 11.215 2.854 ;
      RECT 11.195 2.605 11.205 2.9 ;
      RECT 11.145 2.552 11.195 3.039 ;
      RECT 11.135 2.501 11.145 3.23 ;
      RECT 11.095 2.459 11.135 3.335 ;
      RECT 11.075 2.405 11.095 3.472 ;
      RECT 11.065 2.38 11.075 2.688 ;
      RECT 11.065 2.77 11.075 3.542 ;
      RECT 11.055 2.366 11.065 2.673 ;
      RECT 11.055 2.825 11.065 3.825 ;
      RECT 11.035 2.341 11.055 2.655 ;
      RECT 11.015 3 11.055 3.825 ;
      RECT 11.025 2.315 11.035 2.635 ;
      RECT 10.995 2.28 11.025 2.589 ;
      RECT 11.005 3.125 11.015 3.825 ;
      RECT 10.995 3.205 11.005 3.825 ;
      RECT 10.985 2.245 10.995 2.554 ;
      RECT 10.945 3.275 10.995 3.825 ;
      RECT 10.975 2.225 10.985 2.53 ;
      RECT 10.945 2.095 10.975 2.495 ;
      RECT 10.935 2.095 10.945 2.46 ;
      RECT 10.915 3.375 10.945 3.825 ;
      RECT 10.915 2.095 10.935 2.435 ;
      RECT 10.905 2.095 10.915 2.41 ;
      RECT 10.865 3.475 10.915 3.825 ;
      RECT 10.885 2.095 10.905 2.38 ;
      RECT 10.855 2.095 10.885 2.365 ;
      RECT 10.855 3.55 10.865 3.825 ;
      RECT 10.775 2.635 10.815 2.895 ;
      RECT 6.505 2.055 6.765 2.315 ;
      RECT 6.505 2.085 6.785 2.295 ;
      RECT 8.715 1.905 8.895 2.055 ;
      RECT 10.765 2.63 10.775 2.895 ;
      RECT 10.745 2.62 10.765 2.895 ;
      RECT 10.727 2.613 10.745 2.895 ;
      RECT 10.641 2.602 10.727 2.895 ;
      RECT 10.555 2.585 10.641 2.895 ;
      RECT 10.505 2.572 10.555 2.82 ;
      RECT 10.471 2.564 10.505 2.795 ;
      RECT 10.385 2.553 10.471 2.76 ;
      RECT 10.345 2.53 10.385 2.723 ;
      RECT 10.335 2.495 10.345 2.708 ;
      RECT 10.325 2.455 10.335 2.703 ;
      RECT 10.315 2.435 10.325 2.698 ;
      RECT 10.3 2.395 10.315 2.693 ;
      RECT 10.285 2.347 10.3 2.689 ;
      RECT 10.275 2.306 10.285 2.686 ;
      RECT 10.265 2.268 10.275 2.675 ;
      RECT 10.245 2.212 10.265 2.655 ;
      RECT 10.225 2.16 10.245 2.591 ;
      RECT 10.205 2.11 10.225 2.543 ;
      RECT 10.195 2.08 10.205 2.507 ;
      RECT 10.19 2.062 10.195 2.493 ;
      RECT 10.175 2.053 10.19 2.475 ;
      RECT 10.145 2.034 10.175 2.415 ;
      RECT 10.135 2.017 10.145 2.37 ;
      RECT 10.125 2.009 10.135 2.34 ;
      RECT 10.095 1.997 10.125 2.29 ;
      RECT 10.075 1.985 10.095 2.225 ;
      RECT 10.065 1.977 10.075 2.185 ;
      RECT 10.045 1.974 10.065 2.175 ;
      RECT 10.03 1.972 10.045 2.17 ;
      RECT 10.01 1.971 10.03 2.16 ;
      RECT 9.995 1.97 10.01 2.15 ;
      RECT 9.975 1.969 9.995 2.145 ;
      RECT 9.973 1.969 9.975 2.145 ;
      RECT 9.887 1.966 9.973 2.142 ;
      RECT 9.801 1.961 9.887 2.135 ;
      RECT 9.715 1.956 9.801 2.129 ;
      RECT 9.665 1.953 9.715 2.12 ;
      RECT 9.621 1.951 9.665 2.114 ;
      RECT 9.535 1.947 9.621 2.109 ;
      RECT 9.531 1.945 9.535 2.105 ;
      RECT 9.445 1.942 9.531 2.1 ;
      RECT 9.391 1.938 9.445 2.093 ;
      RECT 9.305 1.935 9.391 2.088 ;
      RECT 9.281 1.932 9.305 2.084 ;
      RECT 9.195 1.93 9.281 2.079 ;
      RECT 9.135 1.926 9.195 2.073 ;
      RECT 9.127 1.924 9.135 2.07 ;
      RECT 9.041 1.92 9.127 2.066 ;
      RECT 8.955 1.913 9.041 2.059 ;
      RECT 8.895 1.907 8.955 2.055 ;
      RECT 8.695 1.905 8.715 2.058 ;
      RECT 8.645 1.915 8.695 2.068 ;
      RECT 8.615 1.925 8.645 2.08 ;
      RECT 8.591 1.927 8.615 2.086 ;
      RECT 8.505 1.93 8.591 2.091 ;
      RECT 8.435 1.935 8.505 2.1 ;
      RECT 8.421 1.937 8.435 2.106 ;
      RECT 8.335 1.941 8.421 2.111 ;
      RECT 8.295 1.945 8.335 2.12 ;
      RECT 8.281 1.947 8.295 2.126 ;
      RECT 8.195 1.951 8.281 2.131 ;
      RECT 8.111 1.957 8.195 2.138 ;
      RECT 8.025 1.963 8.111 2.143 ;
      RECT 8.001 1.967 8.025 2.146 ;
      RECT 7.915 1.971 8.001 2.151 ;
      RECT 7.865 1.976 7.915 2.16 ;
      RECT 7.785 1.981 7.865 2.17 ;
      RECT 7.705 1.987 7.785 2.185 ;
      RECT 7.685 1.991 7.705 2.195 ;
      RECT 7.615 1.994 7.685 2.205 ;
      RECT 7.565 1.999 7.615 2.22 ;
      RECT 7.535 2.002 7.565 2.24 ;
      RECT 7.525 2.004 7.535 2.256 ;
      RECT 7.465 2.016 7.525 2.266 ;
      RECT 7.445 2.031 7.465 2.275 ;
      RECT 7.435 2.05 7.445 2.275 ;
      RECT 7.425 2.07 7.435 2.275 ;
      RECT 7.405 2.08 7.425 2.275 ;
      RECT 7.355 2.09 7.405 2.275 ;
      RECT 7.325 2.096 7.355 2.275 ;
      RECT 7.255 2.101 7.325 2.277 ;
      RECT 7.175 2.102 7.255 2.282 ;
      RECT 7.171 2.1 7.175 2.285 ;
      RECT 7.085 2.097 7.171 2.286 ;
      RECT 7.043 2.094 7.085 2.288 ;
      RECT 6.957 2.092 7.043 2.289 ;
      RECT 6.871 2.089 6.957 2.292 ;
      RECT 6.785 2.086 6.871 2.294 ;
      RECT 8.715 3.145 8.995 3.425 ;
      RECT 8.745 3.125 9.015 3.385 ;
      RECT 8.745 3.075 8.975 3.425 ;
      RECT 8.815 3.065 8.975 3.425 ;
      RECT 8.815 2.775 8.965 3.425 ;
      RECT 8.805 2.455 8.955 2.825 ;
      RECT 8.795 2.455 8.955 2.695 ;
      RECT 8.775 2.165 8.945 2.5 ;
      RECT 8.755 2.165 8.945 2.45 ;
      RECT 8.715 2.165 8.975 2.425 ;
      RECT 8.625 3.635 8.705 3.895 ;
      RECT 7.915 2.355 8.035 2.615 ;
      RECT 8.6 3.615 8.625 3.895 ;
      RECT 8.585 3.577 8.6 3.895 ;
      RECT 8.545 3.52 8.585 3.895 ;
      RECT 8.515 3.43 8.545 3.895 ;
      RECT 8.475 3.33 8.515 3.895 ;
      RECT 8.445 3.23 8.475 3.895 ;
      RECT 8.44 3.177 8.445 3.718 ;
      RECT 8.425 3.147 8.44 3.684 ;
      RECT 8.415 3.108 8.425 3.649 ;
      RECT 8.405 3.075 8.415 3.605 ;
      RECT 8.395 3.042 8.405 3.57 ;
      RECT 8.365 2.976 8.395 3.505 ;
      RECT 8.355 2.911 8.365 3.43 ;
      RECT 8.345 2.881 8.355 3.4 ;
      RECT 8.305 2.811 8.345 3.33 ;
      RECT 8.295 2.746 8.305 3.245 ;
      RECT 8.285 2.728 8.295 3.23 ;
      RECT 8.275 2.711 8.285 3.195 ;
      RECT 8.265 2.694 8.275 3.165 ;
      RECT 8.255 2.677 8.265 3.135 ;
      RECT 8.235 2.652 8.255 3.075 ;
      RECT 8.225 2.626 8.235 3.02 ;
      RECT 8.205 2.601 8.225 2.98 ;
      RECT 8.195 2.57 8.205 2.945 ;
      RECT 8.185 2.557 8.195 2.9 ;
      RECT 8.175 2.542 8.185 2.875 ;
      RECT 8.165 2.355 8.175 2.835 ;
      RECT 8.155 2.355 8.165 2.805 ;
      RECT 8.15 2.355 8.155 2.788 ;
      RECT 8.145 2.355 8.15 2.77 ;
      RECT 8.075 2.355 8.145 2.71 ;
      RECT 8.035 2.355 8.075 2.645 ;
      RECT 7.865 3.225 8.125 3.485 ;
      RECT 6.035 3.145 6.115 3.465 ;
      RECT 5.855 3.205 6.005 3.465 ;
      RECT 6.035 3.145 6.145 3.425 ;
      RECT 7.855 3.317 7.865 3.48 ;
      RECT 7.825 3.327 7.855 3.488 ;
      RECT 7.805 3.335 7.825 3.493 ;
      RECT 7.737 3.343 7.805 3.503 ;
      RECT 7.651 3.363 7.737 3.52 ;
      RECT 7.565 3.384 7.651 3.539 ;
      RECT 7.555 3.4 7.565 3.55 ;
      RECT 7.515 3.41 7.555 3.556 ;
      RECT 7.495 3.415 7.515 3.563 ;
      RECT 7.457 3.416 7.495 3.566 ;
      RECT 7.371 3.419 7.457 3.567 ;
      RECT 7.285 3.423 7.371 3.568 ;
      RECT 7.231 3.425 7.285 3.57 ;
      RECT 7.145 3.425 7.231 3.572 ;
      RECT 7.105 3.42 7.145 3.574 ;
      RECT 7.095 3.414 7.105 3.575 ;
      RECT 7.055 3.409 7.095 3.571 ;
      RECT 7.045 3.4 7.055 3.567 ;
      RECT 7.013 3.391 7.045 3.564 ;
      RECT 6.927 3.379 7.013 3.554 ;
      RECT 6.841 3.362 6.927 3.539 ;
      RECT 6.755 3.344 6.841 3.525 ;
      RECT 6.735 3.335 6.755 3.516 ;
      RECT 6.665 3.325 6.735 3.509 ;
      RECT 6.615 3.31 6.665 3.499 ;
      RECT 6.555 3.3 6.615 3.49 ;
      RECT 6.515 3.29 6.555 3.485 ;
      RECT 6.465 3.28 6.515 3.479 ;
      RECT 6.425 3.268 6.465 3.469 ;
      RECT 6.405 3.258 6.425 3.465 ;
      RECT 6.385 3.248 6.405 3.465 ;
      RECT 6.375 3.238 6.385 3.464 ;
      RECT 6.355 3.23 6.375 3.46 ;
      RECT 6.315 3.205 6.355 3.454 ;
      RECT 6.295 3.145 6.315 3.447 ;
      RECT 6.271 3.145 6.295 3.444 ;
      RECT 6.185 3.145 6.271 3.439 ;
      RECT 6.145 3.145 6.185 3.43 ;
      RECT 6.005 3.195 6.035 3.465 ;
      RECT 7.685 2.775 7.945 3.035 ;
      RECT 7.645 2.775 7.945 2.915 ;
      RECT 7.615 2.775 7.945 2.9 ;
      RECT 7.555 2.775 7.945 2.88 ;
      RECT 7.475 2.585 7.755 2.865 ;
      RECT 7.475 2.77 7.825 2.865 ;
      RECT 7.475 2.71 7.815 2.865 ;
      RECT 7.475 2.66 7.765 2.865 ;
      RECT 5.245 3.115 5.505 3.375 ;
      RECT 5.39 1.205 5.505 3.375 ;
      RECT 5.305 2.585 5.505 3.375 ;
      RECT 6.615 2.635 6.875 2.895 ;
      RECT 5.3 2.585 5.505 2.87 ;
      RECT 5.295 2.585 5.505 2.865 ;
      RECT 6.595 2.645 6.875 2.825 ;
      RECT 6.185 2.615 6.325 2.765 ;
      RECT 5.56 1.205 5.64 1.55 ;
      RECT 5.295 1.205 5.505 1.55 ;
      RECT 6.585 2.644 6.595 2.825 ;
      RECT 6.581 2.644 6.585 2.825 ;
      RECT 6.495 2.639 6.581 2.814 ;
      RECT 6.421 2.63 6.495 2.794 ;
      RECT 6.335 2.621 6.421 2.775 ;
      RECT 6.325 2.615 6.335 2.765 ;
      RECT 6.145 2.615 6.185 2.768 ;
      RECT 6.059 2.615 6.145 2.776 ;
      RECT 5.973 2.615 6.059 2.787 ;
      RECT 5.887 2.615 5.973 2.798 ;
      RECT 5.801 2.615 5.887 2.809 ;
      RECT 5.715 2.615 5.801 2.82 ;
      RECT 5.685 2.615 5.715 2.86 ;
      RECT 5.655 2.615 5.685 2.91 ;
      RECT 5.58 2.615 5.655 2.93 ;
      RECT 5.575 2.59 5.58 2.935 ;
      RECT 5.56 2.585 5.575 2.943 ;
      RECT 5.555 1.205 5.56 2.953 ;
      RECT 5.525 1.205 5.555 2.995 ;
      RECT 5.505 1.205 5.525 3.075 ;
      RECT 4.635 2.965 4.655 3.404 ;
      RECT 4.635 2.965 4.741 3.401 ;
      RECT 4.625 3.08 4.741 3.4 ;
      RECT 4.655 2.115 4.785 3.397 ;
      RECT 4.635 2.985 4.795 3.395 ;
      RECT 4.635 3.07 4.805 3.39 ;
      RECT 4.605 3.115 4.805 3.385 ;
      RECT 4.605 3.115 4.815 3.38 ;
      RECT 4.585 3.115 4.845 3.375 ;
      RECT 4.655 2.115 4.815 2.765 ;
      RECT 4.645 2.115 4.815 2.74 ;
      RECT 4.645 2.115 4.835 2.505 ;
      RECT 4.595 2.115 4.855 2.375 ;
      RECT 4.065 2.605 4.355 2.865 ;
      RECT 4.075 2.585 4.355 2.865 ;
      RECT 4.025 2.665 4.355 2.86 ;
      RECT 4.095 2.578 4.265 2.865 ;
      RECT 4.095 2.565 4.221 2.865 ;
      RECT 4.135 2.558 4.221 2.865 ;
      RECT 3.595 3.705 3.875 3.985 ;
      RECT 3.555 3.67 3.855 3.78 ;
      RECT 3.545 3.62 3.835 3.675 ;
      RECT 3.485 3.385 3.745 3.645 ;
      RECT 3.485 3.525 3.825 3.645 ;
      RECT 3.485 3.475 3.805 3.645 ;
      RECT 3.485 3.43 3.795 3.645 ;
      RECT 3.485 3.415 3.765 3.645 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 75.715 0.93 76.09 1.3 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 57.79 0.93 58.165 1.3 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 39.865 0.93 40.24 1.3 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 21.94 0.93 22.315 1.3 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 4.015 0.93 4.39 1.3 ;
      RECT 0.215 8.5 0.595 8.88 ;
    LAYER via1 ;
      RECT 92.1 7.375 92.25 7.525 ;
      RECT 89.735 6.74 89.885 6.89 ;
      RECT 89.72 2.065 89.87 2.215 ;
      RECT 88.93 2.45 89.08 2.6 ;
      RECT 88.93 6.325 89.08 6.475 ;
      RECT 87.325 3.53 87.475 3.68 ;
      RECT 87.315 1.25 87.465 1.4 ;
      RECT 85.63 2.21 85.78 2.36 ;
      RECT 85.4 6.71 85.55 6.86 ;
      RECT 84.68 3.72 84.83 3.87 ;
      RECT 84.495 7.165 84.645 7.315 ;
      RECT 84.23 2.22 84.38 2.37 ;
      RECT 84.05 3.21 84.2 3.36 ;
      RECT 83.65 3.72 83.8 3.87 ;
      RECT 83.29 3.68 83.44 3.83 ;
      RECT 83.15 2.17 83.3 2.32 ;
      RECT 82.56 3.62 82.71 3.77 ;
      RECT 82.47 2.15 82.62 2.3 ;
      RECT 82.31 2.69 82.46 2.84 ;
      RECT 81.63 3.65 81.78 3.8 ;
      RECT 81.23 2.28 81.38 2.43 ;
      RECT 80.51 3.18 80.66 3.33 ;
      RECT 80.47 2.22 80.62 2.37 ;
      RECT 80.2 3.69 80.35 3.84 ;
      RECT 79.67 2.41 79.82 2.56 ;
      RECT 79.62 3.28 79.77 3.43 ;
      RECT 79.44 2.83 79.59 2.98 ;
      RECT 78.37 2.69 78.52 2.84 ;
      RECT 78.26 2.11 78.41 2.26 ;
      RECT 77.61 3.26 77.76 3.41 ;
      RECT 77.09 1.3 77.24 1.45 ;
      RECT 77 3.17 77.15 3.32 ;
      RECT 76.35 2.17 76.5 2.32 ;
      RECT 76.34 3.17 76.49 3.32 ;
      RECT 75.82 2.66 75.97 2.81 ;
      RECT 75.24 3.44 75.39 3.59 ;
      RECT 74.155 6.755 74.305 6.905 ;
      RECT 71.81 6.74 71.96 6.89 ;
      RECT 71.795 2.065 71.945 2.215 ;
      RECT 71.005 2.45 71.155 2.6 ;
      RECT 71.005 6.325 71.155 6.475 ;
      RECT 69.4 3.53 69.55 3.68 ;
      RECT 69.39 1.25 69.54 1.4 ;
      RECT 67.705 2.21 67.855 2.36 ;
      RECT 67.195 6.71 67.345 6.86 ;
      RECT 66.755 3.72 66.905 3.87 ;
      RECT 66.57 7.165 66.72 7.315 ;
      RECT 66.305 2.22 66.455 2.37 ;
      RECT 66.125 3.21 66.275 3.36 ;
      RECT 65.725 3.72 65.875 3.87 ;
      RECT 65.365 3.68 65.515 3.83 ;
      RECT 65.225 2.17 65.375 2.32 ;
      RECT 64.635 3.62 64.785 3.77 ;
      RECT 64.545 2.15 64.695 2.3 ;
      RECT 64.385 2.69 64.535 2.84 ;
      RECT 63.705 3.65 63.855 3.8 ;
      RECT 63.305 2.28 63.455 2.43 ;
      RECT 62.585 3.18 62.735 3.33 ;
      RECT 62.545 2.22 62.695 2.37 ;
      RECT 62.275 3.69 62.425 3.84 ;
      RECT 61.745 2.41 61.895 2.56 ;
      RECT 61.695 3.28 61.845 3.43 ;
      RECT 61.515 2.83 61.665 2.98 ;
      RECT 60.445 2.69 60.595 2.84 ;
      RECT 60.335 2.11 60.485 2.26 ;
      RECT 59.685 3.26 59.835 3.41 ;
      RECT 59.165 1.3 59.315 1.45 ;
      RECT 59.075 3.17 59.225 3.32 ;
      RECT 58.425 2.17 58.575 2.32 ;
      RECT 58.415 3.17 58.565 3.32 ;
      RECT 57.895 2.66 58.045 2.81 ;
      RECT 57.315 3.44 57.465 3.59 ;
      RECT 56.23 6.755 56.38 6.905 ;
      RECT 53.885 6.74 54.035 6.89 ;
      RECT 53.87 2.065 54.02 2.215 ;
      RECT 53.08 2.45 53.23 2.6 ;
      RECT 53.08 6.325 53.23 6.475 ;
      RECT 51.475 3.53 51.625 3.68 ;
      RECT 51.465 1.25 51.615 1.4 ;
      RECT 49.78 2.21 49.93 2.36 ;
      RECT 49.325 6.715 49.475 6.865 ;
      RECT 48.83 3.72 48.98 3.87 ;
      RECT 48.645 7.165 48.795 7.315 ;
      RECT 48.38 2.22 48.53 2.37 ;
      RECT 48.2 3.21 48.35 3.36 ;
      RECT 47.8 3.72 47.95 3.87 ;
      RECT 47.44 3.68 47.59 3.83 ;
      RECT 47.3 2.17 47.45 2.32 ;
      RECT 46.71 3.62 46.86 3.77 ;
      RECT 46.62 2.15 46.77 2.3 ;
      RECT 46.46 2.69 46.61 2.84 ;
      RECT 45.78 3.65 45.93 3.8 ;
      RECT 45.38 2.28 45.53 2.43 ;
      RECT 44.66 3.18 44.81 3.33 ;
      RECT 44.62 2.22 44.77 2.37 ;
      RECT 44.35 3.69 44.5 3.84 ;
      RECT 43.82 2.41 43.97 2.56 ;
      RECT 43.77 3.28 43.92 3.43 ;
      RECT 43.59 2.83 43.74 2.98 ;
      RECT 42.52 2.69 42.67 2.84 ;
      RECT 42.41 2.11 42.56 2.26 ;
      RECT 41.76 3.26 41.91 3.41 ;
      RECT 41.24 1.3 41.39 1.45 ;
      RECT 41.15 3.17 41.3 3.32 ;
      RECT 40.5 2.17 40.65 2.32 ;
      RECT 40.49 3.17 40.64 3.32 ;
      RECT 39.97 2.66 40.12 2.81 ;
      RECT 39.39 3.44 39.54 3.59 ;
      RECT 38.35 6.76 38.5 6.91 ;
      RECT 35.96 6.74 36.11 6.89 ;
      RECT 35.945 2.065 36.095 2.215 ;
      RECT 35.155 2.45 35.305 2.6 ;
      RECT 35.155 6.325 35.305 6.475 ;
      RECT 33.55 3.53 33.7 3.68 ;
      RECT 33.54 1.25 33.69 1.4 ;
      RECT 31.855 2.21 32.005 2.36 ;
      RECT 31.395 6.71 31.545 6.86 ;
      RECT 30.905 3.72 31.055 3.87 ;
      RECT 30.72 7.165 30.87 7.315 ;
      RECT 30.455 2.22 30.605 2.37 ;
      RECT 30.275 3.21 30.425 3.36 ;
      RECT 29.875 3.72 30.025 3.87 ;
      RECT 29.515 3.68 29.665 3.83 ;
      RECT 29.375 2.17 29.525 2.32 ;
      RECT 28.785 3.62 28.935 3.77 ;
      RECT 28.695 2.15 28.845 2.3 ;
      RECT 28.535 2.69 28.685 2.84 ;
      RECT 27.855 3.65 28.005 3.8 ;
      RECT 27.455 2.28 27.605 2.43 ;
      RECT 26.735 3.18 26.885 3.33 ;
      RECT 26.695 2.22 26.845 2.37 ;
      RECT 26.425 3.69 26.575 3.84 ;
      RECT 25.895 2.41 26.045 2.56 ;
      RECT 25.845 3.28 25.995 3.43 ;
      RECT 25.665 2.83 25.815 2.98 ;
      RECT 24.595 2.69 24.745 2.84 ;
      RECT 24.485 2.11 24.635 2.26 ;
      RECT 23.835 3.26 23.985 3.41 ;
      RECT 23.315 1.3 23.465 1.45 ;
      RECT 23.225 3.17 23.375 3.32 ;
      RECT 22.575 2.17 22.725 2.32 ;
      RECT 22.565 3.17 22.715 3.32 ;
      RECT 22.045 2.66 22.195 2.81 ;
      RECT 21.465 3.44 21.615 3.59 ;
      RECT 20.425 6.755 20.575 6.905 ;
      RECT 18.035 6.74 18.185 6.89 ;
      RECT 18.02 2.065 18.17 2.215 ;
      RECT 17.23 2.45 17.38 2.6 ;
      RECT 17.23 6.325 17.38 6.475 ;
      RECT 15.625 3.53 15.775 3.68 ;
      RECT 15.615 1.25 15.765 1.4 ;
      RECT 13.93 2.21 14.08 2.36 ;
      RECT 13.44 6.705 13.59 6.855 ;
      RECT 12.98 3.72 13.13 3.87 ;
      RECT 12.795 7.165 12.945 7.315 ;
      RECT 12.53 2.22 12.68 2.37 ;
      RECT 12.35 3.21 12.5 3.36 ;
      RECT 11.95 3.72 12.1 3.87 ;
      RECT 11.59 3.68 11.74 3.83 ;
      RECT 11.45 2.17 11.6 2.32 ;
      RECT 10.86 3.62 11.01 3.77 ;
      RECT 10.77 2.15 10.92 2.3 ;
      RECT 10.61 2.69 10.76 2.84 ;
      RECT 9.93 3.65 10.08 3.8 ;
      RECT 9.53 2.28 9.68 2.43 ;
      RECT 8.81 3.18 8.96 3.33 ;
      RECT 8.77 2.22 8.92 2.37 ;
      RECT 8.5 3.69 8.65 3.84 ;
      RECT 7.97 2.41 8.12 2.56 ;
      RECT 7.92 3.28 8.07 3.43 ;
      RECT 7.74 2.83 7.89 2.98 ;
      RECT 6.67 2.69 6.82 2.84 ;
      RECT 6.56 2.11 6.71 2.26 ;
      RECT 5.91 3.26 6.06 3.41 ;
      RECT 5.39 1.3 5.54 1.45 ;
      RECT 5.3 3.17 5.45 3.32 ;
      RECT 4.65 2.17 4.8 2.32 ;
      RECT 4.64 3.17 4.79 3.32 ;
      RECT 4.12 2.66 4.27 2.81 ;
      RECT 3.54 3.44 3.69 3.59 ;
      RECT 1.77 7.095 1.92 7.245 ;
      RECT 1.395 6.355 1.545 6.505 ;
      RECT 0.33 8.615 0.48 8.765 ;
    LAYER met1 ;
      RECT 75.025 1.285 86.985 1.885 ;
      RECT 79.45 0 86.985 1.885 ;
      RECT 57.1 1.285 69.06 1.885 ;
      RECT 61.525 0 69.06 1.885 ;
      RECT 39.175 1.285 51.135 1.885 ;
      RECT 43.6 0 51.135 1.885 ;
      RECT 21.25 1.285 33.21 1.885 ;
      RECT 25.675 0 33.21 1.885 ;
      RECT 3.325 1.285 15.285 1.885 ;
      RECT 7.75 0 15.285 1.885 ;
      RECT 75.02 0 75.765 1.68 ;
      RECT 57.095 0 57.84 1.68 ;
      RECT 39.17 0 39.915 1.68 ;
      RECT 21.245 0 21.99 1.68 ;
      RECT 3.32 0 4.065 1.68 ;
      RECT 78.015 0 79.17 1.885 ;
      RECT 75.02 1.255 77.735 1.68 ;
      RECT 76.045 0 77.735 1.885 ;
      RECT 60.09 0 61.245 1.885 ;
      RECT 57.095 1.255 59.81 1.68 ;
      RECT 58.12 0 59.81 1.885 ;
      RECT 42.165 0 43.32 1.885 ;
      RECT 39.17 1.255 41.885 1.68 ;
      RECT 40.195 0 41.885 1.885 ;
      RECT 24.24 0 25.395 1.885 ;
      RECT 21.245 1.255 23.96 1.68 ;
      RECT 22.27 0 23.96 1.885 ;
      RECT 6.315 0 7.47 1.885 ;
      RECT 3.32 1.255 6.035 1.68 ;
      RECT 4.345 0 6.035 1.885 ;
      RECT 76.045 0 86.985 1.005 ;
      RECT 58.12 0 69.06 1.005 ;
      RECT 40.195 0 51.135 1.005 ;
      RECT 22.27 0 33.21 1.005 ;
      RECT 4.345 0 15.285 1.005 ;
      RECT 75.02 0 86.985 0.975 ;
      RECT 57.095 0 69.06 0.975 ;
      RECT 39.17 0 51.135 0.975 ;
      RECT 21.245 0 33.21 0.975 ;
      RECT 3.32 0 15.285 0.975 ;
      RECT 92.395 0 92.575 0.305 ;
      RECT 74.47 0 90.445 0.305 ;
      RECT 56.545 0 72.52 0.305 ;
      RECT 38.62 0 54.595 0.305 ;
      RECT 20.695 0 36.67 0.305 ;
      RECT 0 0 18.745 0.305 ;
      RECT 0 0 92.575 0.3 ;
      RECT 0.025 8.58 92.575 8.88 ;
      RECT 92.395 8.575 92.575 8.88 ;
      RECT 74.47 8.575 90.445 8.88 ;
      RECT 56.545 8.575 72.52 8.88 ;
      RECT 38.62 8.575 54.595 8.88 ;
      RECT 20.695 8.575 36.67 8.88 ;
      RECT 0.025 8.575 18.745 8.88 ;
      RECT 83.72 6.315 83.89 8.88 ;
      RECT 65.795 6.315 65.965 8.88 ;
      RECT 47.87 6.315 48.04 8.88 ;
      RECT 29.945 6.315 30.115 8.88 ;
      RECT 12.02 6.315 12.19 8.88 ;
      RECT 0.025 8.565 0.83 8.88 ;
      RECT 0.23 8.545 0.58 8.88 ;
      RECT 84.055 6.285 84.345 6.515 ;
      RECT 66.13 6.285 66.42 6.515 ;
      RECT 48.205 6.285 48.495 6.515 ;
      RECT 30.28 6.285 30.57 6.515 ;
      RECT 12.355 6.285 12.645 6.515 ;
      RECT 83.72 6.315 84.345 6.485 ;
      RECT 65.795 6.315 66.42 6.485 ;
      RECT 47.87 6.315 48.495 6.485 ;
      RECT 29.945 6.315 30.57 6.485 ;
      RECT 12.02 6.315 12.645 6.485 ;
      RECT 91.97 7.77 92.26 8 ;
      RECT 92.03 6.29 92.2 8 ;
      RECT 92 7.275 92.35 7.625 ;
      RECT 91.97 6.29 92.26 6.52 ;
      RECT 91.565 2.395 91.67 2.965 ;
      RECT 91.565 2.73 91.89 2.96 ;
      RECT 91.565 2.76 92.06 2.93 ;
      RECT 91.565 2.395 91.755 2.96 ;
      RECT 90.98 2.36 91.27 2.59 ;
      RECT 90.98 2.395 91.755 2.565 ;
      RECT 91.04 0.88 91.21 2.59 ;
      RECT 90.98 0.88 91.27 1.11 ;
      RECT 90.98 7.77 91.27 8 ;
      RECT 91.04 6.29 91.21 8 ;
      RECT 90.98 6.29 91.27 6.52 ;
      RECT 90.98 6.325 91.835 6.485 ;
      RECT 91.665 5.92 91.835 6.485 ;
      RECT 90.98 6.32 91.375 6.485 ;
      RECT 91.6 5.92 91.89 6.15 ;
      RECT 91.6 5.95 92.06 6.12 ;
      RECT 90.61 2.73 90.9 2.96 ;
      RECT 90.61 2.76 91.07 2.93 ;
      RECT 90.675 1.655 90.84 2.96 ;
      RECT 89.19 1.625 89.48 1.855 ;
      RECT 89.19 1.655 90.84 1.825 ;
      RECT 89.25 0.885 89.42 1.855 ;
      RECT 89.19 0.885 89.48 1.115 ;
      RECT 89.19 7.765 89.48 7.995 ;
      RECT 89.25 7.025 89.42 7.995 ;
      RECT 89.25 7.12 90.84 7.29 ;
      RECT 90.67 5.92 90.84 7.29 ;
      RECT 89.19 7.025 89.48 7.255 ;
      RECT 90.61 5.92 90.9 6.15 ;
      RECT 90.61 5.95 91.07 6.12 ;
      RECT 87.225 3.43 87.575 3.78 ;
      RECT 87.315 2.025 87.485 3.78 ;
      RECT 89.62 1.965 89.97 2.315 ;
      RECT 87.315 2.025 88.935 2.2 ;
      RECT 87.315 2.025 89.97 2.195 ;
      RECT 89.645 6.655 89.97 6.98 ;
      RECT 85.3 6.61 85.65 6.96 ;
      RECT 89.62 6.655 89.97 6.885 ;
      RECT 84.86 6.655 85.15 6.885 ;
      RECT 84.69 6.685 89.97 6.855 ;
      RECT 88.845 2.365 89.165 2.685 ;
      RECT 88.815 2.365 89.165 2.595 ;
      RECT 88.645 2.395 89.165 2.565 ;
      RECT 88.845 6.225 89.165 6.545 ;
      RECT 88.815 6.285 89.165 6.515 ;
      RECT 88.645 6.315 89.165 6.485 ;
      RECT 84.685 3.255 84.875 3.925 ;
      RECT 84.625 3.665 84.665 3.925 ;
      RECT 85.995 2.89 86.005 3.111 ;
      RECT 85.925 2.885 85.995 3.236 ;
      RECT 85.915 2.885 85.925 3.36 ;
      RECT 85.885 2.885 85.915 3.41 ;
      RECT 85.865 2.885 85.885 3.485 ;
      RECT 85.845 2.885 85.865 3.555 ;
      RECT 85.815 2.885 85.845 3.595 ;
      RECT 85.805 2.885 85.815 3.615 ;
      RECT 85.795 2.885 85.805 3.626 ;
      RECT 85.785 3.135 85.795 3.628 ;
      RECT 85.775 3.2 85.785 3.63 ;
      RECT 85.765 3.295 85.775 3.632 ;
      RECT 85.755 3.37 85.765 3.634 ;
      RECT 85.705 3.394 85.755 3.64 ;
      RECT 85.665 3.429 85.705 3.649 ;
      RECT 85.655 3.445 85.665 3.654 ;
      RECT 85.641 3.45 85.655 3.657 ;
      RECT 85.555 3.49 85.641 3.668 ;
      RECT 85.475 3.533 85.555 3.686 ;
      RECT 85.455 3.543 85.475 3.697 ;
      RECT 85.425 3.551 85.455 3.702 ;
      RECT 85.405 3.561 85.425 3.707 ;
      RECT 85.381 3.567 85.405 3.712 ;
      RECT 85.295 3.577 85.381 3.725 ;
      RECT 85.217 3.583 85.295 3.745 ;
      RECT 85.131 3.578 85.217 3.764 ;
      RECT 85.045 3.574 85.131 3.785 ;
      RECT 84.965 3.57 85.045 3.8 ;
      RECT 84.895 3.566 84.965 3.831 ;
      RECT 84.885 3.277 84.895 3.345 ;
      RECT 84.885 3.555 84.895 3.861 ;
      RECT 84.875 3.262 84.885 3.49 ;
      RECT 84.875 3.535 84.885 3.925 ;
      RECT 84.665 3.285 84.685 3.925 ;
      RECT 85.465 2.605 85.475 3.345 ;
      RECT 85.285 3.125 85.305 3.345 ;
      RECT 85.295 3.115 85.305 3.345 ;
      RECT 85.795 2.155 85.835 2.415 ;
      RECT 85.785 2.155 85.795 2.425 ;
      RECT 85.751 2.155 85.785 2.452 ;
      RECT 85.665 2.155 85.751 2.512 ;
      RECT 85.645 2.155 85.665 2.575 ;
      RECT 85.585 2.155 85.645 2.74 ;
      RECT 85.575 2.155 85.585 2.9 ;
      RECT 85.545 2.346 85.575 2.995 ;
      RECT 85.535 2.401 85.545 3.095 ;
      RECT 85.525 2.43 85.535 3.14 ;
      RECT 85.515 2.455 85.525 3.173 ;
      RECT 85.505 2.49 85.515 3.228 ;
      RECT 85.485 2.535 85.505 3.29 ;
      RECT 85.475 2.58 85.485 3.34 ;
      RECT 85.455 2.64 85.465 3.345 ;
      RECT 85.445 2.67 85.455 3.345 ;
      RECT 85.425 2.7 85.445 3.345 ;
      RECT 85.375 2.805 85.425 3.345 ;
      RECT 85.365 2.9 85.375 3.345 ;
      RECT 85.355 2.93 85.365 3.345 ;
      RECT 85.33 2.98 85.355 3.345 ;
      RECT 85.325 3.035 85.33 3.345 ;
      RECT 85.305 3.06 85.325 3.345 ;
      RECT 85.265 3.14 85.285 3.335 ;
      RECT 85.015 2.725 85.085 2.935 ;
      RECT 82.255 2.635 82.515 2.895 ;
      RECT 85.085 2.73 85.095 2.93 ;
      RECT 84.971 2.723 85.015 2.935 ;
      RECT 84.885 2.716 84.971 2.935 ;
      RECT 84.865 2.711 84.885 2.925 ;
      RECT 84.855 2.709 84.865 2.905 ;
      RECT 84.805 2.706 84.855 2.9 ;
      RECT 84.775 2.702 84.805 2.895 ;
      RECT 84.755 2.7 84.775 2.89 ;
      RECT 84.715 2.697 84.755 2.885 ;
      RECT 84.645 2.691 84.715 2.88 ;
      RECT 84.615 2.686 84.645 2.875 ;
      RECT 84.595 2.684 84.615 2.87 ;
      RECT 84.565 2.681 84.595 2.865 ;
      RECT 84.505 2.677 84.565 2.86 ;
      RECT 84.435 2.675 84.505 2.85 ;
      RECT 84.401 2.673 84.435 2.843 ;
      RECT 84.315 2.668 84.401 2.835 ;
      RECT 84.281 2.662 84.315 2.827 ;
      RECT 84.195 2.652 84.281 2.819 ;
      RECT 84.161 2.643 84.195 2.811 ;
      RECT 84.075 2.638 84.161 2.803 ;
      RECT 84.005 2.635 84.075 2.793 ;
      RECT 83.985 2.63 84.005 2.787 ;
      RECT 83.981 2.625 83.985 2.786 ;
      RECT 83.895 2.621 83.981 2.781 ;
      RECT 83.855 2.616 83.895 2.774 ;
      RECT 83.775 2.615 83.855 2.769 ;
      RECT 83.755 2.615 83.775 2.766 ;
      RECT 83.729 2.615 83.755 2.766 ;
      RECT 83.643 2.617 83.729 2.77 ;
      RECT 83.557 2.619 83.643 2.777 ;
      RECT 83.471 2.621 83.557 2.783 ;
      RECT 83.385 2.624 83.471 2.79 ;
      RECT 83.351 2.626 83.385 2.795 ;
      RECT 83.265 2.631 83.351 2.8 ;
      RECT 83.241 2.626 83.265 2.804 ;
      RECT 83.155 2.631 83.241 2.809 ;
      RECT 83.117 2.636 83.155 2.814 ;
      RECT 83.031 2.639 83.117 2.819 ;
      RECT 82.945 2.643 83.031 2.826 ;
      RECT 82.881 2.645 82.945 2.832 ;
      RECT 82.795 2.645 82.881 2.838 ;
      RECT 82.711 2.646 82.795 2.845 ;
      RECT 82.625 2.649 82.711 2.852 ;
      RECT 82.601 2.651 82.625 2.856 ;
      RECT 82.515 2.653 82.601 2.861 ;
      RECT 82.245 2.67 82.255 2.865 ;
      RECT 84.43 7.765 84.72 7.995 ;
      RECT 84.49 7.025 84.66 7.995 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 84.43 7.025 84.72 7.425 ;
      RECT 84.485 2.247 84.675 2.455 ;
      RECT 84.475 2.252 84.685 2.45 ;
      RECT 84.465 2.233 84.475 2.445 ;
      RECT 84.435 2.228 84.465 2.44 ;
      RECT 84.395 2.252 84.685 2.43 ;
      RECT 84.175 2.165 84.435 2.425 ;
      RECT 84.475 2.236 84.485 2.45 ;
      RECT 84.175 2.245 84.665 2.425 ;
      RECT 84.175 2.241 84.525 2.425 ;
      RECT 84.125 3.155 84.175 3.435 ;
      RECT 84.055 3.125 84.085 3.435 ;
      RECT 84.195 3.155 84.255 3.415 ;
      RECT 84.055 3.115 84.075 3.435 ;
      RECT 84.175 3.155 84.195 3.425 ;
      RECT 84.095 3.145 84.125 3.435 ;
      RECT 84.085 3.13 84.095 3.435 ;
      RECT 84.035 3.105 84.055 3.435 ;
      RECT 84.005 3.09 84.035 3.435 ;
      RECT 83.995 3.08 84.005 3.435 ;
      RECT 83.975 3.069 83.995 3.43 ;
      RECT 83.955 3.057 83.975 3.4 ;
      RECT 83.945 3.048 83.955 3.383 ;
      RECT 83.915 3.03 83.945 3.375 ;
      RECT 83.905 2.995 83.915 3.367 ;
      RECT 83.895 2.975 83.905 3.36 ;
      RECT 83.885 2.955 83.895 3.353 ;
      RECT 83.875 2.94 83.885 3.348 ;
      RECT 83.865 2.92 83.875 3.343 ;
      RECT 83.855 2.915 83.865 3.338 ;
      RECT 83.851 2.905 83.855 3.334 ;
      RECT 83.765 2.905 83.851 3.309 ;
      RECT 83.735 2.905 83.765 3.275 ;
      RECT 83.725 2.905 83.735 3.255 ;
      RECT 83.665 2.905 83.725 3.2 ;
      RECT 83.655 2.92 83.665 3.145 ;
      RECT 83.645 2.93 83.655 3.125 ;
      RECT 83.595 3.665 83.855 3.925 ;
      RECT 83.515 3.685 83.855 3.901 ;
      RECT 83.495 3.685 83.855 3.896 ;
      RECT 83.471 3.685 83.855 3.894 ;
      RECT 83.385 3.685 83.855 3.889 ;
      RECT 83.235 3.625 83.495 3.885 ;
      RECT 83.195 3.68 83.515 3.88 ;
      RECT 83.185 3.69 83.855 3.875 ;
      RECT 83.205 3.675 83.495 3.885 ;
      RECT 83.095 2.115 83.355 2.375 ;
      RECT 83.095 2.2 83.365 2.3 ;
      RECT 82.265 3.63 82.285 3.874 ;
      RECT 82.265 3.63 82.335 3.869 ;
      RECT 82.245 3.635 82.335 3.868 ;
      RECT 82.235 3.65 82.421 3.858 ;
      RECT 82.235 3.65 82.495 3.855 ;
      RECT 82.23 3.687 82.505 3.845 ;
      RECT 82.23 3.687 82.591 3.841 ;
      RECT 82.23 3.687 82.605 3.827 ;
      RECT 82.505 3.565 82.765 3.825 ;
      RECT 82.225 3.692 82.765 3.82 ;
      RECT 82.215 3.74 82.765 3.795 ;
      RECT 82.485 3.605 82.505 3.854 ;
      RECT 82.421 3.609 82.485 3.857 ;
      RECT 82.285 3.622 82.765 3.825 ;
      RECT 82.335 3.616 82.421 3.862 ;
      RECT 81.735 2.475 81.745 2.645 ;
      RECT 81.795 2.435 81.805 2.615 ;
      RECT 82.095 2.245 82.105 2.455 ;
      RECT 82.425 2.095 82.675 2.355 ;
      RECT 82.415 2.095 82.425 2.357 ;
      RECT 82.405 2.155 82.415 2.361 ;
      RECT 82.375 2.157 82.405 2.369 ;
      RECT 82.345 2.162 82.375 2.383 ;
      RECT 82.335 2.166 82.345 2.393 ;
      RECT 82.305 2.171 82.335 2.405 ;
      RECT 82.275 2.18 82.305 2.406 ;
      RECT 82.205 2.19 82.275 2.41 ;
      RECT 82.165 2.195 82.205 2.414 ;
      RECT 82.145 2.195 82.165 2.425 ;
      RECT 82.135 2.2 82.145 2.435 ;
      RECT 82.125 2.21 82.135 2.438 ;
      RECT 82.115 2.23 82.125 2.443 ;
      RECT 82.105 2.24 82.115 2.445 ;
      RECT 82.075 2.255 82.095 2.462 ;
      RECT 82.065 2.267 82.075 2.472 ;
      RECT 82.055 2.273 82.065 2.475 ;
      RECT 82.021 2.286 82.055 2.485 ;
      RECT 81.935 2.32 82.021 2.518 ;
      RECT 81.915 2.355 81.935 2.547 ;
      RECT 81.895 2.37 81.915 2.559 ;
      RECT 81.875 2.38 81.895 2.571 ;
      RECT 81.825 2.399 81.875 2.591 ;
      RECT 81.815 2.416 81.825 2.605 ;
      RECT 81.805 2.422 81.815 2.61 ;
      RECT 81.785 2.44 81.795 2.618 ;
      RECT 81.775 2.445 81.785 2.625 ;
      RECT 81.765 2.456 81.775 2.632 ;
      RECT 81.745 2.461 81.765 2.64 ;
      RECT 81.725 2.475 81.735 2.65 ;
      RECT 81.715 2.48 81.725 2.66 ;
      RECT 81.685 2.494 81.715 2.67 ;
      RECT 81.675 2.507 81.685 2.68 ;
      RECT 81.595 2.538 81.675 2.705 ;
      RECT 81.575 2.568 81.595 2.73 ;
      RECT 81.565 2.573 81.575 2.737 ;
      RECT 81.535 2.585 81.565 2.743 ;
      RECT 81.525 2.6 81.535 2.749 ;
      RECT 81.515 2.605 81.525 2.752 ;
      RECT 81.495 2.615 81.515 2.756 ;
      RECT 81.475 2.62 81.495 2.762 ;
      RECT 81.445 2.625 81.475 2.77 ;
      RECT 81.415 2.63 81.445 2.78 ;
      RECT 81.385 2.64 81.415 2.789 ;
      RECT 81.345 2.645 81.385 2.797 ;
      RECT 81.295 2.638 81.345 2.809 ;
      RECT 81.275 2.629 81.295 2.82 ;
      RECT 81.265 2.626 81.275 2.825 ;
      RECT 81.225 2.625 81.265 2.826 ;
      RECT 81.215 2.61 81.225 2.827 ;
      RECT 81.187 2.595 81.215 2.828 ;
      RECT 81.101 2.595 81.187 2.83 ;
      RECT 81.015 2.595 81.101 2.834 ;
      RECT 80.995 2.595 81.015 2.83 ;
      RECT 80.985 2.605 80.995 2.823 ;
      RECT 80.975 2.62 80.985 2.818 ;
      RECT 80.965 2.625 80.975 2.795 ;
      RECT 82.445 3.13 82.455 3.33 ;
      RECT 82.395 3.125 82.445 3.35 ;
      RECT 82.385 3.125 82.395 3.37 ;
      RECT 82.341 3.125 82.385 3.374 ;
      RECT 82.255 3.125 82.341 3.371 ;
      RECT 82.195 3.135 82.255 3.368 ;
      RECT 82.135 3.149 82.195 3.366 ;
      RECT 82.125 3.154 82.135 3.364 ;
      RECT 82.115 3.16 82.125 3.363 ;
      RECT 82.045 3.173 82.115 3.359 ;
      RECT 81.997 3.187 82.045 3.36 ;
      RECT 81.911 3.203 81.997 3.372 ;
      RECT 81.825 3.224 81.911 3.388 ;
      RECT 81.805 3.235 81.825 3.398 ;
      RECT 81.725 3.245 81.805 3.408 ;
      RECT 81.691 3.259 81.725 3.42 ;
      RECT 81.605 3.274 81.691 3.435 ;
      RECT 81.575 3.29 81.605 3.445 ;
      RECT 81.52 3.305 81.575 3.456 ;
      RECT 81.475 3.323 81.52 3.476 ;
      RECT 81.421 3.342 81.475 3.496 ;
      RECT 81.335 3.368 81.421 3.523 ;
      RECT 81.315 3.39 81.335 3.543 ;
      RECT 81.255 3.405 81.315 3.559 ;
      RECT 81.245 3.42 81.255 3.573 ;
      RECT 81.225 3.425 81.245 3.579 ;
      RECT 81.195 3.438 81.225 3.589 ;
      RECT 81.175 3.443 81.195 3.598 ;
      RECT 81.165 3.45 81.175 3.603 ;
      RECT 81.155 3.455 81.165 3.606 ;
      RECT 81.115 3.465 81.155 3.615 ;
      RECT 81.09 3.48 81.115 3.627 ;
      RECT 81.045 3.495 81.09 3.639 ;
      RECT 81.025 3.507 81.045 3.651 ;
      RECT 80.995 3.512 81.025 3.661 ;
      RECT 80.975 3.519 80.995 3.671 ;
      RECT 80.965 3.525 80.975 3.68 ;
      RECT 80.941 3.532 80.965 3.69 ;
      RECT 80.855 3.554 80.941 3.71 ;
      RECT 80.845 3.573 80.855 3.725 ;
      RECT 80.821 3.58 80.845 3.731 ;
      RECT 80.735 3.602 80.821 3.756 ;
      RECT 80.695 3.627 80.735 3.783 ;
      RECT 80.685 3.636 80.695 3.793 ;
      RECT 80.635 3.646 80.685 3.802 ;
      RECT 80.615 3.66 80.635 3.812 ;
      RECT 80.585 3.67 80.615 3.817 ;
      RECT 80.575 3.675 80.585 3.82 ;
      RECT 80.501 3.677 80.575 3.827 ;
      RECT 80.415 3.681 80.501 3.839 ;
      RECT 80.405 3.684 80.415 3.845 ;
      RECT 80.145 3.635 80.405 3.895 ;
      RECT 81.675 3.705 81.865 3.915 ;
      RECT 81.665 3.71 81.875 3.91 ;
      RECT 81.655 3.71 81.875 3.875 ;
      RECT 81.575 3.595 81.835 3.855 ;
      RECT 80.485 3.125 80.675 3.425 ;
      RECT 80.475 3.125 80.675 3.42 ;
      RECT 80.465 3.125 80.685 3.415 ;
      RECT 80.455 3.125 80.685 3.41 ;
      RECT 80.455 3.125 80.715 3.385 ;
      RECT 80.415 2.165 80.675 2.425 ;
      RECT 80.225 2.09 80.311 2.423 ;
      RECT 80.225 2.09 80.355 2.419 ;
      RECT 80.205 2.094 80.365 2.418 ;
      RECT 80.355 2.085 80.365 2.418 ;
      RECT 80.225 2.09 80.375 2.417 ;
      RECT 80.205 2.1 80.415 2.416 ;
      RECT 80.195 2.095 80.375 2.408 ;
      RECT 80.185 2.11 80.415 2.315 ;
      RECT 80.185 2.16 80.615 2.315 ;
      RECT 80.185 2.15 80.595 2.315 ;
      RECT 80.185 2.14 80.565 2.315 ;
      RECT 80.185 2.13 80.505 2.315 ;
      RECT 80.185 2.115 80.485 2.315 ;
      RECT 80.311 2.086 80.365 2.418 ;
      RECT 79.385 2.745 79.525 3.035 ;
      RECT 79.645 2.768 79.655 2.955 ;
      RECT 80.345 2.665 80.525 2.895 ;
      RECT 80.345 2.665 80.535 2.885 ;
      RECT 80.555 2.67 80.565 2.875 ;
      RECT 80.535 2.665 80.555 2.88 ;
      RECT 80.295 2.669 80.345 2.895 ;
      RECT 80.285 2.674 80.295 2.895 ;
      RECT 80.251 2.679 80.285 2.896 ;
      RECT 80.165 2.694 80.251 2.898 ;
      RECT 80.151 2.706 80.165 2.901 ;
      RECT 80.065 2.716 80.151 2.903 ;
      RECT 80.041 2.726 80.065 2.905 ;
      RECT 79.955 2.737 80.041 2.905 ;
      RECT 79.925 2.747 79.955 2.905 ;
      RECT 79.895 2.752 79.925 2.908 ;
      RECT 79.875 2.757 79.895 2.913 ;
      RECT 79.855 2.762 79.875 2.915 ;
      RECT 79.805 2.77 79.855 2.915 ;
      RECT 79.785 2.774 79.805 2.915 ;
      RECT 79.765 2.773 79.785 2.92 ;
      RECT 79.705 2.771 79.765 2.935 ;
      RECT 79.655 2.769 79.705 2.95 ;
      RECT 79.565 2.766 79.645 3.035 ;
      RECT 79.535 2.76 79.565 3.035 ;
      RECT 79.525 2.75 79.535 3.035 ;
      RECT 79.335 2.745 79.385 2.96 ;
      RECT 79.325 2.75 79.335 2.95 ;
      RECT 79.565 3.225 79.825 3.485 ;
      RECT 79.565 3.225 79.855 3.375 ;
      RECT 79.565 3.225 79.895 3.36 ;
      RECT 79.825 3.145 80.015 3.355 ;
      RECT 79.825 3.15 80.025 3.345 ;
      RECT 79.775 3.22 80.025 3.345 ;
      RECT 79.805 3.155 79.825 3.485 ;
      RECT 79.795 3.18 80.025 3.345 ;
      RECT 78.975 3.125 78.985 3.355 ;
      RECT 78.875 2.245 78.945 3.355 ;
      RECT 79.615 2.355 79.875 2.615 ;
      RECT 79.315 2.405 79.445 2.565 ;
      RECT 79.531 2.412 79.615 2.565 ;
      RECT 79.445 2.407 79.531 2.565 ;
      RECT 79.255 2.405 79.315 2.575 ;
      RECT 79.225 2.403 79.255 2.59 ;
      RECT 79.205 2.401 79.225 2.6 ;
      RECT 79.195 2.399 79.205 2.605 ;
      RECT 79.175 2.398 79.195 2.615 ;
      RECT 79.165 2.396 79.175 2.62 ;
      RECT 79.145 2.395 79.165 2.625 ;
      RECT 79.125 2.39 79.145 2.63 ;
      RECT 79.095 2.376 79.125 2.64 ;
      RECT 79.055 2.355 79.095 2.655 ;
      RECT 79.045 2.34 79.055 2.665 ;
      RECT 79.025 2.331 79.045 2.675 ;
      RECT 79.015 2.322 79.025 2.695 ;
      RECT 79.005 2.317 79.015 2.755 ;
      RECT 78.985 2.311 79.005 2.84 ;
      RECT 78.985 3.15 78.995 3.35 ;
      RECT 78.975 2.306 78.985 3.07 ;
      RECT 78.965 2.28 78.975 3.355 ;
      RECT 78.945 2.25 78.965 3.355 ;
      RECT 78.855 2.245 78.875 2.58 ;
      RECT 78.865 2.68 78.875 3.355 ;
      RECT 78.855 2.72 78.865 3.355 ;
      RECT 78.825 2.245 78.855 2.525 ;
      RECT 78.835 2.81 78.855 3.355 ;
      RECT 78.82 2.915 78.835 3.355 ;
      RECT 78.795 2.245 78.825 2.48 ;
      RECT 78.815 2.947 78.82 3.355 ;
      RECT 78.795 3.05 78.815 3.355 ;
      RECT 78.785 2.245 78.795 2.47 ;
      RECT 78.785 3.12 78.795 3.35 ;
      RECT 78.765 2.245 78.785 2.46 ;
      RECT 78.755 2.25 78.765 2.45 ;
      RECT 78.965 3.525 78.985 3.765 ;
      RECT 78.285 3.455 78.365 3.725 ;
      RECT 78.195 3.455 78.205 3.665 ;
      RECT 79.475 3.525 79.485 3.725 ;
      RECT 79.395 3.515 79.475 3.75 ;
      RECT 79.391 3.515 79.395 3.776 ;
      RECT 79.305 3.515 79.391 3.786 ;
      RECT 79.285 3.515 79.305 3.794 ;
      RECT 79.261 3.516 79.285 3.792 ;
      RECT 79.175 3.521 79.261 3.787 ;
      RECT 79.157 3.525 79.175 3.781 ;
      RECT 79.071 3.525 79.157 3.777 ;
      RECT 78.985 3.525 79.071 3.769 ;
      RECT 78.881 3.525 78.965 3.762 ;
      RECT 78.795 3.525 78.881 3.756 ;
      RECT 78.735 3.52 78.795 3.75 ;
      RECT 78.707 3.514 78.735 3.747 ;
      RECT 78.621 3.511 78.707 3.744 ;
      RECT 78.535 3.507 78.621 3.738 ;
      RECT 78.49 3.495 78.535 3.734 ;
      RECT 78.465 3.48 78.49 3.732 ;
      RECT 78.425 3.465 78.465 3.73 ;
      RECT 78.365 3.455 78.425 3.727 ;
      RECT 78.275 3.455 78.285 3.72 ;
      RECT 78.26 3.455 78.275 3.71 ;
      RECT 78.205 3.455 78.26 3.685 ;
      RECT 78.185 3.47 78.195 3.66 ;
      RECT 78.315 2.635 78.575 2.895 ;
      RECT 78.315 2.645 78.595 2.855 ;
      RECT 78.315 2.65 78.605 2.85 ;
      RECT 76.295 2.115 76.555 2.375 ;
      RECT 76.285 2.145 76.555 2.355 ;
      RECT 78.215 2.055 78.465 2.315 ;
      RECT 78.205 2.055 78.215 2.316 ;
      RECT 78.175 2.14 78.205 2.318 ;
      RECT 78.165 2.145 78.175 2.32 ;
      RECT 78.105 2.16 78.165 2.326 ;
      RECT 78.075 2.18 78.105 2.333 ;
      RECT 78.045 2.191 78.075 2.34 ;
      RECT 78.025 2.201 78.045 2.345 ;
      RECT 78.007 2.204 78.025 2.344 ;
      RECT 77.921 2.203 78.007 2.344 ;
      RECT 77.835 2.2 77.921 2.343 ;
      RECT 77.749 2.197 77.835 2.342 ;
      RECT 77.663 2.194 77.749 2.342 ;
      RECT 77.577 2.192 77.663 2.341 ;
      RECT 77.491 2.189 77.577 2.34 ;
      RECT 77.405 2.186 77.491 2.34 ;
      RECT 77.387 2.185 77.405 2.339 ;
      RECT 77.301 2.184 77.387 2.339 ;
      RECT 77.215 2.182 77.301 2.338 ;
      RECT 77.129 2.181 77.215 2.338 ;
      RECT 77.043 2.18 77.129 2.337 ;
      RECT 76.957 2.178 77.043 2.337 ;
      RECT 76.871 2.177 76.957 2.336 ;
      RECT 76.785 2.175 76.871 2.336 ;
      RECT 76.761 2.174 76.785 2.335 ;
      RECT 76.675 2.169 76.761 2.335 ;
      RECT 76.641 2.162 76.675 2.335 ;
      RECT 76.555 2.152 76.641 2.335 ;
      RECT 76.275 2.15 76.285 2.35 ;
      RECT 77.555 3.205 77.815 3.465 ;
      RECT 77.555 3.205 77.895 3.251 ;
      RECT 77.695 3.185 77.905 3.24 ;
      RECT 77.755 3.16 77.965 3.2 ;
      RECT 77.765 3.155 77.965 3.2 ;
      RECT 77.775 3.13 77.965 3.2 ;
      RECT 77.835 2.96 77.885 3.29 ;
      RECT 77.785 3.09 77.975 3.15 ;
      RECT 77.825 3.016 77.835 3.329 ;
      RECT 77.785 3.09 78.005 3.125 ;
      RECT 77.785 3.09 78.025 3.1 ;
      RECT 77.895 2.89 78.085 3.095 ;
      RECT 77.885 2.9 78.095 3.09 ;
      RECT 77.805 3.063 78.095 3.09 ;
      RECT 77.815 3.039 77.825 3.345 ;
      RECT 77.905 2.885 78.075 3.095 ;
      RECT 77.195 2.675 77.385 2.885 ;
      RECT 75.765 2.605 76.025 2.865 ;
      RECT 76.115 2.595 76.215 2.805 ;
      RECT 76.065 2.615 76.105 2.805 ;
      RECT 77.385 2.685 77.395 2.88 ;
      RECT 77.185 2.685 77.195 2.88 ;
      RECT 77.165 2.7 77.185 2.87 ;
      RECT 77.155 2.71 77.165 2.865 ;
      RECT 77.115 2.71 77.155 2.863 ;
      RECT 77.091 2.704 77.115 2.86 ;
      RECT 77.005 2.699 77.091 2.857 ;
      RECT 76.945 2.695 77.005 2.852 ;
      RECT 76.911 2.692 76.945 2.849 ;
      RECT 76.825 2.682 76.911 2.845 ;
      RECT 76.821 2.675 76.825 2.842 ;
      RECT 76.735 2.67 76.821 2.84 ;
      RECT 76.707 2.663 76.735 2.836 ;
      RECT 76.621 2.658 76.707 2.833 ;
      RECT 76.535 2.649 76.621 2.828 ;
      RECT 76.525 2.644 76.535 2.825 ;
      RECT 76.511 2.643 76.525 2.825 ;
      RECT 76.425 2.639 76.511 2.82 ;
      RECT 76.405 2.633 76.425 2.816 ;
      RECT 76.345 2.628 76.405 2.815 ;
      RECT 76.315 2.62 76.345 2.815 ;
      RECT 76.305 2.605 76.315 2.815 ;
      RECT 76.301 2.595 76.305 2.814 ;
      RECT 76.215 2.595 76.301 2.81 ;
      RECT 76.105 2.605 76.115 2.805 ;
      RECT 76.035 2.615 76.065 2.8 ;
      RECT 76.025 2.615 76.035 2.8 ;
      RECT 76.945 3.115 77.205 3.375 ;
      RECT 76.875 3.125 77.205 3.335 ;
      RECT 76.865 3.13 77.205 3.33 ;
      RECT 76.285 3.115 76.545 3.375 ;
      RECT 76.285 3.16 76.655 3.365 ;
      RECT 76.285 3.155 76.645 3.365 ;
      RECT 75.195 3.322 75.375 3.765 ;
      RECT 75.185 3.322 75.375 3.763 ;
      RECT 75.185 3.337 75.385 3.76 ;
      RECT 75.175 2.26 75.305 3.758 ;
      RECT 75.175 3.385 75.445 3.645 ;
      RECT 75.175 3.36 75.395 3.645 ;
      RECT 75.175 3.295 75.365 3.758 ;
      RECT 75.175 3.255 75.335 3.758 ;
      RECT 75.175 3.21 75.325 3.758 ;
      RECT 75.175 3.15 75.315 3.758 ;
      RECT 75.165 2.545 75.305 3.2 ;
      RECT 75.205 2.245 75.315 3.065 ;
      RECT 75.175 2.26 75.355 2.52 ;
      RECT 75.175 2.26 75.365 2.47 ;
      RECT 75.205 2.245 75.375 2.463 ;
      RECT 75.195 2.247 75.385 2.458 ;
      RECT 75.185 2.252 75.395 2.45 ;
      RECT 74.045 7.77 74.335 8 ;
      RECT 74.105 6.29 74.275 8 ;
      RECT 74.055 6.655 74.405 7.005 ;
      RECT 74.045 6.29 74.335 6.52 ;
      RECT 73.64 2.395 73.745 2.965 ;
      RECT 73.64 2.73 73.965 2.96 ;
      RECT 73.64 2.76 74.135 2.93 ;
      RECT 73.64 2.395 73.83 2.96 ;
      RECT 73.055 2.36 73.345 2.59 ;
      RECT 73.055 2.395 73.83 2.565 ;
      RECT 73.115 0.88 73.285 2.59 ;
      RECT 73.055 0.88 73.345 1.11 ;
      RECT 73.055 7.77 73.345 8 ;
      RECT 73.115 6.29 73.285 8 ;
      RECT 73.055 6.29 73.345 6.52 ;
      RECT 73.055 6.325 73.91 6.485 ;
      RECT 73.74 5.92 73.91 6.485 ;
      RECT 73.055 6.32 73.45 6.485 ;
      RECT 73.675 5.92 73.965 6.15 ;
      RECT 73.675 5.95 74.135 6.12 ;
      RECT 72.685 2.73 72.975 2.96 ;
      RECT 72.685 2.76 73.145 2.93 ;
      RECT 72.75 1.655 72.915 2.96 ;
      RECT 71.265 1.625 71.555 1.855 ;
      RECT 71.265 1.655 72.915 1.825 ;
      RECT 71.325 0.885 71.495 1.855 ;
      RECT 71.265 0.885 71.555 1.115 ;
      RECT 71.265 7.765 71.555 7.995 ;
      RECT 71.325 7.025 71.495 7.995 ;
      RECT 71.325 7.12 72.915 7.29 ;
      RECT 72.745 5.92 72.915 7.29 ;
      RECT 71.265 7.025 71.555 7.255 ;
      RECT 72.685 5.92 72.975 6.15 ;
      RECT 72.685 5.95 73.145 6.12 ;
      RECT 69.3 3.43 69.65 3.78 ;
      RECT 69.39 2.025 69.56 3.78 ;
      RECT 71.695 1.965 72.045 2.315 ;
      RECT 69.39 2.025 71.01 2.2 ;
      RECT 69.39 2.025 72.045 2.195 ;
      RECT 71.72 6.655 72.045 6.98 ;
      RECT 67.095 6.61 67.445 6.96 ;
      RECT 71.695 6.655 72.045 6.885 ;
      RECT 66.935 6.655 67.445 6.885 ;
      RECT 66.765 6.685 72.045 6.855 ;
      RECT 70.92 2.365 71.24 2.685 ;
      RECT 70.89 2.365 71.24 2.595 ;
      RECT 70.72 2.395 71.24 2.565 ;
      RECT 70.92 6.225 71.24 6.545 ;
      RECT 70.89 6.285 71.24 6.515 ;
      RECT 70.72 6.315 71.24 6.485 ;
      RECT 66.76 3.255 66.95 3.925 ;
      RECT 66.7 3.665 66.74 3.925 ;
      RECT 68.07 2.89 68.08 3.111 ;
      RECT 68 2.885 68.07 3.236 ;
      RECT 67.99 2.885 68 3.36 ;
      RECT 67.96 2.885 67.99 3.41 ;
      RECT 67.94 2.885 67.96 3.485 ;
      RECT 67.92 2.885 67.94 3.555 ;
      RECT 67.89 2.885 67.92 3.595 ;
      RECT 67.88 2.885 67.89 3.615 ;
      RECT 67.87 2.885 67.88 3.626 ;
      RECT 67.86 3.135 67.87 3.628 ;
      RECT 67.85 3.2 67.86 3.63 ;
      RECT 67.84 3.295 67.85 3.632 ;
      RECT 67.83 3.37 67.84 3.634 ;
      RECT 67.78 3.394 67.83 3.64 ;
      RECT 67.74 3.429 67.78 3.649 ;
      RECT 67.73 3.445 67.74 3.654 ;
      RECT 67.716 3.45 67.73 3.657 ;
      RECT 67.63 3.49 67.716 3.668 ;
      RECT 67.55 3.533 67.63 3.686 ;
      RECT 67.53 3.543 67.55 3.697 ;
      RECT 67.5 3.551 67.53 3.702 ;
      RECT 67.48 3.561 67.5 3.707 ;
      RECT 67.456 3.567 67.48 3.712 ;
      RECT 67.37 3.577 67.456 3.725 ;
      RECT 67.292 3.583 67.37 3.745 ;
      RECT 67.206 3.578 67.292 3.764 ;
      RECT 67.12 3.574 67.206 3.785 ;
      RECT 67.04 3.57 67.12 3.8 ;
      RECT 66.97 3.566 67.04 3.831 ;
      RECT 66.96 3.277 66.97 3.345 ;
      RECT 66.96 3.555 66.97 3.861 ;
      RECT 66.95 3.262 66.96 3.49 ;
      RECT 66.95 3.535 66.96 3.925 ;
      RECT 66.74 3.285 66.76 3.925 ;
      RECT 67.54 2.605 67.55 3.345 ;
      RECT 67.36 3.125 67.38 3.345 ;
      RECT 67.37 3.115 67.38 3.345 ;
      RECT 67.87 2.155 67.91 2.415 ;
      RECT 67.86 2.155 67.87 2.425 ;
      RECT 67.826 2.155 67.86 2.452 ;
      RECT 67.74 2.155 67.826 2.512 ;
      RECT 67.72 2.155 67.74 2.575 ;
      RECT 67.66 2.155 67.72 2.74 ;
      RECT 67.65 2.155 67.66 2.9 ;
      RECT 67.62 2.346 67.65 2.995 ;
      RECT 67.61 2.401 67.62 3.095 ;
      RECT 67.6 2.43 67.61 3.14 ;
      RECT 67.59 2.455 67.6 3.173 ;
      RECT 67.58 2.49 67.59 3.228 ;
      RECT 67.56 2.535 67.58 3.29 ;
      RECT 67.55 2.58 67.56 3.34 ;
      RECT 67.53 2.64 67.54 3.345 ;
      RECT 67.52 2.67 67.53 3.345 ;
      RECT 67.5 2.7 67.52 3.345 ;
      RECT 67.45 2.805 67.5 3.345 ;
      RECT 67.44 2.9 67.45 3.345 ;
      RECT 67.43 2.93 67.44 3.345 ;
      RECT 67.405 2.98 67.43 3.345 ;
      RECT 67.4 3.035 67.405 3.345 ;
      RECT 67.38 3.06 67.4 3.345 ;
      RECT 67.34 3.14 67.36 3.335 ;
      RECT 67.09 2.725 67.16 2.935 ;
      RECT 64.33 2.635 64.59 2.895 ;
      RECT 67.16 2.73 67.17 2.93 ;
      RECT 67.046 2.723 67.09 2.935 ;
      RECT 66.96 2.716 67.046 2.935 ;
      RECT 66.94 2.711 66.96 2.925 ;
      RECT 66.93 2.709 66.94 2.905 ;
      RECT 66.88 2.706 66.93 2.9 ;
      RECT 66.85 2.702 66.88 2.895 ;
      RECT 66.83 2.7 66.85 2.89 ;
      RECT 66.79 2.697 66.83 2.885 ;
      RECT 66.72 2.691 66.79 2.88 ;
      RECT 66.69 2.686 66.72 2.875 ;
      RECT 66.67 2.684 66.69 2.87 ;
      RECT 66.64 2.681 66.67 2.865 ;
      RECT 66.58 2.677 66.64 2.86 ;
      RECT 66.51 2.675 66.58 2.85 ;
      RECT 66.476 2.673 66.51 2.843 ;
      RECT 66.39 2.668 66.476 2.835 ;
      RECT 66.356 2.662 66.39 2.827 ;
      RECT 66.27 2.652 66.356 2.819 ;
      RECT 66.236 2.643 66.27 2.811 ;
      RECT 66.15 2.638 66.236 2.803 ;
      RECT 66.08 2.635 66.15 2.793 ;
      RECT 66.06 2.63 66.08 2.787 ;
      RECT 66.056 2.625 66.06 2.786 ;
      RECT 65.97 2.621 66.056 2.781 ;
      RECT 65.93 2.616 65.97 2.774 ;
      RECT 65.85 2.615 65.93 2.769 ;
      RECT 65.83 2.615 65.85 2.766 ;
      RECT 65.804 2.615 65.83 2.766 ;
      RECT 65.718 2.617 65.804 2.77 ;
      RECT 65.632 2.619 65.718 2.777 ;
      RECT 65.546 2.621 65.632 2.783 ;
      RECT 65.46 2.624 65.546 2.79 ;
      RECT 65.426 2.626 65.46 2.795 ;
      RECT 65.34 2.631 65.426 2.8 ;
      RECT 65.316 2.626 65.34 2.804 ;
      RECT 65.23 2.631 65.316 2.809 ;
      RECT 65.192 2.636 65.23 2.814 ;
      RECT 65.106 2.639 65.192 2.819 ;
      RECT 65.02 2.643 65.106 2.826 ;
      RECT 64.956 2.645 65.02 2.832 ;
      RECT 64.87 2.645 64.956 2.838 ;
      RECT 64.786 2.646 64.87 2.845 ;
      RECT 64.7 2.649 64.786 2.852 ;
      RECT 64.676 2.651 64.7 2.856 ;
      RECT 64.59 2.653 64.676 2.861 ;
      RECT 64.32 2.67 64.33 2.865 ;
      RECT 66.505 7.765 66.795 7.995 ;
      RECT 66.565 7.025 66.735 7.995 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 66.505 7.025 66.795 7.425 ;
      RECT 66.56 2.247 66.75 2.455 ;
      RECT 66.55 2.252 66.76 2.45 ;
      RECT 66.54 2.233 66.55 2.445 ;
      RECT 66.51 2.228 66.54 2.44 ;
      RECT 66.47 2.252 66.76 2.43 ;
      RECT 66.25 2.165 66.51 2.425 ;
      RECT 66.55 2.236 66.56 2.45 ;
      RECT 66.25 2.245 66.74 2.425 ;
      RECT 66.25 2.241 66.6 2.425 ;
      RECT 66.2 3.155 66.25 3.435 ;
      RECT 66.13 3.125 66.16 3.435 ;
      RECT 66.27 3.155 66.33 3.415 ;
      RECT 66.13 3.115 66.15 3.435 ;
      RECT 66.25 3.155 66.27 3.425 ;
      RECT 66.17 3.145 66.2 3.435 ;
      RECT 66.16 3.13 66.17 3.435 ;
      RECT 66.11 3.105 66.13 3.435 ;
      RECT 66.08 3.09 66.11 3.435 ;
      RECT 66.07 3.08 66.08 3.435 ;
      RECT 66.05 3.069 66.07 3.43 ;
      RECT 66.03 3.057 66.05 3.4 ;
      RECT 66.02 3.048 66.03 3.383 ;
      RECT 65.99 3.03 66.02 3.375 ;
      RECT 65.98 2.995 65.99 3.367 ;
      RECT 65.97 2.975 65.98 3.36 ;
      RECT 65.96 2.955 65.97 3.353 ;
      RECT 65.95 2.94 65.96 3.348 ;
      RECT 65.94 2.92 65.95 3.343 ;
      RECT 65.93 2.915 65.94 3.338 ;
      RECT 65.926 2.905 65.93 3.334 ;
      RECT 65.84 2.905 65.926 3.309 ;
      RECT 65.81 2.905 65.84 3.275 ;
      RECT 65.8 2.905 65.81 3.255 ;
      RECT 65.74 2.905 65.8 3.2 ;
      RECT 65.73 2.92 65.74 3.145 ;
      RECT 65.72 2.93 65.73 3.125 ;
      RECT 65.67 3.665 65.93 3.925 ;
      RECT 65.59 3.685 65.93 3.901 ;
      RECT 65.57 3.685 65.93 3.896 ;
      RECT 65.546 3.685 65.93 3.894 ;
      RECT 65.46 3.685 65.93 3.889 ;
      RECT 65.31 3.625 65.57 3.885 ;
      RECT 65.27 3.68 65.59 3.88 ;
      RECT 65.26 3.69 65.93 3.875 ;
      RECT 65.28 3.675 65.57 3.885 ;
      RECT 65.17 2.115 65.43 2.375 ;
      RECT 65.17 2.2 65.44 2.3 ;
      RECT 64.34 3.63 64.36 3.874 ;
      RECT 64.34 3.63 64.41 3.869 ;
      RECT 64.32 3.635 64.41 3.868 ;
      RECT 64.31 3.65 64.496 3.858 ;
      RECT 64.31 3.65 64.57 3.855 ;
      RECT 64.305 3.687 64.58 3.845 ;
      RECT 64.305 3.687 64.666 3.841 ;
      RECT 64.305 3.687 64.68 3.827 ;
      RECT 64.58 3.565 64.84 3.825 ;
      RECT 64.3 3.692 64.84 3.82 ;
      RECT 64.29 3.74 64.84 3.795 ;
      RECT 64.56 3.605 64.58 3.854 ;
      RECT 64.496 3.609 64.56 3.857 ;
      RECT 64.36 3.622 64.84 3.825 ;
      RECT 64.41 3.616 64.496 3.862 ;
      RECT 63.81 2.475 63.82 2.645 ;
      RECT 63.87 2.435 63.88 2.615 ;
      RECT 64.17 2.245 64.18 2.455 ;
      RECT 64.5 2.095 64.75 2.355 ;
      RECT 64.49 2.095 64.5 2.357 ;
      RECT 64.48 2.155 64.49 2.361 ;
      RECT 64.45 2.157 64.48 2.369 ;
      RECT 64.42 2.162 64.45 2.383 ;
      RECT 64.41 2.166 64.42 2.393 ;
      RECT 64.38 2.171 64.41 2.405 ;
      RECT 64.35 2.18 64.38 2.406 ;
      RECT 64.28 2.19 64.35 2.41 ;
      RECT 64.24 2.195 64.28 2.414 ;
      RECT 64.22 2.195 64.24 2.425 ;
      RECT 64.21 2.2 64.22 2.435 ;
      RECT 64.2 2.21 64.21 2.438 ;
      RECT 64.19 2.23 64.2 2.443 ;
      RECT 64.18 2.24 64.19 2.445 ;
      RECT 64.15 2.255 64.17 2.462 ;
      RECT 64.14 2.267 64.15 2.472 ;
      RECT 64.13 2.273 64.14 2.475 ;
      RECT 64.096 2.286 64.13 2.485 ;
      RECT 64.01 2.32 64.096 2.518 ;
      RECT 63.99 2.355 64.01 2.547 ;
      RECT 63.97 2.37 63.99 2.559 ;
      RECT 63.95 2.38 63.97 2.571 ;
      RECT 63.9 2.399 63.95 2.591 ;
      RECT 63.89 2.416 63.9 2.605 ;
      RECT 63.88 2.422 63.89 2.61 ;
      RECT 63.86 2.44 63.87 2.618 ;
      RECT 63.85 2.445 63.86 2.625 ;
      RECT 63.84 2.456 63.85 2.632 ;
      RECT 63.82 2.461 63.84 2.64 ;
      RECT 63.8 2.475 63.81 2.65 ;
      RECT 63.79 2.48 63.8 2.66 ;
      RECT 63.76 2.494 63.79 2.67 ;
      RECT 63.75 2.507 63.76 2.68 ;
      RECT 63.67 2.538 63.75 2.705 ;
      RECT 63.65 2.568 63.67 2.73 ;
      RECT 63.64 2.573 63.65 2.737 ;
      RECT 63.61 2.585 63.64 2.743 ;
      RECT 63.6 2.6 63.61 2.749 ;
      RECT 63.59 2.605 63.6 2.752 ;
      RECT 63.57 2.615 63.59 2.756 ;
      RECT 63.55 2.62 63.57 2.762 ;
      RECT 63.52 2.625 63.55 2.77 ;
      RECT 63.49 2.63 63.52 2.78 ;
      RECT 63.46 2.64 63.49 2.789 ;
      RECT 63.42 2.645 63.46 2.797 ;
      RECT 63.37 2.638 63.42 2.809 ;
      RECT 63.35 2.629 63.37 2.82 ;
      RECT 63.34 2.626 63.35 2.825 ;
      RECT 63.3 2.625 63.34 2.826 ;
      RECT 63.29 2.61 63.3 2.827 ;
      RECT 63.262 2.595 63.29 2.828 ;
      RECT 63.176 2.595 63.262 2.83 ;
      RECT 63.09 2.595 63.176 2.834 ;
      RECT 63.07 2.595 63.09 2.83 ;
      RECT 63.06 2.605 63.07 2.823 ;
      RECT 63.05 2.62 63.06 2.818 ;
      RECT 63.04 2.625 63.05 2.795 ;
      RECT 64.52 3.13 64.53 3.33 ;
      RECT 64.47 3.125 64.52 3.35 ;
      RECT 64.46 3.125 64.47 3.37 ;
      RECT 64.416 3.125 64.46 3.374 ;
      RECT 64.33 3.125 64.416 3.371 ;
      RECT 64.27 3.135 64.33 3.368 ;
      RECT 64.21 3.149 64.27 3.366 ;
      RECT 64.2 3.154 64.21 3.364 ;
      RECT 64.19 3.16 64.2 3.363 ;
      RECT 64.12 3.173 64.19 3.359 ;
      RECT 64.072 3.187 64.12 3.36 ;
      RECT 63.986 3.203 64.072 3.372 ;
      RECT 63.9 3.224 63.986 3.388 ;
      RECT 63.88 3.235 63.9 3.398 ;
      RECT 63.8 3.245 63.88 3.408 ;
      RECT 63.766 3.259 63.8 3.42 ;
      RECT 63.68 3.274 63.766 3.435 ;
      RECT 63.65 3.29 63.68 3.445 ;
      RECT 63.595 3.305 63.65 3.456 ;
      RECT 63.55 3.323 63.595 3.476 ;
      RECT 63.496 3.342 63.55 3.496 ;
      RECT 63.41 3.368 63.496 3.523 ;
      RECT 63.39 3.39 63.41 3.543 ;
      RECT 63.33 3.405 63.39 3.559 ;
      RECT 63.32 3.42 63.33 3.573 ;
      RECT 63.3 3.425 63.32 3.579 ;
      RECT 63.27 3.438 63.3 3.589 ;
      RECT 63.25 3.443 63.27 3.598 ;
      RECT 63.24 3.45 63.25 3.603 ;
      RECT 63.23 3.455 63.24 3.606 ;
      RECT 63.19 3.465 63.23 3.615 ;
      RECT 63.165 3.48 63.19 3.627 ;
      RECT 63.12 3.495 63.165 3.639 ;
      RECT 63.1 3.507 63.12 3.651 ;
      RECT 63.07 3.512 63.1 3.661 ;
      RECT 63.05 3.519 63.07 3.671 ;
      RECT 63.04 3.525 63.05 3.68 ;
      RECT 63.016 3.532 63.04 3.69 ;
      RECT 62.93 3.554 63.016 3.71 ;
      RECT 62.92 3.573 62.93 3.725 ;
      RECT 62.896 3.58 62.92 3.731 ;
      RECT 62.81 3.602 62.896 3.756 ;
      RECT 62.77 3.627 62.81 3.783 ;
      RECT 62.76 3.636 62.77 3.793 ;
      RECT 62.71 3.646 62.76 3.802 ;
      RECT 62.69 3.66 62.71 3.812 ;
      RECT 62.66 3.67 62.69 3.817 ;
      RECT 62.65 3.675 62.66 3.82 ;
      RECT 62.576 3.677 62.65 3.827 ;
      RECT 62.49 3.681 62.576 3.839 ;
      RECT 62.48 3.684 62.49 3.845 ;
      RECT 62.22 3.635 62.48 3.895 ;
      RECT 63.75 3.705 63.94 3.915 ;
      RECT 63.74 3.71 63.95 3.91 ;
      RECT 63.73 3.71 63.95 3.875 ;
      RECT 63.65 3.595 63.91 3.855 ;
      RECT 62.56 3.125 62.75 3.425 ;
      RECT 62.55 3.125 62.75 3.42 ;
      RECT 62.54 3.125 62.76 3.415 ;
      RECT 62.53 3.125 62.76 3.41 ;
      RECT 62.53 3.125 62.79 3.385 ;
      RECT 62.49 2.165 62.75 2.425 ;
      RECT 62.3 2.09 62.386 2.423 ;
      RECT 62.3 2.09 62.43 2.419 ;
      RECT 62.28 2.094 62.44 2.418 ;
      RECT 62.43 2.085 62.44 2.418 ;
      RECT 62.3 2.09 62.45 2.417 ;
      RECT 62.28 2.1 62.49 2.416 ;
      RECT 62.27 2.095 62.45 2.408 ;
      RECT 62.26 2.11 62.49 2.315 ;
      RECT 62.26 2.16 62.69 2.315 ;
      RECT 62.26 2.15 62.67 2.315 ;
      RECT 62.26 2.14 62.64 2.315 ;
      RECT 62.26 2.13 62.58 2.315 ;
      RECT 62.26 2.115 62.56 2.315 ;
      RECT 62.386 2.086 62.44 2.418 ;
      RECT 61.46 2.745 61.6 3.035 ;
      RECT 61.72 2.768 61.73 2.955 ;
      RECT 62.42 2.665 62.6 2.895 ;
      RECT 62.42 2.665 62.61 2.885 ;
      RECT 62.63 2.67 62.64 2.875 ;
      RECT 62.61 2.665 62.63 2.88 ;
      RECT 62.37 2.669 62.42 2.895 ;
      RECT 62.36 2.674 62.37 2.895 ;
      RECT 62.326 2.679 62.36 2.896 ;
      RECT 62.24 2.694 62.326 2.898 ;
      RECT 62.226 2.706 62.24 2.901 ;
      RECT 62.14 2.716 62.226 2.903 ;
      RECT 62.116 2.726 62.14 2.905 ;
      RECT 62.03 2.737 62.116 2.905 ;
      RECT 62 2.747 62.03 2.905 ;
      RECT 61.97 2.752 62 2.908 ;
      RECT 61.95 2.757 61.97 2.913 ;
      RECT 61.93 2.762 61.95 2.915 ;
      RECT 61.88 2.77 61.93 2.915 ;
      RECT 61.86 2.774 61.88 2.915 ;
      RECT 61.84 2.773 61.86 2.92 ;
      RECT 61.78 2.771 61.84 2.935 ;
      RECT 61.73 2.769 61.78 2.95 ;
      RECT 61.64 2.766 61.72 3.035 ;
      RECT 61.61 2.76 61.64 3.035 ;
      RECT 61.6 2.75 61.61 3.035 ;
      RECT 61.41 2.745 61.46 2.96 ;
      RECT 61.4 2.75 61.41 2.95 ;
      RECT 61.64 3.225 61.9 3.485 ;
      RECT 61.64 3.225 61.93 3.375 ;
      RECT 61.64 3.225 61.97 3.36 ;
      RECT 61.9 3.145 62.09 3.355 ;
      RECT 61.9 3.15 62.1 3.345 ;
      RECT 61.85 3.22 62.1 3.345 ;
      RECT 61.88 3.155 61.9 3.485 ;
      RECT 61.87 3.18 62.1 3.345 ;
      RECT 61.05 3.125 61.06 3.355 ;
      RECT 60.95 2.245 61.02 3.355 ;
      RECT 61.69 2.355 61.95 2.615 ;
      RECT 61.39 2.405 61.52 2.565 ;
      RECT 61.606 2.412 61.69 2.565 ;
      RECT 61.52 2.407 61.606 2.565 ;
      RECT 61.33 2.405 61.39 2.575 ;
      RECT 61.3 2.403 61.33 2.59 ;
      RECT 61.28 2.401 61.3 2.6 ;
      RECT 61.27 2.399 61.28 2.605 ;
      RECT 61.25 2.398 61.27 2.615 ;
      RECT 61.24 2.396 61.25 2.62 ;
      RECT 61.22 2.395 61.24 2.625 ;
      RECT 61.2 2.39 61.22 2.63 ;
      RECT 61.17 2.376 61.2 2.64 ;
      RECT 61.13 2.355 61.17 2.655 ;
      RECT 61.12 2.34 61.13 2.665 ;
      RECT 61.1 2.331 61.12 2.675 ;
      RECT 61.09 2.322 61.1 2.695 ;
      RECT 61.08 2.317 61.09 2.755 ;
      RECT 61.06 2.311 61.08 2.84 ;
      RECT 61.06 3.15 61.07 3.35 ;
      RECT 61.05 2.306 61.06 3.07 ;
      RECT 61.04 2.28 61.05 3.355 ;
      RECT 61.02 2.25 61.04 3.355 ;
      RECT 60.93 2.245 60.95 2.58 ;
      RECT 60.94 2.68 60.95 3.355 ;
      RECT 60.93 2.72 60.94 3.355 ;
      RECT 60.9 2.245 60.93 2.525 ;
      RECT 60.91 2.81 60.93 3.355 ;
      RECT 60.895 2.915 60.91 3.355 ;
      RECT 60.87 2.245 60.9 2.48 ;
      RECT 60.89 2.947 60.895 3.355 ;
      RECT 60.87 3.05 60.89 3.355 ;
      RECT 60.86 2.245 60.87 2.47 ;
      RECT 60.86 3.12 60.87 3.35 ;
      RECT 60.84 2.245 60.86 2.46 ;
      RECT 60.83 2.25 60.84 2.45 ;
      RECT 61.04 3.525 61.06 3.765 ;
      RECT 60.36 3.455 60.44 3.725 ;
      RECT 60.27 3.455 60.28 3.665 ;
      RECT 61.55 3.525 61.56 3.725 ;
      RECT 61.47 3.515 61.55 3.75 ;
      RECT 61.466 3.515 61.47 3.776 ;
      RECT 61.38 3.515 61.466 3.786 ;
      RECT 61.36 3.515 61.38 3.794 ;
      RECT 61.336 3.516 61.36 3.792 ;
      RECT 61.25 3.521 61.336 3.787 ;
      RECT 61.232 3.525 61.25 3.781 ;
      RECT 61.146 3.525 61.232 3.777 ;
      RECT 61.06 3.525 61.146 3.769 ;
      RECT 60.956 3.525 61.04 3.762 ;
      RECT 60.87 3.525 60.956 3.756 ;
      RECT 60.81 3.52 60.87 3.75 ;
      RECT 60.782 3.514 60.81 3.747 ;
      RECT 60.696 3.511 60.782 3.744 ;
      RECT 60.61 3.507 60.696 3.738 ;
      RECT 60.565 3.495 60.61 3.734 ;
      RECT 60.54 3.48 60.565 3.732 ;
      RECT 60.5 3.465 60.54 3.73 ;
      RECT 60.44 3.455 60.5 3.727 ;
      RECT 60.35 3.455 60.36 3.72 ;
      RECT 60.335 3.455 60.35 3.71 ;
      RECT 60.28 3.455 60.335 3.685 ;
      RECT 60.26 3.47 60.27 3.66 ;
      RECT 60.39 2.635 60.65 2.895 ;
      RECT 60.39 2.645 60.67 2.855 ;
      RECT 60.39 2.65 60.68 2.85 ;
      RECT 58.37 2.115 58.63 2.375 ;
      RECT 58.36 2.145 58.63 2.355 ;
      RECT 60.29 2.055 60.54 2.315 ;
      RECT 60.28 2.055 60.29 2.316 ;
      RECT 60.25 2.14 60.28 2.318 ;
      RECT 60.24 2.145 60.25 2.32 ;
      RECT 60.18 2.16 60.24 2.326 ;
      RECT 60.15 2.18 60.18 2.333 ;
      RECT 60.12 2.191 60.15 2.34 ;
      RECT 60.1 2.201 60.12 2.345 ;
      RECT 60.082 2.204 60.1 2.344 ;
      RECT 59.996 2.203 60.082 2.344 ;
      RECT 59.91 2.2 59.996 2.343 ;
      RECT 59.824 2.197 59.91 2.342 ;
      RECT 59.738 2.194 59.824 2.342 ;
      RECT 59.652 2.192 59.738 2.341 ;
      RECT 59.566 2.189 59.652 2.34 ;
      RECT 59.48 2.186 59.566 2.34 ;
      RECT 59.462 2.185 59.48 2.339 ;
      RECT 59.376 2.184 59.462 2.339 ;
      RECT 59.29 2.182 59.376 2.338 ;
      RECT 59.204 2.181 59.29 2.338 ;
      RECT 59.118 2.18 59.204 2.337 ;
      RECT 59.032 2.178 59.118 2.337 ;
      RECT 58.946 2.177 59.032 2.336 ;
      RECT 58.86 2.175 58.946 2.336 ;
      RECT 58.836 2.174 58.86 2.335 ;
      RECT 58.75 2.169 58.836 2.335 ;
      RECT 58.716 2.162 58.75 2.335 ;
      RECT 58.63 2.152 58.716 2.335 ;
      RECT 58.35 2.15 58.36 2.35 ;
      RECT 59.63 3.205 59.89 3.465 ;
      RECT 59.63 3.205 59.97 3.251 ;
      RECT 59.77 3.185 59.98 3.24 ;
      RECT 59.83 3.16 60.04 3.2 ;
      RECT 59.84 3.155 60.04 3.2 ;
      RECT 59.85 3.13 60.04 3.2 ;
      RECT 59.91 2.96 59.96 3.29 ;
      RECT 59.86 3.09 60.05 3.15 ;
      RECT 59.9 3.016 59.91 3.329 ;
      RECT 59.86 3.09 60.08 3.125 ;
      RECT 59.86 3.09 60.1 3.1 ;
      RECT 59.97 2.89 60.16 3.095 ;
      RECT 59.96 2.9 60.17 3.09 ;
      RECT 59.88 3.063 60.17 3.09 ;
      RECT 59.89 3.039 59.9 3.345 ;
      RECT 59.98 2.885 60.15 3.095 ;
      RECT 59.27 2.675 59.46 2.885 ;
      RECT 57.84 2.605 58.1 2.865 ;
      RECT 58.19 2.595 58.29 2.805 ;
      RECT 58.14 2.615 58.18 2.805 ;
      RECT 59.46 2.685 59.47 2.88 ;
      RECT 59.26 2.685 59.27 2.88 ;
      RECT 59.24 2.7 59.26 2.87 ;
      RECT 59.23 2.71 59.24 2.865 ;
      RECT 59.19 2.71 59.23 2.863 ;
      RECT 59.166 2.704 59.19 2.86 ;
      RECT 59.08 2.699 59.166 2.857 ;
      RECT 59.02 2.695 59.08 2.852 ;
      RECT 58.986 2.692 59.02 2.849 ;
      RECT 58.9 2.682 58.986 2.845 ;
      RECT 58.896 2.675 58.9 2.842 ;
      RECT 58.81 2.67 58.896 2.84 ;
      RECT 58.782 2.663 58.81 2.836 ;
      RECT 58.696 2.658 58.782 2.833 ;
      RECT 58.61 2.649 58.696 2.828 ;
      RECT 58.6 2.644 58.61 2.825 ;
      RECT 58.586 2.643 58.6 2.825 ;
      RECT 58.5 2.639 58.586 2.82 ;
      RECT 58.48 2.633 58.5 2.816 ;
      RECT 58.42 2.628 58.48 2.815 ;
      RECT 58.39 2.62 58.42 2.815 ;
      RECT 58.38 2.605 58.39 2.815 ;
      RECT 58.376 2.595 58.38 2.814 ;
      RECT 58.29 2.595 58.376 2.81 ;
      RECT 58.18 2.605 58.19 2.805 ;
      RECT 58.11 2.615 58.14 2.8 ;
      RECT 58.1 2.615 58.11 2.8 ;
      RECT 59.02 3.115 59.28 3.375 ;
      RECT 58.95 3.125 59.28 3.335 ;
      RECT 58.94 3.13 59.28 3.33 ;
      RECT 58.36 3.115 58.62 3.375 ;
      RECT 58.36 3.16 58.73 3.365 ;
      RECT 58.36 3.155 58.72 3.365 ;
      RECT 57.27 3.322 57.45 3.765 ;
      RECT 57.26 3.322 57.45 3.763 ;
      RECT 57.26 3.337 57.46 3.76 ;
      RECT 57.25 2.26 57.38 3.758 ;
      RECT 57.25 3.385 57.52 3.645 ;
      RECT 57.25 3.36 57.47 3.645 ;
      RECT 57.25 3.295 57.44 3.758 ;
      RECT 57.25 3.255 57.41 3.758 ;
      RECT 57.25 3.21 57.4 3.758 ;
      RECT 57.25 3.15 57.39 3.758 ;
      RECT 57.24 2.545 57.38 3.2 ;
      RECT 57.28 2.245 57.39 3.065 ;
      RECT 57.25 2.26 57.43 2.52 ;
      RECT 57.25 2.26 57.44 2.47 ;
      RECT 57.28 2.245 57.45 2.463 ;
      RECT 57.27 2.247 57.46 2.458 ;
      RECT 57.26 2.252 57.47 2.45 ;
      RECT 56.12 7.77 56.41 8 ;
      RECT 56.18 6.29 56.35 8 ;
      RECT 56.13 6.655 56.48 7.005 ;
      RECT 56.12 6.29 56.41 6.52 ;
      RECT 55.715 2.395 55.82 2.965 ;
      RECT 55.715 2.73 56.04 2.96 ;
      RECT 55.715 2.76 56.21 2.93 ;
      RECT 55.715 2.395 55.905 2.96 ;
      RECT 55.13 2.36 55.42 2.59 ;
      RECT 55.13 2.395 55.905 2.565 ;
      RECT 55.19 0.88 55.36 2.59 ;
      RECT 55.13 0.88 55.42 1.11 ;
      RECT 55.13 7.77 55.42 8 ;
      RECT 55.19 6.29 55.36 8 ;
      RECT 55.13 6.29 55.42 6.52 ;
      RECT 55.13 6.325 55.985 6.485 ;
      RECT 55.815 5.92 55.985 6.485 ;
      RECT 55.13 6.32 55.525 6.485 ;
      RECT 55.75 5.92 56.04 6.15 ;
      RECT 55.75 5.95 56.21 6.12 ;
      RECT 54.76 2.73 55.05 2.96 ;
      RECT 54.76 2.76 55.22 2.93 ;
      RECT 54.825 1.655 54.99 2.96 ;
      RECT 53.34 1.625 53.63 1.855 ;
      RECT 53.34 1.655 54.99 1.825 ;
      RECT 53.4 0.885 53.57 1.855 ;
      RECT 53.34 0.885 53.63 1.115 ;
      RECT 53.34 7.765 53.63 7.995 ;
      RECT 53.4 7.025 53.57 7.995 ;
      RECT 53.4 7.12 54.99 7.29 ;
      RECT 54.82 5.92 54.99 7.29 ;
      RECT 53.34 7.025 53.63 7.255 ;
      RECT 54.76 5.92 55.05 6.15 ;
      RECT 54.76 5.95 55.22 6.12 ;
      RECT 51.375 3.43 51.725 3.78 ;
      RECT 51.465 2.025 51.635 3.78 ;
      RECT 53.77 1.965 54.12 2.315 ;
      RECT 51.465 2.025 53.085 2.2 ;
      RECT 51.465 2.025 54.12 2.195 ;
      RECT 53.795 6.655 54.12 6.98 ;
      RECT 49.225 6.615 49.575 6.965 ;
      RECT 53.77 6.655 54.12 6.885 ;
      RECT 49.01 6.655 49.575 6.885 ;
      RECT 48.84 6.685 54.12 6.855 ;
      RECT 52.995 2.365 53.315 2.685 ;
      RECT 52.965 2.365 53.315 2.595 ;
      RECT 52.795 2.395 53.315 2.565 ;
      RECT 52.995 6.225 53.315 6.545 ;
      RECT 52.965 6.285 53.315 6.515 ;
      RECT 52.795 6.315 53.315 6.485 ;
      RECT 48.835 3.255 49.025 3.925 ;
      RECT 48.775 3.665 48.815 3.925 ;
      RECT 50.145 2.89 50.155 3.111 ;
      RECT 50.075 2.885 50.145 3.236 ;
      RECT 50.065 2.885 50.075 3.36 ;
      RECT 50.035 2.885 50.065 3.41 ;
      RECT 50.015 2.885 50.035 3.485 ;
      RECT 49.995 2.885 50.015 3.555 ;
      RECT 49.965 2.885 49.995 3.595 ;
      RECT 49.955 2.885 49.965 3.615 ;
      RECT 49.945 2.885 49.955 3.626 ;
      RECT 49.935 3.135 49.945 3.628 ;
      RECT 49.925 3.2 49.935 3.63 ;
      RECT 49.915 3.295 49.925 3.632 ;
      RECT 49.905 3.37 49.915 3.634 ;
      RECT 49.855 3.394 49.905 3.64 ;
      RECT 49.815 3.429 49.855 3.649 ;
      RECT 49.805 3.445 49.815 3.654 ;
      RECT 49.791 3.45 49.805 3.657 ;
      RECT 49.705 3.49 49.791 3.668 ;
      RECT 49.625 3.533 49.705 3.686 ;
      RECT 49.605 3.543 49.625 3.697 ;
      RECT 49.575 3.551 49.605 3.702 ;
      RECT 49.555 3.561 49.575 3.707 ;
      RECT 49.531 3.567 49.555 3.712 ;
      RECT 49.445 3.577 49.531 3.725 ;
      RECT 49.367 3.583 49.445 3.745 ;
      RECT 49.281 3.578 49.367 3.764 ;
      RECT 49.195 3.574 49.281 3.785 ;
      RECT 49.115 3.57 49.195 3.8 ;
      RECT 49.045 3.566 49.115 3.831 ;
      RECT 49.035 3.277 49.045 3.345 ;
      RECT 49.035 3.555 49.045 3.861 ;
      RECT 49.025 3.262 49.035 3.49 ;
      RECT 49.025 3.535 49.035 3.925 ;
      RECT 48.815 3.285 48.835 3.925 ;
      RECT 49.615 2.605 49.625 3.345 ;
      RECT 49.435 3.125 49.455 3.345 ;
      RECT 49.445 3.115 49.455 3.345 ;
      RECT 49.945 2.155 49.985 2.415 ;
      RECT 49.935 2.155 49.945 2.425 ;
      RECT 49.901 2.155 49.935 2.452 ;
      RECT 49.815 2.155 49.901 2.512 ;
      RECT 49.795 2.155 49.815 2.575 ;
      RECT 49.735 2.155 49.795 2.74 ;
      RECT 49.725 2.155 49.735 2.9 ;
      RECT 49.695 2.346 49.725 2.995 ;
      RECT 49.685 2.401 49.695 3.095 ;
      RECT 49.675 2.43 49.685 3.14 ;
      RECT 49.665 2.455 49.675 3.173 ;
      RECT 49.655 2.49 49.665 3.228 ;
      RECT 49.635 2.535 49.655 3.29 ;
      RECT 49.625 2.58 49.635 3.34 ;
      RECT 49.605 2.64 49.615 3.345 ;
      RECT 49.595 2.67 49.605 3.345 ;
      RECT 49.575 2.7 49.595 3.345 ;
      RECT 49.525 2.805 49.575 3.345 ;
      RECT 49.515 2.9 49.525 3.345 ;
      RECT 49.505 2.93 49.515 3.345 ;
      RECT 49.48 2.98 49.505 3.345 ;
      RECT 49.475 3.035 49.48 3.345 ;
      RECT 49.455 3.06 49.475 3.345 ;
      RECT 49.415 3.14 49.435 3.335 ;
      RECT 49.165 2.725 49.235 2.935 ;
      RECT 46.405 2.635 46.665 2.895 ;
      RECT 49.235 2.73 49.245 2.93 ;
      RECT 49.121 2.723 49.165 2.935 ;
      RECT 49.035 2.716 49.121 2.935 ;
      RECT 49.015 2.711 49.035 2.925 ;
      RECT 49.005 2.709 49.015 2.905 ;
      RECT 48.955 2.706 49.005 2.9 ;
      RECT 48.925 2.702 48.955 2.895 ;
      RECT 48.905 2.7 48.925 2.89 ;
      RECT 48.865 2.697 48.905 2.885 ;
      RECT 48.795 2.691 48.865 2.88 ;
      RECT 48.765 2.686 48.795 2.875 ;
      RECT 48.745 2.684 48.765 2.87 ;
      RECT 48.715 2.681 48.745 2.865 ;
      RECT 48.655 2.677 48.715 2.86 ;
      RECT 48.585 2.675 48.655 2.85 ;
      RECT 48.551 2.673 48.585 2.843 ;
      RECT 48.465 2.668 48.551 2.835 ;
      RECT 48.431 2.662 48.465 2.827 ;
      RECT 48.345 2.652 48.431 2.819 ;
      RECT 48.311 2.643 48.345 2.811 ;
      RECT 48.225 2.638 48.311 2.803 ;
      RECT 48.155 2.635 48.225 2.793 ;
      RECT 48.135 2.63 48.155 2.787 ;
      RECT 48.131 2.625 48.135 2.786 ;
      RECT 48.045 2.621 48.131 2.781 ;
      RECT 48.005 2.616 48.045 2.774 ;
      RECT 47.925 2.615 48.005 2.769 ;
      RECT 47.905 2.615 47.925 2.766 ;
      RECT 47.879 2.615 47.905 2.766 ;
      RECT 47.793 2.617 47.879 2.77 ;
      RECT 47.707 2.619 47.793 2.777 ;
      RECT 47.621 2.621 47.707 2.783 ;
      RECT 47.535 2.624 47.621 2.79 ;
      RECT 47.501 2.626 47.535 2.795 ;
      RECT 47.415 2.631 47.501 2.8 ;
      RECT 47.391 2.626 47.415 2.804 ;
      RECT 47.305 2.631 47.391 2.809 ;
      RECT 47.267 2.636 47.305 2.814 ;
      RECT 47.181 2.639 47.267 2.819 ;
      RECT 47.095 2.643 47.181 2.826 ;
      RECT 47.031 2.645 47.095 2.832 ;
      RECT 46.945 2.645 47.031 2.838 ;
      RECT 46.861 2.646 46.945 2.845 ;
      RECT 46.775 2.649 46.861 2.852 ;
      RECT 46.751 2.651 46.775 2.856 ;
      RECT 46.665 2.653 46.751 2.861 ;
      RECT 46.395 2.67 46.405 2.865 ;
      RECT 48.58 7.765 48.87 7.995 ;
      RECT 48.64 7.025 48.81 7.995 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 48.58 7.025 48.87 7.425 ;
      RECT 48.635 2.247 48.825 2.455 ;
      RECT 48.625 2.252 48.835 2.45 ;
      RECT 48.615 2.233 48.625 2.445 ;
      RECT 48.585 2.228 48.615 2.44 ;
      RECT 48.545 2.252 48.835 2.43 ;
      RECT 48.325 2.165 48.585 2.425 ;
      RECT 48.625 2.236 48.635 2.45 ;
      RECT 48.325 2.245 48.815 2.425 ;
      RECT 48.325 2.241 48.675 2.425 ;
      RECT 48.275 3.155 48.325 3.435 ;
      RECT 48.205 3.125 48.235 3.435 ;
      RECT 48.345 3.155 48.405 3.415 ;
      RECT 48.205 3.115 48.225 3.435 ;
      RECT 48.325 3.155 48.345 3.425 ;
      RECT 48.245 3.145 48.275 3.435 ;
      RECT 48.235 3.13 48.245 3.435 ;
      RECT 48.185 3.105 48.205 3.435 ;
      RECT 48.155 3.09 48.185 3.435 ;
      RECT 48.145 3.08 48.155 3.435 ;
      RECT 48.125 3.069 48.145 3.43 ;
      RECT 48.105 3.057 48.125 3.4 ;
      RECT 48.095 3.048 48.105 3.383 ;
      RECT 48.065 3.03 48.095 3.375 ;
      RECT 48.055 2.995 48.065 3.367 ;
      RECT 48.045 2.975 48.055 3.36 ;
      RECT 48.035 2.955 48.045 3.353 ;
      RECT 48.025 2.94 48.035 3.348 ;
      RECT 48.015 2.92 48.025 3.343 ;
      RECT 48.005 2.915 48.015 3.338 ;
      RECT 48.001 2.905 48.005 3.334 ;
      RECT 47.915 2.905 48.001 3.309 ;
      RECT 47.885 2.905 47.915 3.275 ;
      RECT 47.875 2.905 47.885 3.255 ;
      RECT 47.815 2.905 47.875 3.2 ;
      RECT 47.805 2.92 47.815 3.145 ;
      RECT 47.795 2.93 47.805 3.125 ;
      RECT 47.745 3.665 48.005 3.925 ;
      RECT 47.665 3.685 48.005 3.901 ;
      RECT 47.645 3.685 48.005 3.896 ;
      RECT 47.621 3.685 48.005 3.894 ;
      RECT 47.535 3.685 48.005 3.889 ;
      RECT 47.385 3.625 47.645 3.885 ;
      RECT 47.345 3.68 47.665 3.88 ;
      RECT 47.335 3.69 48.005 3.875 ;
      RECT 47.355 3.675 47.645 3.885 ;
      RECT 47.245 2.115 47.505 2.375 ;
      RECT 47.245 2.2 47.515 2.3 ;
      RECT 46.415 3.63 46.435 3.874 ;
      RECT 46.415 3.63 46.485 3.869 ;
      RECT 46.395 3.635 46.485 3.868 ;
      RECT 46.385 3.65 46.571 3.858 ;
      RECT 46.385 3.65 46.645 3.855 ;
      RECT 46.38 3.687 46.655 3.845 ;
      RECT 46.38 3.687 46.741 3.841 ;
      RECT 46.38 3.687 46.755 3.827 ;
      RECT 46.655 3.565 46.915 3.825 ;
      RECT 46.375 3.692 46.915 3.82 ;
      RECT 46.365 3.74 46.915 3.795 ;
      RECT 46.635 3.605 46.655 3.854 ;
      RECT 46.571 3.609 46.635 3.857 ;
      RECT 46.435 3.622 46.915 3.825 ;
      RECT 46.485 3.616 46.571 3.862 ;
      RECT 45.885 2.475 45.895 2.645 ;
      RECT 45.945 2.435 45.955 2.615 ;
      RECT 46.245 2.245 46.255 2.455 ;
      RECT 46.575 2.095 46.825 2.355 ;
      RECT 46.565 2.095 46.575 2.357 ;
      RECT 46.555 2.155 46.565 2.361 ;
      RECT 46.525 2.157 46.555 2.369 ;
      RECT 46.495 2.162 46.525 2.383 ;
      RECT 46.485 2.166 46.495 2.393 ;
      RECT 46.455 2.171 46.485 2.405 ;
      RECT 46.425 2.18 46.455 2.406 ;
      RECT 46.355 2.19 46.425 2.41 ;
      RECT 46.315 2.195 46.355 2.414 ;
      RECT 46.295 2.195 46.315 2.425 ;
      RECT 46.285 2.2 46.295 2.435 ;
      RECT 46.275 2.21 46.285 2.438 ;
      RECT 46.265 2.23 46.275 2.443 ;
      RECT 46.255 2.24 46.265 2.445 ;
      RECT 46.225 2.255 46.245 2.462 ;
      RECT 46.215 2.267 46.225 2.472 ;
      RECT 46.205 2.273 46.215 2.475 ;
      RECT 46.171 2.286 46.205 2.485 ;
      RECT 46.085 2.32 46.171 2.518 ;
      RECT 46.065 2.355 46.085 2.547 ;
      RECT 46.045 2.37 46.065 2.559 ;
      RECT 46.025 2.38 46.045 2.571 ;
      RECT 45.975 2.399 46.025 2.591 ;
      RECT 45.965 2.416 45.975 2.605 ;
      RECT 45.955 2.422 45.965 2.61 ;
      RECT 45.935 2.44 45.945 2.618 ;
      RECT 45.925 2.445 45.935 2.625 ;
      RECT 45.915 2.456 45.925 2.632 ;
      RECT 45.895 2.461 45.915 2.64 ;
      RECT 45.875 2.475 45.885 2.65 ;
      RECT 45.865 2.48 45.875 2.66 ;
      RECT 45.835 2.494 45.865 2.67 ;
      RECT 45.825 2.507 45.835 2.68 ;
      RECT 45.745 2.538 45.825 2.705 ;
      RECT 45.725 2.568 45.745 2.73 ;
      RECT 45.715 2.573 45.725 2.737 ;
      RECT 45.685 2.585 45.715 2.743 ;
      RECT 45.675 2.6 45.685 2.749 ;
      RECT 45.665 2.605 45.675 2.752 ;
      RECT 45.645 2.615 45.665 2.756 ;
      RECT 45.625 2.62 45.645 2.762 ;
      RECT 45.595 2.625 45.625 2.77 ;
      RECT 45.565 2.63 45.595 2.78 ;
      RECT 45.535 2.64 45.565 2.789 ;
      RECT 45.495 2.645 45.535 2.797 ;
      RECT 45.445 2.638 45.495 2.809 ;
      RECT 45.425 2.629 45.445 2.82 ;
      RECT 45.415 2.626 45.425 2.825 ;
      RECT 45.375 2.625 45.415 2.826 ;
      RECT 45.365 2.61 45.375 2.827 ;
      RECT 45.337 2.595 45.365 2.828 ;
      RECT 45.251 2.595 45.337 2.83 ;
      RECT 45.165 2.595 45.251 2.834 ;
      RECT 45.145 2.595 45.165 2.83 ;
      RECT 45.135 2.605 45.145 2.823 ;
      RECT 45.125 2.62 45.135 2.818 ;
      RECT 45.115 2.625 45.125 2.795 ;
      RECT 46.595 3.13 46.605 3.33 ;
      RECT 46.545 3.125 46.595 3.35 ;
      RECT 46.535 3.125 46.545 3.37 ;
      RECT 46.491 3.125 46.535 3.374 ;
      RECT 46.405 3.125 46.491 3.371 ;
      RECT 46.345 3.135 46.405 3.368 ;
      RECT 46.285 3.149 46.345 3.366 ;
      RECT 46.275 3.154 46.285 3.364 ;
      RECT 46.265 3.16 46.275 3.363 ;
      RECT 46.195 3.173 46.265 3.359 ;
      RECT 46.147 3.187 46.195 3.36 ;
      RECT 46.061 3.203 46.147 3.372 ;
      RECT 45.975 3.224 46.061 3.388 ;
      RECT 45.955 3.235 45.975 3.398 ;
      RECT 45.875 3.245 45.955 3.408 ;
      RECT 45.841 3.259 45.875 3.42 ;
      RECT 45.755 3.274 45.841 3.435 ;
      RECT 45.725 3.29 45.755 3.445 ;
      RECT 45.67 3.305 45.725 3.456 ;
      RECT 45.625 3.323 45.67 3.476 ;
      RECT 45.571 3.342 45.625 3.496 ;
      RECT 45.485 3.368 45.571 3.523 ;
      RECT 45.465 3.39 45.485 3.543 ;
      RECT 45.405 3.405 45.465 3.559 ;
      RECT 45.395 3.42 45.405 3.573 ;
      RECT 45.375 3.425 45.395 3.579 ;
      RECT 45.345 3.438 45.375 3.589 ;
      RECT 45.325 3.443 45.345 3.598 ;
      RECT 45.315 3.45 45.325 3.603 ;
      RECT 45.305 3.455 45.315 3.606 ;
      RECT 45.265 3.465 45.305 3.615 ;
      RECT 45.24 3.48 45.265 3.627 ;
      RECT 45.195 3.495 45.24 3.639 ;
      RECT 45.175 3.507 45.195 3.651 ;
      RECT 45.145 3.512 45.175 3.661 ;
      RECT 45.125 3.519 45.145 3.671 ;
      RECT 45.115 3.525 45.125 3.68 ;
      RECT 45.091 3.532 45.115 3.69 ;
      RECT 45.005 3.554 45.091 3.71 ;
      RECT 44.995 3.573 45.005 3.725 ;
      RECT 44.971 3.58 44.995 3.731 ;
      RECT 44.885 3.602 44.971 3.756 ;
      RECT 44.845 3.627 44.885 3.783 ;
      RECT 44.835 3.636 44.845 3.793 ;
      RECT 44.785 3.646 44.835 3.802 ;
      RECT 44.765 3.66 44.785 3.812 ;
      RECT 44.735 3.67 44.765 3.817 ;
      RECT 44.725 3.675 44.735 3.82 ;
      RECT 44.651 3.677 44.725 3.827 ;
      RECT 44.565 3.681 44.651 3.839 ;
      RECT 44.555 3.684 44.565 3.845 ;
      RECT 44.295 3.635 44.555 3.895 ;
      RECT 45.825 3.705 46.015 3.915 ;
      RECT 45.815 3.71 46.025 3.91 ;
      RECT 45.805 3.71 46.025 3.875 ;
      RECT 45.725 3.595 45.985 3.855 ;
      RECT 44.635 3.125 44.825 3.425 ;
      RECT 44.625 3.125 44.825 3.42 ;
      RECT 44.615 3.125 44.835 3.415 ;
      RECT 44.605 3.125 44.835 3.41 ;
      RECT 44.605 3.125 44.865 3.385 ;
      RECT 44.565 2.165 44.825 2.425 ;
      RECT 44.375 2.09 44.461 2.423 ;
      RECT 44.375 2.09 44.505 2.419 ;
      RECT 44.355 2.094 44.515 2.418 ;
      RECT 44.505 2.085 44.515 2.418 ;
      RECT 44.375 2.09 44.525 2.417 ;
      RECT 44.355 2.1 44.565 2.416 ;
      RECT 44.345 2.095 44.525 2.408 ;
      RECT 44.335 2.11 44.565 2.315 ;
      RECT 44.335 2.16 44.765 2.315 ;
      RECT 44.335 2.15 44.745 2.315 ;
      RECT 44.335 2.14 44.715 2.315 ;
      RECT 44.335 2.13 44.655 2.315 ;
      RECT 44.335 2.115 44.635 2.315 ;
      RECT 44.461 2.086 44.515 2.418 ;
      RECT 43.535 2.745 43.675 3.035 ;
      RECT 43.795 2.768 43.805 2.955 ;
      RECT 44.495 2.665 44.675 2.895 ;
      RECT 44.495 2.665 44.685 2.885 ;
      RECT 44.705 2.67 44.715 2.875 ;
      RECT 44.685 2.665 44.705 2.88 ;
      RECT 44.445 2.669 44.495 2.895 ;
      RECT 44.435 2.674 44.445 2.895 ;
      RECT 44.401 2.679 44.435 2.896 ;
      RECT 44.315 2.694 44.401 2.898 ;
      RECT 44.301 2.706 44.315 2.901 ;
      RECT 44.215 2.716 44.301 2.903 ;
      RECT 44.191 2.726 44.215 2.905 ;
      RECT 44.105 2.737 44.191 2.905 ;
      RECT 44.075 2.747 44.105 2.905 ;
      RECT 44.045 2.752 44.075 2.908 ;
      RECT 44.025 2.757 44.045 2.913 ;
      RECT 44.005 2.762 44.025 2.915 ;
      RECT 43.955 2.77 44.005 2.915 ;
      RECT 43.935 2.774 43.955 2.915 ;
      RECT 43.915 2.773 43.935 2.92 ;
      RECT 43.855 2.771 43.915 2.935 ;
      RECT 43.805 2.769 43.855 2.95 ;
      RECT 43.715 2.766 43.795 3.035 ;
      RECT 43.685 2.76 43.715 3.035 ;
      RECT 43.675 2.75 43.685 3.035 ;
      RECT 43.485 2.745 43.535 2.96 ;
      RECT 43.475 2.75 43.485 2.95 ;
      RECT 43.715 3.225 43.975 3.485 ;
      RECT 43.715 3.225 44.005 3.375 ;
      RECT 43.715 3.225 44.045 3.36 ;
      RECT 43.975 3.145 44.165 3.355 ;
      RECT 43.975 3.15 44.175 3.345 ;
      RECT 43.925 3.22 44.175 3.345 ;
      RECT 43.955 3.155 43.975 3.485 ;
      RECT 43.945 3.18 44.175 3.345 ;
      RECT 43.125 3.125 43.135 3.355 ;
      RECT 43.025 2.245 43.095 3.355 ;
      RECT 43.765 2.355 44.025 2.615 ;
      RECT 43.465 2.405 43.595 2.565 ;
      RECT 43.681 2.412 43.765 2.565 ;
      RECT 43.595 2.407 43.681 2.565 ;
      RECT 43.405 2.405 43.465 2.575 ;
      RECT 43.375 2.403 43.405 2.59 ;
      RECT 43.355 2.401 43.375 2.6 ;
      RECT 43.345 2.399 43.355 2.605 ;
      RECT 43.325 2.398 43.345 2.615 ;
      RECT 43.315 2.396 43.325 2.62 ;
      RECT 43.295 2.395 43.315 2.625 ;
      RECT 43.275 2.39 43.295 2.63 ;
      RECT 43.245 2.376 43.275 2.64 ;
      RECT 43.205 2.355 43.245 2.655 ;
      RECT 43.195 2.34 43.205 2.665 ;
      RECT 43.175 2.331 43.195 2.675 ;
      RECT 43.165 2.322 43.175 2.695 ;
      RECT 43.155 2.317 43.165 2.755 ;
      RECT 43.135 2.311 43.155 2.84 ;
      RECT 43.135 3.15 43.145 3.35 ;
      RECT 43.125 2.306 43.135 3.07 ;
      RECT 43.115 2.28 43.125 3.355 ;
      RECT 43.095 2.25 43.115 3.355 ;
      RECT 43.005 2.245 43.025 2.58 ;
      RECT 43.015 2.68 43.025 3.355 ;
      RECT 43.005 2.72 43.015 3.355 ;
      RECT 42.975 2.245 43.005 2.525 ;
      RECT 42.985 2.81 43.005 3.355 ;
      RECT 42.97 2.915 42.985 3.355 ;
      RECT 42.945 2.245 42.975 2.48 ;
      RECT 42.965 2.947 42.97 3.355 ;
      RECT 42.945 3.05 42.965 3.355 ;
      RECT 42.935 2.245 42.945 2.47 ;
      RECT 42.935 3.12 42.945 3.35 ;
      RECT 42.915 2.245 42.935 2.46 ;
      RECT 42.905 2.25 42.915 2.45 ;
      RECT 43.115 3.525 43.135 3.765 ;
      RECT 42.435 3.455 42.515 3.725 ;
      RECT 42.345 3.455 42.355 3.665 ;
      RECT 43.625 3.525 43.635 3.725 ;
      RECT 43.545 3.515 43.625 3.75 ;
      RECT 43.541 3.515 43.545 3.776 ;
      RECT 43.455 3.515 43.541 3.786 ;
      RECT 43.435 3.515 43.455 3.794 ;
      RECT 43.411 3.516 43.435 3.792 ;
      RECT 43.325 3.521 43.411 3.787 ;
      RECT 43.307 3.525 43.325 3.781 ;
      RECT 43.221 3.525 43.307 3.777 ;
      RECT 43.135 3.525 43.221 3.769 ;
      RECT 43.031 3.525 43.115 3.762 ;
      RECT 42.945 3.525 43.031 3.756 ;
      RECT 42.885 3.52 42.945 3.75 ;
      RECT 42.857 3.514 42.885 3.747 ;
      RECT 42.771 3.511 42.857 3.744 ;
      RECT 42.685 3.507 42.771 3.738 ;
      RECT 42.64 3.495 42.685 3.734 ;
      RECT 42.615 3.48 42.64 3.732 ;
      RECT 42.575 3.465 42.615 3.73 ;
      RECT 42.515 3.455 42.575 3.727 ;
      RECT 42.425 3.455 42.435 3.72 ;
      RECT 42.41 3.455 42.425 3.71 ;
      RECT 42.355 3.455 42.41 3.685 ;
      RECT 42.335 3.47 42.345 3.66 ;
      RECT 42.465 2.635 42.725 2.895 ;
      RECT 42.465 2.645 42.745 2.855 ;
      RECT 42.465 2.65 42.755 2.85 ;
      RECT 40.445 2.115 40.705 2.375 ;
      RECT 40.435 2.145 40.705 2.355 ;
      RECT 42.365 2.055 42.615 2.315 ;
      RECT 42.355 2.055 42.365 2.316 ;
      RECT 42.325 2.14 42.355 2.318 ;
      RECT 42.315 2.145 42.325 2.32 ;
      RECT 42.255 2.16 42.315 2.326 ;
      RECT 42.225 2.18 42.255 2.333 ;
      RECT 42.195 2.191 42.225 2.34 ;
      RECT 42.175 2.201 42.195 2.345 ;
      RECT 42.157 2.204 42.175 2.344 ;
      RECT 42.071 2.203 42.157 2.344 ;
      RECT 41.985 2.2 42.071 2.343 ;
      RECT 41.899 2.197 41.985 2.342 ;
      RECT 41.813 2.194 41.899 2.342 ;
      RECT 41.727 2.192 41.813 2.341 ;
      RECT 41.641 2.189 41.727 2.34 ;
      RECT 41.555 2.186 41.641 2.34 ;
      RECT 41.537 2.185 41.555 2.339 ;
      RECT 41.451 2.184 41.537 2.339 ;
      RECT 41.365 2.182 41.451 2.338 ;
      RECT 41.279 2.181 41.365 2.338 ;
      RECT 41.193 2.18 41.279 2.337 ;
      RECT 41.107 2.178 41.193 2.337 ;
      RECT 41.021 2.177 41.107 2.336 ;
      RECT 40.935 2.175 41.021 2.336 ;
      RECT 40.911 2.174 40.935 2.335 ;
      RECT 40.825 2.169 40.911 2.335 ;
      RECT 40.791 2.162 40.825 2.335 ;
      RECT 40.705 2.152 40.791 2.335 ;
      RECT 40.425 2.15 40.435 2.35 ;
      RECT 41.705 3.205 41.965 3.465 ;
      RECT 41.705 3.205 42.045 3.251 ;
      RECT 41.845 3.185 42.055 3.24 ;
      RECT 41.905 3.16 42.115 3.2 ;
      RECT 41.915 3.155 42.115 3.2 ;
      RECT 41.925 3.13 42.115 3.2 ;
      RECT 41.985 2.96 42.035 3.29 ;
      RECT 41.935 3.09 42.125 3.15 ;
      RECT 41.975 3.016 41.985 3.329 ;
      RECT 41.935 3.09 42.155 3.125 ;
      RECT 41.935 3.09 42.175 3.1 ;
      RECT 42.045 2.89 42.235 3.095 ;
      RECT 42.035 2.9 42.245 3.09 ;
      RECT 41.955 3.063 42.245 3.09 ;
      RECT 41.965 3.039 41.975 3.345 ;
      RECT 42.055 2.885 42.225 3.095 ;
      RECT 41.345 2.675 41.535 2.885 ;
      RECT 39.915 2.605 40.175 2.865 ;
      RECT 40.265 2.595 40.365 2.805 ;
      RECT 40.215 2.615 40.255 2.805 ;
      RECT 41.535 2.685 41.545 2.88 ;
      RECT 41.335 2.685 41.345 2.88 ;
      RECT 41.315 2.7 41.335 2.87 ;
      RECT 41.305 2.71 41.315 2.865 ;
      RECT 41.265 2.71 41.305 2.863 ;
      RECT 41.241 2.704 41.265 2.86 ;
      RECT 41.155 2.699 41.241 2.857 ;
      RECT 41.095 2.695 41.155 2.852 ;
      RECT 41.061 2.692 41.095 2.849 ;
      RECT 40.975 2.682 41.061 2.845 ;
      RECT 40.971 2.675 40.975 2.842 ;
      RECT 40.885 2.67 40.971 2.84 ;
      RECT 40.857 2.663 40.885 2.836 ;
      RECT 40.771 2.658 40.857 2.833 ;
      RECT 40.685 2.649 40.771 2.828 ;
      RECT 40.675 2.644 40.685 2.825 ;
      RECT 40.661 2.643 40.675 2.825 ;
      RECT 40.575 2.639 40.661 2.82 ;
      RECT 40.555 2.633 40.575 2.816 ;
      RECT 40.495 2.628 40.555 2.815 ;
      RECT 40.465 2.62 40.495 2.815 ;
      RECT 40.455 2.605 40.465 2.815 ;
      RECT 40.451 2.595 40.455 2.814 ;
      RECT 40.365 2.595 40.451 2.81 ;
      RECT 40.255 2.605 40.265 2.805 ;
      RECT 40.185 2.615 40.215 2.8 ;
      RECT 40.175 2.615 40.185 2.8 ;
      RECT 41.095 3.115 41.355 3.375 ;
      RECT 41.025 3.125 41.355 3.335 ;
      RECT 41.015 3.13 41.355 3.33 ;
      RECT 40.435 3.115 40.695 3.375 ;
      RECT 40.435 3.16 40.805 3.365 ;
      RECT 40.435 3.155 40.795 3.365 ;
      RECT 39.345 3.322 39.525 3.765 ;
      RECT 39.335 3.322 39.525 3.763 ;
      RECT 39.335 3.337 39.535 3.76 ;
      RECT 39.325 2.26 39.455 3.758 ;
      RECT 39.325 3.385 39.595 3.645 ;
      RECT 39.325 3.36 39.545 3.645 ;
      RECT 39.325 3.295 39.515 3.758 ;
      RECT 39.325 3.255 39.485 3.758 ;
      RECT 39.325 3.21 39.475 3.758 ;
      RECT 39.325 3.15 39.465 3.758 ;
      RECT 39.315 2.545 39.455 3.2 ;
      RECT 39.355 2.245 39.465 3.065 ;
      RECT 39.325 2.26 39.505 2.52 ;
      RECT 39.325 2.26 39.515 2.47 ;
      RECT 39.355 2.245 39.525 2.463 ;
      RECT 39.345 2.247 39.535 2.458 ;
      RECT 39.335 2.252 39.545 2.45 ;
      RECT 38.195 7.77 38.485 8 ;
      RECT 38.255 6.29 38.425 8 ;
      RECT 38.245 6.66 38.6 7.015 ;
      RECT 38.195 6.29 38.485 6.52 ;
      RECT 37.79 2.395 37.895 2.965 ;
      RECT 37.79 2.73 38.115 2.96 ;
      RECT 37.79 2.76 38.285 2.93 ;
      RECT 37.79 2.395 37.98 2.96 ;
      RECT 37.205 2.36 37.495 2.59 ;
      RECT 37.205 2.395 37.98 2.565 ;
      RECT 37.265 0.88 37.435 2.59 ;
      RECT 37.205 0.88 37.495 1.11 ;
      RECT 37.205 7.77 37.495 8 ;
      RECT 37.265 6.29 37.435 8 ;
      RECT 37.205 6.29 37.495 6.52 ;
      RECT 37.205 6.325 38.06 6.485 ;
      RECT 37.89 5.92 38.06 6.485 ;
      RECT 37.205 6.32 37.6 6.485 ;
      RECT 37.825 5.92 38.115 6.15 ;
      RECT 37.825 5.95 38.285 6.12 ;
      RECT 36.835 2.73 37.125 2.96 ;
      RECT 36.835 2.76 37.295 2.93 ;
      RECT 36.9 1.655 37.065 2.96 ;
      RECT 35.415 1.625 35.705 1.855 ;
      RECT 35.415 1.655 37.065 1.825 ;
      RECT 35.475 0.885 35.645 1.855 ;
      RECT 35.415 0.885 35.705 1.115 ;
      RECT 35.415 7.765 35.705 7.995 ;
      RECT 35.475 7.025 35.645 7.995 ;
      RECT 35.475 7.12 37.065 7.29 ;
      RECT 36.895 5.92 37.065 7.29 ;
      RECT 35.415 7.025 35.705 7.255 ;
      RECT 36.835 5.92 37.125 6.15 ;
      RECT 36.835 5.95 37.295 6.12 ;
      RECT 33.45 3.43 33.8 3.78 ;
      RECT 33.54 2.025 33.71 3.78 ;
      RECT 35.845 1.965 36.195 2.315 ;
      RECT 33.54 2.025 35.16 2.2 ;
      RECT 33.54 2.025 36.195 2.195 ;
      RECT 35.87 6.655 36.195 6.98 ;
      RECT 31.295 6.61 31.645 6.96 ;
      RECT 35.845 6.655 36.195 6.885 ;
      RECT 31.085 6.655 31.645 6.885 ;
      RECT 30.915 6.685 36.195 6.855 ;
      RECT 35.07 2.365 35.39 2.685 ;
      RECT 35.04 2.365 35.39 2.595 ;
      RECT 34.87 2.395 35.39 2.565 ;
      RECT 35.07 6.225 35.39 6.545 ;
      RECT 35.04 6.285 35.39 6.515 ;
      RECT 34.87 6.315 35.39 6.485 ;
      RECT 30.91 3.255 31.1 3.925 ;
      RECT 30.85 3.665 30.89 3.925 ;
      RECT 32.22 2.89 32.23 3.111 ;
      RECT 32.15 2.885 32.22 3.236 ;
      RECT 32.14 2.885 32.15 3.36 ;
      RECT 32.11 2.885 32.14 3.41 ;
      RECT 32.09 2.885 32.11 3.485 ;
      RECT 32.07 2.885 32.09 3.555 ;
      RECT 32.04 2.885 32.07 3.595 ;
      RECT 32.03 2.885 32.04 3.615 ;
      RECT 32.02 2.885 32.03 3.626 ;
      RECT 32.01 3.135 32.02 3.628 ;
      RECT 32 3.2 32.01 3.63 ;
      RECT 31.99 3.295 32 3.632 ;
      RECT 31.98 3.37 31.99 3.634 ;
      RECT 31.93 3.394 31.98 3.64 ;
      RECT 31.89 3.429 31.93 3.649 ;
      RECT 31.88 3.445 31.89 3.654 ;
      RECT 31.866 3.45 31.88 3.657 ;
      RECT 31.78 3.49 31.866 3.668 ;
      RECT 31.7 3.533 31.78 3.686 ;
      RECT 31.68 3.543 31.7 3.697 ;
      RECT 31.65 3.551 31.68 3.702 ;
      RECT 31.63 3.561 31.65 3.707 ;
      RECT 31.606 3.567 31.63 3.712 ;
      RECT 31.52 3.577 31.606 3.725 ;
      RECT 31.442 3.583 31.52 3.745 ;
      RECT 31.356 3.578 31.442 3.764 ;
      RECT 31.27 3.574 31.356 3.785 ;
      RECT 31.19 3.57 31.27 3.8 ;
      RECT 31.12 3.566 31.19 3.831 ;
      RECT 31.11 3.277 31.12 3.345 ;
      RECT 31.11 3.555 31.12 3.861 ;
      RECT 31.1 3.262 31.11 3.49 ;
      RECT 31.1 3.535 31.11 3.925 ;
      RECT 30.89 3.285 30.91 3.925 ;
      RECT 31.69 2.605 31.7 3.345 ;
      RECT 31.51 3.125 31.53 3.345 ;
      RECT 31.52 3.115 31.53 3.345 ;
      RECT 32.02 2.155 32.06 2.415 ;
      RECT 32.01 2.155 32.02 2.425 ;
      RECT 31.976 2.155 32.01 2.452 ;
      RECT 31.89 2.155 31.976 2.512 ;
      RECT 31.87 2.155 31.89 2.575 ;
      RECT 31.81 2.155 31.87 2.74 ;
      RECT 31.8 2.155 31.81 2.9 ;
      RECT 31.77 2.346 31.8 2.995 ;
      RECT 31.76 2.401 31.77 3.095 ;
      RECT 31.75 2.43 31.76 3.14 ;
      RECT 31.74 2.455 31.75 3.173 ;
      RECT 31.73 2.49 31.74 3.228 ;
      RECT 31.71 2.535 31.73 3.29 ;
      RECT 31.7 2.58 31.71 3.34 ;
      RECT 31.68 2.64 31.69 3.345 ;
      RECT 31.67 2.67 31.68 3.345 ;
      RECT 31.65 2.7 31.67 3.345 ;
      RECT 31.6 2.805 31.65 3.345 ;
      RECT 31.59 2.9 31.6 3.345 ;
      RECT 31.58 2.93 31.59 3.345 ;
      RECT 31.555 2.98 31.58 3.345 ;
      RECT 31.55 3.035 31.555 3.345 ;
      RECT 31.53 3.06 31.55 3.345 ;
      RECT 31.49 3.14 31.51 3.335 ;
      RECT 31.24 2.725 31.31 2.935 ;
      RECT 28.48 2.635 28.74 2.895 ;
      RECT 31.31 2.73 31.32 2.93 ;
      RECT 31.196 2.723 31.24 2.935 ;
      RECT 31.11 2.716 31.196 2.935 ;
      RECT 31.09 2.711 31.11 2.925 ;
      RECT 31.08 2.709 31.09 2.905 ;
      RECT 31.03 2.706 31.08 2.9 ;
      RECT 31 2.702 31.03 2.895 ;
      RECT 30.98 2.7 31 2.89 ;
      RECT 30.94 2.697 30.98 2.885 ;
      RECT 30.87 2.691 30.94 2.88 ;
      RECT 30.84 2.686 30.87 2.875 ;
      RECT 30.82 2.684 30.84 2.87 ;
      RECT 30.79 2.681 30.82 2.865 ;
      RECT 30.73 2.677 30.79 2.86 ;
      RECT 30.66 2.675 30.73 2.85 ;
      RECT 30.626 2.673 30.66 2.843 ;
      RECT 30.54 2.668 30.626 2.835 ;
      RECT 30.506 2.662 30.54 2.827 ;
      RECT 30.42 2.652 30.506 2.819 ;
      RECT 30.386 2.643 30.42 2.811 ;
      RECT 30.3 2.638 30.386 2.803 ;
      RECT 30.23 2.635 30.3 2.793 ;
      RECT 30.21 2.63 30.23 2.787 ;
      RECT 30.206 2.625 30.21 2.786 ;
      RECT 30.12 2.621 30.206 2.781 ;
      RECT 30.08 2.616 30.12 2.774 ;
      RECT 30 2.615 30.08 2.769 ;
      RECT 29.98 2.615 30 2.766 ;
      RECT 29.954 2.615 29.98 2.766 ;
      RECT 29.868 2.617 29.954 2.77 ;
      RECT 29.782 2.619 29.868 2.777 ;
      RECT 29.696 2.621 29.782 2.783 ;
      RECT 29.61 2.624 29.696 2.79 ;
      RECT 29.576 2.626 29.61 2.795 ;
      RECT 29.49 2.631 29.576 2.8 ;
      RECT 29.466 2.626 29.49 2.804 ;
      RECT 29.38 2.631 29.466 2.809 ;
      RECT 29.342 2.636 29.38 2.814 ;
      RECT 29.256 2.639 29.342 2.819 ;
      RECT 29.17 2.643 29.256 2.826 ;
      RECT 29.106 2.645 29.17 2.832 ;
      RECT 29.02 2.645 29.106 2.838 ;
      RECT 28.936 2.646 29.02 2.845 ;
      RECT 28.85 2.649 28.936 2.852 ;
      RECT 28.826 2.651 28.85 2.856 ;
      RECT 28.74 2.653 28.826 2.861 ;
      RECT 28.47 2.67 28.48 2.865 ;
      RECT 30.655 7.765 30.945 7.995 ;
      RECT 30.715 7.025 30.885 7.995 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 30.655 7.025 30.945 7.425 ;
      RECT 30.71 2.247 30.9 2.455 ;
      RECT 30.7 2.252 30.91 2.45 ;
      RECT 30.69 2.233 30.7 2.445 ;
      RECT 30.66 2.228 30.69 2.44 ;
      RECT 30.62 2.252 30.91 2.43 ;
      RECT 30.4 2.165 30.66 2.425 ;
      RECT 30.7 2.236 30.71 2.45 ;
      RECT 30.4 2.245 30.89 2.425 ;
      RECT 30.4 2.241 30.75 2.425 ;
      RECT 30.35 3.155 30.4 3.435 ;
      RECT 30.28 3.125 30.31 3.435 ;
      RECT 30.42 3.155 30.48 3.415 ;
      RECT 30.28 3.115 30.3 3.435 ;
      RECT 30.4 3.155 30.42 3.425 ;
      RECT 30.32 3.145 30.35 3.435 ;
      RECT 30.31 3.13 30.32 3.435 ;
      RECT 30.26 3.105 30.28 3.435 ;
      RECT 30.23 3.09 30.26 3.435 ;
      RECT 30.22 3.08 30.23 3.435 ;
      RECT 30.2 3.069 30.22 3.43 ;
      RECT 30.18 3.057 30.2 3.4 ;
      RECT 30.17 3.048 30.18 3.383 ;
      RECT 30.14 3.03 30.17 3.375 ;
      RECT 30.13 2.995 30.14 3.367 ;
      RECT 30.12 2.975 30.13 3.36 ;
      RECT 30.11 2.955 30.12 3.353 ;
      RECT 30.1 2.94 30.11 3.348 ;
      RECT 30.09 2.92 30.1 3.343 ;
      RECT 30.08 2.915 30.09 3.338 ;
      RECT 30.076 2.905 30.08 3.334 ;
      RECT 29.99 2.905 30.076 3.309 ;
      RECT 29.96 2.905 29.99 3.275 ;
      RECT 29.95 2.905 29.96 3.255 ;
      RECT 29.89 2.905 29.95 3.2 ;
      RECT 29.88 2.92 29.89 3.145 ;
      RECT 29.87 2.93 29.88 3.125 ;
      RECT 29.82 3.665 30.08 3.925 ;
      RECT 29.74 3.685 30.08 3.901 ;
      RECT 29.72 3.685 30.08 3.896 ;
      RECT 29.696 3.685 30.08 3.894 ;
      RECT 29.61 3.685 30.08 3.889 ;
      RECT 29.46 3.625 29.72 3.885 ;
      RECT 29.42 3.68 29.74 3.88 ;
      RECT 29.41 3.69 30.08 3.875 ;
      RECT 29.43 3.675 29.72 3.885 ;
      RECT 29.32 2.115 29.58 2.375 ;
      RECT 29.32 2.2 29.59 2.3 ;
      RECT 28.49 3.63 28.51 3.874 ;
      RECT 28.49 3.63 28.56 3.869 ;
      RECT 28.47 3.635 28.56 3.868 ;
      RECT 28.46 3.65 28.646 3.858 ;
      RECT 28.46 3.65 28.72 3.855 ;
      RECT 28.455 3.687 28.73 3.845 ;
      RECT 28.455 3.687 28.816 3.841 ;
      RECT 28.455 3.687 28.83 3.827 ;
      RECT 28.73 3.565 28.99 3.825 ;
      RECT 28.45 3.692 28.99 3.82 ;
      RECT 28.44 3.74 28.99 3.795 ;
      RECT 28.71 3.605 28.73 3.854 ;
      RECT 28.646 3.609 28.71 3.857 ;
      RECT 28.51 3.622 28.99 3.825 ;
      RECT 28.56 3.616 28.646 3.862 ;
      RECT 27.96 2.475 27.97 2.645 ;
      RECT 28.02 2.435 28.03 2.615 ;
      RECT 28.32 2.245 28.33 2.455 ;
      RECT 28.65 2.095 28.9 2.355 ;
      RECT 28.64 2.095 28.65 2.357 ;
      RECT 28.63 2.155 28.64 2.361 ;
      RECT 28.6 2.157 28.63 2.369 ;
      RECT 28.57 2.162 28.6 2.383 ;
      RECT 28.56 2.166 28.57 2.393 ;
      RECT 28.53 2.171 28.56 2.405 ;
      RECT 28.5 2.18 28.53 2.406 ;
      RECT 28.43 2.19 28.5 2.41 ;
      RECT 28.39 2.195 28.43 2.414 ;
      RECT 28.37 2.195 28.39 2.425 ;
      RECT 28.36 2.2 28.37 2.435 ;
      RECT 28.35 2.21 28.36 2.438 ;
      RECT 28.34 2.23 28.35 2.443 ;
      RECT 28.33 2.24 28.34 2.445 ;
      RECT 28.3 2.255 28.32 2.462 ;
      RECT 28.29 2.267 28.3 2.472 ;
      RECT 28.28 2.273 28.29 2.475 ;
      RECT 28.246 2.286 28.28 2.485 ;
      RECT 28.16 2.32 28.246 2.518 ;
      RECT 28.14 2.355 28.16 2.547 ;
      RECT 28.12 2.37 28.14 2.559 ;
      RECT 28.1 2.38 28.12 2.571 ;
      RECT 28.05 2.399 28.1 2.591 ;
      RECT 28.04 2.416 28.05 2.605 ;
      RECT 28.03 2.422 28.04 2.61 ;
      RECT 28.01 2.44 28.02 2.618 ;
      RECT 28 2.445 28.01 2.625 ;
      RECT 27.99 2.456 28 2.632 ;
      RECT 27.97 2.461 27.99 2.64 ;
      RECT 27.95 2.475 27.96 2.65 ;
      RECT 27.94 2.48 27.95 2.66 ;
      RECT 27.91 2.494 27.94 2.67 ;
      RECT 27.9 2.507 27.91 2.68 ;
      RECT 27.82 2.538 27.9 2.705 ;
      RECT 27.8 2.568 27.82 2.73 ;
      RECT 27.79 2.573 27.8 2.737 ;
      RECT 27.76 2.585 27.79 2.743 ;
      RECT 27.75 2.6 27.76 2.749 ;
      RECT 27.74 2.605 27.75 2.752 ;
      RECT 27.72 2.615 27.74 2.756 ;
      RECT 27.7 2.62 27.72 2.762 ;
      RECT 27.67 2.625 27.7 2.77 ;
      RECT 27.64 2.63 27.67 2.78 ;
      RECT 27.61 2.64 27.64 2.789 ;
      RECT 27.57 2.645 27.61 2.797 ;
      RECT 27.52 2.638 27.57 2.809 ;
      RECT 27.5 2.629 27.52 2.82 ;
      RECT 27.49 2.626 27.5 2.825 ;
      RECT 27.45 2.625 27.49 2.826 ;
      RECT 27.44 2.61 27.45 2.827 ;
      RECT 27.412 2.595 27.44 2.828 ;
      RECT 27.326 2.595 27.412 2.83 ;
      RECT 27.24 2.595 27.326 2.834 ;
      RECT 27.22 2.595 27.24 2.83 ;
      RECT 27.21 2.605 27.22 2.823 ;
      RECT 27.2 2.62 27.21 2.818 ;
      RECT 27.19 2.625 27.2 2.795 ;
      RECT 28.67 3.13 28.68 3.33 ;
      RECT 28.62 3.125 28.67 3.35 ;
      RECT 28.61 3.125 28.62 3.37 ;
      RECT 28.566 3.125 28.61 3.374 ;
      RECT 28.48 3.125 28.566 3.371 ;
      RECT 28.42 3.135 28.48 3.368 ;
      RECT 28.36 3.149 28.42 3.366 ;
      RECT 28.35 3.154 28.36 3.364 ;
      RECT 28.34 3.16 28.35 3.363 ;
      RECT 28.27 3.173 28.34 3.359 ;
      RECT 28.222 3.187 28.27 3.36 ;
      RECT 28.136 3.203 28.222 3.372 ;
      RECT 28.05 3.224 28.136 3.388 ;
      RECT 28.03 3.235 28.05 3.398 ;
      RECT 27.95 3.245 28.03 3.408 ;
      RECT 27.916 3.259 27.95 3.42 ;
      RECT 27.83 3.274 27.916 3.435 ;
      RECT 27.8 3.29 27.83 3.445 ;
      RECT 27.745 3.305 27.8 3.456 ;
      RECT 27.7 3.323 27.745 3.476 ;
      RECT 27.646 3.342 27.7 3.496 ;
      RECT 27.56 3.368 27.646 3.523 ;
      RECT 27.54 3.39 27.56 3.543 ;
      RECT 27.48 3.405 27.54 3.559 ;
      RECT 27.47 3.42 27.48 3.573 ;
      RECT 27.45 3.425 27.47 3.579 ;
      RECT 27.42 3.438 27.45 3.589 ;
      RECT 27.4 3.443 27.42 3.598 ;
      RECT 27.39 3.45 27.4 3.603 ;
      RECT 27.38 3.455 27.39 3.606 ;
      RECT 27.34 3.465 27.38 3.615 ;
      RECT 27.315 3.48 27.34 3.627 ;
      RECT 27.27 3.495 27.315 3.639 ;
      RECT 27.25 3.507 27.27 3.651 ;
      RECT 27.22 3.512 27.25 3.661 ;
      RECT 27.2 3.519 27.22 3.671 ;
      RECT 27.19 3.525 27.2 3.68 ;
      RECT 27.166 3.532 27.19 3.69 ;
      RECT 27.08 3.554 27.166 3.71 ;
      RECT 27.07 3.573 27.08 3.725 ;
      RECT 27.046 3.58 27.07 3.731 ;
      RECT 26.96 3.602 27.046 3.756 ;
      RECT 26.92 3.627 26.96 3.783 ;
      RECT 26.91 3.636 26.92 3.793 ;
      RECT 26.86 3.646 26.91 3.802 ;
      RECT 26.84 3.66 26.86 3.812 ;
      RECT 26.81 3.67 26.84 3.817 ;
      RECT 26.8 3.675 26.81 3.82 ;
      RECT 26.726 3.677 26.8 3.827 ;
      RECT 26.64 3.681 26.726 3.839 ;
      RECT 26.63 3.684 26.64 3.845 ;
      RECT 26.37 3.635 26.63 3.895 ;
      RECT 27.9 3.705 28.09 3.915 ;
      RECT 27.89 3.71 28.1 3.91 ;
      RECT 27.88 3.71 28.1 3.875 ;
      RECT 27.8 3.595 28.06 3.855 ;
      RECT 26.71 3.125 26.9 3.425 ;
      RECT 26.7 3.125 26.9 3.42 ;
      RECT 26.69 3.125 26.91 3.415 ;
      RECT 26.68 3.125 26.91 3.41 ;
      RECT 26.68 3.125 26.94 3.385 ;
      RECT 26.64 2.165 26.9 2.425 ;
      RECT 26.45 2.09 26.536 2.423 ;
      RECT 26.45 2.09 26.58 2.419 ;
      RECT 26.43 2.094 26.59 2.418 ;
      RECT 26.58 2.085 26.59 2.418 ;
      RECT 26.45 2.09 26.6 2.417 ;
      RECT 26.43 2.1 26.64 2.416 ;
      RECT 26.42 2.095 26.6 2.408 ;
      RECT 26.41 2.11 26.64 2.315 ;
      RECT 26.41 2.16 26.84 2.315 ;
      RECT 26.41 2.15 26.82 2.315 ;
      RECT 26.41 2.14 26.79 2.315 ;
      RECT 26.41 2.13 26.73 2.315 ;
      RECT 26.41 2.115 26.71 2.315 ;
      RECT 26.536 2.086 26.59 2.418 ;
      RECT 25.61 2.745 25.75 3.035 ;
      RECT 25.87 2.768 25.88 2.955 ;
      RECT 26.57 2.665 26.75 2.895 ;
      RECT 26.57 2.665 26.76 2.885 ;
      RECT 26.78 2.67 26.79 2.875 ;
      RECT 26.76 2.665 26.78 2.88 ;
      RECT 26.52 2.669 26.57 2.895 ;
      RECT 26.51 2.674 26.52 2.895 ;
      RECT 26.476 2.679 26.51 2.896 ;
      RECT 26.39 2.694 26.476 2.898 ;
      RECT 26.376 2.706 26.39 2.901 ;
      RECT 26.29 2.716 26.376 2.903 ;
      RECT 26.266 2.726 26.29 2.905 ;
      RECT 26.18 2.737 26.266 2.905 ;
      RECT 26.15 2.747 26.18 2.905 ;
      RECT 26.12 2.752 26.15 2.908 ;
      RECT 26.1 2.757 26.12 2.913 ;
      RECT 26.08 2.762 26.1 2.915 ;
      RECT 26.03 2.77 26.08 2.915 ;
      RECT 26.01 2.774 26.03 2.915 ;
      RECT 25.99 2.773 26.01 2.92 ;
      RECT 25.93 2.771 25.99 2.935 ;
      RECT 25.88 2.769 25.93 2.95 ;
      RECT 25.79 2.766 25.87 3.035 ;
      RECT 25.76 2.76 25.79 3.035 ;
      RECT 25.75 2.75 25.76 3.035 ;
      RECT 25.56 2.745 25.61 2.96 ;
      RECT 25.55 2.75 25.56 2.95 ;
      RECT 25.79 3.225 26.05 3.485 ;
      RECT 25.79 3.225 26.08 3.375 ;
      RECT 25.79 3.225 26.12 3.36 ;
      RECT 26.05 3.145 26.24 3.355 ;
      RECT 26.05 3.15 26.25 3.345 ;
      RECT 26 3.22 26.25 3.345 ;
      RECT 26.03 3.155 26.05 3.485 ;
      RECT 26.02 3.18 26.25 3.345 ;
      RECT 25.2 3.125 25.21 3.355 ;
      RECT 25.1 2.245 25.17 3.355 ;
      RECT 25.84 2.355 26.1 2.615 ;
      RECT 25.54 2.405 25.67 2.565 ;
      RECT 25.756 2.412 25.84 2.565 ;
      RECT 25.67 2.407 25.756 2.565 ;
      RECT 25.48 2.405 25.54 2.575 ;
      RECT 25.45 2.403 25.48 2.59 ;
      RECT 25.43 2.401 25.45 2.6 ;
      RECT 25.42 2.399 25.43 2.605 ;
      RECT 25.4 2.398 25.42 2.615 ;
      RECT 25.39 2.396 25.4 2.62 ;
      RECT 25.37 2.395 25.39 2.625 ;
      RECT 25.35 2.39 25.37 2.63 ;
      RECT 25.32 2.376 25.35 2.64 ;
      RECT 25.28 2.355 25.32 2.655 ;
      RECT 25.27 2.34 25.28 2.665 ;
      RECT 25.25 2.331 25.27 2.675 ;
      RECT 25.24 2.322 25.25 2.695 ;
      RECT 25.23 2.317 25.24 2.755 ;
      RECT 25.21 2.311 25.23 2.84 ;
      RECT 25.21 3.15 25.22 3.35 ;
      RECT 25.2 2.306 25.21 3.07 ;
      RECT 25.19 2.28 25.2 3.355 ;
      RECT 25.17 2.25 25.19 3.355 ;
      RECT 25.08 2.245 25.1 2.58 ;
      RECT 25.09 2.68 25.1 3.355 ;
      RECT 25.08 2.72 25.09 3.355 ;
      RECT 25.05 2.245 25.08 2.525 ;
      RECT 25.06 2.81 25.08 3.355 ;
      RECT 25.045 2.915 25.06 3.355 ;
      RECT 25.02 2.245 25.05 2.48 ;
      RECT 25.04 2.947 25.045 3.355 ;
      RECT 25.02 3.05 25.04 3.355 ;
      RECT 25.01 2.245 25.02 2.47 ;
      RECT 25.01 3.12 25.02 3.35 ;
      RECT 24.99 2.245 25.01 2.46 ;
      RECT 24.98 2.25 24.99 2.45 ;
      RECT 25.19 3.525 25.21 3.765 ;
      RECT 24.51 3.455 24.59 3.725 ;
      RECT 24.42 3.455 24.43 3.665 ;
      RECT 25.7 3.525 25.71 3.725 ;
      RECT 25.62 3.515 25.7 3.75 ;
      RECT 25.616 3.515 25.62 3.776 ;
      RECT 25.53 3.515 25.616 3.786 ;
      RECT 25.51 3.515 25.53 3.794 ;
      RECT 25.486 3.516 25.51 3.792 ;
      RECT 25.4 3.521 25.486 3.787 ;
      RECT 25.382 3.525 25.4 3.781 ;
      RECT 25.296 3.525 25.382 3.777 ;
      RECT 25.21 3.525 25.296 3.769 ;
      RECT 25.106 3.525 25.19 3.762 ;
      RECT 25.02 3.525 25.106 3.756 ;
      RECT 24.96 3.52 25.02 3.75 ;
      RECT 24.932 3.514 24.96 3.747 ;
      RECT 24.846 3.511 24.932 3.744 ;
      RECT 24.76 3.507 24.846 3.738 ;
      RECT 24.715 3.495 24.76 3.734 ;
      RECT 24.69 3.48 24.715 3.732 ;
      RECT 24.65 3.465 24.69 3.73 ;
      RECT 24.59 3.455 24.65 3.727 ;
      RECT 24.5 3.455 24.51 3.72 ;
      RECT 24.485 3.455 24.5 3.71 ;
      RECT 24.43 3.455 24.485 3.685 ;
      RECT 24.41 3.47 24.42 3.66 ;
      RECT 24.54 2.635 24.8 2.895 ;
      RECT 24.54 2.645 24.82 2.855 ;
      RECT 24.54 2.65 24.83 2.85 ;
      RECT 22.52 2.115 22.78 2.375 ;
      RECT 22.51 2.145 22.78 2.355 ;
      RECT 24.44 2.055 24.69 2.315 ;
      RECT 24.43 2.055 24.44 2.316 ;
      RECT 24.4 2.14 24.43 2.318 ;
      RECT 24.39 2.145 24.4 2.32 ;
      RECT 24.33 2.16 24.39 2.326 ;
      RECT 24.3 2.18 24.33 2.333 ;
      RECT 24.27 2.191 24.3 2.34 ;
      RECT 24.25 2.201 24.27 2.345 ;
      RECT 24.232 2.204 24.25 2.344 ;
      RECT 24.146 2.203 24.232 2.344 ;
      RECT 24.06 2.2 24.146 2.343 ;
      RECT 23.974 2.197 24.06 2.342 ;
      RECT 23.888 2.194 23.974 2.342 ;
      RECT 23.802 2.192 23.888 2.341 ;
      RECT 23.716 2.189 23.802 2.34 ;
      RECT 23.63 2.186 23.716 2.34 ;
      RECT 23.612 2.185 23.63 2.339 ;
      RECT 23.526 2.184 23.612 2.339 ;
      RECT 23.44 2.182 23.526 2.338 ;
      RECT 23.354 2.181 23.44 2.338 ;
      RECT 23.268 2.18 23.354 2.337 ;
      RECT 23.182 2.178 23.268 2.337 ;
      RECT 23.096 2.177 23.182 2.336 ;
      RECT 23.01 2.175 23.096 2.336 ;
      RECT 22.986 2.174 23.01 2.335 ;
      RECT 22.9 2.169 22.986 2.335 ;
      RECT 22.866 2.162 22.9 2.335 ;
      RECT 22.78 2.152 22.866 2.335 ;
      RECT 22.5 2.15 22.51 2.35 ;
      RECT 23.78 3.205 24.04 3.465 ;
      RECT 23.78 3.205 24.12 3.251 ;
      RECT 23.92 3.185 24.13 3.24 ;
      RECT 23.98 3.16 24.19 3.2 ;
      RECT 23.99 3.155 24.19 3.2 ;
      RECT 24 3.13 24.19 3.2 ;
      RECT 24.06 2.96 24.11 3.29 ;
      RECT 24.01 3.09 24.2 3.15 ;
      RECT 24.05 3.016 24.06 3.329 ;
      RECT 24.01 3.09 24.23 3.125 ;
      RECT 24.01 3.09 24.25 3.1 ;
      RECT 24.12 2.89 24.31 3.095 ;
      RECT 24.11 2.9 24.32 3.09 ;
      RECT 24.03 3.063 24.32 3.09 ;
      RECT 24.04 3.039 24.05 3.345 ;
      RECT 24.13 2.885 24.3 3.095 ;
      RECT 23.42 2.675 23.61 2.885 ;
      RECT 21.99 2.605 22.25 2.865 ;
      RECT 22.34 2.595 22.44 2.805 ;
      RECT 22.29 2.615 22.33 2.805 ;
      RECT 23.61 2.685 23.62 2.88 ;
      RECT 23.41 2.685 23.42 2.88 ;
      RECT 23.39 2.7 23.41 2.87 ;
      RECT 23.38 2.71 23.39 2.865 ;
      RECT 23.34 2.71 23.38 2.863 ;
      RECT 23.316 2.704 23.34 2.86 ;
      RECT 23.23 2.699 23.316 2.857 ;
      RECT 23.17 2.695 23.23 2.852 ;
      RECT 23.136 2.692 23.17 2.849 ;
      RECT 23.05 2.682 23.136 2.845 ;
      RECT 23.046 2.675 23.05 2.842 ;
      RECT 22.96 2.67 23.046 2.84 ;
      RECT 22.932 2.663 22.96 2.836 ;
      RECT 22.846 2.658 22.932 2.833 ;
      RECT 22.76 2.649 22.846 2.828 ;
      RECT 22.75 2.644 22.76 2.825 ;
      RECT 22.736 2.643 22.75 2.825 ;
      RECT 22.65 2.639 22.736 2.82 ;
      RECT 22.63 2.633 22.65 2.816 ;
      RECT 22.57 2.628 22.63 2.815 ;
      RECT 22.54 2.62 22.57 2.815 ;
      RECT 22.53 2.605 22.54 2.815 ;
      RECT 22.526 2.595 22.53 2.814 ;
      RECT 22.44 2.595 22.526 2.81 ;
      RECT 22.33 2.605 22.34 2.805 ;
      RECT 22.26 2.615 22.29 2.8 ;
      RECT 22.25 2.615 22.26 2.8 ;
      RECT 23.17 3.115 23.43 3.375 ;
      RECT 23.1 3.125 23.43 3.335 ;
      RECT 23.09 3.13 23.43 3.33 ;
      RECT 22.51 3.115 22.77 3.375 ;
      RECT 22.51 3.16 22.88 3.365 ;
      RECT 22.51 3.155 22.87 3.365 ;
      RECT 21.42 3.322 21.6 3.765 ;
      RECT 21.41 3.322 21.6 3.763 ;
      RECT 21.41 3.337 21.61 3.76 ;
      RECT 21.4 2.26 21.53 3.758 ;
      RECT 21.4 3.385 21.67 3.645 ;
      RECT 21.4 3.36 21.62 3.645 ;
      RECT 21.4 3.295 21.59 3.758 ;
      RECT 21.4 3.255 21.56 3.758 ;
      RECT 21.4 3.21 21.55 3.758 ;
      RECT 21.4 3.15 21.54 3.758 ;
      RECT 21.39 2.545 21.53 3.2 ;
      RECT 21.43 2.245 21.54 3.065 ;
      RECT 21.4 2.26 21.58 2.52 ;
      RECT 21.4 2.26 21.59 2.47 ;
      RECT 21.43 2.245 21.6 2.463 ;
      RECT 21.42 2.247 21.61 2.458 ;
      RECT 21.41 2.252 21.62 2.45 ;
      RECT 20.27 7.77 20.56 8 ;
      RECT 20.33 6.29 20.5 8 ;
      RECT 20.325 6.655 20.675 7.005 ;
      RECT 20.27 6.29 20.56 6.52 ;
      RECT 19.865 2.395 19.97 2.965 ;
      RECT 19.865 2.73 20.19 2.96 ;
      RECT 19.865 2.76 20.36 2.93 ;
      RECT 19.865 2.395 20.055 2.96 ;
      RECT 19.28 2.36 19.57 2.59 ;
      RECT 19.28 2.395 20.055 2.565 ;
      RECT 19.34 0.88 19.51 2.59 ;
      RECT 19.28 0.88 19.57 1.11 ;
      RECT 19.28 7.77 19.57 8 ;
      RECT 19.34 6.29 19.51 8 ;
      RECT 19.28 6.29 19.57 6.52 ;
      RECT 19.28 6.325 20.135 6.485 ;
      RECT 19.965 5.92 20.135 6.485 ;
      RECT 19.28 6.32 19.675 6.485 ;
      RECT 19.9 5.92 20.19 6.15 ;
      RECT 19.9 5.95 20.36 6.12 ;
      RECT 18.91 2.73 19.2 2.96 ;
      RECT 18.91 2.76 19.37 2.93 ;
      RECT 18.975 1.655 19.14 2.96 ;
      RECT 17.49 1.625 17.78 1.855 ;
      RECT 17.49 1.655 19.14 1.825 ;
      RECT 17.55 0.885 17.72 1.855 ;
      RECT 17.49 0.885 17.78 1.115 ;
      RECT 17.49 7.765 17.78 7.995 ;
      RECT 17.55 7.025 17.72 7.995 ;
      RECT 17.55 7.12 19.14 7.29 ;
      RECT 18.97 5.92 19.14 7.29 ;
      RECT 17.49 7.025 17.78 7.255 ;
      RECT 18.91 5.92 19.2 6.15 ;
      RECT 18.91 5.95 19.37 6.12 ;
      RECT 15.525 3.43 15.875 3.78 ;
      RECT 15.615 2.025 15.785 3.78 ;
      RECT 17.92 1.965 18.27 2.315 ;
      RECT 15.615 2.025 17.235 2.2 ;
      RECT 15.615 2.025 18.27 2.195 ;
      RECT 17.945 6.655 18.27 6.98 ;
      RECT 13.34 6.605 13.69 6.955 ;
      RECT 17.92 6.655 18.27 6.885 ;
      RECT 13.16 6.655 13.69 6.885 ;
      RECT 12.99 6.685 18.27 6.855 ;
      RECT 17.145 2.365 17.465 2.685 ;
      RECT 17.115 2.365 17.465 2.595 ;
      RECT 16.945 2.395 17.465 2.565 ;
      RECT 17.145 6.225 17.465 6.545 ;
      RECT 17.115 6.285 17.465 6.515 ;
      RECT 16.945 6.315 17.465 6.485 ;
      RECT 12.985 3.255 13.175 3.925 ;
      RECT 12.925 3.665 12.965 3.925 ;
      RECT 14.295 2.89 14.305 3.111 ;
      RECT 14.225 2.885 14.295 3.236 ;
      RECT 14.215 2.885 14.225 3.36 ;
      RECT 14.185 2.885 14.215 3.41 ;
      RECT 14.165 2.885 14.185 3.485 ;
      RECT 14.145 2.885 14.165 3.555 ;
      RECT 14.115 2.885 14.145 3.595 ;
      RECT 14.105 2.885 14.115 3.615 ;
      RECT 14.095 2.885 14.105 3.626 ;
      RECT 14.085 3.135 14.095 3.628 ;
      RECT 14.075 3.2 14.085 3.63 ;
      RECT 14.065 3.295 14.075 3.632 ;
      RECT 14.055 3.37 14.065 3.634 ;
      RECT 14.005 3.394 14.055 3.64 ;
      RECT 13.965 3.429 14.005 3.649 ;
      RECT 13.955 3.445 13.965 3.654 ;
      RECT 13.941 3.45 13.955 3.657 ;
      RECT 13.855 3.49 13.941 3.668 ;
      RECT 13.775 3.533 13.855 3.686 ;
      RECT 13.755 3.543 13.775 3.697 ;
      RECT 13.725 3.551 13.755 3.702 ;
      RECT 13.705 3.561 13.725 3.707 ;
      RECT 13.681 3.567 13.705 3.712 ;
      RECT 13.595 3.577 13.681 3.725 ;
      RECT 13.517 3.583 13.595 3.745 ;
      RECT 13.431 3.578 13.517 3.764 ;
      RECT 13.345 3.574 13.431 3.785 ;
      RECT 13.265 3.57 13.345 3.8 ;
      RECT 13.195 3.566 13.265 3.831 ;
      RECT 13.185 3.277 13.195 3.345 ;
      RECT 13.185 3.555 13.195 3.861 ;
      RECT 13.175 3.262 13.185 3.49 ;
      RECT 13.175 3.535 13.185 3.925 ;
      RECT 12.965 3.285 12.985 3.925 ;
      RECT 13.765 2.605 13.775 3.345 ;
      RECT 13.585 3.125 13.605 3.345 ;
      RECT 13.595 3.115 13.605 3.345 ;
      RECT 14.095 2.155 14.135 2.415 ;
      RECT 14.085 2.155 14.095 2.425 ;
      RECT 14.051 2.155 14.085 2.452 ;
      RECT 13.965 2.155 14.051 2.512 ;
      RECT 13.945 2.155 13.965 2.575 ;
      RECT 13.885 2.155 13.945 2.74 ;
      RECT 13.875 2.155 13.885 2.9 ;
      RECT 13.845 2.346 13.875 2.995 ;
      RECT 13.835 2.401 13.845 3.095 ;
      RECT 13.825 2.43 13.835 3.14 ;
      RECT 13.815 2.455 13.825 3.173 ;
      RECT 13.805 2.49 13.815 3.228 ;
      RECT 13.785 2.535 13.805 3.29 ;
      RECT 13.775 2.58 13.785 3.34 ;
      RECT 13.755 2.64 13.765 3.345 ;
      RECT 13.745 2.67 13.755 3.345 ;
      RECT 13.725 2.7 13.745 3.345 ;
      RECT 13.675 2.805 13.725 3.345 ;
      RECT 13.665 2.9 13.675 3.345 ;
      RECT 13.655 2.93 13.665 3.345 ;
      RECT 13.63 2.98 13.655 3.345 ;
      RECT 13.625 3.035 13.63 3.345 ;
      RECT 13.605 3.06 13.625 3.345 ;
      RECT 13.565 3.14 13.585 3.335 ;
      RECT 13.315 2.725 13.385 2.935 ;
      RECT 10.555 2.635 10.815 2.895 ;
      RECT 13.385 2.73 13.395 2.93 ;
      RECT 13.271 2.723 13.315 2.935 ;
      RECT 13.185 2.716 13.271 2.935 ;
      RECT 13.165 2.711 13.185 2.925 ;
      RECT 13.155 2.709 13.165 2.905 ;
      RECT 13.105 2.706 13.155 2.9 ;
      RECT 13.075 2.702 13.105 2.895 ;
      RECT 13.055 2.7 13.075 2.89 ;
      RECT 13.015 2.697 13.055 2.885 ;
      RECT 12.945 2.691 13.015 2.88 ;
      RECT 12.915 2.686 12.945 2.875 ;
      RECT 12.895 2.684 12.915 2.87 ;
      RECT 12.865 2.681 12.895 2.865 ;
      RECT 12.805 2.677 12.865 2.86 ;
      RECT 12.735 2.675 12.805 2.85 ;
      RECT 12.701 2.673 12.735 2.843 ;
      RECT 12.615 2.668 12.701 2.835 ;
      RECT 12.581 2.662 12.615 2.827 ;
      RECT 12.495 2.652 12.581 2.819 ;
      RECT 12.461 2.643 12.495 2.811 ;
      RECT 12.375 2.638 12.461 2.803 ;
      RECT 12.305 2.635 12.375 2.793 ;
      RECT 12.285 2.63 12.305 2.787 ;
      RECT 12.281 2.625 12.285 2.786 ;
      RECT 12.195 2.621 12.281 2.781 ;
      RECT 12.155 2.616 12.195 2.774 ;
      RECT 12.075 2.615 12.155 2.769 ;
      RECT 12.055 2.615 12.075 2.766 ;
      RECT 12.029 2.615 12.055 2.766 ;
      RECT 11.943 2.617 12.029 2.77 ;
      RECT 11.857 2.619 11.943 2.777 ;
      RECT 11.771 2.621 11.857 2.783 ;
      RECT 11.685 2.624 11.771 2.79 ;
      RECT 11.651 2.626 11.685 2.795 ;
      RECT 11.565 2.631 11.651 2.8 ;
      RECT 11.541 2.626 11.565 2.804 ;
      RECT 11.455 2.631 11.541 2.809 ;
      RECT 11.417 2.636 11.455 2.814 ;
      RECT 11.331 2.639 11.417 2.819 ;
      RECT 11.245 2.643 11.331 2.826 ;
      RECT 11.181 2.645 11.245 2.832 ;
      RECT 11.095 2.645 11.181 2.838 ;
      RECT 11.011 2.646 11.095 2.845 ;
      RECT 10.925 2.649 11.011 2.852 ;
      RECT 10.901 2.651 10.925 2.856 ;
      RECT 10.815 2.653 10.901 2.861 ;
      RECT 10.545 2.67 10.555 2.865 ;
      RECT 12.73 7.765 13.02 7.995 ;
      RECT 12.79 7.025 12.96 7.995 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 12.73 7.025 13.02 7.425 ;
      RECT 12.785 2.247 12.975 2.455 ;
      RECT 12.775 2.252 12.985 2.45 ;
      RECT 12.765 2.233 12.775 2.445 ;
      RECT 12.735 2.228 12.765 2.44 ;
      RECT 12.695 2.252 12.985 2.43 ;
      RECT 12.475 2.165 12.735 2.425 ;
      RECT 12.775 2.236 12.785 2.45 ;
      RECT 12.475 2.245 12.965 2.425 ;
      RECT 12.475 2.241 12.825 2.425 ;
      RECT 12.425 3.155 12.475 3.435 ;
      RECT 12.355 3.125 12.385 3.435 ;
      RECT 12.495 3.155 12.555 3.415 ;
      RECT 12.355 3.115 12.375 3.435 ;
      RECT 12.475 3.155 12.495 3.425 ;
      RECT 12.395 3.145 12.425 3.435 ;
      RECT 12.385 3.13 12.395 3.435 ;
      RECT 12.335 3.105 12.355 3.435 ;
      RECT 12.305 3.09 12.335 3.435 ;
      RECT 12.295 3.08 12.305 3.435 ;
      RECT 12.275 3.069 12.295 3.43 ;
      RECT 12.255 3.057 12.275 3.4 ;
      RECT 12.245 3.048 12.255 3.383 ;
      RECT 12.215 3.03 12.245 3.375 ;
      RECT 12.205 2.995 12.215 3.367 ;
      RECT 12.195 2.975 12.205 3.36 ;
      RECT 12.185 2.955 12.195 3.353 ;
      RECT 12.175 2.94 12.185 3.348 ;
      RECT 12.165 2.92 12.175 3.343 ;
      RECT 12.155 2.915 12.165 3.338 ;
      RECT 12.151 2.905 12.155 3.334 ;
      RECT 12.065 2.905 12.151 3.309 ;
      RECT 12.035 2.905 12.065 3.275 ;
      RECT 12.025 2.905 12.035 3.255 ;
      RECT 11.965 2.905 12.025 3.2 ;
      RECT 11.955 2.92 11.965 3.145 ;
      RECT 11.945 2.93 11.955 3.125 ;
      RECT 11.895 3.665 12.155 3.925 ;
      RECT 11.815 3.685 12.155 3.901 ;
      RECT 11.795 3.685 12.155 3.896 ;
      RECT 11.771 3.685 12.155 3.894 ;
      RECT 11.685 3.685 12.155 3.889 ;
      RECT 11.535 3.625 11.795 3.885 ;
      RECT 11.495 3.68 11.815 3.88 ;
      RECT 11.485 3.69 12.155 3.875 ;
      RECT 11.505 3.675 11.795 3.885 ;
      RECT 11.395 2.115 11.655 2.375 ;
      RECT 11.395 2.2 11.665 2.3 ;
      RECT 10.565 3.63 10.585 3.874 ;
      RECT 10.565 3.63 10.635 3.869 ;
      RECT 10.545 3.635 10.635 3.868 ;
      RECT 10.535 3.65 10.721 3.858 ;
      RECT 10.535 3.65 10.795 3.855 ;
      RECT 10.53 3.687 10.805 3.845 ;
      RECT 10.53 3.687 10.891 3.841 ;
      RECT 10.53 3.687 10.905 3.827 ;
      RECT 10.805 3.565 11.065 3.825 ;
      RECT 10.525 3.692 11.065 3.82 ;
      RECT 10.515 3.74 11.065 3.795 ;
      RECT 10.785 3.605 10.805 3.854 ;
      RECT 10.721 3.609 10.785 3.857 ;
      RECT 10.585 3.622 11.065 3.825 ;
      RECT 10.635 3.616 10.721 3.862 ;
      RECT 10.035 2.475 10.045 2.645 ;
      RECT 10.095 2.435 10.105 2.615 ;
      RECT 10.395 2.245 10.405 2.455 ;
      RECT 10.725 2.095 10.975 2.355 ;
      RECT 10.715 2.095 10.725 2.357 ;
      RECT 10.705 2.155 10.715 2.361 ;
      RECT 10.675 2.157 10.705 2.369 ;
      RECT 10.645 2.162 10.675 2.383 ;
      RECT 10.635 2.166 10.645 2.393 ;
      RECT 10.605 2.171 10.635 2.405 ;
      RECT 10.575 2.18 10.605 2.406 ;
      RECT 10.505 2.19 10.575 2.41 ;
      RECT 10.465 2.195 10.505 2.414 ;
      RECT 10.445 2.195 10.465 2.425 ;
      RECT 10.435 2.2 10.445 2.435 ;
      RECT 10.425 2.21 10.435 2.438 ;
      RECT 10.415 2.23 10.425 2.443 ;
      RECT 10.405 2.24 10.415 2.445 ;
      RECT 10.375 2.255 10.395 2.462 ;
      RECT 10.365 2.267 10.375 2.472 ;
      RECT 10.355 2.273 10.365 2.475 ;
      RECT 10.321 2.286 10.355 2.485 ;
      RECT 10.235 2.32 10.321 2.518 ;
      RECT 10.215 2.355 10.235 2.547 ;
      RECT 10.195 2.37 10.215 2.559 ;
      RECT 10.175 2.38 10.195 2.571 ;
      RECT 10.125 2.399 10.175 2.591 ;
      RECT 10.115 2.416 10.125 2.605 ;
      RECT 10.105 2.422 10.115 2.61 ;
      RECT 10.085 2.44 10.095 2.618 ;
      RECT 10.075 2.445 10.085 2.625 ;
      RECT 10.065 2.456 10.075 2.632 ;
      RECT 10.045 2.461 10.065 2.64 ;
      RECT 10.025 2.475 10.035 2.65 ;
      RECT 10.015 2.48 10.025 2.66 ;
      RECT 9.985 2.494 10.015 2.67 ;
      RECT 9.975 2.507 9.985 2.68 ;
      RECT 9.895 2.538 9.975 2.705 ;
      RECT 9.875 2.568 9.895 2.73 ;
      RECT 9.865 2.573 9.875 2.737 ;
      RECT 9.835 2.585 9.865 2.743 ;
      RECT 9.825 2.6 9.835 2.749 ;
      RECT 9.815 2.605 9.825 2.752 ;
      RECT 9.795 2.615 9.815 2.756 ;
      RECT 9.775 2.62 9.795 2.762 ;
      RECT 9.745 2.625 9.775 2.77 ;
      RECT 9.715 2.63 9.745 2.78 ;
      RECT 9.685 2.64 9.715 2.789 ;
      RECT 9.645 2.645 9.685 2.797 ;
      RECT 9.595 2.638 9.645 2.809 ;
      RECT 9.575 2.629 9.595 2.82 ;
      RECT 9.565 2.626 9.575 2.825 ;
      RECT 9.525 2.625 9.565 2.826 ;
      RECT 9.515 2.61 9.525 2.827 ;
      RECT 9.487 2.595 9.515 2.828 ;
      RECT 9.401 2.595 9.487 2.83 ;
      RECT 9.315 2.595 9.401 2.834 ;
      RECT 9.295 2.595 9.315 2.83 ;
      RECT 9.285 2.605 9.295 2.823 ;
      RECT 9.275 2.62 9.285 2.818 ;
      RECT 9.265 2.625 9.275 2.795 ;
      RECT 10.745 3.13 10.755 3.33 ;
      RECT 10.695 3.125 10.745 3.35 ;
      RECT 10.685 3.125 10.695 3.37 ;
      RECT 10.641 3.125 10.685 3.374 ;
      RECT 10.555 3.125 10.641 3.371 ;
      RECT 10.495 3.135 10.555 3.368 ;
      RECT 10.435 3.149 10.495 3.366 ;
      RECT 10.425 3.154 10.435 3.364 ;
      RECT 10.415 3.16 10.425 3.363 ;
      RECT 10.345 3.173 10.415 3.359 ;
      RECT 10.297 3.187 10.345 3.36 ;
      RECT 10.211 3.203 10.297 3.372 ;
      RECT 10.125 3.224 10.211 3.388 ;
      RECT 10.105 3.235 10.125 3.398 ;
      RECT 10.025 3.245 10.105 3.408 ;
      RECT 9.991 3.259 10.025 3.42 ;
      RECT 9.905 3.274 9.991 3.435 ;
      RECT 9.875 3.29 9.905 3.445 ;
      RECT 9.82 3.305 9.875 3.456 ;
      RECT 9.775 3.323 9.82 3.476 ;
      RECT 9.721 3.342 9.775 3.496 ;
      RECT 9.635 3.368 9.721 3.523 ;
      RECT 9.615 3.39 9.635 3.543 ;
      RECT 9.555 3.405 9.615 3.559 ;
      RECT 9.545 3.42 9.555 3.573 ;
      RECT 9.525 3.425 9.545 3.579 ;
      RECT 9.495 3.438 9.525 3.589 ;
      RECT 9.475 3.443 9.495 3.598 ;
      RECT 9.465 3.45 9.475 3.603 ;
      RECT 9.455 3.455 9.465 3.606 ;
      RECT 9.415 3.465 9.455 3.615 ;
      RECT 9.39 3.48 9.415 3.627 ;
      RECT 9.345 3.495 9.39 3.639 ;
      RECT 9.325 3.507 9.345 3.651 ;
      RECT 9.295 3.512 9.325 3.661 ;
      RECT 9.275 3.519 9.295 3.671 ;
      RECT 9.265 3.525 9.275 3.68 ;
      RECT 9.241 3.532 9.265 3.69 ;
      RECT 9.155 3.554 9.241 3.71 ;
      RECT 9.145 3.573 9.155 3.725 ;
      RECT 9.121 3.58 9.145 3.731 ;
      RECT 9.035 3.602 9.121 3.756 ;
      RECT 8.995 3.627 9.035 3.783 ;
      RECT 8.985 3.636 8.995 3.793 ;
      RECT 8.935 3.646 8.985 3.802 ;
      RECT 8.915 3.66 8.935 3.812 ;
      RECT 8.885 3.67 8.915 3.817 ;
      RECT 8.875 3.675 8.885 3.82 ;
      RECT 8.801 3.677 8.875 3.827 ;
      RECT 8.715 3.681 8.801 3.839 ;
      RECT 8.705 3.684 8.715 3.845 ;
      RECT 8.445 3.635 8.705 3.895 ;
      RECT 9.975 3.705 10.165 3.915 ;
      RECT 9.965 3.71 10.175 3.91 ;
      RECT 9.955 3.71 10.175 3.875 ;
      RECT 9.875 3.595 10.135 3.855 ;
      RECT 8.785 3.125 8.975 3.425 ;
      RECT 8.775 3.125 8.975 3.42 ;
      RECT 8.765 3.125 8.985 3.415 ;
      RECT 8.755 3.125 8.985 3.41 ;
      RECT 8.755 3.125 9.015 3.385 ;
      RECT 8.715 2.165 8.975 2.425 ;
      RECT 8.525 2.09 8.611 2.423 ;
      RECT 8.525 2.09 8.655 2.419 ;
      RECT 8.505 2.094 8.665 2.418 ;
      RECT 8.655 2.085 8.665 2.418 ;
      RECT 8.525 2.09 8.675 2.417 ;
      RECT 8.505 2.1 8.715 2.416 ;
      RECT 8.495 2.095 8.675 2.408 ;
      RECT 8.485 2.11 8.715 2.315 ;
      RECT 8.485 2.16 8.915 2.315 ;
      RECT 8.485 2.15 8.895 2.315 ;
      RECT 8.485 2.14 8.865 2.315 ;
      RECT 8.485 2.13 8.805 2.315 ;
      RECT 8.485 2.115 8.785 2.315 ;
      RECT 8.611 2.086 8.665 2.418 ;
      RECT 7.685 2.745 7.825 3.035 ;
      RECT 7.945 2.768 7.955 2.955 ;
      RECT 8.645 2.665 8.825 2.895 ;
      RECT 8.645 2.665 8.835 2.885 ;
      RECT 8.855 2.67 8.865 2.875 ;
      RECT 8.835 2.665 8.855 2.88 ;
      RECT 8.595 2.669 8.645 2.895 ;
      RECT 8.585 2.674 8.595 2.895 ;
      RECT 8.551 2.679 8.585 2.896 ;
      RECT 8.465 2.694 8.551 2.898 ;
      RECT 8.451 2.706 8.465 2.901 ;
      RECT 8.365 2.716 8.451 2.903 ;
      RECT 8.341 2.726 8.365 2.905 ;
      RECT 8.255 2.737 8.341 2.905 ;
      RECT 8.225 2.747 8.255 2.905 ;
      RECT 8.195 2.752 8.225 2.908 ;
      RECT 8.175 2.757 8.195 2.913 ;
      RECT 8.155 2.762 8.175 2.915 ;
      RECT 8.105 2.77 8.155 2.915 ;
      RECT 8.085 2.774 8.105 2.915 ;
      RECT 8.065 2.773 8.085 2.92 ;
      RECT 8.005 2.771 8.065 2.935 ;
      RECT 7.955 2.769 8.005 2.95 ;
      RECT 7.865 2.766 7.945 3.035 ;
      RECT 7.835 2.76 7.865 3.035 ;
      RECT 7.825 2.75 7.835 3.035 ;
      RECT 7.635 2.745 7.685 2.96 ;
      RECT 7.625 2.75 7.635 2.95 ;
      RECT 7.865 3.225 8.125 3.485 ;
      RECT 7.865 3.225 8.155 3.375 ;
      RECT 7.865 3.225 8.195 3.36 ;
      RECT 8.125 3.145 8.315 3.355 ;
      RECT 8.125 3.15 8.325 3.345 ;
      RECT 8.075 3.22 8.325 3.345 ;
      RECT 8.105 3.155 8.125 3.485 ;
      RECT 8.095 3.18 8.325 3.345 ;
      RECT 7.275 3.125 7.285 3.355 ;
      RECT 7.175 2.245 7.245 3.355 ;
      RECT 7.915 2.355 8.175 2.615 ;
      RECT 7.615 2.405 7.745 2.565 ;
      RECT 7.831 2.412 7.915 2.565 ;
      RECT 7.745 2.407 7.831 2.565 ;
      RECT 7.555 2.405 7.615 2.575 ;
      RECT 7.525 2.403 7.555 2.59 ;
      RECT 7.505 2.401 7.525 2.6 ;
      RECT 7.495 2.399 7.505 2.605 ;
      RECT 7.475 2.398 7.495 2.615 ;
      RECT 7.465 2.396 7.475 2.62 ;
      RECT 7.445 2.395 7.465 2.625 ;
      RECT 7.425 2.39 7.445 2.63 ;
      RECT 7.395 2.376 7.425 2.64 ;
      RECT 7.355 2.355 7.395 2.655 ;
      RECT 7.345 2.34 7.355 2.665 ;
      RECT 7.325 2.331 7.345 2.675 ;
      RECT 7.315 2.322 7.325 2.695 ;
      RECT 7.305 2.317 7.315 2.755 ;
      RECT 7.285 2.311 7.305 2.84 ;
      RECT 7.285 3.15 7.295 3.35 ;
      RECT 7.275 2.306 7.285 3.07 ;
      RECT 7.265 2.28 7.275 3.355 ;
      RECT 7.245 2.25 7.265 3.355 ;
      RECT 7.155 2.245 7.175 2.58 ;
      RECT 7.165 2.68 7.175 3.355 ;
      RECT 7.155 2.72 7.165 3.355 ;
      RECT 7.125 2.245 7.155 2.525 ;
      RECT 7.135 2.81 7.155 3.355 ;
      RECT 7.12 2.915 7.135 3.355 ;
      RECT 7.095 2.245 7.125 2.48 ;
      RECT 7.115 2.947 7.12 3.355 ;
      RECT 7.095 3.05 7.115 3.355 ;
      RECT 7.085 2.245 7.095 2.47 ;
      RECT 7.085 3.12 7.095 3.35 ;
      RECT 7.065 2.245 7.085 2.46 ;
      RECT 7.055 2.25 7.065 2.45 ;
      RECT 7.265 3.525 7.285 3.765 ;
      RECT 6.585 3.455 6.665 3.725 ;
      RECT 6.495 3.455 6.505 3.665 ;
      RECT 7.775 3.525 7.785 3.725 ;
      RECT 7.695 3.515 7.775 3.75 ;
      RECT 7.691 3.515 7.695 3.776 ;
      RECT 7.605 3.515 7.691 3.786 ;
      RECT 7.585 3.515 7.605 3.794 ;
      RECT 7.561 3.516 7.585 3.792 ;
      RECT 7.475 3.521 7.561 3.787 ;
      RECT 7.457 3.525 7.475 3.781 ;
      RECT 7.371 3.525 7.457 3.777 ;
      RECT 7.285 3.525 7.371 3.769 ;
      RECT 7.181 3.525 7.265 3.762 ;
      RECT 7.095 3.525 7.181 3.756 ;
      RECT 7.035 3.52 7.095 3.75 ;
      RECT 7.007 3.514 7.035 3.747 ;
      RECT 6.921 3.511 7.007 3.744 ;
      RECT 6.835 3.507 6.921 3.738 ;
      RECT 6.79 3.495 6.835 3.734 ;
      RECT 6.765 3.48 6.79 3.732 ;
      RECT 6.725 3.465 6.765 3.73 ;
      RECT 6.665 3.455 6.725 3.727 ;
      RECT 6.575 3.455 6.585 3.72 ;
      RECT 6.56 3.455 6.575 3.71 ;
      RECT 6.505 3.455 6.56 3.685 ;
      RECT 6.485 3.47 6.495 3.66 ;
      RECT 6.615 2.635 6.875 2.895 ;
      RECT 6.615 2.645 6.895 2.855 ;
      RECT 6.615 2.65 6.905 2.85 ;
      RECT 4.595 2.115 4.855 2.375 ;
      RECT 4.585 2.145 4.855 2.355 ;
      RECT 6.515 2.055 6.765 2.315 ;
      RECT 6.505 2.055 6.515 2.316 ;
      RECT 6.475 2.14 6.505 2.318 ;
      RECT 6.465 2.145 6.475 2.32 ;
      RECT 6.405 2.16 6.465 2.326 ;
      RECT 6.375 2.18 6.405 2.333 ;
      RECT 6.345 2.191 6.375 2.34 ;
      RECT 6.325 2.201 6.345 2.345 ;
      RECT 6.307 2.204 6.325 2.344 ;
      RECT 6.221 2.203 6.307 2.344 ;
      RECT 6.135 2.2 6.221 2.343 ;
      RECT 6.049 2.197 6.135 2.342 ;
      RECT 5.963 2.194 6.049 2.342 ;
      RECT 5.877 2.192 5.963 2.341 ;
      RECT 5.791 2.189 5.877 2.34 ;
      RECT 5.705 2.186 5.791 2.34 ;
      RECT 5.687 2.185 5.705 2.339 ;
      RECT 5.601 2.184 5.687 2.339 ;
      RECT 5.515 2.182 5.601 2.338 ;
      RECT 5.429 2.181 5.515 2.338 ;
      RECT 5.343 2.18 5.429 2.337 ;
      RECT 5.257 2.178 5.343 2.337 ;
      RECT 5.171 2.177 5.257 2.336 ;
      RECT 5.085 2.175 5.171 2.336 ;
      RECT 5.061 2.174 5.085 2.335 ;
      RECT 4.975 2.169 5.061 2.335 ;
      RECT 4.941 2.162 4.975 2.335 ;
      RECT 4.855 2.152 4.941 2.335 ;
      RECT 4.575 2.15 4.585 2.35 ;
      RECT 5.855 3.205 6.115 3.465 ;
      RECT 5.855 3.205 6.195 3.251 ;
      RECT 5.995 3.185 6.205 3.24 ;
      RECT 6.055 3.16 6.265 3.2 ;
      RECT 6.065 3.155 6.265 3.2 ;
      RECT 6.075 3.13 6.265 3.2 ;
      RECT 6.135 2.96 6.185 3.29 ;
      RECT 6.085 3.09 6.275 3.15 ;
      RECT 6.125 3.016 6.135 3.329 ;
      RECT 6.085 3.09 6.305 3.125 ;
      RECT 6.085 3.09 6.325 3.1 ;
      RECT 6.195 2.89 6.385 3.095 ;
      RECT 6.185 2.9 6.395 3.09 ;
      RECT 6.105 3.063 6.395 3.09 ;
      RECT 6.115 3.039 6.125 3.345 ;
      RECT 6.205 2.885 6.375 3.095 ;
      RECT 5.495 2.675 5.685 2.885 ;
      RECT 4.065 2.605 4.325 2.865 ;
      RECT 4.415 2.595 4.515 2.805 ;
      RECT 4.365 2.615 4.405 2.805 ;
      RECT 5.685 2.685 5.695 2.88 ;
      RECT 5.485 2.685 5.495 2.88 ;
      RECT 5.465 2.7 5.485 2.87 ;
      RECT 5.455 2.71 5.465 2.865 ;
      RECT 5.415 2.71 5.455 2.863 ;
      RECT 5.391 2.704 5.415 2.86 ;
      RECT 5.305 2.699 5.391 2.857 ;
      RECT 5.245 2.695 5.305 2.852 ;
      RECT 5.211 2.692 5.245 2.849 ;
      RECT 5.125 2.682 5.211 2.845 ;
      RECT 5.121 2.675 5.125 2.842 ;
      RECT 5.035 2.67 5.121 2.84 ;
      RECT 5.007 2.663 5.035 2.836 ;
      RECT 4.921 2.658 5.007 2.833 ;
      RECT 4.835 2.649 4.921 2.828 ;
      RECT 4.825 2.644 4.835 2.825 ;
      RECT 4.811 2.643 4.825 2.825 ;
      RECT 4.725 2.639 4.811 2.82 ;
      RECT 4.705 2.633 4.725 2.816 ;
      RECT 4.645 2.628 4.705 2.815 ;
      RECT 4.615 2.62 4.645 2.815 ;
      RECT 4.605 2.605 4.615 2.815 ;
      RECT 4.601 2.595 4.605 2.814 ;
      RECT 4.515 2.595 4.601 2.81 ;
      RECT 4.405 2.605 4.415 2.805 ;
      RECT 4.335 2.615 4.365 2.8 ;
      RECT 4.325 2.615 4.335 2.8 ;
      RECT 5.245 3.115 5.505 3.375 ;
      RECT 5.175 3.125 5.505 3.335 ;
      RECT 5.165 3.13 5.505 3.33 ;
      RECT 4.585 3.115 4.845 3.375 ;
      RECT 4.585 3.16 4.955 3.365 ;
      RECT 4.585 3.155 4.945 3.365 ;
      RECT 3.495 3.322 3.675 3.765 ;
      RECT 3.485 3.322 3.675 3.763 ;
      RECT 3.485 3.337 3.685 3.76 ;
      RECT 3.475 2.26 3.605 3.758 ;
      RECT 3.475 3.385 3.745 3.645 ;
      RECT 3.475 3.36 3.695 3.645 ;
      RECT 3.475 3.295 3.665 3.758 ;
      RECT 3.475 3.255 3.635 3.758 ;
      RECT 3.475 3.21 3.625 3.758 ;
      RECT 3.475 3.15 3.615 3.758 ;
      RECT 3.465 2.545 3.605 3.2 ;
      RECT 3.505 2.245 3.615 3.065 ;
      RECT 3.475 2.26 3.655 2.52 ;
      RECT 3.475 2.26 3.665 2.47 ;
      RECT 3.505 2.245 3.675 2.463 ;
      RECT 3.495 2.247 3.685 2.458 ;
      RECT 3.485 2.252 3.695 2.45 ;
      RECT 1.7 7.765 1.99 7.995 ;
      RECT 1.76 7.025 1.93 7.995 ;
      RECT 1.67 7.025 2.02 7.315 ;
      RECT 1.295 6.285 1.645 6.575 ;
      RECT 1.155 6.315 1.645 6.485 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 81.175 2.225 81.435 2.485 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 63.25 2.225 63.51 2.485 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 45.325 2.225 45.585 2.485 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 27.4 2.225 27.66 2.485 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 9.475 2.225 9.735 2.485 ;
    LAYER mcon ;
      RECT 92.03 6.32 92.2 6.49 ;
      RECT 92.035 6.315 92.205 6.485 ;
      RECT 74.105 6.32 74.275 6.49 ;
      RECT 74.11 6.315 74.28 6.485 ;
      RECT 56.18 6.32 56.35 6.49 ;
      RECT 56.185 6.315 56.355 6.485 ;
      RECT 38.255 6.32 38.425 6.49 ;
      RECT 38.26 6.315 38.43 6.485 ;
      RECT 20.33 6.32 20.5 6.49 ;
      RECT 20.335 6.315 20.505 6.485 ;
      RECT 92.03 7.8 92.2 7.97 ;
      RECT 91.68 0.1 91.85 0.27 ;
      RECT 91.68 8.61 91.85 8.78 ;
      RECT 91.66 2.76 91.83 2.93 ;
      RECT 91.66 5.95 91.83 6.12 ;
      RECT 91.04 0.91 91.21 1.08 ;
      RECT 91.04 2.39 91.21 2.56 ;
      RECT 91.04 6.32 91.21 6.49 ;
      RECT 91.04 7.8 91.21 7.97 ;
      RECT 90.69 0.1 90.86 0.27 ;
      RECT 90.69 8.61 90.86 8.78 ;
      RECT 90.67 2.76 90.84 2.93 ;
      RECT 90.67 5.95 90.84 6.12 ;
      RECT 89.99 0.105 90.16 0.275 ;
      RECT 89.99 8.605 90.16 8.775 ;
      RECT 89.68 2.025 89.85 2.195 ;
      RECT 89.68 6.685 89.85 6.855 ;
      RECT 89.31 0.105 89.48 0.275 ;
      RECT 89.31 8.605 89.48 8.775 ;
      RECT 89.25 0.915 89.42 1.085 ;
      RECT 89.25 1.655 89.42 1.825 ;
      RECT 89.25 7.055 89.42 7.225 ;
      RECT 89.25 7.795 89.42 7.965 ;
      RECT 88.875 2.395 89.045 2.565 ;
      RECT 88.875 6.315 89.045 6.485 ;
      RECT 88.63 0.105 88.8 0.275 ;
      RECT 88.63 8.605 88.8 8.775 ;
      RECT 87.95 0.105 88.12 0.275 ;
      RECT 87.95 8.605 88.12 8.775 ;
      RECT 86.665 1.565 86.835 1.735 ;
      RECT 86.205 1.565 86.375 1.735 ;
      RECT 85.815 2.905 85.985 3.075 ;
      RECT 85.745 1.565 85.915 1.735 ;
      RECT 85.605 2.245 85.775 2.415 ;
      RECT 85.285 1.565 85.455 1.735 ;
      RECT 85.285 3.155 85.455 3.325 ;
      RECT 85.23 8.605 85.4 8.775 ;
      RECT 84.92 6.685 85.09 6.855 ;
      RECT 84.905 2.745 85.075 2.915 ;
      RECT 84.825 1.565 84.995 1.735 ;
      RECT 84.685 3.315 84.855 3.485 ;
      RECT 84.665 3.715 84.835 3.885 ;
      RECT 84.55 8.605 84.72 8.775 ;
      RECT 84.495 2.265 84.665 2.435 ;
      RECT 84.49 7.055 84.66 7.225 ;
      RECT 84.49 7.795 84.66 7.965 ;
      RECT 84.365 1.565 84.535 1.735 ;
      RECT 84.115 6.315 84.285 6.485 ;
      RECT 83.995 3.245 84.165 3.415 ;
      RECT 83.905 1.565 84.075 1.735 ;
      RECT 83.87 8.605 84.04 8.775 ;
      RECT 83.675 2.935 83.845 3.105 ;
      RECT 83.605 3.715 83.775 3.885 ;
      RECT 83.445 1.565 83.615 1.735 ;
      RECT 83.205 3.695 83.375 3.865 ;
      RECT 83.19 8.605 83.36 8.775 ;
      RECT 83.165 2.185 83.335 2.355 ;
      RECT 82.985 1.565 83.155 1.735 ;
      RECT 82.525 1.565 82.695 1.735 ;
      RECT 82.265 2.685 82.435 2.855 ;
      RECT 82.265 3.145 82.435 3.315 ;
      RECT 82.265 3.655 82.435 3.825 ;
      RECT 82.155 2.215 82.325 2.385 ;
      RECT 82.065 1.565 82.235 1.735 ;
      RECT 81.685 3.725 81.855 3.895 ;
      RECT 81.605 1.565 81.775 1.735 ;
      RECT 81.205 2.255 81.375 2.425 ;
      RECT 81.145 1.565 81.315 1.735 ;
      RECT 80.995 2.635 81.165 2.805 ;
      RECT 80.685 1.565 80.855 1.735 ;
      RECT 80.495 3.235 80.665 3.405 ;
      RECT 80.375 2.685 80.545 2.855 ;
      RECT 80.225 1.565 80.395 1.735 ;
      RECT 80.205 2.135 80.375 2.305 ;
      RECT 79.835 3.165 80.005 3.335 ;
      RECT 79.765 1.565 79.935 1.735 ;
      RECT 79.345 2.765 79.515 2.935 ;
      RECT 79.305 1.565 79.475 1.735 ;
      RECT 79.295 3.535 79.465 3.705 ;
      RECT 78.845 1.565 79.015 1.735 ;
      RECT 78.805 3.165 78.975 3.335 ;
      RECT 78.775 2.265 78.945 2.435 ;
      RECT 78.415 2.665 78.585 2.835 ;
      RECT 78.385 1.565 78.555 1.735 ;
      RECT 78.205 3.475 78.375 3.645 ;
      RECT 77.925 1.565 78.095 1.735 ;
      RECT 77.905 2.905 78.075 3.075 ;
      RECT 77.465 1.565 77.635 1.735 ;
      RECT 77.205 2.695 77.375 2.865 ;
      RECT 77.005 1.565 77.175 1.735 ;
      RECT 76.885 3.145 77.055 3.315 ;
      RECT 76.545 1.565 76.715 1.735 ;
      RECT 76.465 3.175 76.635 3.345 ;
      RECT 76.295 2.165 76.465 2.335 ;
      RECT 76.125 2.615 76.295 2.785 ;
      RECT 76.085 1.565 76.255 1.735 ;
      RECT 75.625 1.565 75.795 1.735 ;
      RECT 75.205 2.265 75.375 2.435 ;
      RECT 75.195 3.585 75.365 3.755 ;
      RECT 75.165 1.565 75.335 1.735 ;
      RECT 74.105 7.8 74.275 7.97 ;
      RECT 73.755 0.1 73.925 0.27 ;
      RECT 73.755 8.61 73.925 8.78 ;
      RECT 73.735 2.76 73.905 2.93 ;
      RECT 73.735 5.95 73.905 6.12 ;
      RECT 73.115 0.91 73.285 1.08 ;
      RECT 73.115 2.39 73.285 2.56 ;
      RECT 73.115 6.32 73.285 6.49 ;
      RECT 73.115 7.8 73.285 7.97 ;
      RECT 72.765 0.1 72.935 0.27 ;
      RECT 72.765 8.61 72.935 8.78 ;
      RECT 72.745 2.76 72.915 2.93 ;
      RECT 72.745 5.95 72.915 6.12 ;
      RECT 72.065 0.105 72.235 0.275 ;
      RECT 72.065 8.605 72.235 8.775 ;
      RECT 71.755 2.025 71.925 2.195 ;
      RECT 71.755 6.685 71.925 6.855 ;
      RECT 71.385 0.105 71.555 0.275 ;
      RECT 71.385 8.605 71.555 8.775 ;
      RECT 71.325 0.915 71.495 1.085 ;
      RECT 71.325 1.655 71.495 1.825 ;
      RECT 71.325 7.055 71.495 7.225 ;
      RECT 71.325 7.795 71.495 7.965 ;
      RECT 70.95 2.395 71.12 2.565 ;
      RECT 70.95 6.315 71.12 6.485 ;
      RECT 70.705 0.105 70.875 0.275 ;
      RECT 70.705 8.605 70.875 8.775 ;
      RECT 70.025 0.105 70.195 0.275 ;
      RECT 70.025 8.605 70.195 8.775 ;
      RECT 68.74 1.565 68.91 1.735 ;
      RECT 68.28 1.565 68.45 1.735 ;
      RECT 67.89 2.905 68.06 3.075 ;
      RECT 67.82 1.565 67.99 1.735 ;
      RECT 67.68 2.245 67.85 2.415 ;
      RECT 67.36 1.565 67.53 1.735 ;
      RECT 67.36 3.155 67.53 3.325 ;
      RECT 67.305 8.605 67.475 8.775 ;
      RECT 66.995 6.685 67.165 6.855 ;
      RECT 66.98 2.745 67.15 2.915 ;
      RECT 66.9 1.565 67.07 1.735 ;
      RECT 66.76 3.315 66.93 3.485 ;
      RECT 66.74 3.715 66.91 3.885 ;
      RECT 66.625 8.605 66.795 8.775 ;
      RECT 66.57 2.265 66.74 2.435 ;
      RECT 66.565 7.055 66.735 7.225 ;
      RECT 66.565 7.795 66.735 7.965 ;
      RECT 66.44 1.565 66.61 1.735 ;
      RECT 66.19 6.315 66.36 6.485 ;
      RECT 66.07 3.245 66.24 3.415 ;
      RECT 65.98 1.565 66.15 1.735 ;
      RECT 65.945 8.605 66.115 8.775 ;
      RECT 65.75 2.935 65.92 3.105 ;
      RECT 65.68 3.715 65.85 3.885 ;
      RECT 65.52 1.565 65.69 1.735 ;
      RECT 65.28 3.695 65.45 3.865 ;
      RECT 65.265 8.605 65.435 8.775 ;
      RECT 65.24 2.185 65.41 2.355 ;
      RECT 65.06 1.565 65.23 1.735 ;
      RECT 64.6 1.565 64.77 1.735 ;
      RECT 64.34 2.685 64.51 2.855 ;
      RECT 64.34 3.145 64.51 3.315 ;
      RECT 64.34 3.655 64.51 3.825 ;
      RECT 64.23 2.215 64.4 2.385 ;
      RECT 64.14 1.565 64.31 1.735 ;
      RECT 63.76 3.725 63.93 3.895 ;
      RECT 63.68 1.565 63.85 1.735 ;
      RECT 63.28 2.255 63.45 2.425 ;
      RECT 63.22 1.565 63.39 1.735 ;
      RECT 63.07 2.635 63.24 2.805 ;
      RECT 62.76 1.565 62.93 1.735 ;
      RECT 62.57 3.235 62.74 3.405 ;
      RECT 62.45 2.685 62.62 2.855 ;
      RECT 62.3 1.565 62.47 1.735 ;
      RECT 62.28 2.135 62.45 2.305 ;
      RECT 61.91 3.165 62.08 3.335 ;
      RECT 61.84 1.565 62.01 1.735 ;
      RECT 61.42 2.765 61.59 2.935 ;
      RECT 61.38 1.565 61.55 1.735 ;
      RECT 61.37 3.535 61.54 3.705 ;
      RECT 60.92 1.565 61.09 1.735 ;
      RECT 60.88 3.165 61.05 3.335 ;
      RECT 60.85 2.265 61.02 2.435 ;
      RECT 60.49 2.665 60.66 2.835 ;
      RECT 60.46 1.565 60.63 1.735 ;
      RECT 60.28 3.475 60.45 3.645 ;
      RECT 60 1.565 60.17 1.735 ;
      RECT 59.98 2.905 60.15 3.075 ;
      RECT 59.54 1.565 59.71 1.735 ;
      RECT 59.28 2.695 59.45 2.865 ;
      RECT 59.08 1.565 59.25 1.735 ;
      RECT 58.96 3.145 59.13 3.315 ;
      RECT 58.62 1.565 58.79 1.735 ;
      RECT 58.54 3.175 58.71 3.345 ;
      RECT 58.37 2.165 58.54 2.335 ;
      RECT 58.2 2.615 58.37 2.785 ;
      RECT 58.16 1.565 58.33 1.735 ;
      RECT 57.7 1.565 57.87 1.735 ;
      RECT 57.28 2.265 57.45 2.435 ;
      RECT 57.27 3.585 57.44 3.755 ;
      RECT 57.24 1.565 57.41 1.735 ;
      RECT 56.18 7.8 56.35 7.97 ;
      RECT 55.83 0.1 56 0.27 ;
      RECT 55.83 8.61 56 8.78 ;
      RECT 55.81 2.76 55.98 2.93 ;
      RECT 55.81 5.95 55.98 6.12 ;
      RECT 55.19 0.91 55.36 1.08 ;
      RECT 55.19 2.39 55.36 2.56 ;
      RECT 55.19 6.32 55.36 6.49 ;
      RECT 55.19 7.8 55.36 7.97 ;
      RECT 54.84 0.1 55.01 0.27 ;
      RECT 54.84 8.61 55.01 8.78 ;
      RECT 54.82 2.76 54.99 2.93 ;
      RECT 54.82 5.95 54.99 6.12 ;
      RECT 54.14 0.105 54.31 0.275 ;
      RECT 54.14 8.605 54.31 8.775 ;
      RECT 53.83 2.025 54 2.195 ;
      RECT 53.83 6.685 54 6.855 ;
      RECT 53.46 0.105 53.63 0.275 ;
      RECT 53.46 8.605 53.63 8.775 ;
      RECT 53.4 0.915 53.57 1.085 ;
      RECT 53.4 1.655 53.57 1.825 ;
      RECT 53.4 7.055 53.57 7.225 ;
      RECT 53.4 7.795 53.57 7.965 ;
      RECT 53.025 2.395 53.195 2.565 ;
      RECT 53.025 6.315 53.195 6.485 ;
      RECT 52.78 0.105 52.95 0.275 ;
      RECT 52.78 8.605 52.95 8.775 ;
      RECT 52.1 0.105 52.27 0.275 ;
      RECT 52.1 8.605 52.27 8.775 ;
      RECT 50.815 1.565 50.985 1.735 ;
      RECT 50.355 1.565 50.525 1.735 ;
      RECT 49.965 2.905 50.135 3.075 ;
      RECT 49.895 1.565 50.065 1.735 ;
      RECT 49.755 2.245 49.925 2.415 ;
      RECT 49.435 1.565 49.605 1.735 ;
      RECT 49.435 3.155 49.605 3.325 ;
      RECT 49.38 8.605 49.55 8.775 ;
      RECT 49.07 6.685 49.24 6.855 ;
      RECT 49.055 2.745 49.225 2.915 ;
      RECT 48.975 1.565 49.145 1.735 ;
      RECT 48.835 3.315 49.005 3.485 ;
      RECT 48.815 3.715 48.985 3.885 ;
      RECT 48.7 8.605 48.87 8.775 ;
      RECT 48.645 2.265 48.815 2.435 ;
      RECT 48.64 7.055 48.81 7.225 ;
      RECT 48.64 7.795 48.81 7.965 ;
      RECT 48.515 1.565 48.685 1.735 ;
      RECT 48.265 6.315 48.435 6.485 ;
      RECT 48.145 3.245 48.315 3.415 ;
      RECT 48.055 1.565 48.225 1.735 ;
      RECT 48.02 8.605 48.19 8.775 ;
      RECT 47.825 2.935 47.995 3.105 ;
      RECT 47.755 3.715 47.925 3.885 ;
      RECT 47.595 1.565 47.765 1.735 ;
      RECT 47.355 3.695 47.525 3.865 ;
      RECT 47.34 8.605 47.51 8.775 ;
      RECT 47.315 2.185 47.485 2.355 ;
      RECT 47.135 1.565 47.305 1.735 ;
      RECT 46.675 1.565 46.845 1.735 ;
      RECT 46.415 2.685 46.585 2.855 ;
      RECT 46.415 3.145 46.585 3.315 ;
      RECT 46.415 3.655 46.585 3.825 ;
      RECT 46.305 2.215 46.475 2.385 ;
      RECT 46.215 1.565 46.385 1.735 ;
      RECT 45.835 3.725 46.005 3.895 ;
      RECT 45.755 1.565 45.925 1.735 ;
      RECT 45.355 2.255 45.525 2.425 ;
      RECT 45.295 1.565 45.465 1.735 ;
      RECT 45.145 2.635 45.315 2.805 ;
      RECT 44.835 1.565 45.005 1.735 ;
      RECT 44.645 3.235 44.815 3.405 ;
      RECT 44.525 2.685 44.695 2.855 ;
      RECT 44.375 1.565 44.545 1.735 ;
      RECT 44.355 2.135 44.525 2.305 ;
      RECT 43.985 3.165 44.155 3.335 ;
      RECT 43.915 1.565 44.085 1.735 ;
      RECT 43.495 2.765 43.665 2.935 ;
      RECT 43.455 1.565 43.625 1.735 ;
      RECT 43.445 3.535 43.615 3.705 ;
      RECT 42.995 1.565 43.165 1.735 ;
      RECT 42.955 3.165 43.125 3.335 ;
      RECT 42.925 2.265 43.095 2.435 ;
      RECT 42.565 2.665 42.735 2.835 ;
      RECT 42.535 1.565 42.705 1.735 ;
      RECT 42.355 3.475 42.525 3.645 ;
      RECT 42.075 1.565 42.245 1.735 ;
      RECT 42.055 2.905 42.225 3.075 ;
      RECT 41.615 1.565 41.785 1.735 ;
      RECT 41.355 2.695 41.525 2.865 ;
      RECT 41.155 1.565 41.325 1.735 ;
      RECT 41.035 3.145 41.205 3.315 ;
      RECT 40.695 1.565 40.865 1.735 ;
      RECT 40.615 3.175 40.785 3.345 ;
      RECT 40.445 2.165 40.615 2.335 ;
      RECT 40.275 2.615 40.445 2.785 ;
      RECT 40.235 1.565 40.405 1.735 ;
      RECT 39.775 1.565 39.945 1.735 ;
      RECT 39.355 2.265 39.525 2.435 ;
      RECT 39.345 3.585 39.515 3.755 ;
      RECT 39.315 1.565 39.485 1.735 ;
      RECT 38.255 7.8 38.425 7.97 ;
      RECT 37.905 0.1 38.075 0.27 ;
      RECT 37.905 8.61 38.075 8.78 ;
      RECT 37.885 2.76 38.055 2.93 ;
      RECT 37.885 5.95 38.055 6.12 ;
      RECT 37.265 0.91 37.435 1.08 ;
      RECT 37.265 2.39 37.435 2.56 ;
      RECT 37.265 6.32 37.435 6.49 ;
      RECT 37.265 7.8 37.435 7.97 ;
      RECT 36.915 0.1 37.085 0.27 ;
      RECT 36.915 8.61 37.085 8.78 ;
      RECT 36.895 2.76 37.065 2.93 ;
      RECT 36.895 5.95 37.065 6.12 ;
      RECT 36.215 0.105 36.385 0.275 ;
      RECT 36.215 8.605 36.385 8.775 ;
      RECT 35.905 2.025 36.075 2.195 ;
      RECT 35.905 6.685 36.075 6.855 ;
      RECT 35.535 0.105 35.705 0.275 ;
      RECT 35.535 8.605 35.705 8.775 ;
      RECT 35.475 0.915 35.645 1.085 ;
      RECT 35.475 1.655 35.645 1.825 ;
      RECT 35.475 7.055 35.645 7.225 ;
      RECT 35.475 7.795 35.645 7.965 ;
      RECT 35.1 2.395 35.27 2.565 ;
      RECT 35.1 6.315 35.27 6.485 ;
      RECT 34.855 0.105 35.025 0.275 ;
      RECT 34.855 8.605 35.025 8.775 ;
      RECT 34.175 0.105 34.345 0.275 ;
      RECT 34.175 8.605 34.345 8.775 ;
      RECT 32.89 1.565 33.06 1.735 ;
      RECT 32.43 1.565 32.6 1.735 ;
      RECT 32.04 2.905 32.21 3.075 ;
      RECT 31.97 1.565 32.14 1.735 ;
      RECT 31.83 2.245 32 2.415 ;
      RECT 31.51 1.565 31.68 1.735 ;
      RECT 31.51 3.155 31.68 3.325 ;
      RECT 31.455 8.605 31.625 8.775 ;
      RECT 31.145 6.685 31.315 6.855 ;
      RECT 31.13 2.745 31.3 2.915 ;
      RECT 31.05 1.565 31.22 1.735 ;
      RECT 30.91 3.315 31.08 3.485 ;
      RECT 30.89 3.715 31.06 3.885 ;
      RECT 30.775 8.605 30.945 8.775 ;
      RECT 30.72 2.265 30.89 2.435 ;
      RECT 30.715 7.055 30.885 7.225 ;
      RECT 30.715 7.795 30.885 7.965 ;
      RECT 30.59 1.565 30.76 1.735 ;
      RECT 30.34 6.315 30.51 6.485 ;
      RECT 30.22 3.245 30.39 3.415 ;
      RECT 30.13 1.565 30.3 1.735 ;
      RECT 30.095 8.605 30.265 8.775 ;
      RECT 29.9 2.935 30.07 3.105 ;
      RECT 29.83 3.715 30 3.885 ;
      RECT 29.67 1.565 29.84 1.735 ;
      RECT 29.43 3.695 29.6 3.865 ;
      RECT 29.415 8.605 29.585 8.775 ;
      RECT 29.39 2.185 29.56 2.355 ;
      RECT 29.21 1.565 29.38 1.735 ;
      RECT 28.75 1.565 28.92 1.735 ;
      RECT 28.49 2.685 28.66 2.855 ;
      RECT 28.49 3.145 28.66 3.315 ;
      RECT 28.49 3.655 28.66 3.825 ;
      RECT 28.38 2.215 28.55 2.385 ;
      RECT 28.29 1.565 28.46 1.735 ;
      RECT 27.91 3.725 28.08 3.895 ;
      RECT 27.83 1.565 28 1.735 ;
      RECT 27.43 2.255 27.6 2.425 ;
      RECT 27.37 1.565 27.54 1.735 ;
      RECT 27.22 2.635 27.39 2.805 ;
      RECT 26.91 1.565 27.08 1.735 ;
      RECT 26.72 3.235 26.89 3.405 ;
      RECT 26.6 2.685 26.77 2.855 ;
      RECT 26.45 1.565 26.62 1.735 ;
      RECT 26.43 2.135 26.6 2.305 ;
      RECT 26.06 3.165 26.23 3.335 ;
      RECT 25.99 1.565 26.16 1.735 ;
      RECT 25.57 2.765 25.74 2.935 ;
      RECT 25.53 1.565 25.7 1.735 ;
      RECT 25.52 3.535 25.69 3.705 ;
      RECT 25.07 1.565 25.24 1.735 ;
      RECT 25.03 3.165 25.2 3.335 ;
      RECT 25 2.265 25.17 2.435 ;
      RECT 24.64 2.665 24.81 2.835 ;
      RECT 24.61 1.565 24.78 1.735 ;
      RECT 24.43 3.475 24.6 3.645 ;
      RECT 24.15 1.565 24.32 1.735 ;
      RECT 24.13 2.905 24.3 3.075 ;
      RECT 23.69 1.565 23.86 1.735 ;
      RECT 23.43 2.695 23.6 2.865 ;
      RECT 23.23 1.565 23.4 1.735 ;
      RECT 23.11 3.145 23.28 3.315 ;
      RECT 22.77 1.565 22.94 1.735 ;
      RECT 22.69 3.175 22.86 3.345 ;
      RECT 22.52 2.165 22.69 2.335 ;
      RECT 22.35 2.615 22.52 2.785 ;
      RECT 22.31 1.565 22.48 1.735 ;
      RECT 21.85 1.565 22.02 1.735 ;
      RECT 21.43 2.265 21.6 2.435 ;
      RECT 21.42 3.585 21.59 3.755 ;
      RECT 21.39 1.565 21.56 1.735 ;
      RECT 20.33 7.8 20.5 7.97 ;
      RECT 19.98 0.1 20.15 0.27 ;
      RECT 19.98 8.61 20.15 8.78 ;
      RECT 19.96 2.76 20.13 2.93 ;
      RECT 19.96 5.95 20.13 6.12 ;
      RECT 19.34 0.91 19.51 1.08 ;
      RECT 19.34 2.39 19.51 2.56 ;
      RECT 19.34 6.32 19.51 6.49 ;
      RECT 19.34 7.8 19.51 7.97 ;
      RECT 18.99 0.1 19.16 0.27 ;
      RECT 18.99 8.61 19.16 8.78 ;
      RECT 18.97 2.76 19.14 2.93 ;
      RECT 18.97 5.95 19.14 6.12 ;
      RECT 18.29 0.105 18.46 0.275 ;
      RECT 18.29 8.605 18.46 8.775 ;
      RECT 17.98 2.025 18.15 2.195 ;
      RECT 17.98 6.685 18.15 6.855 ;
      RECT 17.61 0.105 17.78 0.275 ;
      RECT 17.61 8.605 17.78 8.775 ;
      RECT 17.55 0.915 17.72 1.085 ;
      RECT 17.55 1.655 17.72 1.825 ;
      RECT 17.55 7.055 17.72 7.225 ;
      RECT 17.55 7.795 17.72 7.965 ;
      RECT 17.175 2.395 17.345 2.565 ;
      RECT 17.175 6.315 17.345 6.485 ;
      RECT 16.93 0.105 17.1 0.275 ;
      RECT 16.93 8.605 17.1 8.775 ;
      RECT 16.25 0.105 16.42 0.275 ;
      RECT 16.25 8.605 16.42 8.775 ;
      RECT 14.965 1.565 15.135 1.735 ;
      RECT 14.505 1.565 14.675 1.735 ;
      RECT 14.115 2.905 14.285 3.075 ;
      RECT 14.045 1.565 14.215 1.735 ;
      RECT 13.905 2.245 14.075 2.415 ;
      RECT 13.585 1.565 13.755 1.735 ;
      RECT 13.585 3.155 13.755 3.325 ;
      RECT 13.53 8.605 13.7 8.775 ;
      RECT 13.22 6.685 13.39 6.855 ;
      RECT 13.205 2.745 13.375 2.915 ;
      RECT 13.125 1.565 13.295 1.735 ;
      RECT 12.985 3.315 13.155 3.485 ;
      RECT 12.965 3.715 13.135 3.885 ;
      RECT 12.85 8.605 13.02 8.775 ;
      RECT 12.795 2.265 12.965 2.435 ;
      RECT 12.79 7.055 12.96 7.225 ;
      RECT 12.79 7.795 12.96 7.965 ;
      RECT 12.665 1.565 12.835 1.735 ;
      RECT 12.415 6.315 12.585 6.485 ;
      RECT 12.295 3.245 12.465 3.415 ;
      RECT 12.205 1.565 12.375 1.735 ;
      RECT 12.17 8.605 12.34 8.775 ;
      RECT 11.975 2.935 12.145 3.105 ;
      RECT 11.905 3.715 12.075 3.885 ;
      RECT 11.745 1.565 11.915 1.735 ;
      RECT 11.505 3.695 11.675 3.865 ;
      RECT 11.49 8.605 11.66 8.775 ;
      RECT 11.465 2.185 11.635 2.355 ;
      RECT 11.285 1.565 11.455 1.735 ;
      RECT 10.825 1.565 10.995 1.735 ;
      RECT 10.565 2.685 10.735 2.855 ;
      RECT 10.565 3.145 10.735 3.315 ;
      RECT 10.565 3.655 10.735 3.825 ;
      RECT 10.455 2.215 10.625 2.385 ;
      RECT 10.365 1.565 10.535 1.735 ;
      RECT 9.985 3.725 10.155 3.895 ;
      RECT 9.905 1.565 10.075 1.735 ;
      RECT 9.505 2.255 9.675 2.425 ;
      RECT 9.445 1.565 9.615 1.735 ;
      RECT 9.295 2.635 9.465 2.805 ;
      RECT 8.985 1.565 9.155 1.735 ;
      RECT 8.795 3.235 8.965 3.405 ;
      RECT 8.675 2.685 8.845 2.855 ;
      RECT 8.525 1.565 8.695 1.735 ;
      RECT 8.505 2.135 8.675 2.305 ;
      RECT 8.135 3.165 8.305 3.335 ;
      RECT 8.065 1.565 8.235 1.735 ;
      RECT 7.645 2.765 7.815 2.935 ;
      RECT 7.605 1.565 7.775 1.735 ;
      RECT 7.595 3.535 7.765 3.705 ;
      RECT 7.145 1.565 7.315 1.735 ;
      RECT 7.105 3.165 7.275 3.335 ;
      RECT 7.075 2.265 7.245 2.435 ;
      RECT 6.715 2.665 6.885 2.835 ;
      RECT 6.685 1.565 6.855 1.735 ;
      RECT 6.505 3.475 6.675 3.645 ;
      RECT 6.225 1.565 6.395 1.735 ;
      RECT 6.205 2.905 6.375 3.075 ;
      RECT 5.765 1.565 5.935 1.735 ;
      RECT 5.505 2.695 5.675 2.865 ;
      RECT 5.305 1.565 5.475 1.735 ;
      RECT 5.185 3.145 5.355 3.315 ;
      RECT 4.845 1.565 5.015 1.735 ;
      RECT 4.765 3.175 4.935 3.345 ;
      RECT 4.595 2.165 4.765 2.335 ;
      RECT 4.425 2.615 4.595 2.785 ;
      RECT 4.385 1.565 4.555 1.735 ;
      RECT 3.925 1.565 4.095 1.735 ;
      RECT 3.505 2.265 3.675 2.435 ;
      RECT 3.495 3.585 3.665 3.755 ;
      RECT 3.465 1.565 3.635 1.735 ;
      RECT 2.5 8.605 2.67 8.775 ;
      RECT 1.82 8.605 1.99 8.775 ;
      RECT 1.76 7.055 1.93 7.225 ;
      RECT 1.76 7.795 1.93 7.965 ;
      RECT 1.385 6.315 1.555 6.485 ;
      RECT 1.14 8.605 1.31 8.775 ;
      RECT 0.46 8.605 0.63 8.775 ;
    LAYER li1 ;
      RECT 86.075 0 86.245 2.235 ;
      RECT 85.115 0 85.285 2.235 ;
      RECT 84.155 0 84.325 2.235 ;
      RECT 83.635 0 83.805 2.235 ;
      RECT 82.675 0 82.845 2.235 ;
      RECT 81.675 0 81.845 2.235 ;
      RECT 80.715 0 80.885 2.235 ;
      RECT 79.235 0 79.405 2.235 ;
      RECT 77.315 0 77.485 2.235 ;
      RECT 75.835 0 76.005 2.235 ;
      RECT 68.15 0 68.32 2.235 ;
      RECT 67.19 0 67.36 2.235 ;
      RECT 66.23 0 66.4 2.235 ;
      RECT 65.71 0 65.88 2.235 ;
      RECT 64.75 0 64.92 2.235 ;
      RECT 63.75 0 63.92 2.235 ;
      RECT 62.79 0 62.96 2.235 ;
      RECT 61.31 0 61.48 2.235 ;
      RECT 59.39 0 59.56 2.235 ;
      RECT 57.91 0 58.08 2.235 ;
      RECT 50.225 0 50.395 2.235 ;
      RECT 49.265 0 49.435 2.235 ;
      RECT 48.305 0 48.475 2.235 ;
      RECT 47.785 0 47.955 2.235 ;
      RECT 46.825 0 46.995 2.235 ;
      RECT 45.825 0 45.995 2.235 ;
      RECT 44.865 0 45.035 2.235 ;
      RECT 43.385 0 43.555 2.235 ;
      RECT 41.465 0 41.635 2.235 ;
      RECT 39.985 0 40.155 2.235 ;
      RECT 32.3 0 32.47 2.235 ;
      RECT 31.34 0 31.51 2.235 ;
      RECT 30.38 0 30.55 2.235 ;
      RECT 29.86 0 30.03 2.235 ;
      RECT 28.9 0 29.07 2.235 ;
      RECT 27.9 0 28.07 2.235 ;
      RECT 26.94 0 27.11 2.235 ;
      RECT 25.46 0 25.63 2.235 ;
      RECT 23.54 0 23.71 2.235 ;
      RECT 22.06 0 22.23 2.235 ;
      RECT 14.375 0 14.545 2.235 ;
      RECT 13.415 0 13.585 2.235 ;
      RECT 12.455 0 12.625 2.235 ;
      RECT 11.935 0 12.105 2.235 ;
      RECT 10.975 0 11.145 2.235 ;
      RECT 9.975 0 10.145 2.235 ;
      RECT 9.015 0 9.185 2.235 ;
      RECT 7.535 0 7.705 2.235 ;
      RECT 5.615 0 5.785 2.235 ;
      RECT 4.135 0 4.305 2.235 ;
      RECT 75.025 0 86.985 1.735 ;
      RECT 57.1 0 69.06 1.735 ;
      RECT 39.175 0 51.135 1.735 ;
      RECT 21.25 0 33.21 1.735 ;
      RECT 3.325 0 15.285 1.735 ;
      RECT 75.02 0 86.985 1.68 ;
      RECT 57.095 0 69.06 1.68 ;
      RECT 39.17 0 51.135 1.68 ;
      RECT 21.245 0 33.21 1.68 ;
      RECT 3.32 0 15.285 1.68 ;
      RECT 87.87 0 88.04 0.935 ;
      RECT 69.945 0 70.115 0.935 ;
      RECT 52.02 0 52.19 0.935 ;
      RECT 34.095 0 34.265 0.935 ;
      RECT 16.17 0 16.34 0.935 ;
      RECT 91.6 0 91.77 0.93 ;
      RECT 90.61 0 90.78 0.93 ;
      RECT 73.675 0 73.845 0.93 ;
      RECT 72.685 0 72.855 0.93 ;
      RECT 55.75 0 55.92 0.93 ;
      RECT 54.76 0 54.93 0.93 ;
      RECT 37.825 0 37.995 0.93 ;
      RECT 36.835 0 37.005 0.93 ;
      RECT 19.9 0 20.07 0.93 ;
      RECT 18.91 0 19.08 0.93 ;
      RECT 92.395 0 92.575 0.305 ;
      RECT 74.47 0 90.445 0.305 ;
      RECT 56.545 0 72.52 0.305 ;
      RECT 38.62 0 54.595 0.305 ;
      RECT 20.695 0 36.67 0.305 ;
      RECT 0 0 18.745 0.305 ;
      RECT 0 0 92.575 0.3 ;
      RECT 0.025 8.58 92.575 8.88 ;
      RECT 92.395 8.575 92.575 8.88 ;
      RECT 91.6 7.95 91.77 8.88 ;
      RECT 90.61 7.95 90.78 8.88 ;
      RECT 74.47 8.575 90.445 8.88 ;
      RECT 73.675 7.95 73.845 8.88 ;
      RECT 72.685 7.95 72.855 8.88 ;
      RECT 56.545 8.575 72.52 8.88 ;
      RECT 55.75 7.95 55.92 8.88 ;
      RECT 54.76 7.95 54.93 8.88 ;
      RECT 38.62 8.575 54.595 8.88 ;
      RECT 37.825 7.95 37.995 8.88 ;
      RECT 36.835 7.95 37.005 8.88 ;
      RECT 20.695 8.575 36.67 8.88 ;
      RECT 19.9 7.95 20.07 8.88 ;
      RECT 18.91 7.95 19.08 8.88 ;
      RECT 0.025 8.575 18.745 8.88 ;
      RECT 87.87 7.945 88.04 8.88 ;
      RECT 83.11 7.945 83.28 8.88 ;
      RECT 69.945 7.945 70.115 8.88 ;
      RECT 65.185 7.945 65.355 8.88 ;
      RECT 52.02 7.945 52.19 8.88 ;
      RECT 47.26 7.945 47.43 8.88 ;
      RECT 34.095 7.945 34.265 8.88 ;
      RECT 29.335 7.945 29.505 8.88 ;
      RECT 16.17 7.945 16.34 8.88 ;
      RECT 11.41 7.945 11.58 8.88 ;
      RECT 0.025 8.565 0.83 8.88 ;
      RECT 0.32 8.545 0.55 8.88 ;
      RECT 0.38 7.945 0.55 8.88 ;
      RECT 92.03 5.02 92.2 6.49 ;
      RECT 92.03 6.315 92.205 6.485 ;
      RECT 91.66 1.74 91.83 2.93 ;
      RECT 91.66 1.74 92.13 1.91 ;
      RECT 91.66 6.97 92.13 7.14 ;
      RECT 91.66 5.95 91.83 7.14 ;
      RECT 90.67 1.74 90.84 2.93 ;
      RECT 90.67 1.74 91.14 1.91 ;
      RECT 90.67 6.97 91.14 7.14 ;
      RECT 90.67 5.95 90.84 7.14 ;
      RECT 88.82 2.635 88.99 3.865 ;
      RECT 88.875 0.855 89.045 2.805 ;
      RECT 88.82 0.575 88.99 1.025 ;
      RECT 88.82 7.855 88.99 8.305 ;
      RECT 88.875 6.075 89.045 8.025 ;
      RECT 88.82 5.015 88.99 6.245 ;
      RECT 88.3 0.575 88.47 3.865 ;
      RECT 88.3 2.075 88.705 2.405 ;
      RECT 88.3 1.235 88.705 1.565 ;
      RECT 88.3 5.015 88.47 8.305 ;
      RECT 88.3 7.315 88.705 7.645 ;
      RECT 88.3 6.475 88.705 6.805 ;
      RECT 86.395 3.39 86.415 3.44 ;
      RECT 86.375 3.362 86.395 3.555 ;
      RECT 86.355 3.337 86.375 3.611 ;
      RECT 86.315 3.325 86.355 3.63 ;
      RECT 86.265 3.32 86.315 3.659 ;
      RECT 86.261 3.314 86.265 3.675 ;
      RECT 86.175 3.306 86.261 3.675 ;
      RECT 86.115 3.294 86.175 3.67 ;
      RECT 86.061 3.284 86.115 3.659 ;
      RECT 85.975 3.272 86.061 3.642 ;
      RECT 85.953 3.263 85.975 3.629 ;
      RECT 85.867 3.256 85.953 3.616 ;
      RECT 85.781 3.243 85.867 3.595 ;
      RECT 85.695 3.231 85.781 3.575 ;
      RECT 85.665 3.22 85.695 3.561 ;
      RECT 85.615 3.207 85.665 3.551 ;
      RECT 85.595 3.197 85.615 3.545 ;
      RECT 85.541 3.187 85.595 3.539 ;
      RECT 85.455 3.167 85.541 3.523 ;
      RECT 85.415 3.155 85.455 3.509 ;
      RECT 85.38 3.155 85.415 3.495 ;
      RECT 85.365 3.155 85.38 3.48 ;
      RECT 85.315 3.155 85.365 3.425 ;
      RECT 85.285 3.155 85.315 3.345 ;
      RECT 85.815 2.825 85.985 3.075 ;
      RECT 85.815 2.825 85.995 3.03 ;
      RECT 85.875 2.655 86.005 2.975 ;
      RECT 85.875 2.662 86.015 2.94 ;
      RECT 85.835 2.677 86.025 2.875 ;
      RECT 85.825 2.76 86.025 2.875 ;
      RECT 85.835 2.695 86.035 2.785 ;
      RECT 85.835 2.675 86.015 2.94 ;
      RECT 85.605 1.93 85.775 2.415 ;
      RECT 85.595 1.93 85.775 2.405 ;
      RECT 85.595 1.945 85.795 2.35 ;
      RECT 85.555 1.925 85.745 2.315 ;
      RECT 85.555 1.96 85.805 2.235 ;
      RECT 85.505 1.945 85.795 2.135 ;
      RECT 85.505 1.975 85.815 2.095 ;
      RECT 85.505 1.99 85.825 2.015 ;
      RECT 85.101 2.688 85.115 2.944 ;
      RECT 85.101 2.689 85.201 2.939 ;
      RECT 85.015 2.686 85.101 2.936 ;
      RECT 85.005 2.685 85.015 2.929 ;
      RECT 85.005 2.692 85.287 2.926 ;
      RECT 84.925 2.695 85.287 2.922 ;
      RECT 85.005 2.694 85.305 2.919 ;
      RECT 84.915 2.707 85.325 2.916 ;
      RECT 84.925 2.695 85.325 2.916 ;
      RECT 84.905 2.712 85.325 2.915 ;
      RECT 84.925 2.697 85.411 2.911 ;
      RECT 84.885 2.715 85.411 2.908 ;
      RECT 84.925 2.701 85.497 2.902 ;
      RECT 84.875 2.72 85.497 2.898 ;
      RECT 84.925 2.704 85.525 2.897 ;
      RECT 84.925 2.705 85.565 2.891 ;
      RECT 84.915 2.71 85.575 2.886 ;
      RECT 84.875 2.73 85.585 2.875 ;
      RECT 84.875 2.75 85.595 2.86 ;
      RECT 84.835 3.298 84.855 3.605 ;
      RECT 84.825 3.273 84.835 3.885 ;
      RECT 84.785 3.24 84.825 3.885 ;
      RECT 84.781 3.21 84.785 3.885 ;
      RECT 84.695 3.095 84.781 3.885 ;
      RECT 84.685 2.97 84.695 3.885 ;
      RECT 84.675 2.935 84.685 3.885 ;
      RECT 84.665 2.905 84.675 3.885 ;
      RECT 84.645 2.875 84.665 3.77 ;
      RECT 84.635 2.845 84.645 3.645 ;
      RECT 84.625 2.825 84.635 3.595 ;
      RECT 84.605 2.795 84.625 3.503 ;
      RECT 84.585 2.761 84.605 3.418 ;
      RECT 84.58 2.744 84.585 3.353 ;
      RECT 84.575 2.738 84.58 3.325 ;
      RECT 84.565 2.73 84.575 3.29 ;
      RECT 84.545 2.725 84.555 3.19 ;
      RECT 84.535 2.725 84.545 3.165 ;
      RECT 84.53 2.725 84.535 3.128 ;
      RECT 84.515 2.725 84.53 3.06 ;
      RECT 84.505 2.724 84.515 2.99 ;
      RECT 84.495 2.722 84.505 2.97 ;
      RECT 84.435 2.718 84.495 2.943 ;
      RECT 84.395 2.72 84.435 2.923 ;
      RECT 84.375 2.75 84.395 2.905 ;
      RECT 84.555 2.725 84.565 3.245 ;
      RECT 84.495 2.08 84.665 2.435 ;
      RECT 84.525 1.966 84.665 2.435 ;
      RECT 84.525 1.968 84.675 2.43 ;
      RECT 84.525 1.97 84.695 2.42 ;
      RECT 84.525 1.973 84.725 2.405 ;
      RECT 84.525 1.978 84.775 2.375 ;
      RECT 84.525 1.983 84.795 2.338 ;
      RECT 84.505 1.985 84.805 2.313 ;
      RECT 84.525 1.965 84.635 2.435 ;
      RECT 84.535 1.96 84.635 2.435 ;
      RECT 84.055 3.222 84.245 3.585 ;
      RECT 84.055 3.237 84.285 3.583 ;
      RECT 84.055 3.265 84.305 3.579 ;
      RECT 84.055 3.3 84.315 3.577 ;
      RECT 84.055 3.345 84.325 3.576 ;
      RECT 84.045 3.217 84.205 3.565 ;
      RECT 84.025 3.225 84.245 3.515 ;
      RECT 83.995 3.237 84.285 3.45 ;
      RECT 84.055 3.215 84.205 3.585 ;
      RECT 84.06 7.855 84.23 8.305 ;
      RECT 84.115 6.075 84.285 8.025 ;
      RECT 84.06 5.015 84.23 6.245 ;
      RECT 83.54 5.015 83.71 8.305 ;
      RECT 83.54 7.315 83.945 7.645 ;
      RECT 83.54 6.475 83.945 6.805 ;
      RECT 83.641 2.695 83.845 3.105 ;
      RECT 83.555 2.588 83.641 3.09 ;
      RECT 83.551 2.584 83.555 3.074 ;
      RECT 83.465 2.695 83.845 3.054 ;
      RECT 83.445 2.575 83.465 3.015 ;
      RECT 83.435 2.58 83.551 2.99 ;
      RECT 83.425 2.587 83.555 2.97 ;
      RECT 83.415 2.592 83.645 2.945 ;
      RECT 83.405 2.61 83.735 2.925 ;
      RECT 83.395 2.615 83.735 2.905 ;
      RECT 83.385 2.62 83.775 2.77 ;
      RECT 83.385 2.65 83.835 2.77 ;
      RECT 83.385 2.635 83.825 2.77 ;
      RECT 83.415 2.605 83.735 2.945 ;
      RECT 83.415 2.593 83.675 2.945 ;
      RECT 83.565 3.42 83.815 3.885 ;
      RECT 83.485 3.395 83.805 3.88 ;
      RECT 83.415 3.429 83.815 3.87 ;
      RECT 83.205 3.68 83.815 3.865 ;
      RECT 83.385 3.449 83.815 3.865 ;
      RECT 83.225 3.64 83.815 3.865 ;
      RECT 83.375 3.46 83.815 3.865 ;
      RECT 83.265 3.58 83.815 3.865 ;
      RECT 83.315 3.505 83.815 3.865 ;
      RECT 83.565 3.37 83.805 3.885 ;
      RECT 83.585 3.365 83.805 3.885 ;
      RECT 83.595 3.36 83.725 3.885 ;
      RECT 83.681 3.355 83.685 3.885 ;
      RECT 83.155 1.925 83.241 2.362 ;
      RECT 83.145 1.925 83.241 2.358 ;
      RECT 83.145 1.925 83.305 2.357 ;
      RECT 83.145 1.925 83.335 2.355 ;
      RECT 83.145 1.925 83.345 2.345 ;
      RECT 83.135 1.93 83.345 2.343 ;
      RECT 83.125 1.94 83.345 2.335 ;
      RECT 83.125 1.94 83.355 2.295 ;
      RECT 83.145 1.925 83.375 2.21 ;
      RECT 83.115 1.95 83.375 2.205 ;
      RECT 83.125 1.94 83.385 2.135 ;
      RECT 83.105 1.96 83.385 2.08 ;
      RECT 83.095 1.97 83.385 1.98 ;
      RECT 83.175 2.741 83.185 2.82 ;
      RECT 83.165 2.734 83.175 3.005 ;
      RECT 83.155 2.728 83.165 3.03 ;
      RECT 83.145 2.72 83.155 3.06 ;
      RECT 83.105 2.715 83.145 3.11 ;
      RECT 83.085 2.715 83.105 3.165 ;
      RECT 83.075 2.715 83.085 3.19 ;
      RECT 83.065 2.715 83.075 3.205 ;
      RECT 83.035 2.715 83.065 3.25 ;
      RECT 83.025 2.715 83.035 3.29 ;
      RECT 83.005 2.715 83.025 3.315 ;
      RECT 82.985 2.715 83.005 3.35 ;
      RECT 82.905 2.715 82.985 3.395 ;
      RECT 82.895 2.715 82.905 3.415 ;
      RECT 82.855 2.795 82.895 3.412 ;
      RECT 82.835 2.875 82.855 3.409 ;
      RECT 82.815 2.93 82.835 3.407 ;
      RECT 82.795 2.99 82.815 3.405 ;
      RECT 82.755 3.025 82.795 3.403 ;
      RECT 82.751 3.035 82.755 3.401 ;
      RECT 82.665 3.05 82.751 3.397 ;
      RECT 82.645 3.07 82.665 3.393 ;
      RECT 82.575 3.075 82.645 3.389 ;
      RECT 82.555 3.076 82.575 3.386 ;
      RECT 82.551 3.078 82.555 3.385 ;
      RECT 82.465 3.087 82.551 3.38 ;
      RECT 82.455 3.096 82.465 3.375 ;
      RECT 82.415 3.102 82.455 3.37 ;
      RECT 82.365 3.113 82.415 3.355 ;
      RECT 82.345 3.122 82.365 3.34 ;
      RECT 82.265 3.135 82.345 3.325 ;
      RECT 82.435 2.685 82.605 2.895 ;
      RECT 82.551 2.677 82.605 2.895 ;
      RECT 82.351 2.685 82.605 2.885 ;
      RECT 82.265 2.685 82.605 2.865 ;
      RECT 82.265 2.69 82.615 2.81 ;
      RECT 82.265 2.7 82.625 2.72 ;
      RECT 82.465 2.682 82.605 2.895 ;
      RECT 82.215 3.623 82.465 3.955 ;
      RECT 82.185 3.635 82.465 3.937 ;
      RECT 82.165 3.67 82.465 3.907 ;
      RECT 82.215 3.62 82.387 3.955 ;
      RECT 82.215 3.616 82.301 3.955 ;
      RECT 82.145 1.965 82.325 2.385 ;
      RECT 82.145 1.965 82.345 2.375 ;
      RECT 82.145 1.965 82.365 2.35 ;
      RECT 82.145 1.965 82.375 2.335 ;
      RECT 82.145 1.965 82.385 2.33 ;
      RECT 82.145 2.005 82.405 2.315 ;
      RECT 82.145 2.075 82.425 2.295 ;
      RECT 82.125 2.075 82.425 2.29 ;
      RECT 82.125 2.135 82.435 2.265 ;
      RECT 82.125 2.175 82.445 2.215 ;
      RECT 82.105 1.965 82.385 2.195 ;
      RECT 82.095 1.975 82.385 2.118 ;
      RECT 82.085 2.015 82.405 2.063 ;
      RECT 81.685 3.375 81.855 3.895 ;
      RECT 81.675 3.375 81.855 3.855 ;
      RECT 81.665 3.395 81.855 3.83 ;
      RECT 81.675 3.375 81.865 3.825 ;
      RECT 81.655 3.435 81.865 3.795 ;
      RECT 81.645 3.47 81.865 3.775 ;
      RECT 81.635 3.52 81.865 3.735 ;
      RECT 81.675 3.386 81.875 3.725 ;
      RECT 81.625 3.6 81.875 3.675 ;
      RECT 81.665 3.409 81.885 3.605 ;
      RECT 81.665 3.433 81.895 3.5 ;
      RECT 81.605 2.68 81.625 2.955 ;
      RECT 81.565 2.665 81.605 3 ;
      RECT 81.545 2.65 81.565 3.065 ;
      RECT 81.525 2.649 81.545 3.14 ;
      RECT 81.505 2.657 81.525 3.245 ;
      RECT 81.501 2.662 81.505 3.297 ;
      RECT 81.415 2.681 81.501 3.337 ;
      RECT 81.405 2.702 81.415 3.376 ;
      RECT 81.395 2.71 81.405 3.377 ;
      RECT 81.375 2.845 81.395 3.379 ;
      RECT 81.365 2.995 81.375 3.381 ;
      RECT 81.325 3.08 81.365 3.386 ;
      RECT 81.243 3.102 81.325 3.396 ;
      RECT 81.157 3.117 81.243 3.409 ;
      RECT 81.071 3.132 81.157 3.422 ;
      RECT 80.985 3.147 81.071 3.436 ;
      RECT 80.905 3.161 80.985 3.449 ;
      RECT 80.891 3.169 80.905 3.457 ;
      RECT 80.805 3.177 80.891 3.471 ;
      RECT 80.795 3.185 80.805 3.484 ;
      RECT 80.771 3.185 80.795 3.492 ;
      RECT 80.685 3.187 80.771 3.522 ;
      RECT 80.605 3.189 80.685 3.565 ;
      RECT 80.535 3.192 80.605 3.6 ;
      RECT 80.515 3.194 80.535 3.616 ;
      RECT 80.485 3.2 80.515 3.618 ;
      RECT 80.435 3.215 80.485 3.621 ;
      RECT 80.415 3.23 80.435 3.624 ;
      RECT 80.385 3.235 80.415 3.627 ;
      RECT 80.325 3.25 80.385 3.631 ;
      RECT 80.315 3.266 80.325 3.635 ;
      RECT 80.265 3.276 80.315 3.624 ;
      RECT 80.235 3.295 80.265 3.607 ;
      RECT 80.215 3.315 80.235 3.597 ;
      RECT 80.195 3.34 80.215 3.589 ;
      RECT 81.205 1.932 81.375 2.425 ;
      RECT 81.195 1.932 81.375 2.41 ;
      RECT 81.195 1.947 81.405 2.4 ;
      RECT 81.185 1.947 81.405 2.375 ;
      RECT 81.175 1.947 81.405 2.34 ;
      RECT 81.175 1.955 81.415 2.295 ;
      RECT 81.155 1.925 81.345 2.275 ;
      RECT 81.145 1.932 81.375 2.235 ;
      RECT 81.135 1.947 81.405 2.215 ;
      RECT 81.125 1.96 81.415 2.175 ;
      RECT 81.115 1.975 81.415 2.128 ;
      RECT 81.115 1.975 81.425 2.12 ;
      RECT 81.105 1.99 81.425 2.093 ;
      RECT 81.115 1.985 81.435 2.035 ;
      RECT 80.915 2.612 81.185 2.905 ;
      RECT 80.915 2.614 81.195 2.9 ;
      RECT 80.905 2.64 81.195 2.895 ;
      RECT 80.915 2.63 81.205 2.89 ;
      RECT 80.915 2.608 81.151 2.905 ;
      RECT 80.915 2.605 81.065 2.905 ;
      RECT 80.975 2.6 81.061 2.905 ;
      RECT 80.465 2.648 80.535 2.945 ;
      RECT 80.465 2.648 80.545 2.944 ;
      RECT 80.545 2.635 80.555 2.941 ;
      RECT 80.445 2.662 80.555 2.935 ;
      RECT 80.535 2.64 80.625 2.931 ;
      RECT 80.465 2.655 80.645 2.92 ;
      RECT 80.445 2.72 80.655 2.916 ;
      RECT 80.425 2.668 80.645 2.915 ;
      RECT 80.415 2.673 80.645 2.905 ;
      RECT 80.405 2.795 80.665 2.9 ;
      RECT 80.405 2.875 80.675 2.89 ;
      RECT 80.375 2.681 80.645 2.884 ;
      RECT 80.365 2.695 80.645 2.869 ;
      RECT 80.405 2.676 80.645 2.9 ;
      RECT 80.535 2.636 80.555 2.941 ;
      RECT 80.355 2.072 80.375 2.305 ;
      RECT 80.345 2.053 80.355 2.31 ;
      RECT 80.335 2.041 80.345 2.317 ;
      RECT 80.295 2.027 80.335 2.327 ;
      RECT 80.285 2.017 80.295 2.336 ;
      RECT 80.235 2.002 80.285 2.341 ;
      RECT 80.225 1.987 80.235 2.347 ;
      RECT 80.205 1.978 80.225 2.352 ;
      RECT 80.195 1.968 80.205 2.358 ;
      RECT 80.185 1.965 80.195 2.363 ;
      RECT 80.165 1.965 80.185 2.364 ;
      RECT 80.135 1.96 80.165 2.362 ;
      RECT 80.111 1.953 80.135 2.361 ;
      RECT 80.025 1.943 80.111 2.358 ;
      RECT 80.015 1.935 80.025 2.355 ;
      RECT 79.993 1.935 80.015 2.354 ;
      RECT 79.907 1.935 79.993 2.352 ;
      RECT 79.821 1.935 79.907 2.35 ;
      RECT 79.735 1.935 79.821 2.347 ;
      RECT 79.725 1.935 79.735 2.34 ;
      RECT 79.695 1.935 79.725 2.3 ;
      RECT 79.685 1.945 79.695 2.255 ;
      RECT 79.675 1.99 79.685 2.24 ;
      RECT 79.645 2.085 79.675 2.195 ;
      RECT 79.835 2.822 80.005 3.335 ;
      RECT 79.825 2.853 80.005 3.315 ;
      RECT 79.825 2.853 80.025 3.285 ;
      RECT 79.815 2.861 80.025 3.26 ;
      RECT 79.815 2.861 80.035 3.25 ;
      RECT 79.815 2.861 80.045 3.23 ;
      RECT 79.815 2.861 80.095 3.185 ;
      RECT 79.815 2.861 80.105 3.16 ;
      RECT 79.815 2.861 80.115 3.125 ;
      RECT 79.815 2.861 80.125 3.09 ;
      RECT 79.815 2.861 80.135 3.04 ;
      RECT 79.815 2.861 80.155 2.965 ;
      RECT 79.985 2.725 80.165 2.905 ;
      RECT 79.905 2.78 80.165 2.905 ;
      RECT 79.945 2.745 80.005 3.335 ;
      RECT 79.935 2.765 80.165 2.905 ;
      RECT 79.295 3.235 79.381 3.801 ;
      RECT 79.255 3.235 79.381 3.795 ;
      RECT 79.255 3.235 79.467 3.793 ;
      RECT 79.255 3.235 79.505 3.787 ;
      RECT 79.255 3.242 79.515 3.785 ;
      RECT 79.225 3.235 79.505 3.78 ;
      RECT 79.195 3.25 79.515 3.77 ;
      RECT 79.195 3.277 79.555 3.762 ;
      RECT 79.17 3.277 79.555 3.75 ;
      RECT 79.17 3.315 79.565 3.732 ;
      RECT 79.155 3.297 79.555 3.725 ;
      RECT 79.155 3.345 79.575 3.721 ;
      RECT 79.155 3.411 79.595 3.705 ;
      RECT 79.155 3.466 79.605 3.515 ;
      RECT 79.345 2.755 79.515 2.935 ;
      RECT 79.295 2.694 79.345 2.92 ;
      RECT 79.035 2.675 79.295 2.905 ;
      RECT 78.995 2.735 79.465 2.905 ;
      RECT 78.995 2.725 79.425 2.905 ;
      RECT 78.995 2.714 79.405 2.905 ;
      RECT 78.995 2.7 79.345 2.905 ;
      RECT 79.035 2.67 79.231 2.905 ;
      RECT 79.065 2.649 79.231 2.905 ;
      RECT 79.045 2.65 79.231 2.905 ;
      RECT 79.065 2.635 79.145 2.905 ;
      RECT 78.825 3.165 78.945 3.605 ;
      RECT 78.805 3.165 78.945 3.604 ;
      RECT 78.765 3.185 78.945 3.601 ;
      RECT 78.725 3.229 78.945 3.597 ;
      RECT 78.715 3.259 78.965 3.46 ;
      RECT 78.805 3.165 78.975 3.355 ;
      RECT 78.465 1.945 78.475 2.395 ;
      RECT 78.275 1.945 78.295 2.355 ;
      RECT 78.245 1.945 78.255 2.335 ;
      RECT 78.925 2.255 78.945 2.44 ;
      RECT 78.905 2.215 78.925 2.448 ;
      RECT 78.855 2.182 78.905 2.458 ;
      RECT 78.801 2.156 78.855 2.461 ;
      RECT 78.715 2.121 78.801 2.451 ;
      RECT 78.705 2.097 78.715 2.44 ;
      RECT 78.635 2.063 78.705 2.43 ;
      RECT 78.615 2.023 78.635 2.423 ;
      RECT 78.595 2.005 78.615 2.419 ;
      RECT 78.585 1.995 78.595 2.416 ;
      RECT 78.555 1.98 78.585 2.412 ;
      RECT 78.545 1.965 78.555 2.408 ;
      RECT 78.535 1.96 78.545 2.406 ;
      RECT 78.485 1.95 78.535 2.401 ;
      RECT 78.475 1.945 78.485 2.396 ;
      RECT 78.445 1.945 78.465 2.39 ;
      RECT 78.411 1.945 78.445 2.382 ;
      RECT 78.325 1.945 78.411 2.372 ;
      RECT 78.295 1.945 78.325 2.36 ;
      RECT 78.255 1.945 78.275 2.345 ;
      RECT 78.235 1.945 78.245 2.328 ;
      RECT 78.215 1.955 78.235 2.308 ;
      RECT 78.205 1.975 78.215 2.24 ;
      RECT 78.195 1.985 78.205 2 ;
      RECT 78.465 2.665 78.551 2.99 ;
      RECT 78.465 2.665 78.585 2.982 ;
      RECT 78.415 2.665 78.585 2.98 ;
      RECT 78.415 2.669 78.671 2.975 ;
      RECT 78.415 2.674 78.695 2.968 ;
      RECT 78.415 2.68 78.705 2.966 ;
      RECT 78.415 2.69 78.715 2.963 ;
      RECT 78.415 2.83 78.725 2.958 ;
      RECT 78.475 3.34 78.525 3.656 ;
      RECT 78.465 3.32 78.475 3.681 ;
      RECT 78.455 3.31 78.465 3.69 ;
      RECT 78.435 3.304 78.455 3.705 ;
      RECT 78.405 3.302 78.435 3.725 ;
      RECT 78.391 3.3 78.405 3.735 ;
      RECT 78.305 3.296 78.391 3.735 ;
      RECT 78.235 3.29 78.305 3.725 ;
      RECT 78.155 3.285 78.235 3.7 ;
      RECT 78.095 3.281 78.155 3.665 ;
      RECT 78.025 3.277 78.095 3.625 ;
      RECT 77.995 3.275 78.025 3.6 ;
      RECT 77.891 3.273 77.935 3.595 ;
      RECT 77.805 3.268 77.891 3.595 ;
      RECT 77.725 3.265 77.805 3.595 ;
      RECT 77.645 3.266 77.725 3.62 ;
      RECT 77.563 3.268 77.645 3.645 ;
      RECT 77.477 3.269 77.563 3.645 ;
      RECT 77.391 3.271 77.477 3.645 ;
      RECT 77.305 3.273 77.391 3.645 ;
      RECT 77.285 3.274 77.305 3.637 ;
      RECT 77.275 3.28 77.285 3.626 ;
      RECT 77.235 3.3 77.275 3.607 ;
      RECT 77.225 3.32 77.235 3.589 ;
      RECT 77.935 3.275 77.995 3.595 ;
      RECT 77.905 2.82 78.075 3.075 ;
      RECT 77.905 2.82 78.085 3.068 ;
      RECT 77.905 2.82 78.095 3.053 ;
      RECT 77.905 2.82 78.115 3.035 ;
      RECT 77.905 2.82 78.155 2.99 ;
      RECT 78.085 2.585 78.175 2.943 ;
      RECT 78.075 2.59 78.185 2.924 ;
      RECT 78.025 2.605 78.195 2.911 ;
      RECT 78.015 2.62 78.205 2.895 ;
      RECT 77.915 2.785 78.205 2.895 ;
      RECT 77.955 2.645 78.075 3.075 ;
      RECT 77.925 2.755 78.205 2.895 ;
      RECT 77.945 2.68 78.075 3.075 ;
      RECT 77.935 2.705 78.205 2.895 ;
      RECT 78.055 2.591 78.185 2.924 ;
      RECT 78.075 2.586 78.175 2.943 ;
      RECT 77.535 2.72 77.725 2.895 ;
      RECT 77.495 2.638 77.685 2.89 ;
      RECT 77.461 2.643 77.685 2.884 ;
      RECT 77.375 2.65 77.685 2.879 ;
      RECT 77.291 2.665 77.685 2.874 ;
      RECT 77.205 2.685 77.715 2.868 ;
      RECT 77.291 2.675 77.715 2.874 ;
      RECT 77.535 2.635 77.685 2.895 ;
      RECT 77.535 2.631 77.635 2.895 ;
      RECT 77.621 2.626 77.635 2.895 ;
      RECT 76.375 1.954 77.035 2.345 ;
      RECT 76.633 1.948 77.035 2.345 ;
      RECT 76.365 1.96 77.035 2.344 ;
      RECT 76.355 1.975 77.035 2.343 ;
      RECT 76.295 2.015 77.035 2.339 ;
      RECT 76.461 1.953 77.045 2.335 ;
      RECT 76.365 1.96 77.055 2.325 ;
      RECT 76.365 1.968 77.065 2.305 ;
      RECT 76.355 1.978 77.085 2.278 ;
      RECT 76.295 2.015 77.095 2.253 ;
      RECT 76.355 1.985 77.105 2.24 ;
      RECT 76.461 1.951 77.035 2.345 ;
      RECT 76.547 1.949 77.035 2.345 ;
      RECT 76.633 1.947 77.015 2.345 ;
      RECT 76.719 1.945 77.015 2.345 ;
      RECT 76.885 3.12 77.055 3.315 ;
      RECT 76.875 3.12 77.055 3.26 ;
      RECT 76.87 3.12 77.055 3.188 ;
      RECT 76.855 3.06 77.035 3.155 ;
      RECT 76.845 3.06 77.035 3.105 ;
      RECT 76.815 3.035 77.025 3.06 ;
      RECT 76.795 3.035 77.025 3.045 ;
      RECT 76.735 2.725 76.915 3.036 ;
      RECT 76.735 2.96 77.015 3.036 ;
      RECT 76.725 2.724 76.735 3.026 ;
      RECT 76.705 2.723 76.725 3.02 ;
      RECT 76.675 2.722 76.705 3 ;
      RECT 76.625 2.719 76.675 2.965 ;
      RECT 76.625 2.84 76.985 2.965 ;
      RECT 76.555 2.716 76.625 2.92 ;
      RECT 76.555 2.775 76.965 2.92 ;
      RECT 76.555 2.765 76.955 2.92 ;
      RECT 76.555 2.755 76.945 2.92 ;
      RECT 76.555 2.735 76.925 2.92 ;
      RECT 76.635 3.255 76.645 3.512 ;
      RECT 76.615 3.172 76.635 3.532 ;
      RECT 76.595 3.166 76.615 3.56 ;
      RECT 76.535 3.154 76.595 3.58 ;
      RECT 76.495 3.14 76.535 3.581 ;
      RECT 76.411 3.129 76.495 3.569 ;
      RECT 76.325 3.116 76.411 3.553 ;
      RECT 76.315 3.109 76.325 3.545 ;
      RECT 76.265 3.106 76.315 3.485 ;
      RECT 76.245 3.102 76.265 3.4 ;
      RECT 76.235 3.1 76.245 3.35 ;
      RECT 76.205 3.098 76.235 3.32 ;
      RECT 76.165 3.093 76.205 3.3 ;
      RECT 76.127 3.088 76.165 3.288 ;
      RECT 76.041 3.08 76.127 3.297 ;
      RECT 75.955 3.069 76.041 3.309 ;
      RECT 75.885 3.059 75.955 3.319 ;
      RECT 75.865 3.05 75.885 3.324 ;
      RECT 75.805 3.022 75.865 3.32 ;
      RECT 75.785 2.992 75.805 3.308 ;
      RECT 75.765 2.965 75.785 3.295 ;
      RECT 75.685 2.718 75.765 3.262 ;
      RECT 75.671 2.71 75.685 3.224 ;
      RECT 75.585 2.702 75.671 3.145 ;
      RECT 75.565 2.693 75.585 3.061 ;
      RECT 75.535 2.688 75.565 3.041 ;
      RECT 75.465 2.699 75.535 3.026 ;
      RECT 75.445 2.717 75.465 3 ;
      RECT 75.435 2.723 75.445 2.945 ;
      RECT 75.415 2.745 75.435 2.83 ;
      RECT 76.075 2.705 76.245 2.895 ;
      RECT 76.075 2.705 76.275 2.89 ;
      RECT 76.125 2.615 76.295 2.88 ;
      RECT 76.085 2.65 76.295 2.88 ;
      RECT 75.285 3.388 75.355 3.829 ;
      RECT 75.225 3.413 75.355 3.826 ;
      RECT 75.225 3.413 75.405 3.819 ;
      RECT 75.215 3.435 75.405 3.816 ;
      RECT 75.355 3.375 75.425 3.814 ;
      RECT 75.285 3.4 75.505 3.811 ;
      RECT 75.215 3.439 75.555 3.807 ;
      RECT 75.195 3.465 75.555 3.795 ;
      RECT 75.215 3.459 75.575 3.79 ;
      RECT 75.195 2.205 75.235 2.445 ;
      RECT 75.195 2.205 75.265 2.444 ;
      RECT 75.195 2.205 75.375 2.436 ;
      RECT 75.195 2.205 75.435 2.415 ;
      RECT 75.205 2.15 75.485 2.315 ;
      RECT 75.315 1.99 75.345 2.437 ;
      RECT 75.345 1.985 75.525 2.195 ;
      RECT 75.215 2.125 75.525 2.195 ;
      RECT 75.265 2.02 75.315 2.44 ;
      RECT 75.235 2.075 75.525 2.195 ;
      RECT 74.105 5.02 74.275 6.49 ;
      RECT 74.105 6.315 74.28 6.485 ;
      RECT 73.735 1.74 73.905 2.93 ;
      RECT 73.735 1.74 74.205 1.91 ;
      RECT 73.735 6.97 74.205 7.14 ;
      RECT 73.735 5.95 73.905 7.14 ;
      RECT 72.745 1.74 72.915 2.93 ;
      RECT 72.745 1.74 73.215 1.91 ;
      RECT 72.745 6.97 73.215 7.14 ;
      RECT 72.745 5.95 72.915 7.14 ;
      RECT 70.895 2.635 71.065 3.865 ;
      RECT 70.95 0.855 71.12 2.805 ;
      RECT 70.895 0.575 71.065 1.025 ;
      RECT 70.895 7.855 71.065 8.305 ;
      RECT 70.95 6.075 71.12 8.025 ;
      RECT 70.895 5.015 71.065 6.245 ;
      RECT 70.375 0.575 70.545 3.865 ;
      RECT 70.375 2.075 70.78 2.405 ;
      RECT 70.375 1.235 70.78 1.565 ;
      RECT 70.375 5.015 70.545 8.305 ;
      RECT 70.375 7.315 70.78 7.645 ;
      RECT 70.375 6.475 70.78 6.805 ;
      RECT 68.47 3.39 68.49 3.44 ;
      RECT 68.45 3.362 68.47 3.555 ;
      RECT 68.43 3.337 68.45 3.611 ;
      RECT 68.39 3.325 68.43 3.63 ;
      RECT 68.34 3.32 68.39 3.659 ;
      RECT 68.336 3.314 68.34 3.675 ;
      RECT 68.25 3.306 68.336 3.675 ;
      RECT 68.19 3.294 68.25 3.67 ;
      RECT 68.136 3.284 68.19 3.659 ;
      RECT 68.05 3.272 68.136 3.642 ;
      RECT 68.028 3.263 68.05 3.629 ;
      RECT 67.942 3.256 68.028 3.616 ;
      RECT 67.856 3.243 67.942 3.595 ;
      RECT 67.77 3.231 67.856 3.575 ;
      RECT 67.74 3.22 67.77 3.561 ;
      RECT 67.69 3.207 67.74 3.551 ;
      RECT 67.67 3.197 67.69 3.545 ;
      RECT 67.616 3.187 67.67 3.539 ;
      RECT 67.53 3.167 67.616 3.523 ;
      RECT 67.49 3.155 67.53 3.509 ;
      RECT 67.455 3.155 67.49 3.495 ;
      RECT 67.44 3.155 67.455 3.48 ;
      RECT 67.39 3.155 67.44 3.425 ;
      RECT 67.36 3.155 67.39 3.345 ;
      RECT 67.89 2.825 68.06 3.075 ;
      RECT 67.89 2.825 68.07 3.03 ;
      RECT 67.95 2.655 68.08 2.975 ;
      RECT 67.95 2.662 68.09 2.94 ;
      RECT 67.91 2.677 68.1 2.875 ;
      RECT 67.9 2.76 68.1 2.875 ;
      RECT 67.91 2.695 68.11 2.785 ;
      RECT 67.91 2.675 68.09 2.94 ;
      RECT 67.68 1.93 67.85 2.415 ;
      RECT 67.67 1.93 67.85 2.405 ;
      RECT 67.67 1.945 67.87 2.35 ;
      RECT 67.63 1.925 67.82 2.315 ;
      RECT 67.63 1.96 67.88 2.235 ;
      RECT 67.58 1.945 67.87 2.135 ;
      RECT 67.58 1.975 67.89 2.095 ;
      RECT 67.58 1.99 67.9 2.015 ;
      RECT 67.176 2.688 67.19 2.944 ;
      RECT 67.176 2.689 67.276 2.939 ;
      RECT 67.09 2.686 67.176 2.936 ;
      RECT 67.08 2.685 67.09 2.929 ;
      RECT 67.08 2.692 67.362 2.926 ;
      RECT 67 2.695 67.362 2.922 ;
      RECT 67.08 2.694 67.38 2.919 ;
      RECT 66.99 2.707 67.4 2.916 ;
      RECT 67 2.695 67.4 2.916 ;
      RECT 66.98 2.712 67.4 2.915 ;
      RECT 67 2.697 67.486 2.911 ;
      RECT 66.96 2.715 67.486 2.908 ;
      RECT 67 2.701 67.572 2.902 ;
      RECT 66.95 2.72 67.572 2.898 ;
      RECT 67 2.704 67.6 2.897 ;
      RECT 67 2.705 67.64 2.891 ;
      RECT 66.99 2.71 67.65 2.886 ;
      RECT 66.95 2.73 67.66 2.875 ;
      RECT 66.95 2.75 67.67 2.86 ;
      RECT 66.91 3.298 66.93 3.605 ;
      RECT 66.9 3.273 66.91 3.885 ;
      RECT 66.86 3.24 66.9 3.885 ;
      RECT 66.856 3.21 66.86 3.885 ;
      RECT 66.77 3.095 66.856 3.885 ;
      RECT 66.76 2.97 66.77 3.885 ;
      RECT 66.75 2.935 66.76 3.885 ;
      RECT 66.74 2.905 66.75 3.885 ;
      RECT 66.72 2.875 66.74 3.77 ;
      RECT 66.71 2.845 66.72 3.645 ;
      RECT 66.7 2.825 66.71 3.595 ;
      RECT 66.68 2.795 66.7 3.503 ;
      RECT 66.66 2.761 66.68 3.418 ;
      RECT 66.655 2.744 66.66 3.353 ;
      RECT 66.65 2.738 66.655 3.325 ;
      RECT 66.64 2.73 66.65 3.29 ;
      RECT 66.62 2.725 66.63 3.19 ;
      RECT 66.61 2.725 66.62 3.165 ;
      RECT 66.605 2.725 66.61 3.128 ;
      RECT 66.59 2.725 66.605 3.06 ;
      RECT 66.58 2.724 66.59 2.99 ;
      RECT 66.57 2.722 66.58 2.97 ;
      RECT 66.51 2.718 66.57 2.943 ;
      RECT 66.47 2.72 66.51 2.923 ;
      RECT 66.45 2.75 66.47 2.905 ;
      RECT 66.63 2.725 66.64 3.245 ;
      RECT 66.57 2.08 66.74 2.435 ;
      RECT 66.6 1.966 66.74 2.435 ;
      RECT 66.6 1.968 66.75 2.43 ;
      RECT 66.6 1.97 66.77 2.42 ;
      RECT 66.6 1.973 66.8 2.405 ;
      RECT 66.6 1.978 66.85 2.375 ;
      RECT 66.6 1.983 66.87 2.338 ;
      RECT 66.58 1.985 66.88 2.313 ;
      RECT 66.6 1.965 66.71 2.435 ;
      RECT 66.61 1.96 66.71 2.435 ;
      RECT 66.13 3.222 66.32 3.585 ;
      RECT 66.13 3.237 66.36 3.583 ;
      RECT 66.13 3.265 66.38 3.579 ;
      RECT 66.13 3.3 66.39 3.577 ;
      RECT 66.13 3.345 66.4 3.576 ;
      RECT 66.12 3.217 66.28 3.565 ;
      RECT 66.1 3.225 66.32 3.515 ;
      RECT 66.07 3.237 66.36 3.45 ;
      RECT 66.13 3.215 66.28 3.585 ;
      RECT 66.135 7.855 66.305 8.305 ;
      RECT 66.19 6.075 66.36 8.025 ;
      RECT 66.135 5.015 66.305 6.245 ;
      RECT 65.615 5.015 65.785 8.305 ;
      RECT 65.615 7.315 66.02 7.645 ;
      RECT 65.615 6.475 66.02 6.805 ;
      RECT 65.716 2.695 65.92 3.105 ;
      RECT 65.63 2.588 65.716 3.09 ;
      RECT 65.626 2.584 65.63 3.074 ;
      RECT 65.54 2.695 65.92 3.054 ;
      RECT 65.52 2.575 65.54 3.015 ;
      RECT 65.51 2.58 65.626 2.99 ;
      RECT 65.5 2.587 65.63 2.97 ;
      RECT 65.49 2.592 65.72 2.945 ;
      RECT 65.48 2.61 65.81 2.925 ;
      RECT 65.47 2.615 65.81 2.905 ;
      RECT 65.46 2.62 65.85 2.77 ;
      RECT 65.46 2.65 65.91 2.77 ;
      RECT 65.46 2.635 65.9 2.77 ;
      RECT 65.49 2.605 65.81 2.945 ;
      RECT 65.49 2.593 65.75 2.945 ;
      RECT 65.64 3.42 65.89 3.885 ;
      RECT 65.56 3.395 65.88 3.88 ;
      RECT 65.49 3.429 65.89 3.87 ;
      RECT 65.28 3.68 65.89 3.865 ;
      RECT 65.46 3.449 65.89 3.865 ;
      RECT 65.3 3.64 65.89 3.865 ;
      RECT 65.45 3.46 65.89 3.865 ;
      RECT 65.34 3.58 65.89 3.865 ;
      RECT 65.39 3.505 65.89 3.865 ;
      RECT 65.64 3.37 65.88 3.885 ;
      RECT 65.66 3.365 65.88 3.885 ;
      RECT 65.67 3.36 65.8 3.885 ;
      RECT 65.756 3.355 65.76 3.885 ;
      RECT 65.23 1.925 65.316 2.362 ;
      RECT 65.22 1.925 65.316 2.358 ;
      RECT 65.22 1.925 65.38 2.357 ;
      RECT 65.22 1.925 65.41 2.355 ;
      RECT 65.22 1.925 65.42 2.345 ;
      RECT 65.21 1.93 65.42 2.343 ;
      RECT 65.2 1.94 65.42 2.335 ;
      RECT 65.2 1.94 65.43 2.295 ;
      RECT 65.22 1.925 65.45 2.21 ;
      RECT 65.19 1.95 65.45 2.205 ;
      RECT 65.2 1.94 65.46 2.135 ;
      RECT 65.18 1.96 65.46 2.08 ;
      RECT 65.17 1.97 65.46 1.98 ;
      RECT 65.25 2.741 65.26 2.82 ;
      RECT 65.24 2.734 65.25 3.005 ;
      RECT 65.23 2.728 65.24 3.03 ;
      RECT 65.22 2.72 65.23 3.06 ;
      RECT 65.18 2.715 65.22 3.11 ;
      RECT 65.16 2.715 65.18 3.165 ;
      RECT 65.15 2.715 65.16 3.19 ;
      RECT 65.14 2.715 65.15 3.205 ;
      RECT 65.11 2.715 65.14 3.25 ;
      RECT 65.1 2.715 65.11 3.29 ;
      RECT 65.08 2.715 65.1 3.315 ;
      RECT 65.06 2.715 65.08 3.35 ;
      RECT 64.98 2.715 65.06 3.395 ;
      RECT 64.97 2.715 64.98 3.415 ;
      RECT 64.93 2.795 64.97 3.412 ;
      RECT 64.91 2.875 64.93 3.409 ;
      RECT 64.89 2.93 64.91 3.407 ;
      RECT 64.87 2.99 64.89 3.405 ;
      RECT 64.83 3.025 64.87 3.403 ;
      RECT 64.826 3.035 64.83 3.401 ;
      RECT 64.74 3.05 64.826 3.397 ;
      RECT 64.72 3.07 64.74 3.393 ;
      RECT 64.65 3.075 64.72 3.389 ;
      RECT 64.63 3.076 64.65 3.386 ;
      RECT 64.626 3.078 64.63 3.385 ;
      RECT 64.54 3.087 64.626 3.38 ;
      RECT 64.53 3.096 64.54 3.375 ;
      RECT 64.49 3.102 64.53 3.37 ;
      RECT 64.44 3.113 64.49 3.355 ;
      RECT 64.42 3.122 64.44 3.34 ;
      RECT 64.34 3.135 64.42 3.325 ;
      RECT 64.51 2.685 64.68 2.895 ;
      RECT 64.626 2.677 64.68 2.895 ;
      RECT 64.426 2.685 64.68 2.885 ;
      RECT 64.34 2.685 64.68 2.865 ;
      RECT 64.34 2.69 64.69 2.81 ;
      RECT 64.34 2.7 64.7 2.72 ;
      RECT 64.54 2.682 64.68 2.895 ;
      RECT 64.29 3.623 64.54 3.955 ;
      RECT 64.26 3.635 64.54 3.937 ;
      RECT 64.24 3.67 64.54 3.907 ;
      RECT 64.29 3.62 64.462 3.955 ;
      RECT 64.29 3.616 64.376 3.955 ;
      RECT 64.22 1.965 64.4 2.385 ;
      RECT 64.22 1.965 64.42 2.375 ;
      RECT 64.22 1.965 64.44 2.35 ;
      RECT 64.22 1.965 64.45 2.335 ;
      RECT 64.22 1.965 64.46 2.33 ;
      RECT 64.22 2.005 64.48 2.315 ;
      RECT 64.22 2.075 64.5 2.295 ;
      RECT 64.2 2.075 64.5 2.29 ;
      RECT 64.2 2.135 64.51 2.265 ;
      RECT 64.2 2.175 64.52 2.215 ;
      RECT 64.18 1.965 64.46 2.195 ;
      RECT 64.17 1.975 64.46 2.118 ;
      RECT 64.16 2.015 64.48 2.063 ;
      RECT 63.76 3.375 63.93 3.895 ;
      RECT 63.75 3.375 63.93 3.855 ;
      RECT 63.74 3.395 63.93 3.83 ;
      RECT 63.75 3.375 63.94 3.825 ;
      RECT 63.73 3.435 63.94 3.795 ;
      RECT 63.72 3.47 63.94 3.775 ;
      RECT 63.71 3.52 63.94 3.735 ;
      RECT 63.75 3.386 63.95 3.725 ;
      RECT 63.7 3.6 63.95 3.675 ;
      RECT 63.74 3.409 63.96 3.605 ;
      RECT 63.74 3.433 63.97 3.5 ;
      RECT 63.68 2.68 63.7 2.955 ;
      RECT 63.64 2.665 63.68 3 ;
      RECT 63.62 2.65 63.64 3.065 ;
      RECT 63.6 2.649 63.62 3.14 ;
      RECT 63.58 2.657 63.6 3.245 ;
      RECT 63.576 2.662 63.58 3.297 ;
      RECT 63.49 2.681 63.576 3.337 ;
      RECT 63.48 2.702 63.49 3.376 ;
      RECT 63.47 2.71 63.48 3.377 ;
      RECT 63.45 2.845 63.47 3.379 ;
      RECT 63.44 2.995 63.45 3.381 ;
      RECT 63.4 3.08 63.44 3.386 ;
      RECT 63.318 3.102 63.4 3.396 ;
      RECT 63.232 3.117 63.318 3.409 ;
      RECT 63.146 3.132 63.232 3.422 ;
      RECT 63.06 3.147 63.146 3.436 ;
      RECT 62.98 3.161 63.06 3.449 ;
      RECT 62.966 3.169 62.98 3.457 ;
      RECT 62.88 3.177 62.966 3.471 ;
      RECT 62.87 3.185 62.88 3.484 ;
      RECT 62.846 3.185 62.87 3.492 ;
      RECT 62.76 3.187 62.846 3.522 ;
      RECT 62.68 3.189 62.76 3.565 ;
      RECT 62.61 3.192 62.68 3.6 ;
      RECT 62.59 3.194 62.61 3.616 ;
      RECT 62.56 3.2 62.59 3.618 ;
      RECT 62.51 3.215 62.56 3.621 ;
      RECT 62.49 3.23 62.51 3.624 ;
      RECT 62.46 3.235 62.49 3.627 ;
      RECT 62.4 3.25 62.46 3.631 ;
      RECT 62.39 3.266 62.4 3.635 ;
      RECT 62.34 3.276 62.39 3.624 ;
      RECT 62.31 3.295 62.34 3.607 ;
      RECT 62.29 3.315 62.31 3.597 ;
      RECT 62.27 3.34 62.29 3.589 ;
      RECT 63.28 1.932 63.45 2.425 ;
      RECT 63.27 1.932 63.45 2.41 ;
      RECT 63.27 1.947 63.48 2.4 ;
      RECT 63.26 1.947 63.48 2.375 ;
      RECT 63.25 1.947 63.48 2.34 ;
      RECT 63.25 1.955 63.49 2.295 ;
      RECT 63.23 1.925 63.42 2.275 ;
      RECT 63.22 1.932 63.45 2.235 ;
      RECT 63.21 1.947 63.48 2.215 ;
      RECT 63.2 1.96 63.49 2.175 ;
      RECT 63.19 1.975 63.49 2.128 ;
      RECT 63.19 1.975 63.5 2.12 ;
      RECT 63.18 1.99 63.5 2.093 ;
      RECT 63.19 1.985 63.51 2.035 ;
      RECT 62.99 2.612 63.26 2.905 ;
      RECT 62.99 2.614 63.27 2.9 ;
      RECT 62.98 2.64 63.27 2.895 ;
      RECT 62.99 2.63 63.28 2.89 ;
      RECT 62.99 2.608 63.226 2.905 ;
      RECT 62.99 2.605 63.14 2.905 ;
      RECT 63.05 2.6 63.136 2.905 ;
      RECT 62.54 2.648 62.61 2.945 ;
      RECT 62.54 2.648 62.62 2.944 ;
      RECT 62.62 2.635 62.63 2.941 ;
      RECT 62.52 2.662 62.63 2.935 ;
      RECT 62.61 2.64 62.7 2.931 ;
      RECT 62.54 2.655 62.72 2.92 ;
      RECT 62.52 2.72 62.73 2.916 ;
      RECT 62.5 2.668 62.72 2.915 ;
      RECT 62.49 2.673 62.72 2.905 ;
      RECT 62.48 2.795 62.74 2.9 ;
      RECT 62.48 2.875 62.75 2.89 ;
      RECT 62.45 2.681 62.72 2.884 ;
      RECT 62.44 2.695 62.72 2.869 ;
      RECT 62.48 2.676 62.72 2.9 ;
      RECT 62.61 2.636 62.63 2.941 ;
      RECT 62.43 2.072 62.45 2.305 ;
      RECT 62.42 2.053 62.43 2.31 ;
      RECT 62.41 2.041 62.42 2.317 ;
      RECT 62.37 2.027 62.41 2.327 ;
      RECT 62.36 2.017 62.37 2.336 ;
      RECT 62.31 2.002 62.36 2.341 ;
      RECT 62.3 1.987 62.31 2.347 ;
      RECT 62.28 1.978 62.3 2.352 ;
      RECT 62.27 1.968 62.28 2.358 ;
      RECT 62.26 1.965 62.27 2.363 ;
      RECT 62.24 1.965 62.26 2.364 ;
      RECT 62.21 1.96 62.24 2.362 ;
      RECT 62.186 1.953 62.21 2.361 ;
      RECT 62.1 1.943 62.186 2.358 ;
      RECT 62.09 1.935 62.1 2.355 ;
      RECT 62.068 1.935 62.09 2.354 ;
      RECT 61.982 1.935 62.068 2.352 ;
      RECT 61.896 1.935 61.982 2.35 ;
      RECT 61.81 1.935 61.896 2.347 ;
      RECT 61.8 1.935 61.81 2.34 ;
      RECT 61.77 1.935 61.8 2.3 ;
      RECT 61.76 1.945 61.77 2.255 ;
      RECT 61.75 1.99 61.76 2.24 ;
      RECT 61.72 2.085 61.75 2.195 ;
      RECT 61.91 2.822 62.08 3.335 ;
      RECT 61.9 2.853 62.08 3.315 ;
      RECT 61.9 2.853 62.1 3.285 ;
      RECT 61.89 2.861 62.1 3.26 ;
      RECT 61.89 2.861 62.11 3.25 ;
      RECT 61.89 2.861 62.12 3.23 ;
      RECT 61.89 2.861 62.17 3.185 ;
      RECT 61.89 2.861 62.18 3.16 ;
      RECT 61.89 2.861 62.19 3.125 ;
      RECT 61.89 2.861 62.2 3.09 ;
      RECT 61.89 2.861 62.21 3.04 ;
      RECT 61.89 2.861 62.23 2.965 ;
      RECT 62.06 2.725 62.24 2.905 ;
      RECT 61.98 2.78 62.24 2.905 ;
      RECT 62.02 2.745 62.08 3.335 ;
      RECT 62.01 2.765 62.24 2.905 ;
      RECT 61.37 3.235 61.456 3.801 ;
      RECT 61.33 3.235 61.456 3.795 ;
      RECT 61.33 3.235 61.542 3.793 ;
      RECT 61.33 3.235 61.58 3.787 ;
      RECT 61.33 3.242 61.59 3.785 ;
      RECT 61.3 3.235 61.58 3.78 ;
      RECT 61.27 3.25 61.59 3.77 ;
      RECT 61.27 3.277 61.63 3.762 ;
      RECT 61.245 3.277 61.63 3.75 ;
      RECT 61.245 3.315 61.64 3.732 ;
      RECT 61.23 3.297 61.63 3.725 ;
      RECT 61.23 3.345 61.65 3.721 ;
      RECT 61.23 3.411 61.67 3.705 ;
      RECT 61.23 3.466 61.68 3.515 ;
      RECT 61.42 2.755 61.59 2.935 ;
      RECT 61.37 2.694 61.42 2.92 ;
      RECT 61.11 2.675 61.37 2.905 ;
      RECT 61.07 2.735 61.54 2.905 ;
      RECT 61.07 2.725 61.5 2.905 ;
      RECT 61.07 2.714 61.48 2.905 ;
      RECT 61.07 2.7 61.42 2.905 ;
      RECT 61.11 2.67 61.306 2.905 ;
      RECT 61.14 2.649 61.306 2.905 ;
      RECT 61.12 2.65 61.306 2.905 ;
      RECT 61.14 2.635 61.22 2.905 ;
      RECT 60.9 3.165 61.02 3.605 ;
      RECT 60.88 3.165 61.02 3.604 ;
      RECT 60.84 3.185 61.02 3.601 ;
      RECT 60.8 3.229 61.02 3.597 ;
      RECT 60.79 3.259 61.04 3.46 ;
      RECT 60.88 3.165 61.05 3.355 ;
      RECT 60.54 1.945 60.55 2.395 ;
      RECT 60.35 1.945 60.37 2.355 ;
      RECT 60.32 1.945 60.33 2.335 ;
      RECT 61 2.255 61.02 2.44 ;
      RECT 60.98 2.215 61 2.448 ;
      RECT 60.93 2.182 60.98 2.458 ;
      RECT 60.876 2.156 60.93 2.461 ;
      RECT 60.79 2.121 60.876 2.451 ;
      RECT 60.78 2.097 60.79 2.44 ;
      RECT 60.71 2.063 60.78 2.43 ;
      RECT 60.69 2.023 60.71 2.423 ;
      RECT 60.67 2.005 60.69 2.419 ;
      RECT 60.66 1.995 60.67 2.416 ;
      RECT 60.63 1.98 60.66 2.412 ;
      RECT 60.62 1.965 60.63 2.408 ;
      RECT 60.61 1.96 60.62 2.406 ;
      RECT 60.56 1.95 60.61 2.401 ;
      RECT 60.55 1.945 60.56 2.396 ;
      RECT 60.52 1.945 60.54 2.39 ;
      RECT 60.486 1.945 60.52 2.382 ;
      RECT 60.4 1.945 60.486 2.372 ;
      RECT 60.37 1.945 60.4 2.36 ;
      RECT 60.33 1.945 60.35 2.345 ;
      RECT 60.31 1.945 60.32 2.328 ;
      RECT 60.29 1.955 60.31 2.308 ;
      RECT 60.28 1.975 60.29 2.24 ;
      RECT 60.27 1.985 60.28 2 ;
      RECT 60.54 2.665 60.626 2.99 ;
      RECT 60.54 2.665 60.66 2.982 ;
      RECT 60.49 2.665 60.66 2.98 ;
      RECT 60.49 2.669 60.746 2.975 ;
      RECT 60.49 2.674 60.77 2.968 ;
      RECT 60.49 2.68 60.78 2.966 ;
      RECT 60.49 2.69 60.79 2.963 ;
      RECT 60.49 2.83 60.8 2.958 ;
      RECT 60.55 3.34 60.6 3.656 ;
      RECT 60.54 3.32 60.55 3.681 ;
      RECT 60.53 3.31 60.54 3.69 ;
      RECT 60.51 3.304 60.53 3.705 ;
      RECT 60.48 3.302 60.51 3.725 ;
      RECT 60.466 3.3 60.48 3.735 ;
      RECT 60.38 3.296 60.466 3.735 ;
      RECT 60.31 3.29 60.38 3.725 ;
      RECT 60.23 3.285 60.31 3.7 ;
      RECT 60.17 3.281 60.23 3.665 ;
      RECT 60.1 3.277 60.17 3.625 ;
      RECT 60.07 3.275 60.1 3.6 ;
      RECT 59.966 3.273 60.01 3.595 ;
      RECT 59.88 3.268 59.966 3.595 ;
      RECT 59.8 3.265 59.88 3.595 ;
      RECT 59.72 3.266 59.8 3.62 ;
      RECT 59.638 3.268 59.72 3.645 ;
      RECT 59.552 3.269 59.638 3.645 ;
      RECT 59.466 3.271 59.552 3.645 ;
      RECT 59.38 3.273 59.466 3.645 ;
      RECT 59.36 3.274 59.38 3.637 ;
      RECT 59.35 3.28 59.36 3.626 ;
      RECT 59.31 3.3 59.35 3.607 ;
      RECT 59.3 3.32 59.31 3.589 ;
      RECT 60.01 3.275 60.07 3.595 ;
      RECT 59.98 2.82 60.15 3.075 ;
      RECT 59.98 2.82 60.16 3.068 ;
      RECT 59.98 2.82 60.17 3.053 ;
      RECT 59.98 2.82 60.19 3.035 ;
      RECT 59.98 2.82 60.23 2.99 ;
      RECT 60.16 2.585 60.25 2.943 ;
      RECT 60.15 2.59 60.26 2.924 ;
      RECT 60.1 2.605 60.27 2.911 ;
      RECT 60.09 2.62 60.28 2.895 ;
      RECT 59.99 2.785 60.28 2.895 ;
      RECT 60.03 2.645 60.15 3.075 ;
      RECT 60 2.755 60.28 2.895 ;
      RECT 60.02 2.68 60.15 3.075 ;
      RECT 60.01 2.705 60.28 2.895 ;
      RECT 60.13 2.591 60.26 2.924 ;
      RECT 60.15 2.586 60.25 2.943 ;
      RECT 59.61 2.72 59.8 2.895 ;
      RECT 59.57 2.638 59.76 2.89 ;
      RECT 59.536 2.643 59.76 2.884 ;
      RECT 59.45 2.65 59.76 2.879 ;
      RECT 59.366 2.665 59.76 2.874 ;
      RECT 59.28 2.685 59.79 2.868 ;
      RECT 59.366 2.675 59.79 2.874 ;
      RECT 59.61 2.635 59.76 2.895 ;
      RECT 59.61 2.631 59.71 2.895 ;
      RECT 59.696 2.626 59.71 2.895 ;
      RECT 58.45 1.954 59.11 2.345 ;
      RECT 58.708 1.948 59.11 2.345 ;
      RECT 58.44 1.96 59.11 2.344 ;
      RECT 58.43 1.975 59.11 2.343 ;
      RECT 58.37 2.015 59.11 2.339 ;
      RECT 58.536 1.953 59.12 2.335 ;
      RECT 58.44 1.96 59.13 2.325 ;
      RECT 58.44 1.968 59.14 2.305 ;
      RECT 58.43 1.978 59.16 2.278 ;
      RECT 58.37 2.015 59.17 2.253 ;
      RECT 58.43 1.985 59.18 2.24 ;
      RECT 58.536 1.951 59.11 2.345 ;
      RECT 58.622 1.949 59.11 2.345 ;
      RECT 58.708 1.947 59.09 2.345 ;
      RECT 58.794 1.945 59.09 2.345 ;
      RECT 58.96 3.12 59.13 3.315 ;
      RECT 58.95 3.12 59.13 3.26 ;
      RECT 58.945 3.12 59.13 3.188 ;
      RECT 58.93 3.06 59.11 3.155 ;
      RECT 58.92 3.06 59.11 3.105 ;
      RECT 58.89 3.035 59.1 3.06 ;
      RECT 58.87 3.035 59.1 3.045 ;
      RECT 58.81 2.725 58.99 3.036 ;
      RECT 58.81 2.96 59.09 3.036 ;
      RECT 58.8 2.724 58.81 3.026 ;
      RECT 58.78 2.723 58.8 3.02 ;
      RECT 58.75 2.722 58.78 3 ;
      RECT 58.7 2.719 58.75 2.965 ;
      RECT 58.7 2.84 59.06 2.965 ;
      RECT 58.63 2.716 58.7 2.92 ;
      RECT 58.63 2.775 59.04 2.92 ;
      RECT 58.63 2.765 59.03 2.92 ;
      RECT 58.63 2.755 59.02 2.92 ;
      RECT 58.63 2.735 59 2.92 ;
      RECT 58.71 3.255 58.72 3.512 ;
      RECT 58.69 3.172 58.71 3.532 ;
      RECT 58.67 3.166 58.69 3.56 ;
      RECT 58.61 3.154 58.67 3.58 ;
      RECT 58.57 3.14 58.61 3.581 ;
      RECT 58.486 3.129 58.57 3.569 ;
      RECT 58.4 3.116 58.486 3.553 ;
      RECT 58.39 3.109 58.4 3.545 ;
      RECT 58.34 3.106 58.39 3.485 ;
      RECT 58.32 3.102 58.34 3.4 ;
      RECT 58.31 3.1 58.32 3.35 ;
      RECT 58.28 3.098 58.31 3.32 ;
      RECT 58.24 3.093 58.28 3.3 ;
      RECT 58.202 3.088 58.24 3.288 ;
      RECT 58.116 3.08 58.202 3.297 ;
      RECT 58.03 3.069 58.116 3.309 ;
      RECT 57.96 3.059 58.03 3.319 ;
      RECT 57.94 3.05 57.96 3.324 ;
      RECT 57.88 3.022 57.94 3.32 ;
      RECT 57.86 2.992 57.88 3.308 ;
      RECT 57.84 2.965 57.86 3.295 ;
      RECT 57.76 2.718 57.84 3.262 ;
      RECT 57.746 2.71 57.76 3.224 ;
      RECT 57.66 2.702 57.746 3.145 ;
      RECT 57.64 2.693 57.66 3.061 ;
      RECT 57.61 2.688 57.64 3.041 ;
      RECT 57.54 2.699 57.61 3.026 ;
      RECT 57.52 2.717 57.54 3 ;
      RECT 57.51 2.723 57.52 2.945 ;
      RECT 57.49 2.745 57.51 2.83 ;
      RECT 58.15 2.705 58.32 2.895 ;
      RECT 58.15 2.705 58.35 2.89 ;
      RECT 58.2 2.615 58.37 2.88 ;
      RECT 58.16 2.65 58.37 2.88 ;
      RECT 57.36 3.388 57.43 3.829 ;
      RECT 57.3 3.413 57.43 3.826 ;
      RECT 57.3 3.413 57.48 3.819 ;
      RECT 57.29 3.435 57.48 3.816 ;
      RECT 57.43 3.375 57.5 3.814 ;
      RECT 57.36 3.4 57.58 3.811 ;
      RECT 57.29 3.439 57.63 3.807 ;
      RECT 57.27 3.465 57.63 3.795 ;
      RECT 57.29 3.459 57.65 3.79 ;
      RECT 57.27 2.205 57.31 2.445 ;
      RECT 57.27 2.205 57.34 2.444 ;
      RECT 57.27 2.205 57.45 2.436 ;
      RECT 57.27 2.205 57.51 2.415 ;
      RECT 57.28 2.15 57.56 2.315 ;
      RECT 57.39 1.99 57.42 2.437 ;
      RECT 57.42 1.985 57.6 2.195 ;
      RECT 57.29 2.125 57.6 2.195 ;
      RECT 57.34 2.02 57.39 2.44 ;
      RECT 57.31 2.075 57.6 2.195 ;
      RECT 56.18 5.02 56.35 6.49 ;
      RECT 56.18 6.315 56.355 6.485 ;
      RECT 55.81 1.74 55.98 2.93 ;
      RECT 55.81 1.74 56.28 1.91 ;
      RECT 55.81 6.97 56.28 7.14 ;
      RECT 55.81 5.95 55.98 7.14 ;
      RECT 54.82 1.74 54.99 2.93 ;
      RECT 54.82 1.74 55.29 1.91 ;
      RECT 54.82 6.97 55.29 7.14 ;
      RECT 54.82 5.95 54.99 7.14 ;
      RECT 52.97 2.635 53.14 3.865 ;
      RECT 53.025 0.855 53.195 2.805 ;
      RECT 52.97 0.575 53.14 1.025 ;
      RECT 52.97 7.855 53.14 8.305 ;
      RECT 53.025 6.075 53.195 8.025 ;
      RECT 52.97 5.015 53.14 6.245 ;
      RECT 52.45 0.575 52.62 3.865 ;
      RECT 52.45 2.075 52.855 2.405 ;
      RECT 52.45 1.235 52.855 1.565 ;
      RECT 52.45 5.015 52.62 8.305 ;
      RECT 52.45 7.315 52.855 7.645 ;
      RECT 52.45 6.475 52.855 6.805 ;
      RECT 50.545 3.39 50.565 3.44 ;
      RECT 50.525 3.362 50.545 3.555 ;
      RECT 50.505 3.337 50.525 3.611 ;
      RECT 50.465 3.325 50.505 3.63 ;
      RECT 50.415 3.32 50.465 3.659 ;
      RECT 50.411 3.314 50.415 3.675 ;
      RECT 50.325 3.306 50.411 3.675 ;
      RECT 50.265 3.294 50.325 3.67 ;
      RECT 50.211 3.284 50.265 3.659 ;
      RECT 50.125 3.272 50.211 3.642 ;
      RECT 50.103 3.263 50.125 3.629 ;
      RECT 50.017 3.256 50.103 3.616 ;
      RECT 49.931 3.243 50.017 3.595 ;
      RECT 49.845 3.231 49.931 3.575 ;
      RECT 49.815 3.22 49.845 3.561 ;
      RECT 49.765 3.207 49.815 3.551 ;
      RECT 49.745 3.197 49.765 3.545 ;
      RECT 49.691 3.187 49.745 3.539 ;
      RECT 49.605 3.167 49.691 3.523 ;
      RECT 49.565 3.155 49.605 3.509 ;
      RECT 49.53 3.155 49.565 3.495 ;
      RECT 49.515 3.155 49.53 3.48 ;
      RECT 49.465 3.155 49.515 3.425 ;
      RECT 49.435 3.155 49.465 3.345 ;
      RECT 49.965 2.825 50.135 3.075 ;
      RECT 49.965 2.825 50.145 3.03 ;
      RECT 50.025 2.655 50.155 2.975 ;
      RECT 50.025 2.662 50.165 2.94 ;
      RECT 49.985 2.677 50.175 2.875 ;
      RECT 49.975 2.76 50.175 2.875 ;
      RECT 49.985 2.695 50.185 2.785 ;
      RECT 49.985 2.675 50.165 2.94 ;
      RECT 49.755 1.93 49.925 2.415 ;
      RECT 49.745 1.93 49.925 2.405 ;
      RECT 49.745 1.945 49.945 2.35 ;
      RECT 49.705 1.925 49.895 2.315 ;
      RECT 49.705 1.96 49.955 2.235 ;
      RECT 49.655 1.945 49.945 2.135 ;
      RECT 49.655 1.975 49.965 2.095 ;
      RECT 49.655 1.99 49.975 2.015 ;
      RECT 49.251 2.688 49.265 2.944 ;
      RECT 49.251 2.689 49.351 2.939 ;
      RECT 49.165 2.686 49.251 2.936 ;
      RECT 49.155 2.685 49.165 2.929 ;
      RECT 49.155 2.692 49.437 2.926 ;
      RECT 49.075 2.695 49.437 2.922 ;
      RECT 49.155 2.694 49.455 2.919 ;
      RECT 49.065 2.707 49.475 2.916 ;
      RECT 49.075 2.695 49.475 2.916 ;
      RECT 49.055 2.712 49.475 2.915 ;
      RECT 49.075 2.697 49.561 2.911 ;
      RECT 49.035 2.715 49.561 2.908 ;
      RECT 49.075 2.701 49.647 2.902 ;
      RECT 49.025 2.72 49.647 2.898 ;
      RECT 49.075 2.704 49.675 2.897 ;
      RECT 49.075 2.705 49.715 2.891 ;
      RECT 49.065 2.71 49.725 2.886 ;
      RECT 49.025 2.73 49.735 2.875 ;
      RECT 49.025 2.75 49.745 2.86 ;
      RECT 48.985 3.298 49.005 3.605 ;
      RECT 48.975 3.273 48.985 3.885 ;
      RECT 48.935 3.24 48.975 3.885 ;
      RECT 48.931 3.21 48.935 3.885 ;
      RECT 48.845 3.095 48.931 3.885 ;
      RECT 48.835 2.97 48.845 3.885 ;
      RECT 48.825 2.935 48.835 3.885 ;
      RECT 48.815 2.905 48.825 3.885 ;
      RECT 48.795 2.875 48.815 3.77 ;
      RECT 48.785 2.845 48.795 3.645 ;
      RECT 48.775 2.825 48.785 3.595 ;
      RECT 48.755 2.795 48.775 3.503 ;
      RECT 48.735 2.761 48.755 3.418 ;
      RECT 48.73 2.744 48.735 3.353 ;
      RECT 48.725 2.738 48.73 3.325 ;
      RECT 48.715 2.73 48.725 3.29 ;
      RECT 48.695 2.725 48.705 3.19 ;
      RECT 48.685 2.725 48.695 3.165 ;
      RECT 48.68 2.725 48.685 3.128 ;
      RECT 48.665 2.725 48.68 3.06 ;
      RECT 48.655 2.724 48.665 2.99 ;
      RECT 48.645 2.722 48.655 2.97 ;
      RECT 48.585 2.718 48.645 2.943 ;
      RECT 48.545 2.72 48.585 2.923 ;
      RECT 48.525 2.75 48.545 2.905 ;
      RECT 48.705 2.725 48.715 3.245 ;
      RECT 48.645 2.08 48.815 2.435 ;
      RECT 48.675 1.966 48.815 2.435 ;
      RECT 48.675 1.968 48.825 2.43 ;
      RECT 48.675 1.97 48.845 2.42 ;
      RECT 48.675 1.973 48.875 2.405 ;
      RECT 48.675 1.978 48.925 2.375 ;
      RECT 48.675 1.983 48.945 2.338 ;
      RECT 48.655 1.985 48.955 2.313 ;
      RECT 48.675 1.965 48.785 2.435 ;
      RECT 48.685 1.96 48.785 2.435 ;
      RECT 48.205 3.222 48.395 3.585 ;
      RECT 48.205 3.237 48.435 3.583 ;
      RECT 48.205 3.265 48.455 3.579 ;
      RECT 48.205 3.3 48.465 3.577 ;
      RECT 48.205 3.345 48.475 3.576 ;
      RECT 48.195 3.217 48.355 3.565 ;
      RECT 48.175 3.225 48.395 3.515 ;
      RECT 48.145 3.237 48.435 3.45 ;
      RECT 48.205 3.215 48.355 3.585 ;
      RECT 48.21 7.855 48.38 8.305 ;
      RECT 48.265 6.075 48.435 8.025 ;
      RECT 48.21 5.015 48.38 6.245 ;
      RECT 47.69 5.015 47.86 8.305 ;
      RECT 47.69 7.315 48.095 7.645 ;
      RECT 47.69 6.475 48.095 6.805 ;
      RECT 47.791 2.695 47.995 3.105 ;
      RECT 47.705 2.588 47.791 3.09 ;
      RECT 47.701 2.584 47.705 3.074 ;
      RECT 47.615 2.695 47.995 3.054 ;
      RECT 47.595 2.575 47.615 3.015 ;
      RECT 47.585 2.58 47.701 2.99 ;
      RECT 47.575 2.587 47.705 2.97 ;
      RECT 47.565 2.592 47.795 2.945 ;
      RECT 47.555 2.61 47.885 2.925 ;
      RECT 47.545 2.615 47.885 2.905 ;
      RECT 47.535 2.62 47.925 2.77 ;
      RECT 47.535 2.65 47.985 2.77 ;
      RECT 47.535 2.635 47.975 2.77 ;
      RECT 47.565 2.605 47.885 2.945 ;
      RECT 47.565 2.593 47.825 2.945 ;
      RECT 47.715 3.42 47.965 3.885 ;
      RECT 47.635 3.395 47.955 3.88 ;
      RECT 47.565 3.429 47.965 3.87 ;
      RECT 47.355 3.68 47.965 3.865 ;
      RECT 47.535 3.449 47.965 3.865 ;
      RECT 47.375 3.64 47.965 3.865 ;
      RECT 47.525 3.46 47.965 3.865 ;
      RECT 47.415 3.58 47.965 3.865 ;
      RECT 47.465 3.505 47.965 3.865 ;
      RECT 47.715 3.37 47.955 3.885 ;
      RECT 47.735 3.365 47.955 3.885 ;
      RECT 47.745 3.36 47.875 3.885 ;
      RECT 47.831 3.355 47.835 3.885 ;
      RECT 47.305 1.925 47.391 2.362 ;
      RECT 47.295 1.925 47.391 2.358 ;
      RECT 47.295 1.925 47.455 2.357 ;
      RECT 47.295 1.925 47.485 2.355 ;
      RECT 47.295 1.925 47.495 2.345 ;
      RECT 47.285 1.93 47.495 2.343 ;
      RECT 47.275 1.94 47.495 2.335 ;
      RECT 47.275 1.94 47.505 2.295 ;
      RECT 47.295 1.925 47.525 2.21 ;
      RECT 47.265 1.95 47.525 2.205 ;
      RECT 47.275 1.94 47.535 2.135 ;
      RECT 47.255 1.96 47.535 2.08 ;
      RECT 47.245 1.97 47.535 1.98 ;
      RECT 47.325 2.741 47.335 2.82 ;
      RECT 47.315 2.734 47.325 3.005 ;
      RECT 47.305 2.728 47.315 3.03 ;
      RECT 47.295 2.72 47.305 3.06 ;
      RECT 47.255 2.715 47.295 3.11 ;
      RECT 47.235 2.715 47.255 3.165 ;
      RECT 47.225 2.715 47.235 3.19 ;
      RECT 47.215 2.715 47.225 3.205 ;
      RECT 47.185 2.715 47.215 3.25 ;
      RECT 47.175 2.715 47.185 3.29 ;
      RECT 47.155 2.715 47.175 3.315 ;
      RECT 47.135 2.715 47.155 3.35 ;
      RECT 47.055 2.715 47.135 3.395 ;
      RECT 47.045 2.715 47.055 3.415 ;
      RECT 47.005 2.795 47.045 3.412 ;
      RECT 46.985 2.875 47.005 3.409 ;
      RECT 46.965 2.93 46.985 3.407 ;
      RECT 46.945 2.99 46.965 3.405 ;
      RECT 46.905 3.025 46.945 3.403 ;
      RECT 46.901 3.035 46.905 3.401 ;
      RECT 46.815 3.05 46.901 3.397 ;
      RECT 46.795 3.07 46.815 3.393 ;
      RECT 46.725 3.075 46.795 3.389 ;
      RECT 46.705 3.076 46.725 3.386 ;
      RECT 46.701 3.078 46.705 3.385 ;
      RECT 46.615 3.087 46.701 3.38 ;
      RECT 46.605 3.096 46.615 3.375 ;
      RECT 46.565 3.102 46.605 3.37 ;
      RECT 46.515 3.113 46.565 3.355 ;
      RECT 46.495 3.122 46.515 3.34 ;
      RECT 46.415 3.135 46.495 3.325 ;
      RECT 46.585 2.685 46.755 2.895 ;
      RECT 46.701 2.677 46.755 2.895 ;
      RECT 46.501 2.685 46.755 2.885 ;
      RECT 46.415 2.685 46.755 2.865 ;
      RECT 46.415 2.69 46.765 2.81 ;
      RECT 46.415 2.7 46.775 2.72 ;
      RECT 46.615 2.682 46.755 2.895 ;
      RECT 46.365 3.623 46.615 3.955 ;
      RECT 46.335 3.635 46.615 3.937 ;
      RECT 46.315 3.67 46.615 3.907 ;
      RECT 46.365 3.62 46.537 3.955 ;
      RECT 46.365 3.616 46.451 3.955 ;
      RECT 46.295 1.965 46.475 2.385 ;
      RECT 46.295 1.965 46.495 2.375 ;
      RECT 46.295 1.965 46.515 2.35 ;
      RECT 46.295 1.965 46.525 2.335 ;
      RECT 46.295 1.965 46.535 2.33 ;
      RECT 46.295 2.005 46.555 2.315 ;
      RECT 46.295 2.075 46.575 2.295 ;
      RECT 46.275 2.075 46.575 2.29 ;
      RECT 46.275 2.135 46.585 2.265 ;
      RECT 46.275 2.175 46.595 2.215 ;
      RECT 46.255 1.965 46.535 2.195 ;
      RECT 46.245 1.975 46.535 2.118 ;
      RECT 46.235 2.015 46.555 2.063 ;
      RECT 45.835 3.375 46.005 3.895 ;
      RECT 45.825 3.375 46.005 3.855 ;
      RECT 45.815 3.395 46.005 3.83 ;
      RECT 45.825 3.375 46.015 3.825 ;
      RECT 45.805 3.435 46.015 3.795 ;
      RECT 45.795 3.47 46.015 3.775 ;
      RECT 45.785 3.52 46.015 3.735 ;
      RECT 45.825 3.386 46.025 3.725 ;
      RECT 45.775 3.6 46.025 3.675 ;
      RECT 45.815 3.409 46.035 3.605 ;
      RECT 45.815 3.433 46.045 3.5 ;
      RECT 45.755 2.68 45.775 2.955 ;
      RECT 45.715 2.665 45.755 3 ;
      RECT 45.695 2.65 45.715 3.065 ;
      RECT 45.675 2.649 45.695 3.14 ;
      RECT 45.655 2.657 45.675 3.245 ;
      RECT 45.651 2.662 45.655 3.297 ;
      RECT 45.565 2.681 45.651 3.337 ;
      RECT 45.555 2.702 45.565 3.376 ;
      RECT 45.545 2.71 45.555 3.377 ;
      RECT 45.525 2.845 45.545 3.379 ;
      RECT 45.515 2.995 45.525 3.381 ;
      RECT 45.475 3.08 45.515 3.386 ;
      RECT 45.393 3.102 45.475 3.396 ;
      RECT 45.307 3.117 45.393 3.409 ;
      RECT 45.221 3.132 45.307 3.422 ;
      RECT 45.135 3.147 45.221 3.436 ;
      RECT 45.055 3.161 45.135 3.449 ;
      RECT 45.041 3.169 45.055 3.457 ;
      RECT 44.955 3.177 45.041 3.471 ;
      RECT 44.945 3.185 44.955 3.484 ;
      RECT 44.921 3.185 44.945 3.492 ;
      RECT 44.835 3.187 44.921 3.522 ;
      RECT 44.755 3.189 44.835 3.565 ;
      RECT 44.685 3.192 44.755 3.6 ;
      RECT 44.665 3.194 44.685 3.616 ;
      RECT 44.635 3.2 44.665 3.618 ;
      RECT 44.585 3.215 44.635 3.621 ;
      RECT 44.565 3.23 44.585 3.624 ;
      RECT 44.535 3.235 44.565 3.627 ;
      RECT 44.475 3.25 44.535 3.631 ;
      RECT 44.465 3.266 44.475 3.635 ;
      RECT 44.415 3.276 44.465 3.624 ;
      RECT 44.385 3.295 44.415 3.607 ;
      RECT 44.365 3.315 44.385 3.597 ;
      RECT 44.345 3.34 44.365 3.589 ;
      RECT 45.355 1.932 45.525 2.425 ;
      RECT 45.345 1.932 45.525 2.41 ;
      RECT 45.345 1.947 45.555 2.4 ;
      RECT 45.335 1.947 45.555 2.375 ;
      RECT 45.325 1.947 45.555 2.34 ;
      RECT 45.325 1.955 45.565 2.295 ;
      RECT 45.305 1.925 45.495 2.275 ;
      RECT 45.295 1.932 45.525 2.235 ;
      RECT 45.285 1.947 45.555 2.215 ;
      RECT 45.275 1.96 45.565 2.175 ;
      RECT 45.265 1.975 45.565 2.128 ;
      RECT 45.265 1.975 45.575 2.12 ;
      RECT 45.255 1.99 45.575 2.093 ;
      RECT 45.265 1.985 45.585 2.035 ;
      RECT 45.065 2.612 45.335 2.905 ;
      RECT 45.065 2.614 45.345 2.9 ;
      RECT 45.055 2.64 45.345 2.895 ;
      RECT 45.065 2.63 45.355 2.89 ;
      RECT 45.065 2.608 45.301 2.905 ;
      RECT 45.065 2.605 45.215 2.905 ;
      RECT 45.125 2.6 45.211 2.905 ;
      RECT 44.615 2.648 44.685 2.945 ;
      RECT 44.615 2.648 44.695 2.944 ;
      RECT 44.695 2.635 44.705 2.941 ;
      RECT 44.595 2.662 44.705 2.935 ;
      RECT 44.685 2.64 44.775 2.931 ;
      RECT 44.615 2.655 44.795 2.92 ;
      RECT 44.595 2.72 44.805 2.916 ;
      RECT 44.575 2.668 44.795 2.915 ;
      RECT 44.565 2.673 44.795 2.905 ;
      RECT 44.555 2.795 44.815 2.9 ;
      RECT 44.555 2.875 44.825 2.89 ;
      RECT 44.525 2.681 44.795 2.884 ;
      RECT 44.515 2.695 44.795 2.869 ;
      RECT 44.555 2.676 44.795 2.9 ;
      RECT 44.685 2.636 44.705 2.941 ;
      RECT 44.505 2.072 44.525 2.305 ;
      RECT 44.495 2.053 44.505 2.31 ;
      RECT 44.485 2.041 44.495 2.317 ;
      RECT 44.445 2.027 44.485 2.327 ;
      RECT 44.435 2.017 44.445 2.336 ;
      RECT 44.385 2.002 44.435 2.341 ;
      RECT 44.375 1.987 44.385 2.347 ;
      RECT 44.355 1.978 44.375 2.352 ;
      RECT 44.345 1.968 44.355 2.358 ;
      RECT 44.335 1.965 44.345 2.363 ;
      RECT 44.315 1.965 44.335 2.364 ;
      RECT 44.285 1.96 44.315 2.362 ;
      RECT 44.261 1.953 44.285 2.361 ;
      RECT 44.175 1.943 44.261 2.358 ;
      RECT 44.165 1.935 44.175 2.355 ;
      RECT 44.143 1.935 44.165 2.354 ;
      RECT 44.057 1.935 44.143 2.352 ;
      RECT 43.971 1.935 44.057 2.35 ;
      RECT 43.885 1.935 43.971 2.347 ;
      RECT 43.875 1.935 43.885 2.34 ;
      RECT 43.845 1.935 43.875 2.3 ;
      RECT 43.835 1.945 43.845 2.255 ;
      RECT 43.825 1.99 43.835 2.24 ;
      RECT 43.795 2.085 43.825 2.195 ;
      RECT 43.985 2.822 44.155 3.335 ;
      RECT 43.975 2.853 44.155 3.315 ;
      RECT 43.975 2.853 44.175 3.285 ;
      RECT 43.965 2.861 44.175 3.26 ;
      RECT 43.965 2.861 44.185 3.25 ;
      RECT 43.965 2.861 44.195 3.23 ;
      RECT 43.965 2.861 44.245 3.185 ;
      RECT 43.965 2.861 44.255 3.16 ;
      RECT 43.965 2.861 44.265 3.125 ;
      RECT 43.965 2.861 44.275 3.09 ;
      RECT 43.965 2.861 44.285 3.04 ;
      RECT 43.965 2.861 44.305 2.965 ;
      RECT 44.135 2.725 44.315 2.905 ;
      RECT 44.055 2.78 44.315 2.905 ;
      RECT 44.095 2.745 44.155 3.335 ;
      RECT 44.085 2.765 44.315 2.905 ;
      RECT 43.445 3.235 43.531 3.801 ;
      RECT 43.405 3.235 43.531 3.795 ;
      RECT 43.405 3.235 43.617 3.793 ;
      RECT 43.405 3.235 43.655 3.787 ;
      RECT 43.405 3.242 43.665 3.785 ;
      RECT 43.375 3.235 43.655 3.78 ;
      RECT 43.345 3.25 43.665 3.77 ;
      RECT 43.345 3.277 43.705 3.762 ;
      RECT 43.32 3.277 43.705 3.75 ;
      RECT 43.32 3.315 43.715 3.732 ;
      RECT 43.305 3.297 43.705 3.725 ;
      RECT 43.305 3.345 43.725 3.721 ;
      RECT 43.305 3.411 43.745 3.705 ;
      RECT 43.305 3.466 43.755 3.515 ;
      RECT 43.495 2.755 43.665 2.935 ;
      RECT 43.445 2.694 43.495 2.92 ;
      RECT 43.185 2.675 43.445 2.905 ;
      RECT 43.145 2.735 43.615 2.905 ;
      RECT 43.145 2.725 43.575 2.905 ;
      RECT 43.145 2.714 43.555 2.905 ;
      RECT 43.145 2.7 43.495 2.905 ;
      RECT 43.185 2.67 43.381 2.905 ;
      RECT 43.215 2.649 43.381 2.905 ;
      RECT 43.195 2.65 43.381 2.905 ;
      RECT 43.215 2.635 43.295 2.905 ;
      RECT 42.975 3.165 43.095 3.605 ;
      RECT 42.955 3.165 43.095 3.604 ;
      RECT 42.915 3.185 43.095 3.601 ;
      RECT 42.875 3.229 43.095 3.597 ;
      RECT 42.865 3.259 43.115 3.46 ;
      RECT 42.955 3.165 43.125 3.355 ;
      RECT 42.615 1.945 42.625 2.395 ;
      RECT 42.425 1.945 42.445 2.355 ;
      RECT 42.395 1.945 42.405 2.335 ;
      RECT 43.075 2.255 43.095 2.44 ;
      RECT 43.055 2.215 43.075 2.448 ;
      RECT 43.005 2.182 43.055 2.458 ;
      RECT 42.951 2.156 43.005 2.461 ;
      RECT 42.865 2.121 42.951 2.451 ;
      RECT 42.855 2.097 42.865 2.44 ;
      RECT 42.785 2.063 42.855 2.43 ;
      RECT 42.765 2.023 42.785 2.423 ;
      RECT 42.745 2.005 42.765 2.419 ;
      RECT 42.735 1.995 42.745 2.416 ;
      RECT 42.705 1.98 42.735 2.412 ;
      RECT 42.695 1.965 42.705 2.408 ;
      RECT 42.685 1.96 42.695 2.406 ;
      RECT 42.635 1.95 42.685 2.401 ;
      RECT 42.625 1.945 42.635 2.396 ;
      RECT 42.595 1.945 42.615 2.39 ;
      RECT 42.561 1.945 42.595 2.382 ;
      RECT 42.475 1.945 42.561 2.372 ;
      RECT 42.445 1.945 42.475 2.36 ;
      RECT 42.405 1.945 42.425 2.345 ;
      RECT 42.385 1.945 42.395 2.328 ;
      RECT 42.365 1.955 42.385 2.308 ;
      RECT 42.355 1.975 42.365 2.24 ;
      RECT 42.345 1.985 42.355 2 ;
      RECT 42.615 2.665 42.701 2.99 ;
      RECT 42.615 2.665 42.735 2.982 ;
      RECT 42.565 2.665 42.735 2.98 ;
      RECT 42.565 2.669 42.821 2.975 ;
      RECT 42.565 2.674 42.845 2.968 ;
      RECT 42.565 2.68 42.855 2.966 ;
      RECT 42.565 2.69 42.865 2.963 ;
      RECT 42.565 2.83 42.875 2.958 ;
      RECT 42.625 3.34 42.675 3.656 ;
      RECT 42.615 3.32 42.625 3.681 ;
      RECT 42.605 3.31 42.615 3.69 ;
      RECT 42.585 3.304 42.605 3.705 ;
      RECT 42.555 3.302 42.585 3.725 ;
      RECT 42.541 3.3 42.555 3.735 ;
      RECT 42.455 3.296 42.541 3.735 ;
      RECT 42.385 3.29 42.455 3.725 ;
      RECT 42.305 3.285 42.385 3.7 ;
      RECT 42.245 3.281 42.305 3.665 ;
      RECT 42.175 3.277 42.245 3.625 ;
      RECT 42.145 3.275 42.175 3.6 ;
      RECT 42.041 3.273 42.085 3.595 ;
      RECT 41.955 3.268 42.041 3.595 ;
      RECT 41.875 3.265 41.955 3.595 ;
      RECT 41.795 3.266 41.875 3.62 ;
      RECT 41.713 3.268 41.795 3.645 ;
      RECT 41.627 3.269 41.713 3.645 ;
      RECT 41.541 3.271 41.627 3.645 ;
      RECT 41.455 3.273 41.541 3.645 ;
      RECT 41.435 3.274 41.455 3.637 ;
      RECT 41.425 3.28 41.435 3.626 ;
      RECT 41.385 3.3 41.425 3.607 ;
      RECT 41.375 3.32 41.385 3.589 ;
      RECT 42.085 3.275 42.145 3.595 ;
      RECT 42.055 2.82 42.225 3.075 ;
      RECT 42.055 2.82 42.235 3.068 ;
      RECT 42.055 2.82 42.245 3.053 ;
      RECT 42.055 2.82 42.265 3.035 ;
      RECT 42.055 2.82 42.305 2.99 ;
      RECT 42.235 2.585 42.325 2.943 ;
      RECT 42.225 2.59 42.335 2.924 ;
      RECT 42.175 2.605 42.345 2.911 ;
      RECT 42.165 2.62 42.355 2.895 ;
      RECT 42.065 2.785 42.355 2.895 ;
      RECT 42.105 2.645 42.225 3.075 ;
      RECT 42.075 2.755 42.355 2.895 ;
      RECT 42.095 2.68 42.225 3.075 ;
      RECT 42.085 2.705 42.355 2.895 ;
      RECT 42.205 2.591 42.335 2.924 ;
      RECT 42.225 2.586 42.325 2.943 ;
      RECT 41.685 2.72 41.875 2.895 ;
      RECT 41.645 2.638 41.835 2.89 ;
      RECT 41.611 2.643 41.835 2.884 ;
      RECT 41.525 2.65 41.835 2.879 ;
      RECT 41.441 2.665 41.835 2.874 ;
      RECT 41.355 2.685 41.865 2.868 ;
      RECT 41.441 2.675 41.865 2.874 ;
      RECT 41.685 2.635 41.835 2.895 ;
      RECT 41.685 2.631 41.785 2.895 ;
      RECT 41.771 2.626 41.785 2.895 ;
      RECT 40.525 1.954 41.185 2.345 ;
      RECT 40.783 1.948 41.185 2.345 ;
      RECT 40.515 1.96 41.185 2.344 ;
      RECT 40.505 1.975 41.185 2.343 ;
      RECT 40.445 2.015 41.185 2.339 ;
      RECT 40.611 1.953 41.195 2.335 ;
      RECT 40.515 1.96 41.205 2.325 ;
      RECT 40.515 1.968 41.215 2.305 ;
      RECT 40.505 1.978 41.235 2.278 ;
      RECT 40.445 2.015 41.245 2.253 ;
      RECT 40.505 1.985 41.255 2.24 ;
      RECT 40.611 1.951 41.185 2.345 ;
      RECT 40.697 1.949 41.185 2.345 ;
      RECT 40.783 1.947 41.165 2.345 ;
      RECT 40.869 1.945 41.165 2.345 ;
      RECT 41.035 3.12 41.205 3.315 ;
      RECT 41.025 3.12 41.205 3.26 ;
      RECT 41.02 3.12 41.205 3.188 ;
      RECT 41.005 3.06 41.185 3.155 ;
      RECT 40.995 3.06 41.185 3.105 ;
      RECT 40.965 3.035 41.175 3.06 ;
      RECT 40.945 3.035 41.175 3.045 ;
      RECT 40.885 2.725 41.065 3.036 ;
      RECT 40.885 2.96 41.165 3.036 ;
      RECT 40.875 2.724 40.885 3.026 ;
      RECT 40.855 2.723 40.875 3.02 ;
      RECT 40.825 2.722 40.855 3 ;
      RECT 40.775 2.719 40.825 2.965 ;
      RECT 40.775 2.84 41.135 2.965 ;
      RECT 40.705 2.716 40.775 2.92 ;
      RECT 40.705 2.775 41.115 2.92 ;
      RECT 40.705 2.765 41.105 2.92 ;
      RECT 40.705 2.755 41.095 2.92 ;
      RECT 40.705 2.735 41.075 2.92 ;
      RECT 40.785 3.255 40.795 3.512 ;
      RECT 40.765 3.172 40.785 3.532 ;
      RECT 40.745 3.166 40.765 3.56 ;
      RECT 40.685 3.154 40.745 3.58 ;
      RECT 40.645 3.14 40.685 3.581 ;
      RECT 40.561 3.129 40.645 3.569 ;
      RECT 40.475 3.116 40.561 3.553 ;
      RECT 40.465 3.109 40.475 3.545 ;
      RECT 40.415 3.106 40.465 3.485 ;
      RECT 40.395 3.102 40.415 3.4 ;
      RECT 40.385 3.1 40.395 3.35 ;
      RECT 40.355 3.098 40.385 3.32 ;
      RECT 40.315 3.093 40.355 3.3 ;
      RECT 40.277 3.088 40.315 3.288 ;
      RECT 40.191 3.08 40.277 3.297 ;
      RECT 40.105 3.069 40.191 3.309 ;
      RECT 40.035 3.059 40.105 3.319 ;
      RECT 40.015 3.05 40.035 3.324 ;
      RECT 39.955 3.022 40.015 3.32 ;
      RECT 39.935 2.992 39.955 3.308 ;
      RECT 39.915 2.965 39.935 3.295 ;
      RECT 39.835 2.718 39.915 3.262 ;
      RECT 39.821 2.71 39.835 3.224 ;
      RECT 39.735 2.702 39.821 3.145 ;
      RECT 39.715 2.693 39.735 3.061 ;
      RECT 39.685 2.688 39.715 3.041 ;
      RECT 39.615 2.699 39.685 3.026 ;
      RECT 39.595 2.717 39.615 3 ;
      RECT 39.585 2.723 39.595 2.945 ;
      RECT 39.565 2.745 39.585 2.83 ;
      RECT 40.225 2.705 40.395 2.895 ;
      RECT 40.225 2.705 40.425 2.89 ;
      RECT 40.275 2.615 40.445 2.88 ;
      RECT 40.235 2.65 40.445 2.88 ;
      RECT 39.435 3.388 39.505 3.829 ;
      RECT 39.375 3.413 39.505 3.826 ;
      RECT 39.375 3.413 39.555 3.819 ;
      RECT 39.365 3.435 39.555 3.816 ;
      RECT 39.505 3.375 39.575 3.814 ;
      RECT 39.435 3.4 39.655 3.811 ;
      RECT 39.365 3.439 39.705 3.807 ;
      RECT 39.345 3.465 39.705 3.795 ;
      RECT 39.365 3.459 39.725 3.79 ;
      RECT 39.345 2.205 39.385 2.445 ;
      RECT 39.345 2.205 39.415 2.444 ;
      RECT 39.345 2.205 39.525 2.436 ;
      RECT 39.345 2.205 39.585 2.415 ;
      RECT 39.355 2.15 39.635 2.315 ;
      RECT 39.465 1.99 39.495 2.437 ;
      RECT 39.495 1.985 39.675 2.195 ;
      RECT 39.365 2.125 39.675 2.195 ;
      RECT 39.415 2.02 39.465 2.44 ;
      RECT 39.385 2.075 39.675 2.195 ;
      RECT 38.255 5.02 38.425 6.49 ;
      RECT 38.255 6.315 38.43 6.485 ;
      RECT 37.885 1.74 38.055 2.93 ;
      RECT 37.885 1.74 38.355 1.91 ;
      RECT 37.885 6.97 38.355 7.14 ;
      RECT 37.885 5.95 38.055 7.14 ;
      RECT 36.895 1.74 37.065 2.93 ;
      RECT 36.895 1.74 37.365 1.91 ;
      RECT 36.895 6.97 37.365 7.14 ;
      RECT 36.895 5.95 37.065 7.14 ;
      RECT 35.045 2.635 35.215 3.865 ;
      RECT 35.1 0.855 35.27 2.805 ;
      RECT 35.045 0.575 35.215 1.025 ;
      RECT 35.045 7.855 35.215 8.305 ;
      RECT 35.1 6.075 35.27 8.025 ;
      RECT 35.045 5.015 35.215 6.245 ;
      RECT 34.525 0.575 34.695 3.865 ;
      RECT 34.525 2.075 34.93 2.405 ;
      RECT 34.525 1.235 34.93 1.565 ;
      RECT 34.525 5.015 34.695 8.305 ;
      RECT 34.525 7.315 34.93 7.645 ;
      RECT 34.525 6.475 34.93 6.805 ;
      RECT 32.62 3.39 32.64 3.44 ;
      RECT 32.6 3.362 32.62 3.555 ;
      RECT 32.58 3.337 32.6 3.611 ;
      RECT 32.54 3.325 32.58 3.63 ;
      RECT 32.49 3.32 32.54 3.659 ;
      RECT 32.486 3.314 32.49 3.675 ;
      RECT 32.4 3.306 32.486 3.675 ;
      RECT 32.34 3.294 32.4 3.67 ;
      RECT 32.286 3.284 32.34 3.659 ;
      RECT 32.2 3.272 32.286 3.642 ;
      RECT 32.178 3.263 32.2 3.629 ;
      RECT 32.092 3.256 32.178 3.616 ;
      RECT 32.006 3.243 32.092 3.595 ;
      RECT 31.92 3.231 32.006 3.575 ;
      RECT 31.89 3.22 31.92 3.561 ;
      RECT 31.84 3.207 31.89 3.551 ;
      RECT 31.82 3.197 31.84 3.545 ;
      RECT 31.766 3.187 31.82 3.539 ;
      RECT 31.68 3.167 31.766 3.523 ;
      RECT 31.64 3.155 31.68 3.509 ;
      RECT 31.605 3.155 31.64 3.495 ;
      RECT 31.59 3.155 31.605 3.48 ;
      RECT 31.54 3.155 31.59 3.425 ;
      RECT 31.51 3.155 31.54 3.345 ;
      RECT 32.04 2.825 32.21 3.075 ;
      RECT 32.04 2.825 32.22 3.03 ;
      RECT 32.1 2.655 32.23 2.975 ;
      RECT 32.1 2.662 32.24 2.94 ;
      RECT 32.06 2.677 32.25 2.875 ;
      RECT 32.05 2.76 32.25 2.875 ;
      RECT 32.06 2.695 32.26 2.785 ;
      RECT 32.06 2.675 32.24 2.94 ;
      RECT 31.83 1.93 32 2.415 ;
      RECT 31.82 1.93 32 2.405 ;
      RECT 31.82 1.945 32.02 2.35 ;
      RECT 31.78 1.925 31.97 2.315 ;
      RECT 31.78 1.96 32.03 2.235 ;
      RECT 31.73 1.945 32.02 2.135 ;
      RECT 31.73 1.975 32.04 2.095 ;
      RECT 31.73 1.99 32.05 2.015 ;
      RECT 31.326 2.688 31.34 2.944 ;
      RECT 31.326 2.689 31.426 2.939 ;
      RECT 31.24 2.686 31.326 2.936 ;
      RECT 31.23 2.685 31.24 2.929 ;
      RECT 31.23 2.692 31.512 2.926 ;
      RECT 31.15 2.695 31.512 2.922 ;
      RECT 31.23 2.694 31.53 2.919 ;
      RECT 31.14 2.707 31.55 2.916 ;
      RECT 31.15 2.695 31.55 2.916 ;
      RECT 31.13 2.712 31.55 2.915 ;
      RECT 31.15 2.697 31.636 2.911 ;
      RECT 31.11 2.715 31.636 2.908 ;
      RECT 31.15 2.701 31.722 2.902 ;
      RECT 31.1 2.72 31.722 2.898 ;
      RECT 31.15 2.704 31.75 2.897 ;
      RECT 31.15 2.705 31.79 2.891 ;
      RECT 31.14 2.71 31.8 2.886 ;
      RECT 31.1 2.73 31.81 2.875 ;
      RECT 31.1 2.75 31.82 2.86 ;
      RECT 31.06 3.298 31.08 3.605 ;
      RECT 31.05 3.273 31.06 3.885 ;
      RECT 31.01 3.24 31.05 3.885 ;
      RECT 31.006 3.21 31.01 3.885 ;
      RECT 30.92 3.095 31.006 3.885 ;
      RECT 30.91 2.97 30.92 3.885 ;
      RECT 30.9 2.935 30.91 3.885 ;
      RECT 30.89 2.905 30.9 3.885 ;
      RECT 30.87 2.875 30.89 3.77 ;
      RECT 30.86 2.845 30.87 3.645 ;
      RECT 30.85 2.825 30.86 3.595 ;
      RECT 30.83 2.795 30.85 3.503 ;
      RECT 30.81 2.761 30.83 3.418 ;
      RECT 30.805 2.744 30.81 3.353 ;
      RECT 30.8 2.738 30.805 3.325 ;
      RECT 30.79 2.73 30.8 3.29 ;
      RECT 30.77 2.725 30.78 3.19 ;
      RECT 30.76 2.725 30.77 3.165 ;
      RECT 30.755 2.725 30.76 3.128 ;
      RECT 30.74 2.725 30.755 3.06 ;
      RECT 30.73 2.724 30.74 2.99 ;
      RECT 30.72 2.722 30.73 2.97 ;
      RECT 30.66 2.718 30.72 2.943 ;
      RECT 30.62 2.72 30.66 2.923 ;
      RECT 30.6 2.75 30.62 2.905 ;
      RECT 30.78 2.725 30.79 3.245 ;
      RECT 30.72 2.08 30.89 2.435 ;
      RECT 30.75 1.966 30.89 2.435 ;
      RECT 30.75 1.968 30.9 2.43 ;
      RECT 30.75 1.97 30.92 2.42 ;
      RECT 30.75 1.973 30.95 2.405 ;
      RECT 30.75 1.978 31 2.375 ;
      RECT 30.75 1.983 31.02 2.338 ;
      RECT 30.73 1.985 31.03 2.313 ;
      RECT 30.75 1.965 30.86 2.435 ;
      RECT 30.76 1.96 30.86 2.435 ;
      RECT 30.28 3.222 30.47 3.585 ;
      RECT 30.28 3.237 30.51 3.583 ;
      RECT 30.28 3.265 30.53 3.579 ;
      RECT 30.28 3.3 30.54 3.577 ;
      RECT 30.28 3.345 30.55 3.576 ;
      RECT 30.27 3.217 30.43 3.565 ;
      RECT 30.25 3.225 30.47 3.515 ;
      RECT 30.22 3.237 30.51 3.45 ;
      RECT 30.28 3.215 30.43 3.585 ;
      RECT 30.285 7.855 30.455 8.305 ;
      RECT 30.34 6.075 30.51 8.025 ;
      RECT 30.285 5.015 30.455 6.245 ;
      RECT 29.765 5.015 29.935 8.305 ;
      RECT 29.765 7.315 30.17 7.645 ;
      RECT 29.765 6.475 30.17 6.805 ;
      RECT 29.866 2.695 30.07 3.105 ;
      RECT 29.78 2.588 29.866 3.09 ;
      RECT 29.776 2.584 29.78 3.074 ;
      RECT 29.69 2.695 30.07 3.054 ;
      RECT 29.67 2.575 29.69 3.015 ;
      RECT 29.66 2.58 29.776 2.99 ;
      RECT 29.65 2.587 29.78 2.97 ;
      RECT 29.64 2.592 29.87 2.945 ;
      RECT 29.63 2.61 29.96 2.925 ;
      RECT 29.62 2.615 29.96 2.905 ;
      RECT 29.61 2.62 30 2.77 ;
      RECT 29.61 2.65 30.06 2.77 ;
      RECT 29.61 2.635 30.05 2.77 ;
      RECT 29.64 2.605 29.96 2.945 ;
      RECT 29.64 2.593 29.9 2.945 ;
      RECT 29.79 3.42 30.04 3.885 ;
      RECT 29.71 3.395 30.03 3.88 ;
      RECT 29.64 3.429 30.04 3.87 ;
      RECT 29.43 3.68 30.04 3.865 ;
      RECT 29.61 3.449 30.04 3.865 ;
      RECT 29.45 3.64 30.04 3.865 ;
      RECT 29.6 3.46 30.04 3.865 ;
      RECT 29.49 3.58 30.04 3.865 ;
      RECT 29.54 3.505 30.04 3.865 ;
      RECT 29.79 3.37 30.03 3.885 ;
      RECT 29.81 3.365 30.03 3.885 ;
      RECT 29.82 3.36 29.95 3.885 ;
      RECT 29.906 3.355 29.91 3.885 ;
      RECT 29.38 1.925 29.466 2.362 ;
      RECT 29.37 1.925 29.466 2.358 ;
      RECT 29.37 1.925 29.53 2.357 ;
      RECT 29.37 1.925 29.56 2.355 ;
      RECT 29.37 1.925 29.57 2.345 ;
      RECT 29.36 1.93 29.57 2.343 ;
      RECT 29.35 1.94 29.57 2.335 ;
      RECT 29.35 1.94 29.58 2.295 ;
      RECT 29.37 1.925 29.6 2.21 ;
      RECT 29.34 1.95 29.6 2.205 ;
      RECT 29.35 1.94 29.61 2.135 ;
      RECT 29.33 1.96 29.61 2.08 ;
      RECT 29.32 1.97 29.61 1.98 ;
      RECT 29.4 2.741 29.41 2.82 ;
      RECT 29.39 2.734 29.4 3.005 ;
      RECT 29.38 2.728 29.39 3.03 ;
      RECT 29.37 2.72 29.38 3.06 ;
      RECT 29.33 2.715 29.37 3.11 ;
      RECT 29.31 2.715 29.33 3.165 ;
      RECT 29.3 2.715 29.31 3.19 ;
      RECT 29.29 2.715 29.3 3.205 ;
      RECT 29.26 2.715 29.29 3.25 ;
      RECT 29.25 2.715 29.26 3.29 ;
      RECT 29.23 2.715 29.25 3.315 ;
      RECT 29.21 2.715 29.23 3.35 ;
      RECT 29.13 2.715 29.21 3.395 ;
      RECT 29.12 2.715 29.13 3.415 ;
      RECT 29.08 2.795 29.12 3.412 ;
      RECT 29.06 2.875 29.08 3.409 ;
      RECT 29.04 2.93 29.06 3.407 ;
      RECT 29.02 2.99 29.04 3.405 ;
      RECT 28.98 3.025 29.02 3.403 ;
      RECT 28.976 3.035 28.98 3.401 ;
      RECT 28.89 3.05 28.976 3.397 ;
      RECT 28.87 3.07 28.89 3.393 ;
      RECT 28.8 3.075 28.87 3.389 ;
      RECT 28.78 3.076 28.8 3.386 ;
      RECT 28.776 3.078 28.78 3.385 ;
      RECT 28.69 3.087 28.776 3.38 ;
      RECT 28.68 3.096 28.69 3.375 ;
      RECT 28.64 3.102 28.68 3.37 ;
      RECT 28.59 3.113 28.64 3.355 ;
      RECT 28.57 3.122 28.59 3.34 ;
      RECT 28.49 3.135 28.57 3.325 ;
      RECT 28.66 2.685 28.83 2.895 ;
      RECT 28.776 2.677 28.83 2.895 ;
      RECT 28.576 2.685 28.83 2.885 ;
      RECT 28.49 2.685 28.83 2.865 ;
      RECT 28.49 2.69 28.84 2.81 ;
      RECT 28.49 2.7 28.85 2.72 ;
      RECT 28.69 2.682 28.83 2.895 ;
      RECT 28.44 3.623 28.69 3.955 ;
      RECT 28.41 3.635 28.69 3.937 ;
      RECT 28.39 3.67 28.69 3.907 ;
      RECT 28.44 3.62 28.612 3.955 ;
      RECT 28.44 3.616 28.526 3.955 ;
      RECT 28.37 1.965 28.55 2.385 ;
      RECT 28.37 1.965 28.57 2.375 ;
      RECT 28.37 1.965 28.59 2.35 ;
      RECT 28.37 1.965 28.6 2.335 ;
      RECT 28.37 1.965 28.61 2.33 ;
      RECT 28.37 2.005 28.63 2.315 ;
      RECT 28.37 2.075 28.65 2.295 ;
      RECT 28.35 2.075 28.65 2.29 ;
      RECT 28.35 2.135 28.66 2.265 ;
      RECT 28.35 2.175 28.67 2.215 ;
      RECT 28.33 1.965 28.61 2.195 ;
      RECT 28.32 1.975 28.61 2.118 ;
      RECT 28.31 2.015 28.63 2.063 ;
      RECT 27.91 3.375 28.08 3.895 ;
      RECT 27.9 3.375 28.08 3.855 ;
      RECT 27.89 3.395 28.08 3.83 ;
      RECT 27.9 3.375 28.09 3.825 ;
      RECT 27.88 3.435 28.09 3.795 ;
      RECT 27.87 3.47 28.09 3.775 ;
      RECT 27.86 3.52 28.09 3.735 ;
      RECT 27.9 3.386 28.1 3.725 ;
      RECT 27.85 3.6 28.1 3.675 ;
      RECT 27.89 3.409 28.11 3.605 ;
      RECT 27.89 3.433 28.12 3.5 ;
      RECT 27.83 2.68 27.85 2.955 ;
      RECT 27.79 2.665 27.83 3 ;
      RECT 27.77 2.65 27.79 3.065 ;
      RECT 27.75 2.649 27.77 3.14 ;
      RECT 27.73 2.657 27.75 3.245 ;
      RECT 27.726 2.662 27.73 3.297 ;
      RECT 27.64 2.681 27.726 3.337 ;
      RECT 27.63 2.702 27.64 3.376 ;
      RECT 27.62 2.71 27.63 3.377 ;
      RECT 27.6 2.845 27.62 3.379 ;
      RECT 27.59 2.995 27.6 3.381 ;
      RECT 27.55 3.08 27.59 3.386 ;
      RECT 27.468 3.102 27.55 3.396 ;
      RECT 27.382 3.117 27.468 3.409 ;
      RECT 27.296 3.132 27.382 3.422 ;
      RECT 27.21 3.147 27.296 3.436 ;
      RECT 27.13 3.161 27.21 3.449 ;
      RECT 27.116 3.169 27.13 3.457 ;
      RECT 27.03 3.177 27.116 3.471 ;
      RECT 27.02 3.185 27.03 3.484 ;
      RECT 26.996 3.185 27.02 3.492 ;
      RECT 26.91 3.187 26.996 3.522 ;
      RECT 26.83 3.189 26.91 3.565 ;
      RECT 26.76 3.192 26.83 3.6 ;
      RECT 26.74 3.194 26.76 3.616 ;
      RECT 26.71 3.2 26.74 3.618 ;
      RECT 26.66 3.215 26.71 3.621 ;
      RECT 26.64 3.23 26.66 3.624 ;
      RECT 26.61 3.235 26.64 3.627 ;
      RECT 26.55 3.25 26.61 3.631 ;
      RECT 26.54 3.266 26.55 3.635 ;
      RECT 26.49 3.276 26.54 3.624 ;
      RECT 26.46 3.295 26.49 3.607 ;
      RECT 26.44 3.315 26.46 3.597 ;
      RECT 26.42 3.34 26.44 3.589 ;
      RECT 27.43 1.932 27.6 2.425 ;
      RECT 27.42 1.932 27.6 2.41 ;
      RECT 27.42 1.947 27.63 2.4 ;
      RECT 27.41 1.947 27.63 2.375 ;
      RECT 27.4 1.947 27.63 2.34 ;
      RECT 27.4 1.955 27.64 2.295 ;
      RECT 27.38 1.925 27.57 2.275 ;
      RECT 27.37 1.932 27.6 2.235 ;
      RECT 27.36 1.947 27.63 2.215 ;
      RECT 27.35 1.96 27.64 2.175 ;
      RECT 27.34 1.975 27.64 2.128 ;
      RECT 27.34 1.975 27.65 2.12 ;
      RECT 27.33 1.99 27.65 2.093 ;
      RECT 27.34 1.985 27.66 2.035 ;
      RECT 27.14 2.612 27.41 2.905 ;
      RECT 27.14 2.614 27.42 2.9 ;
      RECT 27.13 2.64 27.42 2.895 ;
      RECT 27.14 2.63 27.43 2.89 ;
      RECT 27.14 2.608 27.376 2.905 ;
      RECT 27.14 2.605 27.29 2.905 ;
      RECT 27.2 2.6 27.286 2.905 ;
      RECT 26.69 2.648 26.76 2.945 ;
      RECT 26.69 2.648 26.77 2.944 ;
      RECT 26.77 2.635 26.78 2.941 ;
      RECT 26.67 2.662 26.78 2.935 ;
      RECT 26.76 2.64 26.85 2.931 ;
      RECT 26.69 2.655 26.87 2.92 ;
      RECT 26.67 2.72 26.88 2.916 ;
      RECT 26.65 2.668 26.87 2.915 ;
      RECT 26.64 2.673 26.87 2.905 ;
      RECT 26.63 2.795 26.89 2.9 ;
      RECT 26.63 2.875 26.9 2.89 ;
      RECT 26.6 2.681 26.87 2.884 ;
      RECT 26.59 2.695 26.87 2.869 ;
      RECT 26.63 2.676 26.87 2.9 ;
      RECT 26.76 2.636 26.78 2.941 ;
      RECT 26.58 2.072 26.6 2.305 ;
      RECT 26.57 2.053 26.58 2.31 ;
      RECT 26.56 2.041 26.57 2.317 ;
      RECT 26.52 2.027 26.56 2.327 ;
      RECT 26.51 2.017 26.52 2.336 ;
      RECT 26.46 2.002 26.51 2.341 ;
      RECT 26.45 1.987 26.46 2.347 ;
      RECT 26.43 1.978 26.45 2.352 ;
      RECT 26.42 1.968 26.43 2.358 ;
      RECT 26.41 1.965 26.42 2.363 ;
      RECT 26.39 1.965 26.41 2.364 ;
      RECT 26.36 1.96 26.39 2.362 ;
      RECT 26.336 1.953 26.36 2.361 ;
      RECT 26.25 1.943 26.336 2.358 ;
      RECT 26.24 1.935 26.25 2.355 ;
      RECT 26.218 1.935 26.24 2.354 ;
      RECT 26.132 1.935 26.218 2.352 ;
      RECT 26.046 1.935 26.132 2.35 ;
      RECT 25.96 1.935 26.046 2.347 ;
      RECT 25.95 1.935 25.96 2.34 ;
      RECT 25.92 1.935 25.95 2.3 ;
      RECT 25.91 1.945 25.92 2.255 ;
      RECT 25.9 1.99 25.91 2.24 ;
      RECT 25.87 2.085 25.9 2.195 ;
      RECT 26.06 2.822 26.23 3.335 ;
      RECT 26.05 2.853 26.23 3.315 ;
      RECT 26.05 2.853 26.25 3.285 ;
      RECT 26.04 2.861 26.25 3.26 ;
      RECT 26.04 2.861 26.26 3.25 ;
      RECT 26.04 2.861 26.27 3.23 ;
      RECT 26.04 2.861 26.32 3.185 ;
      RECT 26.04 2.861 26.33 3.16 ;
      RECT 26.04 2.861 26.34 3.125 ;
      RECT 26.04 2.861 26.35 3.09 ;
      RECT 26.04 2.861 26.36 3.04 ;
      RECT 26.04 2.861 26.38 2.965 ;
      RECT 26.21 2.725 26.39 2.905 ;
      RECT 26.13 2.78 26.39 2.905 ;
      RECT 26.17 2.745 26.23 3.335 ;
      RECT 26.16 2.765 26.39 2.905 ;
      RECT 25.52 3.235 25.606 3.801 ;
      RECT 25.48 3.235 25.606 3.795 ;
      RECT 25.48 3.235 25.692 3.793 ;
      RECT 25.48 3.235 25.73 3.787 ;
      RECT 25.48 3.242 25.74 3.785 ;
      RECT 25.45 3.235 25.73 3.78 ;
      RECT 25.42 3.25 25.74 3.77 ;
      RECT 25.42 3.277 25.78 3.762 ;
      RECT 25.395 3.277 25.78 3.75 ;
      RECT 25.395 3.315 25.79 3.732 ;
      RECT 25.38 3.297 25.78 3.725 ;
      RECT 25.38 3.345 25.8 3.721 ;
      RECT 25.38 3.411 25.82 3.705 ;
      RECT 25.38 3.466 25.83 3.515 ;
      RECT 25.57 2.755 25.74 2.935 ;
      RECT 25.52 2.694 25.57 2.92 ;
      RECT 25.26 2.675 25.52 2.905 ;
      RECT 25.22 2.735 25.69 2.905 ;
      RECT 25.22 2.725 25.65 2.905 ;
      RECT 25.22 2.714 25.63 2.905 ;
      RECT 25.22 2.7 25.57 2.905 ;
      RECT 25.26 2.67 25.456 2.905 ;
      RECT 25.29 2.649 25.456 2.905 ;
      RECT 25.27 2.65 25.456 2.905 ;
      RECT 25.29 2.635 25.37 2.905 ;
      RECT 25.05 3.165 25.17 3.605 ;
      RECT 25.03 3.165 25.17 3.604 ;
      RECT 24.99 3.185 25.17 3.601 ;
      RECT 24.95 3.229 25.17 3.597 ;
      RECT 24.94 3.259 25.19 3.46 ;
      RECT 25.03 3.165 25.2 3.355 ;
      RECT 24.69 1.945 24.7 2.395 ;
      RECT 24.5 1.945 24.52 2.355 ;
      RECT 24.47 1.945 24.48 2.335 ;
      RECT 25.15 2.255 25.17 2.44 ;
      RECT 25.13 2.215 25.15 2.448 ;
      RECT 25.08 2.182 25.13 2.458 ;
      RECT 25.026 2.156 25.08 2.461 ;
      RECT 24.94 2.121 25.026 2.451 ;
      RECT 24.93 2.097 24.94 2.44 ;
      RECT 24.86 2.063 24.93 2.43 ;
      RECT 24.84 2.023 24.86 2.423 ;
      RECT 24.82 2.005 24.84 2.419 ;
      RECT 24.81 1.995 24.82 2.416 ;
      RECT 24.78 1.98 24.81 2.412 ;
      RECT 24.77 1.965 24.78 2.408 ;
      RECT 24.76 1.96 24.77 2.406 ;
      RECT 24.71 1.95 24.76 2.401 ;
      RECT 24.7 1.945 24.71 2.396 ;
      RECT 24.67 1.945 24.69 2.39 ;
      RECT 24.636 1.945 24.67 2.382 ;
      RECT 24.55 1.945 24.636 2.372 ;
      RECT 24.52 1.945 24.55 2.36 ;
      RECT 24.48 1.945 24.5 2.345 ;
      RECT 24.46 1.945 24.47 2.328 ;
      RECT 24.44 1.955 24.46 2.308 ;
      RECT 24.43 1.975 24.44 2.24 ;
      RECT 24.42 1.985 24.43 2 ;
      RECT 24.69 2.665 24.776 2.99 ;
      RECT 24.69 2.665 24.81 2.982 ;
      RECT 24.64 2.665 24.81 2.98 ;
      RECT 24.64 2.669 24.896 2.975 ;
      RECT 24.64 2.674 24.92 2.968 ;
      RECT 24.64 2.68 24.93 2.966 ;
      RECT 24.64 2.69 24.94 2.963 ;
      RECT 24.64 2.83 24.95 2.958 ;
      RECT 24.7 3.34 24.75 3.656 ;
      RECT 24.69 3.32 24.7 3.681 ;
      RECT 24.68 3.31 24.69 3.69 ;
      RECT 24.66 3.304 24.68 3.705 ;
      RECT 24.63 3.302 24.66 3.725 ;
      RECT 24.616 3.3 24.63 3.735 ;
      RECT 24.53 3.296 24.616 3.735 ;
      RECT 24.46 3.29 24.53 3.725 ;
      RECT 24.38 3.285 24.46 3.7 ;
      RECT 24.32 3.281 24.38 3.665 ;
      RECT 24.25 3.277 24.32 3.625 ;
      RECT 24.22 3.275 24.25 3.6 ;
      RECT 24.116 3.273 24.16 3.595 ;
      RECT 24.03 3.268 24.116 3.595 ;
      RECT 23.95 3.265 24.03 3.595 ;
      RECT 23.87 3.266 23.95 3.62 ;
      RECT 23.788 3.268 23.87 3.645 ;
      RECT 23.702 3.269 23.788 3.645 ;
      RECT 23.616 3.271 23.702 3.645 ;
      RECT 23.53 3.273 23.616 3.645 ;
      RECT 23.51 3.274 23.53 3.637 ;
      RECT 23.5 3.28 23.51 3.626 ;
      RECT 23.46 3.3 23.5 3.607 ;
      RECT 23.45 3.32 23.46 3.589 ;
      RECT 24.16 3.275 24.22 3.595 ;
      RECT 24.13 2.82 24.3 3.075 ;
      RECT 24.13 2.82 24.31 3.068 ;
      RECT 24.13 2.82 24.32 3.053 ;
      RECT 24.13 2.82 24.34 3.035 ;
      RECT 24.13 2.82 24.38 2.99 ;
      RECT 24.31 2.585 24.4 2.943 ;
      RECT 24.3 2.59 24.41 2.924 ;
      RECT 24.25 2.605 24.42 2.911 ;
      RECT 24.24 2.62 24.43 2.895 ;
      RECT 24.14 2.785 24.43 2.895 ;
      RECT 24.18 2.645 24.3 3.075 ;
      RECT 24.15 2.755 24.43 2.895 ;
      RECT 24.17 2.68 24.3 3.075 ;
      RECT 24.16 2.705 24.43 2.895 ;
      RECT 24.28 2.591 24.41 2.924 ;
      RECT 24.3 2.586 24.4 2.943 ;
      RECT 23.76 2.72 23.95 2.895 ;
      RECT 23.72 2.638 23.91 2.89 ;
      RECT 23.686 2.643 23.91 2.884 ;
      RECT 23.6 2.65 23.91 2.879 ;
      RECT 23.516 2.665 23.91 2.874 ;
      RECT 23.43 2.685 23.94 2.868 ;
      RECT 23.516 2.675 23.94 2.874 ;
      RECT 23.76 2.635 23.91 2.895 ;
      RECT 23.76 2.631 23.86 2.895 ;
      RECT 23.846 2.626 23.86 2.895 ;
      RECT 22.6 1.954 23.26 2.345 ;
      RECT 22.858 1.948 23.26 2.345 ;
      RECT 22.59 1.96 23.26 2.344 ;
      RECT 22.58 1.975 23.26 2.343 ;
      RECT 22.52 2.015 23.26 2.339 ;
      RECT 22.686 1.953 23.27 2.335 ;
      RECT 22.59 1.96 23.28 2.325 ;
      RECT 22.59 1.968 23.29 2.305 ;
      RECT 22.58 1.978 23.31 2.278 ;
      RECT 22.52 2.015 23.32 2.253 ;
      RECT 22.58 1.985 23.33 2.24 ;
      RECT 22.686 1.951 23.26 2.345 ;
      RECT 22.772 1.949 23.26 2.345 ;
      RECT 22.858 1.947 23.24 2.345 ;
      RECT 22.944 1.945 23.24 2.345 ;
      RECT 23.11 3.12 23.28 3.315 ;
      RECT 23.1 3.12 23.28 3.26 ;
      RECT 23.095 3.12 23.28 3.188 ;
      RECT 23.08 3.06 23.26 3.155 ;
      RECT 23.07 3.06 23.26 3.105 ;
      RECT 23.04 3.035 23.25 3.06 ;
      RECT 23.02 3.035 23.25 3.045 ;
      RECT 22.96 2.725 23.14 3.036 ;
      RECT 22.96 2.96 23.24 3.036 ;
      RECT 22.95 2.724 22.96 3.026 ;
      RECT 22.93 2.723 22.95 3.02 ;
      RECT 22.9 2.722 22.93 3 ;
      RECT 22.85 2.719 22.9 2.965 ;
      RECT 22.85 2.84 23.21 2.965 ;
      RECT 22.78 2.716 22.85 2.92 ;
      RECT 22.78 2.775 23.19 2.92 ;
      RECT 22.78 2.765 23.18 2.92 ;
      RECT 22.78 2.755 23.17 2.92 ;
      RECT 22.78 2.735 23.15 2.92 ;
      RECT 22.86 3.255 22.87 3.512 ;
      RECT 22.84 3.172 22.86 3.532 ;
      RECT 22.82 3.166 22.84 3.56 ;
      RECT 22.76 3.154 22.82 3.58 ;
      RECT 22.72 3.14 22.76 3.581 ;
      RECT 22.636 3.129 22.72 3.569 ;
      RECT 22.55 3.116 22.636 3.553 ;
      RECT 22.54 3.109 22.55 3.545 ;
      RECT 22.49 3.106 22.54 3.485 ;
      RECT 22.47 3.102 22.49 3.4 ;
      RECT 22.46 3.1 22.47 3.35 ;
      RECT 22.43 3.098 22.46 3.32 ;
      RECT 22.39 3.093 22.43 3.3 ;
      RECT 22.352 3.088 22.39 3.288 ;
      RECT 22.266 3.08 22.352 3.297 ;
      RECT 22.18 3.069 22.266 3.309 ;
      RECT 22.11 3.059 22.18 3.319 ;
      RECT 22.09 3.05 22.11 3.324 ;
      RECT 22.03 3.022 22.09 3.32 ;
      RECT 22.01 2.992 22.03 3.308 ;
      RECT 21.99 2.965 22.01 3.295 ;
      RECT 21.91 2.718 21.99 3.262 ;
      RECT 21.896 2.71 21.91 3.224 ;
      RECT 21.81 2.702 21.896 3.145 ;
      RECT 21.79 2.693 21.81 3.061 ;
      RECT 21.76 2.688 21.79 3.041 ;
      RECT 21.69 2.699 21.76 3.026 ;
      RECT 21.67 2.717 21.69 3 ;
      RECT 21.66 2.723 21.67 2.945 ;
      RECT 21.64 2.745 21.66 2.83 ;
      RECT 22.3 2.705 22.47 2.895 ;
      RECT 22.3 2.705 22.5 2.89 ;
      RECT 22.35 2.615 22.52 2.88 ;
      RECT 22.31 2.65 22.52 2.88 ;
      RECT 21.51 3.388 21.58 3.829 ;
      RECT 21.45 3.413 21.58 3.826 ;
      RECT 21.45 3.413 21.63 3.819 ;
      RECT 21.44 3.435 21.63 3.816 ;
      RECT 21.58 3.375 21.65 3.814 ;
      RECT 21.51 3.4 21.73 3.811 ;
      RECT 21.44 3.439 21.78 3.807 ;
      RECT 21.42 3.465 21.78 3.795 ;
      RECT 21.44 3.459 21.8 3.79 ;
      RECT 21.42 2.205 21.46 2.445 ;
      RECT 21.42 2.205 21.49 2.444 ;
      RECT 21.42 2.205 21.6 2.436 ;
      RECT 21.42 2.205 21.66 2.415 ;
      RECT 21.43 2.15 21.71 2.315 ;
      RECT 21.54 1.99 21.57 2.437 ;
      RECT 21.57 1.985 21.75 2.195 ;
      RECT 21.44 2.125 21.75 2.195 ;
      RECT 21.49 2.02 21.54 2.44 ;
      RECT 21.46 2.075 21.75 2.195 ;
      RECT 20.33 5.02 20.5 6.49 ;
      RECT 20.33 6.315 20.505 6.485 ;
      RECT 19.96 1.74 20.13 2.93 ;
      RECT 19.96 1.74 20.43 1.91 ;
      RECT 19.96 6.97 20.43 7.14 ;
      RECT 19.96 5.95 20.13 7.14 ;
      RECT 18.97 1.74 19.14 2.93 ;
      RECT 18.97 1.74 19.44 1.91 ;
      RECT 18.97 6.97 19.44 7.14 ;
      RECT 18.97 5.95 19.14 7.14 ;
      RECT 17.12 2.635 17.29 3.865 ;
      RECT 17.175 0.855 17.345 2.805 ;
      RECT 17.12 0.575 17.29 1.025 ;
      RECT 17.12 7.855 17.29 8.305 ;
      RECT 17.175 6.075 17.345 8.025 ;
      RECT 17.12 5.015 17.29 6.245 ;
      RECT 16.6 0.575 16.77 3.865 ;
      RECT 16.6 2.075 17.005 2.405 ;
      RECT 16.6 1.235 17.005 1.565 ;
      RECT 16.6 5.015 16.77 8.305 ;
      RECT 16.6 7.315 17.005 7.645 ;
      RECT 16.6 6.475 17.005 6.805 ;
      RECT 14.695 3.39 14.715 3.44 ;
      RECT 14.675 3.362 14.695 3.555 ;
      RECT 14.655 3.337 14.675 3.611 ;
      RECT 14.615 3.325 14.655 3.63 ;
      RECT 14.565 3.32 14.615 3.659 ;
      RECT 14.561 3.314 14.565 3.675 ;
      RECT 14.475 3.306 14.561 3.675 ;
      RECT 14.415 3.294 14.475 3.67 ;
      RECT 14.361 3.284 14.415 3.659 ;
      RECT 14.275 3.272 14.361 3.642 ;
      RECT 14.253 3.263 14.275 3.629 ;
      RECT 14.167 3.256 14.253 3.616 ;
      RECT 14.081 3.243 14.167 3.595 ;
      RECT 13.995 3.231 14.081 3.575 ;
      RECT 13.965 3.22 13.995 3.561 ;
      RECT 13.915 3.207 13.965 3.551 ;
      RECT 13.895 3.197 13.915 3.545 ;
      RECT 13.841 3.187 13.895 3.539 ;
      RECT 13.755 3.167 13.841 3.523 ;
      RECT 13.715 3.155 13.755 3.509 ;
      RECT 13.68 3.155 13.715 3.495 ;
      RECT 13.665 3.155 13.68 3.48 ;
      RECT 13.615 3.155 13.665 3.425 ;
      RECT 13.585 3.155 13.615 3.345 ;
      RECT 14.115 2.825 14.285 3.075 ;
      RECT 14.115 2.825 14.295 3.03 ;
      RECT 14.175 2.655 14.305 2.975 ;
      RECT 14.175 2.662 14.315 2.94 ;
      RECT 14.135 2.677 14.325 2.875 ;
      RECT 14.125 2.76 14.325 2.875 ;
      RECT 14.135 2.695 14.335 2.785 ;
      RECT 14.135 2.675 14.315 2.94 ;
      RECT 13.905 1.93 14.075 2.415 ;
      RECT 13.895 1.93 14.075 2.405 ;
      RECT 13.895 1.945 14.095 2.35 ;
      RECT 13.855 1.925 14.045 2.315 ;
      RECT 13.855 1.96 14.105 2.235 ;
      RECT 13.805 1.945 14.095 2.135 ;
      RECT 13.805 1.975 14.115 2.095 ;
      RECT 13.805 1.99 14.125 2.015 ;
      RECT 13.401 2.688 13.415 2.944 ;
      RECT 13.401 2.689 13.501 2.939 ;
      RECT 13.315 2.686 13.401 2.936 ;
      RECT 13.305 2.685 13.315 2.929 ;
      RECT 13.305 2.692 13.587 2.926 ;
      RECT 13.225 2.695 13.587 2.922 ;
      RECT 13.305 2.694 13.605 2.919 ;
      RECT 13.215 2.707 13.625 2.916 ;
      RECT 13.225 2.695 13.625 2.916 ;
      RECT 13.205 2.712 13.625 2.915 ;
      RECT 13.225 2.697 13.711 2.911 ;
      RECT 13.185 2.715 13.711 2.908 ;
      RECT 13.225 2.701 13.797 2.902 ;
      RECT 13.175 2.72 13.797 2.898 ;
      RECT 13.225 2.704 13.825 2.897 ;
      RECT 13.225 2.705 13.865 2.891 ;
      RECT 13.215 2.71 13.875 2.886 ;
      RECT 13.175 2.73 13.885 2.875 ;
      RECT 13.175 2.75 13.895 2.86 ;
      RECT 13.135 3.298 13.155 3.605 ;
      RECT 13.125 3.273 13.135 3.885 ;
      RECT 13.085 3.24 13.125 3.885 ;
      RECT 13.081 3.21 13.085 3.885 ;
      RECT 12.995 3.095 13.081 3.885 ;
      RECT 12.985 2.97 12.995 3.885 ;
      RECT 12.975 2.935 12.985 3.885 ;
      RECT 12.965 2.905 12.975 3.885 ;
      RECT 12.945 2.875 12.965 3.77 ;
      RECT 12.935 2.845 12.945 3.645 ;
      RECT 12.925 2.825 12.935 3.595 ;
      RECT 12.905 2.795 12.925 3.503 ;
      RECT 12.885 2.761 12.905 3.418 ;
      RECT 12.88 2.744 12.885 3.353 ;
      RECT 12.875 2.738 12.88 3.325 ;
      RECT 12.865 2.73 12.875 3.29 ;
      RECT 12.845 2.725 12.855 3.19 ;
      RECT 12.835 2.725 12.845 3.165 ;
      RECT 12.83 2.725 12.835 3.128 ;
      RECT 12.815 2.725 12.83 3.06 ;
      RECT 12.805 2.724 12.815 2.99 ;
      RECT 12.795 2.722 12.805 2.97 ;
      RECT 12.735 2.718 12.795 2.943 ;
      RECT 12.695 2.72 12.735 2.923 ;
      RECT 12.675 2.75 12.695 2.905 ;
      RECT 12.855 2.725 12.865 3.245 ;
      RECT 12.795 2.08 12.965 2.435 ;
      RECT 12.825 1.966 12.965 2.435 ;
      RECT 12.825 1.968 12.975 2.43 ;
      RECT 12.825 1.97 12.995 2.42 ;
      RECT 12.825 1.973 13.025 2.405 ;
      RECT 12.825 1.978 13.075 2.375 ;
      RECT 12.825 1.983 13.095 2.338 ;
      RECT 12.805 1.985 13.105 2.313 ;
      RECT 12.825 1.965 12.935 2.435 ;
      RECT 12.835 1.96 12.935 2.435 ;
      RECT 12.355 3.222 12.545 3.585 ;
      RECT 12.355 3.237 12.585 3.583 ;
      RECT 12.355 3.265 12.605 3.579 ;
      RECT 12.355 3.3 12.615 3.577 ;
      RECT 12.355 3.345 12.625 3.576 ;
      RECT 12.345 3.217 12.505 3.565 ;
      RECT 12.325 3.225 12.545 3.515 ;
      RECT 12.295 3.237 12.585 3.45 ;
      RECT 12.355 3.215 12.505 3.585 ;
      RECT 12.36 7.855 12.53 8.305 ;
      RECT 12.415 6.075 12.585 8.025 ;
      RECT 12.36 5.015 12.53 6.245 ;
      RECT 11.84 5.015 12.01 8.305 ;
      RECT 11.84 7.315 12.245 7.645 ;
      RECT 11.84 6.475 12.245 6.805 ;
      RECT 11.941 2.695 12.145 3.105 ;
      RECT 11.855 2.588 11.941 3.09 ;
      RECT 11.851 2.584 11.855 3.074 ;
      RECT 11.765 2.695 12.145 3.054 ;
      RECT 11.745 2.575 11.765 3.015 ;
      RECT 11.735 2.58 11.851 2.99 ;
      RECT 11.725 2.587 11.855 2.97 ;
      RECT 11.715 2.592 11.945 2.945 ;
      RECT 11.705 2.61 12.035 2.925 ;
      RECT 11.695 2.615 12.035 2.905 ;
      RECT 11.685 2.62 12.075 2.77 ;
      RECT 11.685 2.65 12.135 2.77 ;
      RECT 11.685 2.635 12.125 2.77 ;
      RECT 11.715 2.605 12.035 2.945 ;
      RECT 11.715 2.593 11.975 2.945 ;
      RECT 11.865 3.42 12.115 3.885 ;
      RECT 11.785 3.395 12.105 3.88 ;
      RECT 11.715 3.429 12.115 3.87 ;
      RECT 11.505 3.68 12.115 3.865 ;
      RECT 11.685 3.449 12.115 3.865 ;
      RECT 11.525 3.64 12.115 3.865 ;
      RECT 11.675 3.46 12.115 3.865 ;
      RECT 11.565 3.58 12.115 3.865 ;
      RECT 11.615 3.505 12.115 3.865 ;
      RECT 11.865 3.37 12.105 3.885 ;
      RECT 11.885 3.365 12.105 3.885 ;
      RECT 11.895 3.36 12.025 3.885 ;
      RECT 11.981 3.355 11.985 3.885 ;
      RECT 11.455 1.925 11.541 2.362 ;
      RECT 11.445 1.925 11.541 2.358 ;
      RECT 11.445 1.925 11.605 2.357 ;
      RECT 11.445 1.925 11.635 2.355 ;
      RECT 11.445 1.925 11.645 2.345 ;
      RECT 11.435 1.93 11.645 2.343 ;
      RECT 11.425 1.94 11.645 2.335 ;
      RECT 11.425 1.94 11.655 2.295 ;
      RECT 11.445 1.925 11.675 2.21 ;
      RECT 11.415 1.95 11.675 2.205 ;
      RECT 11.425 1.94 11.685 2.135 ;
      RECT 11.405 1.96 11.685 2.08 ;
      RECT 11.395 1.97 11.685 1.98 ;
      RECT 11.475 2.741 11.485 2.82 ;
      RECT 11.465 2.734 11.475 3.005 ;
      RECT 11.455 2.728 11.465 3.03 ;
      RECT 11.445 2.72 11.455 3.06 ;
      RECT 11.405 2.715 11.445 3.11 ;
      RECT 11.385 2.715 11.405 3.165 ;
      RECT 11.375 2.715 11.385 3.19 ;
      RECT 11.365 2.715 11.375 3.205 ;
      RECT 11.335 2.715 11.365 3.25 ;
      RECT 11.325 2.715 11.335 3.29 ;
      RECT 11.305 2.715 11.325 3.315 ;
      RECT 11.285 2.715 11.305 3.35 ;
      RECT 11.205 2.715 11.285 3.395 ;
      RECT 11.195 2.715 11.205 3.415 ;
      RECT 11.155 2.795 11.195 3.412 ;
      RECT 11.135 2.875 11.155 3.409 ;
      RECT 11.115 2.93 11.135 3.407 ;
      RECT 11.095 2.99 11.115 3.405 ;
      RECT 11.055 3.025 11.095 3.403 ;
      RECT 11.051 3.035 11.055 3.401 ;
      RECT 10.965 3.05 11.051 3.397 ;
      RECT 10.945 3.07 10.965 3.393 ;
      RECT 10.875 3.075 10.945 3.389 ;
      RECT 10.855 3.076 10.875 3.386 ;
      RECT 10.851 3.078 10.855 3.385 ;
      RECT 10.765 3.087 10.851 3.38 ;
      RECT 10.755 3.096 10.765 3.375 ;
      RECT 10.715 3.102 10.755 3.37 ;
      RECT 10.665 3.113 10.715 3.355 ;
      RECT 10.645 3.122 10.665 3.34 ;
      RECT 10.565 3.135 10.645 3.325 ;
      RECT 10.735 2.685 10.905 2.895 ;
      RECT 10.851 2.677 10.905 2.895 ;
      RECT 10.651 2.685 10.905 2.885 ;
      RECT 10.565 2.685 10.905 2.865 ;
      RECT 10.565 2.69 10.915 2.81 ;
      RECT 10.565 2.7 10.925 2.72 ;
      RECT 10.765 2.682 10.905 2.895 ;
      RECT 10.515 3.623 10.765 3.955 ;
      RECT 10.485 3.635 10.765 3.937 ;
      RECT 10.465 3.67 10.765 3.907 ;
      RECT 10.515 3.62 10.687 3.955 ;
      RECT 10.515 3.616 10.601 3.955 ;
      RECT 10.445 1.965 10.625 2.385 ;
      RECT 10.445 1.965 10.645 2.375 ;
      RECT 10.445 1.965 10.665 2.35 ;
      RECT 10.445 1.965 10.675 2.335 ;
      RECT 10.445 1.965 10.685 2.33 ;
      RECT 10.445 2.005 10.705 2.315 ;
      RECT 10.445 2.075 10.725 2.295 ;
      RECT 10.425 2.075 10.725 2.29 ;
      RECT 10.425 2.135 10.735 2.265 ;
      RECT 10.425 2.175 10.745 2.215 ;
      RECT 10.405 1.965 10.685 2.195 ;
      RECT 10.395 1.975 10.685 2.118 ;
      RECT 10.385 2.015 10.705 2.063 ;
      RECT 9.985 3.375 10.155 3.895 ;
      RECT 9.975 3.375 10.155 3.855 ;
      RECT 9.965 3.395 10.155 3.83 ;
      RECT 9.975 3.375 10.165 3.825 ;
      RECT 9.955 3.435 10.165 3.795 ;
      RECT 9.945 3.47 10.165 3.775 ;
      RECT 9.935 3.52 10.165 3.735 ;
      RECT 9.975 3.386 10.175 3.725 ;
      RECT 9.925 3.6 10.175 3.675 ;
      RECT 9.965 3.409 10.185 3.605 ;
      RECT 9.965 3.433 10.195 3.5 ;
      RECT 9.905 2.68 9.925 2.955 ;
      RECT 9.865 2.665 9.905 3 ;
      RECT 9.845 2.65 9.865 3.065 ;
      RECT 9.825 2.649 9.845 3.14 ;
      RECT 9.805 2.657 9.825 3.245 ;
      RECT 9.801 2.662 9.805 3.297 ;
      RECT 9.715 2.681 9.801 3.337 ;
      RECT 9.705 2.702 9.715 3.376 ;
      RECT 9.695 2.71 9.705 3.377 ;
      RECT 9.675 2.845 9.695 3.379 ;
      RECT 9.665 2.995 9.675 3.381 ;
      RECT 9.625 3.08 9.665 3.386 ;
      RECT 9.543 3.102 9.625 3.396 ;
      RECT 9.457 3.117 9.543 3.409 ;
      RECT 9.371 3.132 9.457 3.422 ;
      RECT 9.285 3.147 9.371 3.436 ;
      RECT 9.205 3.161 9.285 3.449 ;
      RECT 9.191 3.169 9.205 3.457 ;
      RECT 9.105 3.177 9.191 3.471 ;
      RECT 9.095 3.185 9.105 3.484 ;
      RECT 9.071 3.185 9.095 3.492 ;
      RECT 8.985 3.187 9.071 3.522 ;
      RECT 8.905 3.189 8.985 3.565 ;
      RECT 8.835 3.192 8.905 3.6 ;
      RECT 8.815 3.194 8.835 3.616 ;
      RECT 8.785 3.2 8.815 3.618 ;
      RECT 8.735 3.215 8.785 3.621 ;
      RECT 8.715 3.23 8.735 3.624 ;
      RECT 8.685 3.235 8.715 3.627 ;
      RECT 8.625 3.25 8.685 3.631 ;
      RECT 8.615 3.266 8.625 3.635 ;
      RECT 8.565 3.276 8.615 3.624 ;
      RECT 8.535 3.295 8.565 3.607 ;
      RECT 8.515 3.315 8.535 3.597 ;
      RECT 8.495 3.34 8.515 3.589 ;
      RECT 9.505 1.932 9.675 2.425 ;
      RECT 9.495 1.932 9.675 2.41 ;
      RECT 9.495 1.947 9.705 2.4 ;
      RECT 9.485 1.947 9.705 2.375 ;
      RECT 9.475 1.947 9.705 2.34 ;
      RECT 9.475 1.955 9.715 2.295 ;
      RECT 9.455 1.925 9.645 2.275 ;
      RECT 9.445 1.932 9.675 2.235 ;
      RECT 9.435 1.947 9.705 2.215 ;
      RECT 9.425 1.96 9.715 2.175 ;
      RECT 9.415 1.975 9.715 2.128 ;
      RECT 9.415 1.975 9.725 2.12 ;
      RECT 9.405 1.99 9.725 2.093 ;
      RECT 9.415 1.985 9.735 2.035 ;
      RECT 9.215 2.612 9.485 2.905 ;
      RECT 9.215 2.614 9.495 2.9 ;
      RECT 9.205 2.64 9.495 2.895 ;
      RECT 9.215 2.63 9.505 2.89 ;
      RECT 9.215 2.608 9.451 2.905 ;
      RECT 9.215 2.605 9.365 2.905 ;
      RECT 9.275 2.6 9.361 2.905 ;
      RECT 8.765 2.648 8.835 2.945 ;
      RECT 8.765 2.648 8.845 2.944 ;
      RECT 8.845 2.635 8.855 2.941 ;
      RECT 8.745 2.662 8.855 2.935 ;
      RECT 8.835 2.64 8.925 2.931 ;
      RECT 8.765 2.655 8.945 2.92 ;
      RECT 8.745 2.72 8.955 2.916 ;
      RECT 8.725 2.668 8.945 2.915 ;
      RECT 8.715 2.673 8.945 2.905 ;
      RECT 8.705 2.795 8.965 2.9 ;
      RECT 8.705 2.875 8.975 2.89 ;
      RECT 8.675 2.681 8.945 2.884 ;
      RECT 8.665 2.695 8.945 2.869 ;
      RECT 8.705 2.676 8.945 2.9 ;
      RECT 8.835 2.636 8.855 2.941 ;
      RECT 8.655 2.072 8.675 2.305 ;
      RECT 8.645 2.053 8.655 2.31 ;
      RECT 8.635 2.041 8.645 2.317 ;
      RECT 8.595 2.027 8.635 2.327 ;
      RECT 8.585 2.017 8.595 2.336 ;
      RECT 8.535 2.002 8.585 2.341 ;
      RECT 8.525 1.987 8.535 2.347 ;
      RECT 8.505 1.978 8.525 2.352 ;
      RECT 8.495 1.968 8.505 2.358 ;
      RECT 8.485 1.965 8.495 2.363 ;
      RECT 8.465 1.965 8.485 2.364 ;
      RECT 8.435 1.96 8.465 2.362 ;
      RECT 8.411 1.953 8.435 2.361 ;
      RECT 8.325 1.943 8.411 2.358 ;
      RECT 8.315 1.935 8.325 2.355 ;
      RECT 8.293 1.935 8.315 2.354 ;
      RECT 8.207 1.935 8.293 2.352 ;
      RECT 8.121 1.935 8.207 2.35 ;
      RECT 8.035 1.935 8.121 2.347 ;
      RECT 8.025 1.935 8.035 2.34 ;
      RECT 7.995 1.935 8.025 2.3 ;
      RECT 7.985 1.945 7.995 2.255 ;
      RECT 7.975 1.99 7.985 2.24 ;
      RECT 7.945 2.085 7.975 2.195 ;
      RECT 8.135 2.822 8.305 3.335 ;
      RECT 8.125 2.853 8.305 3.315 ;
      RECT 8.125 2.853 8.325 3.285 ;
      RECT 8.115 2.861 8.325 3.26 ;
      RECT 8.115 2.861 8.335 3.25 ;
      RECT 8.115 2.861 8.345 3.23 ;
      RECT 8.115 2.861 8.395 3.185 ;
      RECT 8.115 2.861 8.405 3.16 ;
      RECT 8.115 2.861 8.415 3.125 ;
      RECT 8.115 2.861 8.425 3.09 ;
      RECT 8.115 2.861 8.435 3.04 ;
      RECT 8.115 2.861 8.455 2.965 ;
      RECT 8.285 2.725 8.465 2.905 ;
      RECT 8.205 2.78 8.465 2.905 ;
      RECT 8.245 2.745 8.305 3.335 ;
      RECT 8.235 2.765 8.465 2.905 ;
      RECT 7.595 3.235 7.681 3.801 ;
      RECT 7.555 3.235 7.681 3.795 ;
      RECT 7.555 3.235 7.767 3.793 ;
      RECT 7.555 3.235 7.805 3.787 ;
      RECT 7.555 3.242 7.815 3.785 ;
      RECT 7.525 3.235 7.805 3.78 ;
      RECT 7.495 3.25 7.815 3.77 ;
      RECT 7.495 3.277 7.855 3.762 ;
      RECT 7.47 3.277 7.855 3.75 ;
      RECT 7.47 3.315 7.865 3.732 ;
      RECT 7.455 3.297 7.855 3.725 ;
      RECT 7.455 3.345 7.875 3.721 ;
      RECT 7.455 3.411 7.895 3.705 ;
      RECT 7.455 3.466 7.905 3.515 ;
      RECT 7.645 2.755 7.815 2.935 ;
      RECT 7.595 2.694 7.645 2.92 ;
      RECT 7.335 2.675 7.595 2.905 ;
      RECT 7.295 2.735 7.765 2.905 ;
      RECT 7.295 2.725 7.725 2.905 ;
      RECT 7.295 2.714 7.705 2.905 ;
      RECT 7.295 2.7 7.645 2.905 ;
      RECT 7.335 2.67 7.531 2.905 ;
      RECT 7.365 2.649 7.531 2.905 ;
      RECT 7.345 2.65 7.531 2.905 ;
      RECT 7.365 2.635 7.445 2.905 ;
      RECT 7.125 3.165 7.245 3.605 ;
      RECT 7.105 3.165 7.245 3.604 ;
      RECT 7.065 3.185 7.245 3.601 ;
      RECT 7.025 3.229 7.245 3.597 ;
      RECT 7.015 3.259 7.265 3.46 ;
      RECT 7.105 3.165 7.275 3.355 ;
      RECT 6.765 1.945 6.775 2.395 ;
      RECT 6.575 1.945 6.595 2.355 ;
      RECT 6.545 1.945 6.555 2.335 ;
      RECT 7.225 2.255 7.245 2.44 ;
      RECT 7.205 2.215 7.225 2.448 ;
      RECT 7.155 2.182 7.205 2.458 ;
      RECT 7.101 2.156 7.155 2.461 ;
      RECT 7.015 2.121 7.101 2.451 ;
      RECT 7.005 2.097 7.015 2.44 ;
      RECT 6.935 2.063 7.005 2.43 ;
      RECT 6.915 2.023 6.935 2.423 ;
      RECT 6.895 2.005 6.915 2.419 ;
      RECT 6.885 1.995 6.895 2.416 ;
      RECT 6.855 1.98 6.885 2.412 ;
      RECT 6.845 1.965 6.855 2.408 ;
      RECT 6.835 1.96 6.845 2.406 ;
      RECT 6.785 1.95 6.835 2.401 ;
      RECT 6.775 1.945 6.785 2.396 ;
      RECT 6.745 1.945 6.765 2.39 ;
      RECT 6.711 1.945 6.745 2.382 ;
      RECT 6.625 1.945 6.711 2.372 ;
      RECT 6.595 1.945 6.625 2.36 ;
      RECT 6.555 1.945 6.575 2.345 ;
      RECT 6.535 1.945 6.545 2.328 ;
      RECT 6.515 1.955 6.535 2.308 ;
      RECT 6.505 1.975 6.515 2.24 ;
      RECT 6.495 1.985 6.505 2 ;
      RECT 6.765 2.665 6.851 2.99 ;
      RECT 6.765 2.665 6.885 2.982 ;
      RECT 6.715 2.665 6.885 2.98 ;
      RECT 6.715 2.669 6.971 2.975 ;
      RECT 6.715 2.674 6.995 2.968 ;
      RECT 6.715 2.68 7.005 2.966 ;
      RECT 6.715 2.69 7.015 2.963 ;
      RECT 6.715 2.83 7.025 2.958 ;
      RECT 6.775 3.34 6.825 3.656 ;
      RECT 6.765 3.32 6.775 3.681 ;
      RECT 6.755 3.31 6.765 3.69 ;
      RECT 6.735 3.304 6.755 3.705 ;
      RECT 6.705 3.302 6.735 3.725 ;
      RECT 6.691 3.3 6.705 3.735 ;
      RECT 6.605 3.296 6.691 3.735 ;
      RECT 6.535 3.29 6.605 3.725 ;
      RECT 6.455 3.285 6.535 3.7 ;
      RECT 6.395 3.281 6.455 3.665 ;
      RECT 6.325 3.277 6.395 3.625 ;
      RECT 6.295 3.275 6.325 3.6 ;
      RECT 6.191 3.273 6.235 3.595 ;
      RECT 6.105 3.268 6.191 3.595 ;
      RECT 6.025 3.265 6.105 3.595 ;
      RECT 5.945 3.266 6.025 3.62 ;
      RECT 5.863 3.268 5.945 3.645 ;
      RECT 5.777 3.269 5.863 3.645 ;
      RECT 5.691 3.271 5.777 3.645 ;
      RECT 5.605 3.273 5.691 3.645 ;
      RECT 5.585 3.274 5.605 3.637 ;
      RECT 5.575 3.28 5.585 3.626 ;
      RECT 5.535 3.3 5.575 3.607 ;
      RECT 5.525 3.32 5.535 3.589 ;
      RECT 6.235 3.275 6.295 3.595 ;
      RECT 6.205 2.82 6.375 3.075 ;
      RECT 6.205 2.82 6.385 3.068 ;
      RECT 6.205 2.82 6.395 3.053 ;
      RECT 6.205 2.82 6.415 3.035 ;
      RECT 6.205 2.82 6.455 2.99 ;
      RECT 6.385 2.585 6.475 2.943 ;
      RECT 6.375 2.59 6.485 2.924 ;
      RECT 6.325 2.605 6.495 2.911 ;
      RECT 6.315 2.62 6.505 2.895 ;
      RECT 6.215 2.785 6.505 2.895 ;
      RECT 6.255 2.645 6.375 3.075 ;
      RECT 6.225 2.755 6.505 2.895 ;
      RECT 6.245 2.68 6.375 3.075 ;
      RECT 6.235 2.705 6.505 2.895 ;
      RECT 6.355 2.591 6.485 2.924 ;
      RECT 6.375 2.586 6.475 2.943 ;
      RECT 5.835 2.72 6.025 2.895 ;
      RECT 5.795 2.638 5.985 2.89 ;
      RECT 5.761 2.643 5.985 2.884 ;
      RECT 5.675 2.65 5.985 2.879 ;
      RECT 5.591 2.665 5.985 2.874 ;
      RECT 5.505 2.685 6.015 2.868 ;
      RECT 5.591 2.675 6.015 2.874 ;
      RECT 5.835 2.635 5.985 2.895 ;
      RECT 5.835 2.631 5.935 2.895 ;
      RECT 5.921 2.626 5.935 2.895 ;
      RECT 4.675 1.954 5.335 2.345 ;
      RECT 4.933 1.948 5.335 2.345 ;
      RECT 4.665 1.96 5.335 2.344 ;
      RECT 4.655 1.975 5.335 2.343 ;
      RECT 4.595 2.015 5.335 2.339 ;
      RECT 4.761 1.953 5.345 2.335 ;
      RECT 4.665 1.96 5.355 2.325 ;
      RECT 4.665 1.968 5.365 2.305 ;
      RECT 4.655 1.978 5.385 2.278 ;
      RECT 4.595 2.015 5.395 2.253 ;
      RECT 4.655 1.985 5.405 2.24 ;
      RECT 4.761 1.951 5.335 2.345 ;
      RECT 4.847 1.949 5.335 2.345 ;
      RECT 4.933 1.947 5.315 2.345 ;
      RECT 5.019 1.945 5.315 2.345 ;
      RECT 5.185 3.12 5.355 3.315 ;
      RECT 5.175 3.12 5.355 3.26 ;
      RECT 5.17 3.12 5.355 3.188 ;
      RECT 5.155 3.06 5.335 3.155 ;
      RECT 5.145 3.06 5.335 3.105 ;
      RECT 5.115 3.035 5.325 3.06 ;
      RECT 5.095 3.035 5.325 3.045 ;
      RECT 5.035 2.725 5.215 3.036 ;
      RECT 5.035 2.96 5.315 3.036 ;
      RECT 5.025 2.724 5.035 3.026 ;
      RECT 5.005 2.723 5.025 3.02 ;
      RECT 4.975 2.722 5.005 3 ;
      RECT 4.925 2.719 4.975 2.965 ;
      RECT 4.925 2.84 5.285 2.965 ;
      RECT 4.855 2.716 4.925 2.92 ;
      RECT 4.855 2.775 5.265 2.92 ;
      RECT 4.855 2.765 5.255 2.92 ;
      RECT 4.855 2.755 5.245 2.92 ;
      RECT 4.855 2.735 5.225 2.92 ;
      RECT 4.935 3.255 4.945 3.512 ;
      RECT 4.915 3.172 4.935 3.532 ;
      RECT 4.895 3.166 4.915 3.56 ;
      RECT 4.835 3.154 4.895 3.58 ;
      RECT 4.795 3.14 4.835 3.581 ;
      RECT 4.711 3.129 4.795 3.569 ;
      RECT 4.625 3.116 4.711 3.553 ;
      RECT 4.615 3.109 4.625 3.545 ;
      RECT 4.565 3.106 4.615 3.485 ;
      RECT 4.545 3.102 4.565 3.4 ;
      RECT 4.535 3.1 4.545 3.35 ;
      RECT 4.505 3.098 4.535 3.32 ;
      RECT 4.465 3.093 4.505 3.3 ;
      RECT 4.427 3.088 4.465 3.288 ;
      RECT 4.341 3.08 4.427 3.297 ;
      RECT 4.255 3.069 4.341 3.309 ;
      RECT 4.185 3.059 4.255 3.319 ;
      RECT 4.165 3.05 4.185 3.324 ;
      RECT 4.105 3.022 4.165 3.32 ;
      RECT 4.085 2.992 4.105 3.308 ;
      RECT 4.065 2.965 4.085 3.295 ;
      RECT 3.985 2.718 4.065 3.262 ;
      RECT 3.971 2.71 3.985 3.224 ;
      RECT 3.885 2.702 3.971 3.145 ;
      RECT 3.865 2.693 3.885 3.061 ;
      RECT 3.835 2.688 3.865 3.041 ;
      RECT 3.765 2.699 3.835 3.026 ;
      RECT 3.745 2.717 3.765 3 ;
      RECT 3.735 2.723 3.745 2.945 ;
      RECT 3.715 2.745 3.735 2.83 ;
      RECT 4.375 2.705 4.545 2.895 ;
      RECT 4.375 2.705 4.575 2.89 ;
      RECT 4.425 2.615 4.595 2.88 ;
      RECT 4.385 2.65 4.595 2.88 ;
      RECT 3.585 3.388 3.655 3.829 ;
      RECT 3.525 3.413 3.655 3.826 ;
      RECT 3.525 3.413 3.705 3.819 ;
      RECT 3.515 3.435 3.705 3.816 ;
      RECT 3.655 3.375 3.725 3.814 ;
      RECT 3.585 3.4 3.805 3.811 ;
      RECT 3.515 3.439 3.855 3.807 ;
      RECT 3.495 3.465 3.855 3.795 ;
      RECT 3.515 3.459 3.875 3.79 ;
      RECT 3.495 2.205 3.535 2.445 ;
      RECT 3.495 2.205 3.565 2.444 ;
      RECT 3.495 2.205 3.675 2.436 ;
      RECT 3.495 2.205 3.735 2.415 ;
      RECT 3.505 2.15 3.785 2.315 ;
      RECT 3.615 1.99 3.645 2.437 ;
      RECT 3.645 1.985 3.825 2.195 ;
      RECT 3.515 2.125 3.825 2.195 ;
      RECT 3.565 2.02 3.615 2.44 ;
      RECT 3.535 2.075 3.825 2.195 ;
      RECT 1.33 7.855 1.5 8.305 ;
      RECT 1.385 6.075 1.555 8.025 ;
      RECT 1.33 5.015 1.5 6.245 ;
      RECT 0.81 5.015 0.98 8.305 ;
      RECT 0.81 7.315 1.215 7.645 ;
      RECT 0.81 6.475 1.215 6.805 ;
      RECT 92.03 7.8 92.2 8.31 ;
      RECT 91.04 0.57 91.21 1.08 ;
      RECT 91.04 2.39 91.21 3.86 ;
      RECT 91.04 5.02 91.21 6.49 ;
      RECT 91.04 7.8 91.21 8.31 ;
      RECT 89.68 0.575 89.85 3.865 ;
      RECT 89.68 5.015 89.85 8.305 ;
      RECT 89.25 0.575 89.42 1.085 ;
      RECT 89.25 1.655 89.42 3.865 ;
      RECT 89.25 5.015 89.42 7.225 ;
      RECT 89.25 7.795 89.42 8.305 ;
      RECT 84.92 5.015 85.09 8.305 ;
      RECT 84.49 5.015 84.66 7.225 ;
      RECT 84.49 7.795 84.66 8.305 ;
      RECT 74.105 7.8 74.275 8.31 ;
      RECT 73.115 0.57 73.285 1.08 ;
      RECT 73.115 2.39 73.285 3.86 ;
      RECT 73.115 5.02 73.285 6.49 ;
      RECT 73.115 7.8 73.285 8.31 ;
      RECT 71.755 0.575 71.925 3.865 ;
      RECT 71.755 5.015 71.925 8.305 ;
      RECT 71.325 0.575 71.495 1.085 ;
      RECT 71.325 1.655 71.495 3.865 ;
      RECT 71.325 5.015 71.495 7.225 ;
      RECT 71.325 7.795 71.495 8.305 ;
      RECT 66.995 5.015 67.165 8.305 ;
      RECT 66.565 5.015 66.735 7.225 ;
      RECT 66.565 7.795 66.735 8.305 ;
      RECT 56.18 7.8 56.35 8.31 ;
      RECT 55.19 0.57 55.36 1.08 ;
      RECT 55.19 2.39 55.36 3.86 ;
      RECT 55.19 5.02 55.36 6.49 ;
      RECT 55.19 7.8 55.36 8.31 ;
      RECT 53.83 0.575 54 3.865 ;
      RECT 53.83 5.015 54 8.305 ;
      RECT 53.4 0.575 53.57 1.085 ;
      RECT 53.4 1.655 53.57 3.865 ;
      RECT 53.4 5.015 53.57 7.225 ;
      RECT 53.4 7.795 53.57 8.305 ;
      RECT 49.07 5.015 49.24 8.305 ;
      RECT 48.64 5.015 48.81 7.225 ;
      RECT 48.64 7.795 48.81 8.305 ;
      RECT 38.255 7.8 38.425 8.31 ;
      RECT 37.265 0.57 37.435 1.08 ;
      RECT 37.265 2.39 37.435 3.86 ;
      RECT 37.265 5.02 37.435 6.49 ;
      RECT 37.265 7.8 37.435 8.31 ;
      RECT 35.905 0.575 36.075 3.865 ;
      RECT 35.905 5.015 36.075 8.305 ;
      RECT 35.475 0.575 35.645 1.085 ;
      RECT 35.475 1.655 35.645 3.865 ;
      RECT 35.475 5.015 35.645 7.225 ;
      RECT 35.475 7.795 35.645 8.305 ;
      RECT 31.145 5.015 31.315 8.305 ;
      RECT 30.715 5.015 30.885 7.225 ;
      RECT 30.715 7.795 30.885 8.305 ;
      RECT 20.33 7.8 20.5 8.31 ;
      RECT 19.34 0.57 19.51 1.08 ;
      RECT 19.34 2.39 19.51 3.86 ;
      RECT 19.34 5.02 19.51 6.49 ;
      RECT 19.34 7.8 19.51 8.31 ;
      RECT 17.98 0.575 18.15 3.865 ;
      RECT 17.98 5.015 18.15 8.305 ;
      RECT 17.55 0.575 17.72 1.085 ;
      RECT 17.55 1.655 17.72 3.865 ;
      RECT 17.55 5.015 17.72 7.225 ;
      RECT 17.55 7.795 17.72 8.305 ;
      RECT 13.22 5.015 13.39 8.305 ;
      RECT 12.79 5.015 12.96 7.225 ;
      RECT 12.79 7.795 12.96 8.305 ;
      RECT 1.76 5.015 1.93 7.225 ;
      RECT 1.76 7.795 1.93 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r1 ;
  SIZE 85.755 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 18.85 2.395 19.02 2.565 ;
        RECT 18.845 2.39 19.015 2.56 ;
        RECT 18.845 0.91 19.015 1.08 ;
      LAYER li1 ;
        RECT 18.845 2.395 19.02 2.565 ;
        RECT 18.845 2.39 19.015 3.86 ;
        RECT 18.845 0.57 19.015 1.08 ;
      LAYER met1 ;
        RECT 18.785 2.36 19.075 2.59 ;
        RECT 18.785 0.88 19.075 1.11 ;
        RECT 18.845 0.88 19.015 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 35.435 2.395 35.605 2.565 ;
        RECT 35.43 2.39 35.6 2.56 ;
        RECT 35.43 0.91 35.6 1.08 ;
      LAYER li1 ;
        RECT 35.43 2.395 35.605 2.565 ;
        RECT 35.43 2.39 35.6 3.86 ;
        RECT 35.43 0.57 35.6 1.08 ;
      LAYER met1 ;
        RECT 35.37 2.36 35.66 2.59 ;
        RECT 35.37 0.88 35.66 1.11 ;
        RECT 35.43 0.88 35.6 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 52.02 2.395 52.19 2.565 ;
        RECT 52.015 2.39 52.185 2.56 ;
        RECT 52.015 0.91 52.185 1.08 ;
      LAYER li1 ;
        RECT 52.015 2.395 52.19 2.565 ;
        RECT 52.015 2.39 52.185 3.86 ;
        RECT 52.015 0.57 52.185 1.08 ;
      LAYER met1 ;
        RECT 51.955 2.36 52.245 2.59 ;
        RECT 51.955 0.88 52.245 1.11 ;
        RECT 52.015 0.88 52.185 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 68.605 2.395 68.775 2.565 ;
        RECT 68.6 2.39 68.77 2.56 ;
        RECT 68.6 0.91 68.77 1.08 ;
      LAYER li1 ;
        RECT 68.6 2.395 68.775 2.565 ;
        RECT 68.6 2.39 68.77 3.86 ;
        RECT 68.6 0.57 68.77 1.08 ;
      LAYER met1 ;
        RECT 68.54 2.36 68.83 2.59 ;
        RECT 68.54 0.88 68.83 1.11 ;
        RECT 68.6 0.88 68.77 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 85.185 2.395 85.355 2.565 ;
        RECT 85.18 2.39 85.35 2.56 ;
        RECT 85.18 0.91 85.35 1.08 ;
      LAYER li1 ;
        RECT 85.18 2.395 85.355 2.565 ;
        RECT 85.18 2.39 85.35 3.86 ;
        RECT 85.18 0.57 85.35 1.08 ;
      LAYER met1 ;
        RECT 85.12 2.36 85.41 2.59 ;
        RECT 85.12 0.88 85.41 1.11 ;
        RECT 85.18 0.88 85.35 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 14.695 1.66 14.865 2.935 ;
        RECT 14.695 5.945 14.865 7.22 ;
        RECT 3.47 5.945 3.64 7.22 ;
      LAYER met2 ;
        RECT 14.62 5.865 14.945 6.19 ;
        RECT 14.615 3.635 14.94 3.96 ;
        RECT 5.775 7.885 14.86 8.055 ;
        RECT 14.685 3.635 14.86 8.055 ;
        RECT 5.72 5.86 6 6.2 ;
        RECT 5.775 5.86 5.945 8.055 ;
      LAYER met1 ;
        RECT 14.635 2.765 15.095 2.935 ;
        RECT 14.615 3.635 14.94 3.96 ;
        RECT 14.635 2.735 14.925 2.965 ;
        RECT 14.69 2.735 14.87 3.96 ;
        RECT 14.62 5.945 15.095 6.115 ;
        RECT 14.62 5.865 14.945 6.19 ;
        RECT 5.69 5.89 6.03 6.17 ;
        RECT 3.41 5.945 6.03 6.115 ;
        RECT 3.41 5.915 3.7 6.145 ;
      LAYER mcon ;
        RECT 3.47 5.945 3.64 6.115 ;
        RECT 14.695 5.945 14.865 6.115 ;
        RECT 14.695 2.765 14.865 2.935 ;
      LAYER via1 ;
        RECT 5.785 5.955 5.935 6.105 ;
        RECT 14.705 3.72 14.855 3.87 ;
        RECT 14.71 5.95 14.86 6.1 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 31.28 1.66 31.45 2.935 ;
        RECT 31.28 5.945 31.45 7.22 ;
        RECT 20.055 5.945 20.225 7.22 ;
      LAYER met2 ;
        RECT 31.205 5.865 31.53 6.19 ;
        RECT 31.2 3.635 31.525 3.96 ;
        RECT 22.36 7.885 31.445 8.055 ;
        RECT 31.27 3.635 31.445 8.055 ;
        RECT 22.305 5.86 22.585 6.2 ;
        RECT 22.36 5.86 22.53 8.055 ;
      LAYER met1 ;
        RECT 31.22 2.765 31.68 2.935 ;
        RECT 31.2 3.635 31.525 3.96 ;
        RECT 31.22 2.735 31.51 2.965 ;
        RECT 31.275 2.735 31.455 3.96 ;
        RECT 31.205 5.945 31.68 6.115 ;
        RECT 31.205 5.865 31.53 6.19 ;
        RECT 22.275 5.89 22.615 6.17 ;
        RECT 19.995 5.945 22.615 6.115 ;
        RECT 19.995 5.915 20.285 6.145 ;
      LAYER mcon ;
        RECT 20.055 5.945 20.225 6.115 ;
        RECT 31.28 5.945 31.45 6.115 ;
        RECT 31.28 2.765 31.45 2.935 ;
      LAYER via1 ;
        RECT 22.37 5.955 22.52 6.105 ;
        RECT 31.29 3.72 31.44 3.87 ;
        RECT 31.295 5.95 31.445 6.1 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 47.865 1.66 48.035 2.935 ;
        RECT 47.865 5.945 48.035 7.22 ;
        RECT 36.64 5.945 36.81 7.22 ;
      LAYER met2 ;
        RECT 47.79 5.865 48.115 6.19 ;
        RECT 47.785 3.635 48.11 3.96 ;
        RECT 38.945 7.885 48.03 8.055 ;
        RECT 47.855 3.635 48.03 8.055 ;
        RECT 38.89 5.86 39.17 6.2 ;
        RECT 38.945 5.86 39.115 8.055 ;
      LAYER met1 ;
        RECT 47.805 2.765 48.265 2.935 ;
        RECT 47.785 3.635 48.11 3.96 ;
        RECT 47.805 2.735 48.095 2.965 ;
        RECT 47.86 2.735 48.04 3.96 ;
        RECT 47.79 5.945 48.265 6.115 ;
        RECT 47.79 5.865 48.115 6.19 ;
        RECT 38.86 5.89 39.2 6.17 ;
        RECT 36.58 5.945 39.2 6.115 ;
        RECT 36.58 5.915 36.87 6.145 ;
      LAYER mcon ;
        RECT 36.64 5.945 36.81 6.115 ;
        RECT 47.865 5.945 48.035 6.115 ;
        RECT 47.865 2.765 48.035 2.935 ;
      LAYER via1 ;
        RECT 38.955 5.955 39.105 6.105 ;
        RECT 47.875 3.72 48.025 3.87 ;
        RECT 47.88 5.95 48.03 6.1 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 64.45 1.66 64.62 2.935 ;
        RECT 64.45 5.945 64.62 7.22 ;
        RECT 53.225 5.945 53.395 7.22 ;
      LAYER met2 ;
        RECT 64.375 5.865 64.7 6.19 ;
        RECT 64.37 3.635 64.695 3.96 ;
        RECT 55.53 7.885 64.615 8.055 ;
        RECT 64.44 3.635 64.615 8.055 ;
        RECT 55.475 5.86 55.755 6.2 ;
        RECT 55.53 5.86 55.7 8.055 ;
      LAYER met1 ;
        RECT 64.39 2.765 64.85 2.935 ;
        RECT 64.37 3.635 64.695 3.96 ;
        RECT 64.39 2.735 64.68 2.965 ;
        RECT 64.445 2.735 64.625 3.96 ;
        RECT 64.375 5.945 64.85 6.115 ;
        RECT 64.375 5.865 64.7 6.19 ;
        RECT 55.445 5.89 55.785 6.17 ;
        RECT 53.165 5.945 55.785 6.115 ;
        RECT 53.165 5.915 53.455 6.145 ;
      LAYER mcon ;
        RECT 53.225 5.945 53.395 6.115 ;
        RECT 64.45 5.945 64.62 6.115 ;
        RECT 64.45 2.765 64.62 2.935 ;
      LAYER via1 ;
        RECT 55.54 5.955 55.69 6.105 ;
        RECT 64.46 3.72 64.61 3.87 ;
        RECT 64.465 5.95 64.615 6.1 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 81.03 1.66 81.2 2.935 ;
        RECT 81.03 5.945 81.2 7.22 ;
        RECT 69.805 5.945 69.975 7.22 ;
      LAYER met2 ;
        RECT 80.955 5.865 81.28 6.19 ;
        RECT 80.95 3.635 81.275 3.96 ;
        RECT 72.11 7.885 81.195 8.055 ;
        RECT 81.02 3.635 81.195 8.055 ;
        RECT 72.055 5.86 72.335 6.2 ;
        RECT 72.11 5.86 72.28 8.055 ;
      LAYER met1 ;
        RECT 80.97 2.765 81.43 2.935 ;
        RECT 80.95 3.635 81.275 3.96 ;
        RECT 80.97 2.735 81.26 2.965 ;
        RECT 81.025 2.735 81.205 3.96 ;
        RECT 80.955 5.945 81.43 6.115 ;
        RECT 80.955 5.865 81.28 6.19 ;
        RECT 72.025 5.89 72.365 6.17 ;
        RECT 69.745 5.945 72.365 6.115 ;
        RECT 69.745 5.915 70.035 6.145 ;
      LAYER mcon ;
        RECT 69.805 5.945 69.975 6.115 ;
        RECT 81.03 5.945 81.2 6.115 ;
        RECT 81.03 2.765 81.2 2.935 ;
      LAYER via1 ;
        RECT 72.12 5.955 72.27 6.105 ;
        RECT 81.04 3.72 81.19 3.87 ;
        RECT 81.045 5.95 81.195 6.1 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.24 5.945 0.41 7.22 ;
      LAYER met1 ;
        RECT 0.18 5.945 0.64 6.115 ;
        RECT 0.18 5.915 0.47 6.145 ;
      LAYER mcon ;
        RECT 0.24 5.945 0.41 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.33 4.255 2.135 4.635 ;
      LAYER li1 ;
        RECT 79.785 4.135 85.725 4.745 ;
        RECT 83.59 4.13 85.57 4.75 ;
        RECT 84.75 3.4 84.92 5.48 ;
        RECT 83.76 3.4 83.93 5.48 ;
        RECT 81.02 3.405 81.19 5.475 ;
        RECT 79.655 4.135 85.725 4.67 ;
        RECT 79.325 3.2 79.655 4.515 ;
        RECT 72.855 4.34 85.725 4.515 ;
        RECT 77.585 3.8 77.845 4.515 ;
        RECT 77.025 4.34 77.395 4.89 ;
        RECT 76.585 3.42 76.915 3.66 ;
        RECT 76.585 3.42 76.775 3.79 ;
        RECT 76.155 3.69 76.765 4.515 ;
        RECT 76.205 3.69 76.475 5.29 ;
        RECT 75.285 3.8 75.505 4.515 ;
        RECT 75.045 4.34 75.325 5.18 ;
        RECT 74.275 3.47 74.605 3.66 ;
        RECT 73.855 3.84 74.475 4.515 ;
        RECT 74.275 3.47 74.475 4.515 ;
        RECT 74.045 3.84 74.375 5.23 ;
        RECT 72.935 3.83 73.195 4.515 ;
        RECT 1.795 4.345 85.725 4.515 ;
        RECT 69.14 4.13 72.715 4.74 ;
        RECT 69.62 4.13 72.37 4.745 ;
        RECT 69.795 4.13 69.965 5.475 ;
        RECT 63.205 4.135 69.145 4.745 ;
        RECT 67.01 4.13 68.99 4.75 ;
        RECT 68.17 3.4 68.34 5.48 ;
        RECT 67.18 3.4 67.35 5.48 ;
        RECT 64.44 3.405 64.61 5.475 ;
        RECT 63.075 4.135 72.715 4.67 ;
        RECT 62.745 3.2 63.075 4.515 ;
        RECT 56.275 4.34 72.715 4.515 ;
        RECT 61.005 3.8 61.265 4.515 ;
        RECT 60.445 4.34 60.815 4.89 ;
        RECT 60.005 3.42 60.335 3.66 ;
        RECT 60.005 3.42 60.195 3.79 ;
        RECT 59.575 3.69 60.185 4.515 ;
        RECT 59.625 3.69 59.895 5.29 ;
        RECT 58.705 3.8 58.925 4.515 ;
        RECT 58.465 4.34 58.745 5.18 ;
        RECT 57.695 3.47 58.025 3.66 ;
        RECT 57.275 3.84 57.895 4.515 ;
        RECT 57.695 3.47 57.895 4.515 ;
        RECT 57.465 3.84 57.795 5.23 ;
        RECT 56.355 3.83 56.615 4.515 ;
        RECT 52.56 4.13 56.135 4.74 ;
        RECT 53.04 4.13 55.79 4.745 ;
        RECT 53.215 4.13 53.385 5.475 ;
        RECT 46.62 4.135 52.56 4.745 ;
        RECT 50.425 4.13 52.405 4.75 ;
        RECT 51.585 3.4 51.755 5.48 ;
        RECT 50.595 3.4 50.765 5.48 ;
        RECT 47.855 3.405 48.025 5.475 ;
        RECT 46.49 4.135 56.135 4.67 ;
        RECT 46.16 3.2 46.49 4.515 ;
        RECT 39.69 4.34 56.135 4.515 ;
        RECT 44.42 3.8 44.68 4.515 ;
        RECT 43.86 4.34 44.23 4.89 ;
        RECT 43.42 3.42 43.75 3.66 ;
        RECT 43.42 3.42 43.61 3.79 ;
        RECT 42.99 3.69 43.6 4.515 ;
        RECT 43.04 3.69 43.31 5.29 ;
        RECT 42.12 3.8 42.34 4.515 ;
        RECT 41.88 4.34 42.16 5.18 ;
        RECT 41.11 3.47 41.44 3.66 ;
        RECT 40.69 3.84 41.31 4.515 ;
        RECT 41.11 3.47 41.31 4.515 ;
        RECT 40.88 3.84 41.21 5.23 ;
        RECT 39.77 3.83 40.03 4.515 ;
        RECT 35.975 4.13 39.55 4.74 ;
        RECT 36.455 4.13 39.205 4.745 ;
        RECT 36.63 4.13 36.8 5.475 ;
        RECT 30.035 4.135 35.975 4.745 ;
        RECT 33.84 4.13 35.82 4.75 ;
        RECT 35 3.4 35.17 5.48 ;
        RECT 34.01 3.4 34.18 5.48 ;
        RECT 31.27 3.405 31.44 5.475 ;
        RECT 29.905 4.135 39.55 4.67 ;
        RECT 29.575 3.2 29.905 4.515 ;
        RECT 23.105 4.34 39.55 4.515 ;
        RECT 27.835 3.8 28.095 4.515 ;
        RECT 27.275 4.34 27.645 4.89 ;
        RECT 26.835 3.42 27.165 3.66 ;
        RECT 26.835 3.42 27.025 3.79 ;
        RECT 26.405 3.69 27.015 4.515 ;
        RECT 26.455 3.69 26.725 5.29 ;
        RECT 25.535 3.8 25.755 4.515 ;
        RECT 25.295 4.34 25.575 5.18 ;
        RECT 24.525 3.47 24.855 3.66 ;
        RECT 24.105 3.84 24.725 4.515 ;
        RECT 24.525 3.47 24.725 4.515 ;
        RECT 24.295 3.84 24.625 5.23 ;
        RECT 23.185 3.83 23.445 4.515 ;
        RECT 19.39 4.13 22.965 4.74 ;
        RECT 19.87 4.13 22.62 4.745 ;
        RECT 20.045 4.13 20.215 5.475 ;
        RECT 13.45 4.135 19.39 4.745 ;
        RECT 17.255 4.13 19.235 4.75 ;
        RECT 18.415 3.4 18.585 5.48 ;
        RECT 17.425 3.4 17.595 5.48 ;
        RECT 14.685 3.405 14.855 5.475 ;
        RECT 13.32 4.135 22.965 4.67 ;
        RECT 12.99 3.2 13.32 4.515 ;
        RECT 6.52 4.34 22.965 4.515 ;
        RECT 11.25 3.8 11.51 4.515 ;
        RECT 10.69 4.34 11.06 4.89 ;
        RECT 10.25 3.42 10.58 3.66 ;
        RECT 10.25 3.42 10.44 3.79 ;
        RECT 9.82 3.69 10.43 4.515 ;
        RECT 9.87 3.69 10.14 5.29 ;
        RECT 8.95 3.8 9.17 4.515 ;
        RECT 8.71 4.34 8.99 5.18 ;
        RECT 7.94 3.47 8.27 3.66 ;
        RECT 7.52 3.84 8.14 4.515 ;
        RECT 7.94 3.47 8.14 4.515 ;
        RECT 7.71 3.84 8.04 5.23 ;
        RECT 6.6 3.83 6.86 4.515 ;
        RECT 1.795 4.13 6.38 4.74 ;
        RECT 3.285 4.13 6.035 4.745 ;
        RECT 3.46 4.13 3.63 5.475 ;
        RECT 0 4.44 2.805 4.745 ;
        RECT 2.04 4.13 2.21 8.305 ;
        RECT 0 4.13 6.38 4.33 ;
        RECT 0 4.13 1.625 4.745 ;
        RECT 0.23 4.13 0.4 5.475 ;
      LAYER met2 ;
        RECT 1.52 4.255 1.9 4.635 ;
      LAYER met1 ;
        RECT 79.785 4.15 85.725 4.745 ;
        RECT 80.245 4.135 85.725 4.745 ;
        RECT 83.59 4.13 85.57 4.75 ;
        RECT 0 4.19 85.725 4.67 ;
        RECT 79.655 4.15 85.725 4.67 ;
        RECT 69.14 4.13 72.715 4.74 ;
        RECT 69.62 4.13 72.37 4.745 ;
        RECT 63.205 4.15 69.145 4.745 ;
        RECT 63.665 4.135 72.715 4.74 ;
        RECT 67.01 4.13 68.99 4.75 ;
        RECT 63.075 4.15 72.715 4.67 ;
        RECT 52.56 4.13 56.135 4.74 ;
        RECT 53.04 4.13 55.79 4.745 ;
        RECT 46.62 4.15 52.56 4.745 ;
        RECT 47.08 4.135 56.135 4.74 ;
        RECT 50.425 4.13 52.405 4.75 ;
        RECT 46.49 4.15 56.135 4.67 ;
        RECT 35.975 4.13 39.55 4.74 ;
        RECT 36.455 4.13 39.205 4.745 ;
        RECT 30.035 4.15 35.975 4.745 ;
        RECT 30.495 4.135 39.55 4.74 ;
        RECT 33.84 4.13 35.82 4.75 ;
        RECT 29.905 4.15 39.55 4.67 ;
        RECT 19.39 4.13 22.965 4.74 ;
        RECT 19.87 4.13 22.62 4.745 ;
        RECT 13.45 4.15 19.39 4.745 ;
        RECT 13.91 4.135 22.965 4.74 ;
        RECT 17.255 4.13 19.235 4.75 ;
        RECT 13.32 4.15 22.965 4.67 ;
        RECT 0 4.13 6.38 4.74 ;
        RECT 3.285 4.13 6.035 4.745 ;
        RECT 0 4.13 2.805 4.745 ;
        RECT 1.98 6.655 2.27 6.885 ;
        RECT 1.81 6.685 2.27 6.855 ;
      LAYER via2 ;
        RECT 1.61 4.345 1.81 4.545 ;
      LAYER mcon ;
        RECT 2.04 6.685 2.21 6.855 ;
        RECT 2.35 4.545 2.52 4.715 ;
        RECT 5.58 4.545 5.75 4.715 ;
        RECT 6.66 4.34 6.83 4.51 ;
        RECT 7.12 4.34 7.29 4.51 ;
        RECT 7.58 4.34 7.75 4.51 ;
        RECT 8.04 4.34 8.21 4.51 ;
        RECT 8.5 4.34 8.67 4.51 ;
        RECT 8.96 4.34 9.13 4.51 ;
        RECT 9.42 4.34 9.59 4.51 ;
        RECT 9.88 4.34 10.05 4.51 ;
        RECT 10.34 4.34 10.51 4.51 ;
        RECT 10.8 4.34 10.97 4.51 ;
        RECT 11.26 4.34 11.43 4.51 ;
        RECT 11.72 4.34 11.89 4.51 ;
        RECT 12.18 4.34 12.35 4.51 ;
        RECT 12.64 4.34 12.81 4.51 ;
        RECT 13.1 4.34 13.27 4.51 ;
        RECT 16.805 4.545 16.975 4.715 ;
        RECT 16.805 4.165 16.975 4.335 ;
        RECT 17.505 4.55 17.675 4.72 ;
        RECT 17.505 4.16 17.675 4.33 ;
        RECT 18.495 4.55 18.665 4.72 ;
        RECT 18.495 4.16 18.665 4.33 ;
        RECT 22.165 4.545 22.335 4.715 ;
        RECT 23.245 4.34 23.415 4.51 ;
        RECT 23.705 4.34 23.875 4.51 ;
        RECT 24.165 4.34 24.335 4.51 ;
        RECT 24.625 4.34 24.795 4.51 ;
        RECT 25.085 4.34 25.255 4.51 ;
        RECT 25.545 4.34 25.715 4.51 ;
        RECT 26.005 4.34 26.175 4.51 ;
        RECT 26.465 4.34 26.635 4.51 ;
        RECT 26.925 4.34 27.095 4.51 ;
        RECT 27.385 4.34 27.555 4.51 ;
        RECT 27.845 4.34 28.015 4.51 ;
        RECT 28.305 4.34 28.475 4.51 ;
        RECT 28.765 4.34 28.935 4.51 ;
        RECT 29.225 4.34 29.395 4.51 ;
        RECT 29.685 4.34 29.855 4.51 ;
        RECT 33.39 4.545 33.56 4.715 ;
        RECT 33.39 4.165 33.56 4.335 ;
        RECT 34.09 4.55 34.26 4.72 ;
        RECT 34.09 4.16 34.26 4.33 ;
        RECT 35.08 4.55 35.25 4.72 ;
        RECT 35.08 4.16 35.25 4.33 ;
        RECT 38.75 4.545 38.92 4.715 ;
        RECT 39.83 4.34 40 4.51 ;
        RECT 40.29 4.34 40.46 4.51 ;
        RECT 40.75 4.34 40.92 4.51 ;
        RECT 41.21 4.34 41.38 4.51 ;
        RECT 41.67 4.34 41.84 4.51 ;
        RECT 42.13 4.34 42.3 4.51 ;
        RECT 42.59 4.34 42.76 4.51 ;
        RECT 43.05 4.34 43.22 4.51 ;
        RECT 43.51 4.34 43.68 4.51 ;
        RECT 43.97 4.34 44.14 4.51 ;
        RECT 44.43 4.34 44.6 4.51 ;
        RECT 44.89 4.34 45.06 4.51 ;
        RECT 45.35 4.34 45.52 4.51 ;
        RECT 45.81 4.34 45.98 4.51 ;
        RECT 46.27 4.34 46.44 4.51 ;
        RECT 49.975 4.545 50.145 4.715 ;
        RECT 49.975 4.165 50.145 4.335 ;
        RECT 50.675 4.55 50.845 4.72 ;
        RECT 50.675 4.16 50.845 4.33 ;
        RECT 51.665 4.55 51.835 4.72 ;
        RECT 51.665 4.16 51.835 4.33 ;
        RECT 55.335 4.545 55.505 4.715 ;
        RECT 56.415 4.34 56.585 4.51 ;
        RECT 56.875 4.34 57.045 4.51 ;
        RECT 57.335 4.34 57.505 4.51 ;
        RECT 57.795 4.34 57.965 4.51 ;
        RECT 58.255 4.34 58.425 4.51 ;
        RECT 58.715 4.34 58.885 4.51 ;
        RECT 59.175 4.34 59.345 4.51 ;
        RECT 59.635 4.34 59.805 4.51 ;
        RECT 60.095 4.34 60.265 4.51 ;
        RECT 60.555 4.34 60.725 4.51 ;
        RECT 61.015 4.34 61.185 4.51 ;
        RECT 61.475 4.34 61.645 4.51 ;
        RECT 61.935 4.34 62.105 4.51 ;
        RECT 62.395 4.34 62.565 4.51 ;
        RECT 62.855 4.34 63.025 4.51 ;
        RECT 66.56 4.545 66.73 4.715 ;
        RECT 66.56 4.165 66.73 4.335 ;
        RECT 67.26 4.55 67.43 4.72 ;
        RECT 67.26 4.16 67.43 4.33 ;
        RECT 68.25 4.55 68.42 4.72 ;
        RECT 68.25 4.16 68.42 4.33 ;
        RECT 71.915 4.545 72.085 4.715 ;
        RECT 72.995 4.34 73.165 4.51 ;
        RECT 73.455 4.34 73.625 4.51 ;
        RECT 73.915 4.34 74.085 4.51 ;
        RECT 74.375 4.34 74.545 4.51 ;
        RECT 74.835 4.34 75.005 4.51 ;
        RECT 75.295 4.34 75.465 4.51 ;
        RECT 75.755 4.34 75.925 4.51 ;
        RECT 76.215 4.34 76.385 4.51 ;
        RECT 76.675 4.34 76.845 4.51 ;
        RECT 77.135 4.34 77.305 4.51 ;
        RECT 77.595 4.34 77.765 4.51 ;
        RECT 78.055 4.34 78.225 4.51 ;
        RECT 78.515 4.34 78.685 4.51 ;
        RECT 78.975 4.34 79.145 4.51 ;
        RECT 79.435 4.34 79.605 4.51 ;
        RECT 83.14 4.545 83.31 4.715 ;
        RECT 83.14 4.165 83.31 4.335 ;
        RECT 83.84 4.55 84.01 4.72 ;
        RECT 83.84 4.16 84.01 4.33 ;
        RECT 84.83 4.55 85 4.72 ;
        RECT 84.83 4.16 85 4.33 ;
      LAYER via1 ;
        RECT 1.635 4.37 1.785 4.52 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 75.225 6.47 75.555 6.8 ;
        RECT 75.195 6.49 75.495 6.9 ;
        RECT 74.755 6.49 75.555 6.79 ;
        RECT 58.645 6.47 58.975 6.8 ;
        RECT 58.615 6.49 58.915 6.9 ;
        RECT 58.175 6.49 58.975 6.79 ;
        RECT 42.06 6.47 42.39 6.8 ;
        RECT 42.03 6.49 42.33 6.9 ;
        RECT 41.59 6.49 42.39 6.79 ;
        RECT 25.475 6.47 25.805 6.8 ;
        RECT 25.445 6.49 25.745 6.9 ;
        RECT 25.005 6.49 25.805 6.79 ;
        RECT 8.89 6.47 9.22 6.8 ;
        RECT 8.86 6.49 9.16 6.9 ;
        RECT 8.42 6.49 9.22 6.79 ;
        RECT 0 0 0.805 0.38 ;
        RECT 0 8.5 0.805 8.88 ;
      LAYER li1 ;
        RECT 0 8.57 85.755 8.88 ;
        RECT 84.75 7.95 84.92 8.88 ;
        RECT 83.76 7.95 83.93 8.88 ;
        RECT 81.02 7.945 81.19 8.88 ;
        RECT 72.56 7.18 79.76 8.88 ;
        RECT 72.855 7.06 79.755 8.88 ;
        RECT 78.285 6.55 78.735 8.88 ;
        RECT 76.195 6.66 76.525 8.88 ;
        RECT 74.125 6.6 74.375 8.88 ;
        RECT 69.795 7.945 69.965 8.88 ;
        RECT 68.17 7.95 68.34 8.88 ;
        RECT 67.18 7.95 67.35 8.88 ;
        RECT 64.44 7.945 64.61 8.88 ;
        RECT 55.98 7.18 63.18 8.88 ;
        RECT 56.275 7.06 63.175 8.88 ;
        RECT 61.705 6.55 62.155 8.88 ;
        RECT 59.615 6.66 59.945 8.88 ;
        RECT 57.545 6.6 57.795 8.88 ;
        RECT 53.215 7.945 53.385 8.88 ;
        RECT 51.585 7.95 51.755 8.88 ;
        RECT 50.595 7.95 50.765 8.88 ;
        RECT 47.855 7.945 48.025 8.88 ;
        RECT 39.395 7.18 46.595 8.88 ;
        RECT 39.69 7.06 46.59 8.88 ;
        RECT 45.12 6.55 45.57 8.88 ;
        RECT 43.03 6.66 43.36 8.88 ;
        RECT 40.96 6.6 41.21 8.88 ;
        RECT 36.63 7.945 36.8 8.88 ;
        RECT 35 7.95 35.17 8.88 ;
        RECT 34.01 7.95 34.18 8.88 ;
        RECT 31.27 7.945 31.44 8.88 ;
        RECT 22.81 7.18 30.01 8.88 ;
        RECT 23.105 7.06 30.005 8.88 ;
        RECT 28.535 6.55 28.985 8.88 ;
        RECT 26.445 6.66 26.775 8.88 ;
        RECT 24.375 6.6 24.625 8.88 ;
        RECT 20.045 7.945 20.215 8.88 ;
        RECT 18.415 7.95 18.585 8.88 ;
        RECT 17.425 7.95 17.595 8.88 ;
        RECT 14.685 7.945 14.855 8.88 ;
        RECT 6.225 7.18 13.425 8.88 ;
        RECT 6.52 7.06 13.42 8.88 ;
        RECT 11.95 6.55 12.4 8.88 ;
        RECT 9.86 6.66 10.19 8.88 ;
        RECT 7.79 6.6 8.04 8.88 ;
        RECT 3.46 7.945 3.63 8.88 ;
        RECT 0 8.565 0.805 8.88 ;
        RECT 0.23 8.545 0.465 8.88 ;
        RECT 0.23 7.945 0.4 8.88 ;
        RECT 0.465 0 85.73 0.31 ;
        RECT 84.75 0 84.92 0.93 ;
        RECT 83.76 0 83.93 0.93 ;
        RECT 81.02 0 81.19 0.935 ;
        RECT 79.75 0 79.945 1.795 ;
        RECT 72.855 0 79.945 1.79 ;
        RECT 79.385 0 79.655 2.6 ;
        RECT 78.475 0 78.715 2.6 ;
        RECT 77.605 0 77.855 2.33 ;
        RECT 75.225 0 75.555 2.25 ;
        RECT 72.935 0 73.195 2.61 ;
        RECT 72.6 0 79.945 1.655 ;
        RECT 68.17 0 68.34 0.93 ;
        RECT 67.18 0 67.35 0.93 ;
        RECT 64.44 0 64.61 0.935 ;
        RECT 63.17 0 63.365 1.795 ;
        RECT 56.275 0 63.365 1.79 ;
        RECT 62.805 0 63.075 2.6 ;
        RECT 61.895 0 62.135 2.6 ;
        RECT 61.025 0 61.275 2.33 ;
        RECT 58.645 0 58.975 2.25 ;
        RECT 56.355 0 56.615 2.61 ;
        RECT 56.02 0 63.365 1.655 ;
        RECT 51.585 0 51.755 0.93 ;
        RECT 50.595 0 50.765 0.93 ;
        RECT 47.855 0 48.025 0.935 ;
        RECT 46.585 0 46.78 1.795 ;
        RECT 39.69 0 46.78 1.79 ;
        RECT 46.22 0 46.49 2.6 ;
        RECT 45.31 0 45.55 2.6 ;
        RECT 44.44 0 44.69 2.33 ;
        RECT 42.06 0 42.39 2.25 ;
        RECT 39.77 0 40.03 2.61 ;
        RECT 39.435 0 46.78 1.655 ;
        RECT 35 0 35.17 0.93 ;
        RECT 34.01 0 34.18 0.93 ;
        RECT 31.27 0 31.44 0.935 ;
        RECT 30 0 30.195 1.795 ;
        RECT 23.105 0 30.195 1.79 ;
        RECT 29.635 0 29.905 2.6 ;
        RECT 28.725 0 28.965 2.6 ;
        RECT 27.855 0 28.105 2.33 ;
        RECT 25.475 0 25.805 2.25 ;
        RECT 23.185 0 23.445 2.61 ;
        RECT 22.85 0 30.195 1.655 ;
        RECT 18.415 0 18.585 0.93 ;
        RECT 17.425 0 17.595 0.93 ;
        RECT 14.685 0 14.855 0.935 ;
        RECT 13.415 0 13.61 1.795 ;
        RECT 6.52 0 13.61 1.79 ;
        RECT 13.05 0 13.32 2.6 ;
        RECT 12.14 0 12.38 2.6 ;
        RECT 11.27 0 11.52 2.33 ;
        RECT 8.89 0 9.22 2.25 ;
        RECT 6.6 0 6.86 2.61 ;
        RECT 6.265 0 13.61 1.655 ;
        RECT 0 0.245 0.805 0.315 ;
        RECT 0.295 0.245 0.465 0.335 ;
        RECT 0 0 85.73 0.075 ;
        RECT 0 0 0.295 0.315 ;
        RECT 76.495 5.82 76.825 6.15 ;
        RECT 74.275 5.82 74.615 6.07 ;
        RECT 70.8 6.075 70.97 8.025 ;
        RECT 70.745 7.855 70.915 8.305 ;
        RECT 70.745 5.015 70.915 6.245 ;
        RECT 59.915 5.82 60.245 6.15 ;
        RECT 57.695 5.82 58.035 6.07 ;
        RECT 54.22 6.075 54.39 8.025 ;
        RECT 54.165 7.855 54.335 8.305 ;
        RECT 54.165 5.015 54.335 6.245 ;
        RECT 43.33 5.82 43.66 6.15 ;
        RECT 41.11 5.82 41.45 6.07 ;
        RECT 37.635 6.075 37.805 8.025 ;
        RECT 37.58 7.855 37.75 8.305 ;
        RECT 37.58 5.015 37.75 6.245 ;
        RECT 26.745 5.82 27.075 6.15 ;
        RECT 24.525 5.82 24.865 6.07 ;
        RECT 21.05 6.075 21.22 8.025 ;
        RECT 20.995 7.855 21.165 8.305 ;
        RECT 20.995 5.015 21.165 6.245 ;
        RECT 10.16 5.82 10.49 6.15 ;
        RECT 7.94 5.82 8.28 6.07 ;
        RECT 4.465 6.075 4.635 8.025 ;
        RECT 4.41 7.855 4.58 8.305 ;
        RECT 4.41 5.015 4.58 6.245 ;
      LAYER met2 ;
        RECT 75.255 6.45 75.535 6.82 ;
        RECT 58.675 6.45 58.955 6.82 ;
        RECT 42.09 6.45 42.37 6.82 ;
        RECT 25.505 6.45 25.785 6.82 ;
        RECT 8.92 6.45 9.2 6.82 ;
        RECT 0.19 8.5 0.57 8.88 ;
        RECT 0.19 0 0.57 0.38 ;
        RECT 0.235 0 0.39 8.88 ;
      LAYER met1 ;
        RECT 0 8.57 85.755 8.88 ;
        RECT 72.56 7.18 79.76 8.88 ;
        RECT 72.855 6.91 79.755 8.88 ;
        RECT 76.445 5.84 76.735 6.07 ;
        RECT 74.315 6.57 76.665 6.71 ;
        RECT 76.525 5.84 76.665 6.71 ;
        RECT 75.245 6.51 75.565 6.77 ;
        RECT 75.28 6.51 75.535 8.88 ;
        RECT 74.235 5.84 74.525 6.07 ;
        RECT 74.315 5.84 74.455 6.71 ;
        RECT 70.74 6.285 71.03 6.515 ;
        RECT 70.58 6.315 70.75 8.88 ;
        RECT 70.57 6.315 71.03 6.485 ;
        RECT 55.98 7.18 63.18 8.88 ;
        RECT 56.275 6.91 63.175 8.88 ;
        RECT 59.865 5.84 60.155 6.07 ;
        RECT 57.735 6.57 60.085 6.71 ;
        RECT 59.945 5.84 60.085 6.71 ;
        RECT 58.665 6.51 58.985 6.77 ;
        RECT 58.7 6.51 58.955 8.88 ;
        RECT 57.655 5.84 57.945 6.07 ;
        RECT 57.735 5.84 57.875 6.71 ;
        RECT 54.16 6.285 54.45 6.515 ;
        RECT 54 6.315 54.17 8.88 ;
        RECT 53.99 6.315 54.45 6.485 ;
        RECT 39.395 7.18 46.595 8.88 ;
        RECT 39.69 6.91 46.59 8.88 ;
        RECT 43.28 5.84 43.57 6.07 ;
        RECT 41.15 6.57 43.5 6.71 ;
        RECT 43.36 5.84 43.5 6.71 ;
        RECT 42.08 6.51 42.4 6.77 ;
        RECT 42.115 6.51 42.37 8.88 ;
        RECT 41.07 5.84 41.36 6.07 ;
        RECT 41.15 5.84 41.29 6.71 ;
        RECT 37.575 6.285 37.865 6.515 ;
        RECT 37.415 6.315 37.585 8.88 ;
        RECT 37.405 6.315 37.865 6.485 ;
        RECT 22.81 7.18 30.01 8.88 ;
        RECT 23.105 6.91 30.005 8.88 ;
        RECT 26.695 5.84 26.985 6.07 ;
        RECT 24.565 6.57 26.915 6.71 ;
        RECT 26.775 5.84 26.915 6.71 ;
        RECT 25.495 6.51 25.815 6.77 ;
        RECT 25.53 6.51 25.785 8.88 ;
        RECT 24.485 5.84 24.775 6.07 ;
        RECT 24.565 5.84 24.705 6.71 ;
        RECT 20.99 6.285 21.28 6.515 ;
        RECT 20.83 6.315 21 8.88 ;
        RECT 20.82 6.315 21.28 6.485 ;
        RECT 6.225 7.18 13.425 8.88 ;
        RECT 6.52 6.91 13.42 8.88 ;
        RECT 10.11 5.84 10.4 6.07 ;
        RECT 7.98 6.57 10.33 6.71 ;
        RECT 10.19 5.84 10.33 6.71 ;
        RECT 8.91 6.51 9.23 6.77 ;
        RECT 8.945 6.51 9.2 8.88 ;
        RECT 7.9 5.84 8.19 6.07 ;
        RECT 7.98 5.84 8.12 6.71 ;
        RECT 4.405 6.285 4.695 6.515 ;
        RECT 4.245 6.315 4.415 8.88 ;
        RECT 4.235 6.315 4.695 6.485 ;
        RECT 0 8.565 0.805 8.88 ;
        RECT 0.205 8.545 0.555 8.88 ;
        RECT 0 0 85.73 0.31 ;
        RECT 72.855 0 79.945 1.795 ;
        RECT 72.855 0 79.755 1.95 ;
        RECT 72.6 0 79.945 1.655 ;
        RECT 56.275 0 63.365 1.795 ;
        RECT 56.275 0 63.175 1.95 ;
        RECT 56.02 0 63.365 1.655 ;
        RECT 39.69 0 46.78 1.795 ;
        RECT 39.69 0 46.59 1.95 ;
        RECT 39.435 0 46.78 1.655 ;
        RECT 23.105 0 30.195 1.795 ;
        RECT 23.105 0 30.005 1.95 ;
        RECT 22.85 0 30.195 1.655 ;
        RECT 6.52 0 13.61 1.795 ;
        RECT 6.52 0 13.42 1.95 ;
        RECT 6.265 0 13.61 1.655 ;
        RECT 0 0 0.805 0.315 ;
        RECT 0.205 0 0.555 0.335 ;
      LAYER via2 ;
        RECT 0.28 8.59 0.48 8.79 ;
        RECT 0.28 0.09 0.48 0.29 ;
        RECT 8.96 6.54 9.16 6.74 ;
        RECT 25.545 6.54 25.745 6.74 ;
        RECT 42.13 6.54 42.33 6.74 ;
        RECT 58.715 6.54 58.915 6.74 ;
        RECT 75.295 6.54 75.495 6.74 ;
      LAYER mcon ;
        RECT 0.31 8.605 0.48 8.775 ;
        RECT 0.99 8.605 1.16 8.775 ;
        RECT 1.67 8.605 1.84 8.775 ;
        RECT 2.35 8.605 2.52 8.775 ;
        RECT 3.54 8.605 3.71 8.775 ;
        RECT 4.22 8.605 4.39 8.775 ;
        RECT 4.465 6.315 4.635 6.485 ;
        RECT 4.9 8.605 5.07 8.775 ;
        RECT 5.58 8.605 5.75 8.775 ;
        RECT 6.66 7.06 6.83 7.23 ;
        RECT 7.12 7.06 7.29 7.23 ;
        RECT 7.58 7.06 7.75 7.23 ;
        RECT 7.96 5.87 8.13 6.04 ;
        RECT 8.04 7.06 8.21 7.23 ;
        RECT 8.5 7.06 8.67 7.23 ;
        RECT 8.96 7.06 9.13 7.23 ;
        RECT 9.42 7.06 9.59 7.23 ;
        RECT 9.88 7.06 10.05 7.23 ;
        RECT 10.17 5.87 10.34 6.04 ;
        RECT 10.34 7.06 10.51 7.23 ;
        RECT 10.8 7.06 10.97 7.23 ;
        RECT 11.26 7.06 11.43 7.23 ;
        RECT 11.72 7.06 11.89 7.23 ;
        RECT 12.18 7.06 12.35 7.23 ;
        RECT 12.64 7.06 12.81 7.23 ;
        RECT 13.1 7.06 13.27 7.23 ;
        RECT 14.765 8.605 14.935 8.775 ;
        RECT 14.765 0.105 14.935 0.275 ;
        RECT 15.445 8.605 15.615 8.775 ;
        RECT 15.445 0.105 15.615 0.275 ;
        RECT 16.125 8.605 16.295 8.775 ;
        RECT 16.125 0.105 16.295 0.275 ;
        RECT 16.805 8.605 16.975 8.775 ;
        RECT 16.805 0.105 16.975 0.275 ;
        RECT 17.505 8.61 17.675 8.78 ;
        RECT 17.505 0.1 17.675 0.27 ;
        RECT 18.495 8.61 18.665 8.78 ;
        RECT 18.495 0.1 18.665 0.27 ;
        RECT 20.125 8.605 20.295 8.775 ;
        RECT 20.805 8.605 20.975 8.775 ;
        RECT 21.05 6.315 21.22 6.485 ;
        RECT 21.485 8.605 21.655 8.775 ;
        RECT 22.165 8.605 22.335 8.775 ;
        RECT 23.245 7.06 23.415 7.23 ;
        RECT 23.705 7.06 23.875 7.23 ;
        RECT 24.165 7.06 24.335 7.23 ;
        RECT 24.545 5.87 24.715 6.04 ;
        RECT 24.625 7.06 24.795 7.23 ;
        RECT 25.085 7.06 25.255 7.23 ;
        RECT 25.545 7.06 25.715 7.23 ;
        RECT 26.005 7.06 26.175 7.23 ;
        RECT 26.465 7.06 26.635 7.23 ;
        RECT 26.755 5.87 26.925 6.04 ;
        RECT 26.925 7.06 27.095 7.23 ;
        RECT 27.385 7.06 27.555 7.23 ;
        RECT 27.845 7.06 28.015 7.23 ;
        RECT 28.305 7.06 28.475 7.23 ;
        RECT 28.765 7.06 28.935 7.23 ;
        RECT 29.225 7.06 29.395 7.23 ;
        RECT 29.685 7.06 29.855 7.23 ;
        RECT 31.35 8.605 31.52 8.775 ;
        RECT 31.35 0.105 31.52 0.275 ;
        RECT 32.03 8.605 32.2 8.775 ;
        RECT 32.03 0.105 32.2 0.275 ;
        RECT 32.71 8.605 32.88 8.775 ;
        RECT 32.71 0.105 32.88 0.275 ;
        RECT 33.39 8.605 33.56 8.775 ;
        RECT 33.39 0.105 33.56 0.275 ;
        RECT 34.09 8.61 34.26 8.78 ;
        RECT 34.09 0.1 34.26 0.27 ;
        RECT 35.08 8.61 35.25 8.78 ;
        RECT 35.08 0.1 35.25 0.27 ;
        RECT 36.71 8.605 36.88 8.775 ;
        RECT 37.39 8.605 37.56 8.775 ;
        RECT 37.635 6.315 37.805 6.485 ;
        RECT 38.07 8.605 38.24 8.775 ;
        RECT 38.75 8.605 38.92 8.775 ;
        RECT 39.83 7.06 40 7.23 ;
        RECT 40.29 7.06 40.46 7.23 ;
        RECT 40.75 7.06 40.92 7.23 ;
        RECT 41.13 5.87 41.3 6.04 ;
        RECT 41.21 7.06 41.38 7.23 ;
        RECT 41.67 7.06 41.84 7.23 ;
        RECT 42.13 7.06 42.3 7.23 ;
        RECT 42.59 7.06 42.76 7.23 ;
        RECT 43.05 7.06 43.22 7.23 ;
        RECT 43.34 5.87 43.51 6.04 ;
        RECT 43.51 7.06 43.68 7.23 ;
        RECT 43.97 7.06 44.14 7.23 ;
        RECT 44.43 7.06 44.6 7.23 ;
        RECT 44.89 7.06 45.06 7.23 ;
        RECT 45.35 7.06 45.52 7.23 ;
        RECT 45.81 7.06 45.98 7.23 ;
        RECT 46.27 7.06 46.44 7.23 ;
        RECT 47.935 8.605 48.105 8.775 ;
        RECT 47.935 0.105 48.105 0.275 ;
        RECT 48.615 8.605 48.785 8.775 ;
        RECT 48.615 0.105 48.785 0.275 ;
        RECT 49.295 8.605 49.465 8.775 ;
        RECT 49.295 0.105 49.465 0.275 ;
        RECT 49.975 8.605 50.145 8.775 ;
        RECT 49.975 0.105 50.145 0.275 ;
        RECT 50.675 8.61 50.845 8.78 ;
        RECT 50.675 0.1 50.845 0.27 ;
        RECT 51.665 8.61 51.835 8.78 ;
        RECT 51.665 0.1 51.835 0.27 ;
        RECT 53.295 8.605 53.465 8.775 ;
        RECT 53.975 8.605 54.145 8.775 ;
        RECT 54.22 6.315 54.39 6.485 ;
        RECT 54.655 8.605 54.825 8.775 ;
        RECT 55.335 8.605 55.505 8.775 ;
        RECT 56.415 7.06 56.585 7.23 ;
        RECT 56.875 7.06 57.045 7.23 ;
        RECT 57.335 7.06 57.505 7.23 ;
        RECT 57.715 5.87 57.885 6.04 ;
        RECT 57.795 7.06 57.965 7.23 ;
        RECT 58.255 7.06 58.425 7.23 ;
        RECT 58.715 7.06 58.885 7.23 ;
        RECT 59.175 7.06 59.345 7.23 ;
        RECT 59.635 7.06 59.805 7.23 ;
        RECT 59.925 5.87 60.095 6.04 ;
        RECT 60.095 7.06 60.265 7.23 ;
        RECT 60.555 7.06 60.725 7.23 ;
        RECT 61.015 7.06 61.185 7.23 ;
        RECT 61.475 7.06 61.645 7.23 ;
        RECT 61.935 7.06 62.105 7.23 ;
        RECT 62.395 7.06 62.565 7.23 ;
        RECT 62.855 7.06 63.025 7.23 ;
        RECT 64.52 8.605 64.69 8.775 ;
        RECT 64.52 0.105 64.69 0.275 ;
        RECT 65.2 8.605 65.37 8.775 ;
        RECT 65.2 0.105 65.37 0.275 ;
        RECT 65.88 8.605 66.05 8.775 ;
        RECT 65.88 0.105 66.05 0.275 ;
        RECT 66.56 8.605 66.73 8.775 ;
        RECT 66.56 0.105 66.73 0.275 ;
        RECT 67.26 8.61 67.43 8.78 ;
        RECT 67.26 0.1 67.43 0.27 ;
        RECT 68.25 8.61 68.42 8.78 ;
        RECT 68.25 0.1 68.42 0.27 ;
        RECT 69.875 8.605 70.045 8.775 ;
        RECT 70.555 8.605 70.725 8.775 ;
        RECT 70.8 6.315 70.97 6.485 ;
        RECT 71.235 8.605 71.405 8.775 ;
        RECT 71.915 8.605 72.085 8.775 ;
        RECT 72.995 7.06 73.165 7.23 ;
        RECT 73.455 7.06 73.625 7.23 ;
        RECT 73.915 7.06 74.085 7.23 ;
        RECT 74.295 5.87 74.465 6.04 ;
        RECT 74.375 7.06 74.545 7.23 ;
        RECT 74.835 7.06 75.005 7.23 ;
        RECT 75.295 7.06 75.465 7.23 ;
        RECT 75.755 7.06 75.925 7.23 ;
        RECT 76.215 7.06 76.385 7.23 ;
        RECT 76.505 5.87 76.675 6.04 ;
        RECT 76.675 7.06 76.845 7.23 ;
        RECT 77.135 7.06 77.305 7.23 ;
        RECT 77.595 7.06 77.765 7.23 ;
        RECT 78.055 7.06 78.225 7.23 ;
        RECT 78.515 7.06 78.685 7.23 ;
        RECT 78.975 7.06 79.145 7.23 ;
        RECT 79.435 7.06 79.605 7.23 ;
        RECT 81.1 8.605 81.27 8.775 ;
        RECT 81.1 0.105 81.27 0.275 ;
        RECT 81.78 8.605 81.95 8.775 ;
        RECT 81.78 0.105 81.95 0.275 ;
        RECT 82.46 8.605 82.63 8.775 ;
        RECT 82.46 0.105 82.63 0.275 ;
        RECT 83.14 8.605 83.31 8.775 ;
        RECT 83.14 0.105 83.31 0.275 ;
        RECT 83.84 8.61 84.01 8.78 ;
        RECT 83.84 0.1 84.01 0.27 ;
        RECT 84.83 8.61 85 8.78 ;
        RECT 84.83 0.1 85 0.27 ;
      LAYER via1 ;
        RECT 0.305 8.615 0.455 8.765 ;
        RECT 0.305 0.115 0.455 0.265 ;
        RECT 8.995 6.565 9.145 6.715 ;
        RECT 25.58 6.565 25.73 6.715 ;
        RECT 42.165 6.565 42.315 6.715 ;
        RECT 58.75 6.565 58.9 6.715 ;
        RECT 75.33 6.565 75.48 6.715 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 77.65 2.73 77.95 3.065 ;
      RECT 77.625 2.73 77.955 3.06 ;
      RECT 77.625 2.75 78.425 3.05 ;
      RECT 71.95 7.97 76.23 8.27 ;
      RECT 75.925 5.79 76.225 8.27 ;
      RECT 71.95 7.03 72.25 8.27 ;
      RECT 71.075 6.995 71.445 7.365 ;
      RECT 71.075 7.03 72.25 7.33 ;
      RECT 75.3 5.795 76.235 6.125 ;
      RECT 75.905 5.79 76.235 6.125 ;
      RECT 76.945 5.79 77.275 6.12 ;
      RECT 75.3 5.81 77.745 6.11 ;
      RECT 75.3 5.795 77.275 6.11 ;
      RECT 75.3 3.765 75.63 6.125 ;
      RECT 75.3 3.765 77.595 4.095 ;
      RECT 75.3 3.765 77.95 4.085 ;
      RECT 77.625 3.75 77.955 4.08 ;
      RECT 75.3 3.77 78.425 4.07 ;
      RECT 77.635 3.7 77.935 4.085 ;
      RECT 76.925 3.07 77.255 3.4 ;
      RECT 76.955 3.06 77.255 3.4 ;
      RECT 76.455 3.09 77.255 3.39 ;
      RECT 76.27 4.77 76.305 5.105 ;
      RECT 76.265 4.77 76.595 5.1 ;
      RECT 76.265 4.79 77.065 5.09 ;
      RECT 76.265 4.785 76.6 5.09 ;
      RECT 75.585 2.39 75.915 2.72 ;
      RECT 75.115 2.41 75.475 2.71 ;
      RECT 75.475 2.4 75.915 2.7 ;
      RECT 61.07 2.73 61.37 3.065 ;
      RECT 61.045 2.73 61.375 3.06 ;
      RECT 61.045 2.75 61.845 3.05 ;
      RECT 55.37 7.97 59.65 8.27 ;
      RECT 59.345 5.79 59.645 8.27 ;
      RECT 55.37 7.03 55.67 8.27 ;
      RECT 54.495 6.995 54.865 7.365 ;
      RECT 54.495 7.03 55.67 7.33 ;
      RECT 58.72 5.795 59.655 6.125 ;
      RECT 59.325 5.79 59.655 6.125 ;
      RECT 60.365 5.79 60.695 6.12 ;
      RECT 58.72 5.81 61.165 6.11 ;
      RECT 58.72 5.795 60.695 6.11 ;
      RECT 58.72 3.765 59.05 6.125 ;
      RECT 58.72 3.765 61.015 4.095 ;
      RECT 58.72 3.765 61.37 4.085 ;
      RECT 61.045 3.75 61.375 4.08 ;
      RECT 58.72 3.77 61.845 4.07 ;
      RECT 61.055 3.7 61.355 4.085 ;
      RECT 60.345 3.07 60.675 3.4 ;
      RECT 60.375 3.06 60.675 3.4 ;
      RECT 59.875 3.09 60.675 3.39 ;
      RECT 59.69 4.77 59.725 5.105 ;
      RECT 59.685 4.77 60.015 5.1 ;
      RECT 59.685 4.79 60.485 5.09 ;
      RECT 59.685 4.785 60.02 5.09 ;
      RECT 59.005 2.39 59.335 2.72 ;
      RECT 58.535 2.41 58.895 2.71 ;
      RECT 58.895 2.4 59.335 2.7 ;
      RECT 44.485 2.73 44.785 3.065 ;
      RECT 44.46 2.73 44.79 3.06 ;
      RECT 44.46 2.75 45.26 3.05 ;
      RECT 38.785 7.97 43.065 8.27 ;
      RECT 42.76 5.79 43.06 8.27 ;
      RECT 38.785 7.03 39.085 8.27 ;
      RECT 37.91 6.995 38.28 7.365 ;
      RECT 37.91 7.03 39.085 7.33 ;
      RECT 42.135 5.795 43.07 6.125 ;
      RECT 42.74 5.79 43.07 6.125 ;
      RECT 43.78 5.79 44.11 6.12 ;
      RECT 42.135 5.81 44.58 6.11 ;
      RECT 42.135 5.795 44.11 6.11 ;
      RECT 42.135 3.765 42.465 6.125 ;
      RECT 42.135 3.765 44.43 4.095 ;
      RECT 42.135 3.765 44.785 4.085 ;
      RECT 44.46 3.75 44.79 4.08 ;
      RECT 42.135 3.77 45.26 4.07 ;
      RECT 44.47 3.7 44.77 4.085 ;
      RECT 43.76 3.07 44.09 3.4 ;
      RECT 43.79 3.06 44.09 3.4 ;
      RECT 43.29 3.09 44.09 3.39 ;
      RECT 43.105 4.77 43.14 5.105 ;
      RECT 43.1 4.77 43.43 5.1 ;
      RECT 43.1 4.79 43.9 5.09 ;
      RECT 43.1 4.785 43.435 5.09 ;
      RECT 42.42 2.39 42.75 2.72 ;
      RECT 41.95 2.41 42.31 2.71 ;
      RECT 42.31 2.4 42.75 2.7 ;
      RECT 27.9 2.73 28.2 3.065 ;
      RECT 27.875 2.73 28.205 3.06 ;
      RECT 27.875 2.75 28.675 3.05 ;
      RECT 22.2 7.97 26.48 8.27 ;
      RECT 26.175 5.79 26.475 8.27 ;
      RECT 22.2 7.03 22.5 8.27 ;
      RECT 21.325 6.995 21.695 7.365 ;
      RECT 21.325 7.03 22.5 7.33 ;
      RECT 25.55 5.795 26.485 6.125 ;
      RECT 26.155 5.79 26.485 6.125 ;
      RECT 27.195 5.79 27.525 6.12 ;
      RECT 25.55 5.81 27.995 6.11 ;
      RECT 25.55 5.795 27.525 6.11 ;
      RECT 25.55 3.765 25.88 6.125 ;
      RECT 25.55 3.765 27.845 4.095 ;
      RECT 25.55 3.765 28.2 4.085 ;
      RECT 27.875 3.75 28.205 4.08 ;
      RECT 25.55 3.77 28.675 4.07 ;
      RECT 27.885 3.7 28.185 4.085 ;
      RECT 27.175 3.07 27.505 3.4 ;
      RECT 27.205 3.06 27.505 3.4 ;
      RECT 26.705 3.09 27.505 3.39 ;
      RECT 26.52 4.77 26.555 5.105 ;
      RECT 26.515 4.77 26.845 5.1 ;
      RECT 26.515 4.79 27.315 5.09 ;
      RECT 26.515 4.785 26.85 5.09 ;
      RECT 25.835 2.39 26.165 2.72 ;
      RECT 25.365 2.41 25.725 2.71 ;
      RECT 25.725 2.4 26.165 2.7 ;
      RECT 11.315 2.73 11.615 3.065 ;
      RECT 11.29 2.73 11.62 3.06 ;
      RECT 11.29 2.75 12.09 3.05 ;
      RECT 5.615 7.97 9.895 8.27 ;
      RECT 9.59 5.79 9.89 8.27 ;
      RECT 5.615 7.03 5.915 8.27 ;
      RECT 4.74 6.995 5.11 7.365 ;
      RECT 4.74 7.03 5.915 7.33 ;
      RECT 8.965 5.795 9.9 6.125 ;
      RECT 9.57 5.79 9.9 6.125 ;
      RECT 10.61 5.79 10.94 6.12 ;
      RECT 8.965 5.81 11.41 6.11 ;
      RECT 8.965 5.795 10.94 6.11 ;
      RECT 8.965 3.765 9.295 6.125 ;
      RECT 8.965 3.765 11.26 4.095 ;
      RECT 8.965 3.765 11.615 4.085 ;
      RECT 11.29 3.75 11.62 4.08 ;
      RECT 8.965 3.77 12.09 4.07 ;
      RECT 11.3 3.7 11.6 4.085 ;
      RECT 10.59 3.07 10.92 3.4 ;
      RECT 10.62 3.06 10.92 3.4 ;
      RECT 10.12 3.09 10.92 3.39 ;
      RECT 9.935 4.77 9.97 5.105 ;
      RECT 9.93 4.77 10.26 5.1 ;
      RECT 9.93 4.79 10.73 5.09 ;
      RECT 9.93 4.785 10.265 5.09 ;
      RECT 9.25 2.39 9.58 2.72 ;
      RECT 8.78 2.41 9.14 2.71 ;
      RECT 9.14 2.4 9.58 2.7 ;
    LAYER via2 ;
      RECT 77.695 2.8 77.895 3 ;
      RECT 77.695 3.82 77.895 4.02 ;
      RECT 77.015 5.86 77.215 6.06 ;
      RECT 76.995 3.14 77.195 3.34 ;
      RECT 76.335 4.84 76.535 5.04 ;
      RECT 75.965 5.86 76.165 6.06 ;
      RECT 75.655 2.45 75.855 2.65 ;
      RECT 71.16 7.08 71.36 7.28 ;
      RECT 61.115 2.8 61.315 3 ;
      RECT 61.115 3.82 61.315 4.02 ;
      RECT 60.435 5.86 60.635 6.06 ;
      RECT 60.415 3.14 60.615 3.34 ;
      RECT 59.755 4.84 59.955 5.04 ;
      RECT 59.385 5.86 59.585 6.06 ;
      RECT 59.075 2.45 59.275 2.65 ;
      RECT 54.58 7.08 54.78 7.28 ;
      RECT 44.53 2.8 44.73 3 ;
      RECT 44.53 3.82 44.73 4.02 ;
      RECT 43.85 5.86 44.05 6.06 ;
      RECT 43.83 3.14 44.03 3.34 ;
      RECT 43.17 4.84 43.37 5.04 ;
      RECT 42.8 5.86 43 6.06 ;
      RECT 42.49 2.45 42.69 2.65 ;
      RECT 37.995 7.08 38.195 7.28 ;
      RECT 27.945 2.8 28.145 3 ;
      RECT 27.945 3.82 28.145 4.02 ;
      RECT 27.265 5.86 27.465 6.06 ;
      RECT 27.245 3.14 27.445 3.34 ;
      RECT 26.585 4.84 26.785 5.04 ;
      RECT 26.215 5.86 26.415 6.06 ;
      RECT 25.905 2.45 26.105 2.65 ;
      RECT 21.41 7.08 21.61 7.28 ;
      RECT 11.36 2.8 11.56 3 ;
      RECT 11.36 3.82 11.56 4.02 ;
      RECT 10.68 5.86 10.88 6.06 ;
      RECT 10.66 3.14 10.86 3.34 ;
      RECT 10 4.84 10.2 5.04 ;
      RECT 9.63 5.86 9.83 6.06 ;
      RECT 9.32 2.45 9.52 2.65 ;
      RECT 4.825 7.08 5.025 7.28 ;
    LAYER met2 ;
      RECT 1.23 8.6 85.355 8.77 ;
      RECT 85.185 7.3 85.355 8.77 ;
      RECT 1.23 6.255 1.4 8.77 ;
      RECT 85.15 7.3 85.475 7.625 ;
      RECT 1.175 6.255 1.455 6.595 ;
      RECT 81.995 6.28 82.315 6.605 ;
      RECT 82.025 5.695 82.195 6.605 ;
      RECT 82.025 5.695 82.2 6.045 ;
      RECT 82.025 5.695 83 5.87 ;
      RECT 82.825 1.965 83 5.87 ;
      RECT 82.77 1.965 83.12 2.315 ;
      RECT 71.66 8.29 81.84 8.46 ;
      RECT 81.68 2.395 81.84 8.46 ;
      RECT 71.66 6.6 71.83 8.46 ;
      RECT 82.795 6.655 83.12 6.98 ;
      RECT 68.605 6.655 68.93 6.98 ;
      RECT 71.605 6.6 71.885 6.94 ;
      RECT 81.68 6.745 83.12 6.915 ;
      RECT 68.605 6.685 71.885 6.855 ;
      RECT 81.995 2.365 82.315 2.685 ;
      RECT 81.68 2.395 82.315 2.565 ;
      RECT 79.74 3.185 80.065 3.51 ;
      RECT 79.74 3.215 80.57 3.4 ;
      RECT 80.4 1.995 80.57 3.4 ;
      RECT 80.325 1.995 80.65 2.32 ;
      RECT 79.355 4.78 79.615 5.1 ;
      RECT 79.415 2.74 79.555 5.1 ;
      RECT 79.355 2.74 79.615 3.06 ;
      RECT 78.335 5.8 78.595 6.12 ;
      RECT 77.715 5.89 78.595 6.03 ;
      RECT 77.715 3.73 77.855 6.03 ;
      RECT 77.655 3.73 77.935 4.1 ;
      RECT 76.975 5.77 77.255 6.14 ;
      RECT 77.035 3.85 77.175 6.14 ;
      RECT 77.035 3.85 77.515 3.99 ;
      RECT 77.375 2.06 77.515 3.99 ;
      RECT 77.315 2.06 77.575 2.38 ;
      RECT 76.295 4.75 76.575 5.12 ;
      RECT 76.355 2.4 76.495 5.12 ;
      RECT 76.295 2.4 76.555 2.72 ;
      RECT 75.925 5.77 76.205 6.14 ;
      RECT 75.925 5.8 76.215 6.12 ;
      RECT 65.415 6.28 65.735 6.605 ;
      RECT 65.445 5.695 65.615 6.605 ;
      RECT 65.445 5.695 65.62 6.045 ;
      RECT 65.445 5.695 66.42 5.87 ;
      RECT 66.245 1.965 66.42 5.87 ;
      RECT 66.19 1.965 66.54 2.315 ;
      RECT 55.08 8.29 65.26 8.46 ;
      RECT 65.1 2.395 65.26 8.46 ;
      RECT 55.08 6.6 55.25 8.46 ;
      RECT 66.215 6.655 66.54 6.98 ;
      RECT 52.02 6.655 52.345 6.98 ;
      RECT 55.025 6.6 55.305 6.94 ;
      RECT 65.1 6.745 66.54 6.915 ;
      RECT 52.02 6.685 55.305 6.855 ;
      RECT 65.415 2.365 65.735 2.685 ;
      RECT 65.1 2.395 65.735 2.565 ;
      RECT 63.16 3.185 63.485 3.51 ;
      RECT 63.16 3.215 63.99 3.4 ;
      RECT 63.82 1.995 63.99 3.4 ;
      RECT 63.745 1.995 64.07 2.32 ;
      RECT 62.775 4.78 63.035 5.1 ;
      RECT 62.835 2.74 62.975 5.1 ;
      RECT 62.775 2.74 63.035 3.06 ;
      RECT 61.755 5.8 62.015 6.12 ;
      RECT 61.135 5.89 62.015 6.03 ;
      RECT 61.135 3.73 61.275 6.03 ;
      RECT 61.075 3.73 61.355 4.1 ;
      RECT 60.395 5.77 60.675 6.14 ;
      RECT 60.455 3.85 60.595 6.14 ;
      RECT 60.455 3.85 60.935 3.99 ;
      RECT 60.795 2.06 60.935 3.99 ;
      RECT 60.735 2.06 60.995 2.38 ;
      RECT 59.715 4.75 59.995 5.12 ;
      RECT 59.775 2.4 59.915 5.12 ;
      RECT 59.715 2.4 59.975 2.72 ;
      RECT 59.345 5.77 59.625 6.14 ;
      RECT 59.345 5.8 59.635 6.12 ;
      RECT 48.83 6.28 49.15 6.605 ;
      RECT 48.86 5.695 49.03 6.605 ;
      RECT 48.86 5.695 49.035 6.045 ;
      RECT 48.86 5.695 49.835 5.87 ;
      RECT 49.66 1.965 49.835 5.87 ;
      RECT 49.605 1.965 49.955 2.315 ;
      RECT 38.495 8.29 48.675 8.46 ;
      RECT 48.515 2.395 48.675 8.46 ;
      RECT 38.495 6.6 38.665 8.46 ;
      RECT 49.63 6.655 49.955 6.98 ;
      RECT 35.435 6.655 35.76 6.98 ;
      RECT 38.44 6.6 38.72 6.94 ;
      RECT 48.515 6.745 49.955 6.915 ;
      RECT 35.435 6.685 38.72 6.855 ;
      RECT 48.83 2.365 49.15 2.685 ;
      RECT 48.515 2.395 49.15 2.565 ;
      RECT 46.575 3.185 46.9 3.51 ;
      RECT 46.575 3.215 47.405 3.4 ;
      RECT 47.235 1.995 47.405 3.4 ;
      RECT 47.16 1.995 47.485 2.32 ;
      RECT 46.19 4.78 46.45 5.1 ;
      RECT 46.25 2.74 46.39 5.1 ;
      RECT 46.19 2.74 46.45 3.06 ;
      RECT 45.17 5.8 45.43 6.12 ;
      RECT 44.55 5.89 45.43 6.03 ;
      RECT 44.55 3.73 44.69 6.03 ;
      RECT 44.49 3.73 44.77 4.1 ;
      RECT 43.81 5.77 44.09 6.14 ;
      RECT 43.87 3.85 44.01 6.14 ;
      RECT 43.87 3.85 44.35 3.99 ;
      RECT 44.21 2.06 44.35 3.99 ;
      RECT 44.15 2.06 44.41 2.38 ;
      RECT 43.13 4.75 43.41 5.12 ;
      RECT 43.19 2.4 43.33 5.12 ;
      RECT 43.13 2.4 43.39 2.72 ;
      RECT 42.76 5.77 43.04 6.14 ;
      RECT 42.76 5.8 43.05 6.12 ;
      RECT 32.245 6.28 32.565 6.605 ;
      RECT 32.275 5.695 32.445 6.605 ;
      RECT 32.275 5.695 32.45 6.045 ;
      RECT 32.275 5.695 33.25 5.87 ;
      RECT 33.075 1.965 33.25 5.87 ;
      RECT 33.02 1.965 33.37 2.315 ;
      RECT 21.91 8.29 32.09 8.46 ;
      RECT 31.93 2.395 32.09 8.46 ;
      RECT 21.91 6.6 22.08 8.46 ;
      RECT 33.045 6.655 33.37 6.98 ;
      RECT 18.85 6.655 19.175 6.98 ;
      RECT 21.855 6.6 22.135 6.94 ;
      RECT 31.93 6.745 33.37 6.915 ;
      RECT 18.85 6.685 22.135 6.855 ;
      RECT 32.245 2.365 32.565 2.685 ;
      RECT 31.93 2.395 32.565 2.565 ;
      RECT 29.99 3.185 30.315 3.51 ;
      RECT 29.99 3.215 30.82 3.4 ;
      RECT 30.65 1.995 30.82 3.4 ;
      RECT 30.575 1.995 30.9 2.32 ;
      RECT 29.605 4.78 29.865 5.1 ;
      RECT 29.665 2.74 29.805 5.1 ;
      RECT 29.605 2.74 29.865 3.06 ;
      RECT 28.585 5.8 28.845 6.12 ;
      RECT 27.965 5.89 28.845 6.03 ;
      RECT 27.965 3.73 28.105 6.03 ;
      RECT 27.905 3.73 28.185 4.1 ;
      RECT 27.225 5.77 27.505 6.14 ;
      RECT 27.285 3.85 27.425 6.14 ;
      RECT 27.285 3.85 27.765 3.99 ;
      RECT 27.625 2.06 27.765 3.99 ;
      RECT 27.565 2.06 27.825 2.38 ;
      RECT 26.545 4.75 26.825 5.12 ;
      RECT 26.605 2.4 26.745 5.12 ;
      RECT 26.545 2.4 26.805 2.72 ;
      RECT 26.175 5.77 26.455 6.14 ;
      RECT 26.175 5.8 26.465 6.12 ;
      RECT 15.66 6.28 15.98 6.605 ;
      RECT 15.69 5.695 15.86 6.605 ;
      RECT 15.69 5.695 15.865 6.045 ;
      RECT 15.69 5.695 16.665 5.87 ;
      RECT 16.49 1.965 16.665 5.87 ;
      RECT 16.435 1.965 16.785 2.315 ;
      RECT 5.325 8.29 15.505 8.46 ;
      RECT 15.345 2.395 15.505 8.46 ;
      RECT 5.325 6.6 5.495 8.46 ;
      RECT 1.55 6.995 1.83 7.335 ;
      RECT 1.55 7.06 2.715 7.23 ;
      RECT 2.545 6.685 2.715 7.23 ;
      RECT 16.46 6.655 16.785 6.98 ;
      RECT 5.27 6.6 5.55 6.94 ;
      RECT 15.345 6.745 16.785 6.915 ;
      RECT 2.545 6.685 5.55 6.855 ;
      RECT 15.66 2.365 15.98 2.685 ;
      RECT 15.345 2.395 15.98 2.565 ;
      RECT 13.405 3.185 13.73 3.51 ;
      RECT 13.405 3.215 14.235 3.4 ;
      RECT 14.065 1.995 14.235 3.4 ;
      RECT 13.99 1.995 14.315 2.32 ;
      RECT 13.02 4.78 13.28 5.1 ;
      RECT 13.08 2.74 13.22 5.1 ;
      RECT 13.02 2.74 13.28 3.06 ;
      RECT 12 5.8 12.26 6.12 ;
      RECT 11.38 5.89 12.26 6.03 ;
      RECT 11.38 3.73 11.52 6.03 ;
      RECT 11.32 3.73 11.6 4.1 ;
      RECT 10.64 5.77 10.92 6.14 ;
      RECT 10.7 3.85 10.84 6.14 ;
      RECT 10.7 3.85 11.18 3.99 ;
      RECT 11.04 2.06 11.18 3.99 ;
      RECT 10.98 2.06 11.24 2.38 ;
      RECT 9.96 4.75 10.24 5.12 ;
      RECT 10.02 2.4 10.16 5.12 ;
      RECT 9.96 2.4 10.22 2.72 ;
      RECT 9.59 5.77 9.87 6.14 ;
      RECT 9.59 5.8 9.88 6.12 ;
      RECT 77.655 2.71 77.935 3.08 ;
      RECT 76.955 3.05 77.235 3.42 ;
      RECT 75.615 2.37 75.895 2.74 ;
      RECT 71.075 6.995 71.45 7.365 ;
      RECT 61.075 2.71 61.355 3.08 ;
      RECT 60.375 3.05 60.655 3.42 ;
      RECT 59.035 2.37 59.315 2.74 ;
      RECT 54.495 6.995 54.865 7.365 ;
      RECT 44.49 2.71 44.77 3.08 ;
      RECT 43.79 3.05 44.07 3.42 ;
      RECT 42.45 2.37 42.73 2.74 ;
      RECT 37.91 6.995 38.28 7.365 ;
      RECT 27.905 2.71 28.185 3.08 ;
      RECT 27.205 3.05 27.485 3.42 ;
      RECT 25.865 2.37 26.145 2.74 ;
      RECT 21.325 6.995 21.695 7.365 ;
      RECT 11.32 2.71 11.6 3.08 ;
      RECT 10.62 3.05 10.9 3.42 ;
      RECT 9.28 2.37 9.56 2.74 ;
      RECT 4.74 6.995 5.11 7.365 ;
    LAYER via1 ;
      RECT 85.24 7.385 85.39 7.535 ;
      RECT 82.885 6.74 83.035 6.89 ;
      RECT 82.87 2.065 83.02 2.215 ;
      RECT 82.08 2.45 82.23 2.6 ;
      RECT 82.08 6.37 82.23 6.52 ;
      RECT 80.415 2.08 80.565 2.23 ;
      RECT 79.83 3.27 79.98 3.42 ;
      RECT 79.41 2.825 79.56 2.975 ;
      RECT 79.41 4.865 79.56 5.015 ;
      RECT 78.39 5.885 78.54 6.035 ;
      RECT 77.71 2.825 77.86 2.975 ;
      RECT 77.71 3.845 77.86 3.995 ;
      RECT 77.37 2.145 77.52 2.295 ;
      RECT 77.03 3.165 77.18 3.315 ;
      RECT 77.03 5.885 77.18 6.035 ;
      RECT 76.35 2.485 76.5 2.635 ;
      RECT 76.35 4.865 76.5 5.015 ;
      RECT 76.01 5.885 76.16 6.035 ;
      RECT 75.67 2.475 75.82 2.625 ;
      RECT 71.67 6.695 71.82 6.845 ;
      RECT 71.185 7.105 71.335 7.255 ;
      RECT 68.695 6.74 68.845 6.89 ;
      RECT 66.305 6.74 66.455 6.89 ;
      RECT 66.29 2.065 66.44 2.215 ;
      RECT 65.5 2.45 65.65 2.6 ;
      RECT 65.5 6.37 65.65 6.52 ;
      RECT 63.835 2.08 63.985 2.23 ;
      RECT 63.25 3.27 63.4 3.42 ;
      RECT 62.83 2.825 62.98 2.975 ;
      RECT 62.83 4.865 62.98 5.015 ;
      RECT 61.81 5.885 61.96 6.035 ;
      RECT 61.13 2.825 61.28 2.975 ;
      RECT 61.13 3.845 61.28 3.995 ;
      RECT 60.79 2.145 60.94 2.295 ;
      RECT 60.45 3.165 60.6 3.315 ;
      RECT 60.45 5.885 60.6 6.035 ;
      RECT 59.77 2.485 59.92 2.635 ;
      RECT 59.77 4.865 59.92 5.015 ;
      RECT 59.43 5.885 59.58 6.035 ;
      RECT 59.09 2.475 59.24 2.625 ;
      RECT 55.09 6.695 55.24 6.845 ;
      RECT 54.605 7.105 54.755 7.255 ;
      RECT 52.11 6.74 52.26 6.89 ;
      RECT 49.72 6.74 49.87 6.89 ;
      RECT 49.705 2.065 49.855 2.215 ;
      RECT 48.915 2.45 49.065 2.6 ;
      RECT 48.915 6.37 49.065 6.52 ;
      RECT 47.25 2.08 47.4 2.23 ;
      RECT 46.665 3.27 46.815 3.42 ;
      RECT 46.245 2.825 46.395 2.975 ;
      RECT 46.245 4.865 46.395 5.015 ;
      RECT 45.225 5.885 45.375 6.035 ;
      RECT 44.545 2.825 44.695 2.975 ;
      RECT 44.545 3.845 44.695 3.995 ;
      RECT 44.205 2.145 44.355 2.295 ;
      RECT 43.865 3.165 44.015 3.315 ;
      RECT 43.865 5.885 44.015 6.035 ;
      RECT 43.185 2.485 43.335 2.635 ;
      RECT 43.185 4.865 43.335 5.015 ;
      RECT 42.845 5.885 42.995 6.035 ;
      RECT 42.505 2.475 42.655 2.625 ;
      RECT 38.505 6.695 38.655 6.845 ;
      RECT 38.02 7.105 38.17 7.255 ;
      RECT 35.525 6.74 35.675 6.89 ;
      RECT 33.135 6.74 33.285 6.89 ;
      RECT 33.12 2.065 33.27 2.215 ;
      RECT 32.33 2.45 32.48 2.6 ;
      RECT 32.33 6.37 32.48 6.52 ;
      RECT 30.665 2.08 30.815 2.23 ;
      RECT 30.08 3.27 30.23 3.42 ;
      RECT 29.66 2.825 29.81 2.975 ;
      RECT 29.66 4.865 29.81 5.015 ;
      RECT 28.64 5.885 28.79 6.035 ;
      RECT 27.96 2.825 28.11 2.975 ;
      RECT 27.96 3.845 28.11 3.995 ;
      RECT 27.62 2.145 27.77 2.295 ;
      RECT 27.28 3.165 27.43 3.315 ;
      RECT 27.28 5.885 27.43 6.035 ;
      RECT 26.6 2.485 26.75 2.635 ;
      RECT 26.6 4.865 26.75 5.015 ;
      RECT 26.26 5.885 26.41 6.035 ;
      RECT 25.92 2.475 26.07 2.625 ;
      RECT 21.92 6.695 22.07 6.845 ;
      RECT 21.435 7.105 21.585 7.255 ;
      RECT 18.94 6.74 19.09 6.89 ;
      RECT 16.55 6.74 16.7 6.89 ;
      RECT 16.535 2.065 16.685 2.215 ;
      RECT 15.745 2.45 15.895 2.6 ;
      RECT 15.745 6.37 15.895 6.52 ;
      RECT 14.08 2.08 14.23 2.23 ;
      RECT 13.495 3.27 13.645 3.42 ;
      RECT 13.075 2.825 13.225 2.975 ;
      RECT 13.075 4.865 13.225 5.015 ;
      RECT 12.055 5.885 12.205 6.035 ;
      RECT 11.375 2.825 11.525 2.975 ;
      RECT 11.375 3.845 11.525 3.995 ;
      RECT 11.035 2.145 11.185 2.295 ;
      RECT 10.695 3.165 10.845 3.315 ;
      RECT 10.695 5.885 10.845 6.035 ;
      RECT 10.015 2.485 10.165 2.635 ;
      RECT 10.015 4.865 10.165 5.015 ;
      RECT 9.675 5.885 9.825 6.035 ;
      RECT 9.335 2.475 9.485 2.625 ;
      RECT 5.335 6.695 5.485 6.845 ;
      RECT 4.85 7.105 5 7.255 ;
      RECT 1.615 7.09 1.765 7.24 ;
      RECT 1.24 6.35 1.39 6.5 ;
    LAYER met1 ;
      RECT 85.12 7.77 85.41 8 ;
      RECT 85.18 6.29 85.35 8 ;
      RECT 85.15 7.3 85.475 7.625 ;
      RECT 85.12 6.29 85.41 6.52 ;
      RECT 84.715 2.395 84.82 2.965 ;
      RECT 84.715 2.73 85.04 2.96 ;
      RECT 84.715 2.76 85.21 2.93 ;
      RECT 84.715 2.395 84.905 2.96 ;
      RECT 84.13 2.36 84.42 2.59 ;
      RECT 84.13 2.395 84.905 2.565 ;
      RECT 84.19 0.88 84.36 2.59 ;
      RECT 84.13 0.88 84.42 1.11 ;
      RECT 84.13 7.77 84.42 8 ;
      RECT 84.19 6.29 84.36 8 ;
      RECT 84.13 6.29 84.42 6.52 ;
      RECT 84.13 6.325 84.985 6.485 ;
      RECT 84.815 5.92 84.985 6.485 ;
      RECT 84.13 6.32 84.525 6.485 ;
      RECT 84.75 5.92 85.04 6.15 ;
      RECT 84.75 5.95 85.21 6.12 ;
      RECT 83.76 2.73 84.05 2.96 ;
      RECT 83.76 2.76 84.22 2.93 ;
      RECT 83.825 1.655 83.99 2.96 ;
      RECT 82.34 1.625 82.63 1.855 ;
      RECT 82.34 1.655 83.99 1.825 ;
      RECT 82.4 0.885 82.57 1.855 ;
      RECT 82.34 0.885 82.63 1.115 ;
      RECT 82.34 7.765 82.63 7.995 ;
      RECT 82.4 7.025 82.57 7.995 ;
      RECT 82.4 7.12 83.99 7.29 ;
      RECT 83.82 5.92 83.99 7.29 ;
      RECT 82.34 7.025 82.63 7.255 ;
      RECT 83.76 5.92 84.05 6.15 ;
      RECT 83.76 5.95 84.22 6.12 ;
      RECT 80.325 1.995 80.65 2.32 ;
      RECT 82.77 1.965 83.12 2.315 ;
      RECT 80.325 2.025 83.12 2.195 ;
      RECT 82.795 6.655 83.12 6.98 ;
      RECT 82.77 6.655 83.12 6.885 ;
      RECT 82.6 6.685 83.12 6.855 ;
      RECT 81.995 2.365 82.315 2.685 ;
      RECT 81.965 2.365 82.315 2.595 ;
      RECT 81.68 2.395 82.315 2.565 ;
      RECT 81.995 6.28 82.315 6.605 ;
      RECT 81.965 6.285 82.315 6.515 ;
      RECT 81.795 6.315 82.315 6.485 ;
      RECT 79.74 3.185 80.065 3.51 ;
      RECT 76.945 3.11 77.265 3.37 ;
      RECT 78.915 3.12 79.205 3.35 ;
      RECT 79.64 3.185 80.065 3.325 ;
      RECT 76.945 3.17 79.78 3.31 ;
      RECT 79.325 2.77 79.645 3.03 ;
      RECT 79.045 2.83 79.645 2.97 ;
      RECT 78.305 5.83 78.625 6.09 ;
      RECT 78.305 5.89 78.895 6.03 ;
      RECT 77.625 2.77 77.945 3.03 ;
      RECT 72.885 2.78 73.175 3.01 ;
      RECT 72.885 2.83 77.945 2.97 ;
      RECT 77.715 2.49 77.855 3.03 ;
      RECT 77.715 2.49 78.195 2.63 ;
      RECT 78.055 2.1 78.195 2.63 ;
      RECT 77.975 2.1 78.265 2.33 ;
      RECT 77.625 3.79 77.945 4.05 ;
      RECT 76.955 3.8 77.245 4.03 ;
      RECT 74.745 3.8 75.035 4.03 ;
      RECT 74.745 3.85 77.945 3.99 ;
      RECT 75.925 5.83 76.245 6.09 ;
      RECT 77.635 5.84 77.925 6.07 ;
      RECT 75.255 5.84 75.545 6.07 ;
      RECT 75.255 5.89 76.245 6.03 ;
      RECT 77.715 5.55 77.855 6.07 ;
      RECT 76.015 5.55 76.155 6.09 ;
      RECT 76.015 5.55 77.855 5.69 ;
      RECT 74.915 2.44 75.205 2.67 ;
      RECT 74.995 2.15 75.135 2.67 ;
      RECT 77.285 2.09 77.605 2.35 ;
      RECT 77.185 2.1 77.605 2.33 ;
      RECT 74.995 2.15 77.605 2.29 ;
      RECT 76.265 2.43 76.585 2.69 ;
      RECT 76.265 2.49 76.855 2.63 ;
      RECT 76.265 4.81 76.585 5.07 ;
      RECT 73.555 4.82 73.845 5.05 ;
      RECT 73.555 4.87 76.585 5.01 ;
      RECT 75.585 2.39 75.915 2.72 ;
      RECT 75.585 2.44 76.045 2.67 ;
      RECT 75.585 2.49 76.065 2.63 ;
      RECT 75.465 2.49 75.475 2.63 ;
      RECT 75.475 2.48 76.045 2.62 ;
      RECT 71.575 6.63 71.915 6.91 ;
      RECT 71.545 6.655 71.915 6.885 ;
      RECT 71.375 6.685 71.915 6.855 ;
      RECT 71.115 7.765 71.405 7.995 ;
      RECT 71.175 6.995 71.345 7.995 ;
      RECT 71.075 6.995 71.445 7.365 ;
      RECT 68.54 7.77 68.83 8 ;
      RECT 68.6 6.29 68.77 8 ;
      RECT 68.6 6.655 68.93 6.98 ;
      RECT 68.54 6.29 68.83 6.52 ;
      RECT 68.135 2.395 68.24 2.965 ;
      RECT 68.135 2.73 68.46 2.96 ;
      RECT 68.135 2.76 68.63 2.93 ;
      RECT 68.135 2.395 68.325 2.96 ;
      RECT 67.55 2.36 67.84 2.59 ;
      RECT 67.55 2.395 68.325 2.565 ;
      RECT 67.61 0.88 67.78 2.59 ;
      RECT 67.55 0.88 67.84 1.11 ;
      RECT 67.55 7.77 67.84 8 ;
      RECT 67.61 6.29 67.78 8 ;
      RECT 67.55 6.29 67.84 6.52 ;
      RECT 67.55 6.325 68.405 6.485 ;
      RECT 68.235 5.92 68.405 6.485 ;
      RECT 67.55 6.32 67.945 6.485 ;
      RECT 68.17 5.92 68.46 6.15 ;
      RECT 68.17 5.95 68.63 6.12 ;
      RECT 67.18 2.73 67.47 2.96 ;
      RECT 67.18 2.76 67.64 2.93 ;
      RECT 67.245 1.655 67.41 2.96 ;
      RECT 65.76 1.625 66.05 1.855 ;
      RECT 65.76 1.655 67.41 1.825 ;
      RECT 65.82 0.885 65.99 1.855 ;
      RECT 65.76 0.885 66.05 1.115 ;
      RECT 65.76 7.765 66.05 7.995 ;
      RECT 65.82 7.025 65.99 7.995 ;
      RECT 65.82 7.12 67.41 7.29 ;
      RECT 67.24 5.92 67.41 7.29 ;
      RECT 65.76 7.025 66.05 7.255 ;
      RECT 67.18 5.92 67.47 6.15 ;
      RECT 67.18 5.95 67.64 6.12 ;
      RECT 63.745 1.995 64.07 2.32 ;
      RECT 66.19 1.965 66.54 2.315 ;
      RECT 63.745 2.025 66.54 2.195 ;
      RECT 66.215 6.655 66.54 6.98 ;
      RECT 66.19 6.655 66.54 6.885 ;
      RECT 66.02 6.685 66.54 6.855 ;
      RECT 65.415 2.365 65.735 2.685 ;
      RECT 65.385 2.365 65.735 2.595 ;
      RECT 65.1 2.395 65.735 2.565 ;
      RECT 65.415 6.28 65.735 6.605 ;
      RECT 65.385 6.285 65.735 6.515 ;
      RECT 65.215 6.315 65.735 6.485 ;
      RECT 63.16 3.185 63.485 3.51 ;
      RECT 60.365 3.11 60.685 3.37 ;
      RECT 62.335 3.12 62.625 3.35 ;
      RECT 63.06 3.185 63.485 3.325 ;
      RECT 60.365 3.17 63.2 3.31 ;
      RECT 62.745 2.77 63.065 3.03 ;
      RECT 62.465 2.83 63.065 2.97 ;
      RECT 61.725 5.83 62.045 6.09 ;
      RECT 61.725 5.89 62.315 6.03 ;
      RECT 61.045 2.77 61.365 3.03 ;
      RECT 56.305 2.78 56.595 3.01 ;
      RECT 56.305 2.83 61.365 2.97 ;
      RECT 61.135 2.49 61.275 3.03 ;
      RECT 61.135 2.49 61.615 2.63 ;
      RECT 61.475 2.1 61.615 2.63 ;
      RECT 61.395 2.1 61.685 2.33 ;
      RECT 61.045 3.79 61.365 4.05 ;
      RECT 60.375 3.8 60.665 4.03 ;
      RECT 58.165 3.8 58.455 4.03 ;
      RECT 58.165 3.85 61.365 3.99 ;
      RECT 59.345 5.83 59.665 6.09 ;
      RECT 61.055 5.84 61.345 6.07 ;
      RECT 58.675 5.84 58.965 6.07 ;
      RECT 58.675 5.89 59.665 6.03 ;
      RECT 61.135 5.55 61.275 6.07 ;
      RECT 59.435 5.55 59.575 6.09 ;
      RECT 59.435 5.55 61.275 5.69 ;
      RECT 58.335 2.44 58.625 2.67 ;
      RECT 58.415 2.15 58.555 2.67 ;
      RECT 60.705 2.09 61.025 2.35 ;
      RECT 60.605 2.1 61.025 2.33 ;
      RECT 58.415 2.15 61.025 2.29 ;
      RECT 59.685 2.43 60.005 2.69 ;
      RECT 59.685 2.49 60.275 2.63 ;
      RECT 59.685 4.81 60.005 5.07 ;
      RECT 56.975 4.82 57.265 5.05 ;
      RECT 56.975 4.87 60.005 5.01 ;
      RECT 59.005 2.39 59.335 2.72 ;
      RECT 59.005 2.44 59.465 2.67 ;
      RECT 59.005 2.49 59.485 2.63 ;
      RECT 58.885 2.49 58.895 2.63 ;
      RECT 58.895 2.48 59.465 2.62 ;
      RECT 54.995 6.63 55.335 6.91 ;
      RECT 54.965 6.655 55.335 6.885 ;
      RECT 54.795 6.685 55.335 6.855 ;
      RECT 54.535 7.765 54.825 7.995 ;
      RECT 54.595 6.995 54.765 7.995 ;
      RECT 54.495 6.995 54.865 7.365 ;
      RECT 51.955 7.77 52.245 8 ;
      RECT 52.015 6.29 52.185 8 ;
      RECT 52.015 6.655 52.345 6.98 ;
      RECT 51.955 6.29 52.245 6.52 ;
      RECT 51.55 2.395 51.655 2.965 ;
      RECT 51.55 2.73 51.875 2.96 ;
      RECT 51.55 2.76 52.045 2.93 ;
      RECT 51.55 2.395 51.74 2.96 ;
      RECT 50.965 2.36 51.255 2.59 ;
      RECT 50.965 2.395 51.74 2.565 ;
      RECT 51.025 0.88 51.195 2.59 ;
      RECT 50.965 0.88 51.255 1.11 ;
      RECT 50.965 7.77 51.255 8 ;
      RECT 51.025 6.29 51.195 8 ;
      RECT 50.965 6.29 51.255 6.52 ;
      RECT 50.965 6.325 51.82 6.485 ;
      RECT 51.65 5.92 51.82 6.485 ;
      RECT 50.965 6.32 51.36 6.485 ;
      RECT 51.585 5.92 51.875 6.15 ;
      RECT 51.585 5.95 52.045 6.12 ;
      RECT 50.595 2.73 50.885 2.96 ;
      RECT 50.595 2.76 51.055 2.93 ;
      RECT 50.66 1.655 50.825 2.96 ;
      RECT 49.175 1.625 49.465 1.855 ;
      RECT 49.175 1.655 50.825 1.825 ;
      RECT 49.235 0.885 49.405 1.855 ;
      RECT 49.175 0.885 49.465 1.115 ;
      RECT 49.175 7.765 49.465 7.995 ;
      RECT 49.235 7.025 49.405 7.995 ;
      RECT 49.235 7.12 50.825 7.29 ;
      RECT 50.655 5.92 50.825 7.29 ;
      RECT 49.175 7.025 49.465 7.255 ;
      RECT 50.595 5.92 50.885 6.15 ;
      RECT 50.595 5.95 51.055 6.12 ;
      RECT 47.16 1.995 47.485 2.32 ;
      RECT 49.605 1.965 49.955 2.315 ;
      RECT 47.16 2.025 49.955 2.195 ;
      RECT 49.63 6.655 49.955 6.98 ;
      RECT 49.605 6.655 49.955 6.885 ;
      RECT 49.435 6.685 49.955 6.855 ;
      RECT 48.83 2.365 49.15 2.685 ;
      RECT 48.8 2.365 49.15 2.595 ;
      RECT 48.515 2.395 49.15 2.565 ;
      RECT 48.83 6.28 49.15 6.605 ;
      RECT 48.8 6.285 49.15 6.515 ;
      RECT 48.63 6.315 49.15 6.485 ;
      RECT 46.575 3.185 46.9 3.51 ;
      RECT 43.78 3.11 44.1 3.37 ;
      RECT 45.75 3.12 46.04 3.35 ;
      RECT 46.475 3.185 46.9 3.325 ;
      RECT 43.78 3.17 46.615 3.31 ;
      RECT 46.16 2.77 46.48 3.03 ;
      RECT 45.88 2.83 46.48 2.97 ;
      RECT 45.14 5.83 45.46 6.09 ;
      RECT 45.14 5.89 45.73 6.03 ;
      RECT 44.46 2.77 44.78 3.03 ;
      RECT 39.72 2.78 40.01 3.01 ;
      RECT 39.72 2.83 44.78 2.97 ;
      RECT 44.55 2.49 44.69 3.03 ;
      RECT 44.55 2.49 45.03 2.63 ;
      RECT 44.89 2.1 45.03 2.63 ;
      RECT 44.81 2.1 45.1 2.33 ;
      RECT 44.46 3.79 44.78 4.05 ;
      RECT 43.79 3.8 44.08 4.03 ;
      RECT 41.58 3.8 41.87 4.03 ;
      RECT 41.58 3.85 44.78 3.99 ;
      RECT 42.76 5.83 43.08 6.09 ;
      RECT 44.47 5.84 44.76 6.07 ;
      RECT 42.09 5.84 42.38 6.07 ;
      RECT 42.09 5.89 43.08 6.03 ;
      RECT 44.55 5.55 44.69 6.07 ;
      RECT 42.85 5.55 42.99 6.09 ;
      RECT 42.85 5.55 44.69 5.69 ;
      RECT 41.75 2.44 42.04 2.67 ;
      RECT 41.83 2.15 41.97 2.67 ;
      RECT 44.12 2.09 44.44 2.35 ;
      RECT 44.02 2.1 44.44 2.33 ;
      RECT 41.83 2.15 44.44 2.29 ;
      RECT 43.1 2.43 43.42 2.69 ;
      RECT 43.1 2.49 43.69 2.63 ;
      RECT 43.1 4.81 43.42 5.07 ;
      RECT 40.39 4.82 40.68 5.05 ;
      RECT 40.39 4.87 43.42 5.01 ;
      RECT 42.42 2.39 42.75 2.72 ;
      RECT 42.42 2.44 42.88 2.67 ;
      RECT 42.42 2.49 42.9 2.63 ;
      RECT 42.3 2.49 42.31 2.63 ;
      RECT 42.31 2.48 42.88 2.62 ;
      RECT 38.41 6.63 38.75 6.91 ;
      RECT 38.38 6.655 38.75 6.885 ;
      RECT 38.21 6.685 38.75 6.855 ;
      RECT 37.95 7.765 38.24 7.995 ;
      RECT 38.01 6.995 38.18 7.995 ;
      RECT 37.91 6.995 38.28 7.365 ;
      RECT 35.37 7.77 35.66 8 ;
      RECT 35.43 6.29 35.6 8 ;
      RECT 35.43 6.655 35.76 6.98 ;
      RECT 35.37 6.29 35.66 6.52 ;
      RECT 34.965 2.395 35.07 2.965 ;
      RECT 34.965 2.73 35.29 2.96 ;
      RECT 34.965 2.76 35.46 2.93 ;
      RECT 34.965 2.395 35.155 2.96 ;
      RECT 34.38 2.36 34.67 2.59 ;
      RECT 34.38 2.395 35.155 2.565 ;
      RECT 34.44 0.88 34.61 2.59 ;
      RECT 34.38 0.88 34.67 1.11 ;
      RECT 34.38 7.77 34.67 8 ;
      RECT 34.44 6.29 34.61 8 ;
      RECT 34.38 6.29 34.67 6.52 ;
      RECT 34.38 6.325 35.235 6.485 ;
      RECT 35.065 5.92 35.235 6.485 ;
      RECT 34.38 6.32 34.775 6.485 ;
      RECT 35 5.92 35.29 6.15 ;
      RECT 35 5.95 35.46 6.12 ;
      RECT 34.01 2.73 34.3 2.96 ;
      RECT 34.01 2.76 34.47 2.93 ;
      RECT 34.075 1.655 34.24 2.96 ;
      RECT 32.59 1.625 32.88 1.855 ;
      RECT 32.59 1.655 34.24 1.825 ;
      RECT 32.65 0.885 32.82 1.855 ;
      RECT 32.59 0.885 32.88 1.115 ;
      RECT 32.59 7.765 32.88 7.995 ;
      RECT 32.65 7.025 32.82 7.995 ;
      RECT 32.65 7.12 34.24 7.29 ;
      RECT 34.07 5.92 34.24 7.29 ;
      RECT 32.59 7.025 32.88 7.255 ;
      RECT 34.01 5.92 34.3 6.15 ;
      RECT 34.01 5.95 34.47 6.12 ;
      RECT 30.575 1.995 30.9 2.32 ;
      RECT 33.02 1.965 33.37 2.315 ;
      RECT 30.575 2.025 33.37 2.195 ;
      RECT 33.045 6.655 33.37 6.98 ;
      RECT 33.02 6.655 33.37 6.885 ;
      RECT 32.85 6.685 33.37 6.855 ;
      RECT 32.245 2.365 32.565 2.685 ;
      RECT 32.215 2.365 32.565 2.595 ;
      RECT 31.93 2.395 32.565 2.565 ;
      RECT 32.245 6.28 32.565 6.605 ;
      RECT 32.215 6.285 32.565 6.515 ;
      RECT 32.045 6.315 32.565 6.485 ;
      RECT 29.99 3.185 30.315 3.51 ;
      RECT 27.195 3.11 27.515 3.37 ;
      RECT 29.165 3.12 29.455 3.35 ;
      RECT 29.89 3.185 30.315 3.325 ;
      RECT 27.195 3.17 30.03 3.31 ;
      RECT 29.575 2.77 29.895 3.03 ;
      RECT 29.295 2.83 29.895 2.97 ;
      RECT 28.555 5.83 28.875 6.09 ;
      RECT 28.555 5.89 29.145 6.03 ;
      RECT 27.875 2.77 28.195 3.03 ;
      RECT 23.135 2.78 23.425 3.01 ;
      RECT 23.135 2.83 28.195 2.97 ;
      RECT 27.965 2.49 28.105 3.03 ;
      RECT 27.965 2.49 28.445 2.63 ;
      RECT 28.305 2.1 28.445 2.63 ;
      RECT 28.225 2.1 28.515 2.33 ;
      RECT 27.875 3.79 28.195 4.05 ;
      RECT 27.205 3.8 27.495 4.03 ;
      RECT 24.995 3.8 25.285 4.03 ;
      RECT 24.995 3.85 28.195 3.99 ;
      RECT 26.175 5.83 26.495 6.09 ;
      RECT 27.885 5.84 28.175 6.07 ;
      RECT 25.505 5.84 25.795 6.07 ;
      RECT 25.505 5.89 26.495 6.03 ;
      RECT 27.965 5.55 28.105 6.07 ;
      RECT 26.265 5.55 26.405 6.09 ;
      RECT 26.265 5.55 28.105 5.69 ;
      RECT 25.165 2.44 25.455 2.67 ;
      RECT 25.245 2.15 25.385 2.67 ;
      RECT 27.535 2.09 27.855 2.35 ;
      RECT 27.435 2.1 27.855 2.33 ;
      RECT 25.245 2.15 27.855 2.29 ;
      RECT 26.515 2.43 26.835 2.69 ;
      RECT 26.515 2.49 27.105 2.63 ;
      RECT 26.515 4.81 26.835 5.07 ;
      RECT 23.805 4.82 24.095 5.05 ;
      RECT 23.805 4.87 26.835 5.01 ;
      RECT 25.835 2.39 26.165 2.72 ;
      RECT 25.835 2.44 26.295 2.67 ;
      RECT 25.835 2.49 26.315 2.63 ;
      RECT 25.715 2.49 25.725 2.63 ;
      RECT 25.725 2.48 26.295 2.62 ;
      RECT 21.825 6.63 22.165 6.91 ;
      RECT 21.795 6.655 22.165 6.885 ;
      RECT 21.625 6.685 22.165 6.855 ;
      RECT 21.365 7.765 21.655 7.995 ;
      RECT 21.425 6.995 21.595 7.995 ;
      RECT 21.325 6.995 21.695 7.365 ;
      RECT 18.785 7.77 19.075 8 ;
      RECT 18.845 6.29 19.015 8 ;
      RECT 18.845 6.655 19.175 6.98 ;
      RECT 18.785 6.29 19.075 6.52 ;
      RECT 18.38 2.395 18.485 2.965 ;
      RECT 18.38 2.73 18.705 2.96 ;
      RECT 18.38 2.76 18.875 2.93 ;
      RECT 18.38 2.395 18.57 2.96 ;
      RECT 17.795 2.36 18.085 2.59 ;
      RECT 17.795 2.395 18.57 2.565 ;
      RECT 17.855 0.88 18.025 2.59 ;
      RECT 17.795 0.88 18.085 1.11 ;
      RECT 17.795 7.77 18.085 8 ;
      RECT 17.855 6.29 18.025 8 ;
      RECT 17.795 6.29 18.085 6.52 ;
      RECT 17.795 6.325 18.65 6.485 ;
      RECT 18.48 5.92 18.65 6.485 ;
      RECT 17.795 6.32 18.19 6.485 ;
      RECT 18.415 5.92 18.705 6.15 ;
      RECT 18.415 5.95 18.875 6.12 ;
      RECT 17.425 2.73 17.715 2.96 ;
      RECT 17.425 2.76 17.885 2.93 ;
      RECT 17.49 1.655 17.655 2.96 ;
      RECT 16.005 1.625 16.295 1.855 ;
      RECT 16.005 1.655 17.655 1.825 ;
      RECT 16.065 0.885 16.235 1.855 ;
      RECT 16.005 0.885 16.295 1.115 ;
      RECT 16.005 7.765 16.295 7.995 ;
      RECT 16.065 7.025 16.235 7.995 ;
      RECT 16.065 7.12 17.655 7.29 ;
      RECT 17.485 5.92 17.655 7.29 ;
      RECT 16.005 7.025 16.295 7.255 ;
      RECT 17.425 5.92 17.715 6.15 ;
      RECT 17.425 5.95 17.885 6.12 ;
      RECT 13.99 1.995 14.315 2.32 ;
      RECT 16.435 1.965 16.785 2.315 ;
      RECT 13.99 2.025 16.785 2.195 ;
      RECT 16.46 6.655 16.785 6.98 ;
      RECT 16.435 6.655 16.785 6.885 ;
      RECT 16.265 6.685 16.785 6.855 ;
      RECT 15.66 2.365 15.98 2.685 ;
      RECT 15.63 2.365 15.98 2.595 ;
      RECT 15.345 2.395 15.98 2.565 ;
      RECT 15.66 6.28 15.98 6.605 ;
      RECT 15.63 6.285 15.98 6.515 ;
      RECT 15.46 6.315 15.98 6.485 ;
      RECT 13.405 3.185 13.73 3.51 ;
      RECT 10.61 3.11 10.93 3.37 ;
      RECT 12.58 3.12 12.87 3.35 ;
      RECT 13.305 3.185 13.73 3.325 ;
      RECT 10.61 3.17 13.445 3.31 ;
      RECT 12.99 2.77 13.31 3.03 ;
      RECT 12.71 2.83 13.31 2.97 ;
      RECT 11.97 5.83 12.29 6.09 ;
      RECT 11.97 5.89 12.56 6.03 ;
      RECT 11.29 2.77 11.61 3.03 ;
      RECT 6.55 2.78 6.84 3.01 ;
      RECT 6.55 2.83 11.61 2.97 ;
      RECT 11.38 2.49 11.52 3.03 ;
      RECT 11.38 2.49 11.86 2.63 ;
      RECT 11.72 2.1 11.86 2.63 ;
      RECT 11.64 2.1 11.93 2.33 ;
      RECT 11.29 3.79 11.61 4.05 ;
      RECT 10.62 3.8 10.91 4.03 ;
      RECT 8.41 3.8 8.7 4.03 ;
      RECT 8.41 3.85 11.61 3.99 ;
      RECT 9.59 5.83 9.91 6.09 ;
      RECT 11.3 5.84 11.59 6.07 ;
      RECT 8.92 5.84 9.21 6.07 ;
      RECT 8.92 5.89 9.91 6.03 ;
      RECT 11.38 5.55 11.52 6.07 ;
      RECT 9.68 5.55 9.82 6.09 ;
      RECT 9.68 5.55 11.52 5.69 ;
      RECT 8.58 2.44 8.87 2.67 ;
      RECT 8.66 2.15 8.8 2.67 ;
      RECT 10.95 2.09 11.27 2.35 ;
      RECT 10.85 2.1 11.27 2.33 ;
      RECT 8.66 2.15 11.27 2.29 ;
      RECT 9.93 2.43 10.25 2.69 ;
      RECT 9.93 2.49 10.52 2.63 ;
      RECT 9.93 4.81 10.25 5.07 ;
      RECT 7.22 4.82 7.51 5.05 ;
      RECT 7.22 4.87 10.25 5.01 ;
      RECT 9.25 2.39 9.58 2.72 ;
      RECT 9.25 2.44 9.71 2.67 ;
      RECT 9.25 2.49 9.73 2.63 ;
      RECT 9.13 2.49 9.14 2.63 ;
      RECT 9.14 2.48 9.71 2.62 ;
      RECT 5.24 6.63 5.58 6.91 ;
      RECT 5.21 6.655 5.58 6.885 ;
      RECT 5.04 6.685 5.58 6.855 ;
      RECT 4.78 7.765 5.07 7.995 ;
      RECT 4.84 6.995 5.01 7.995 ;
      RECT 4.74 6.995 5.11 7.365 ;
      RECT 1.55 7.765 1.84 7.995 ;
      RECT 1.61 7.025 1.78 7.995 ;
      RECT 1.52 7.025 1.86 7.305 ;
      RECT 1.145 6.285 1.485 6.565 ;
      RECT 1.005 6.315 1.485 6.485 ;
      RECT 78.995 4.81 79.645 5.07 ;
      RECT 76.945 5.83 77.265 6.09 ;
      RECT 62.415 4.81 63.065 5.07 ;
      RECT 60.365 5.83 60.685 6.09 ;
      RECT 45.83 4.81 46.48 5.07 ;
      RECT 43.78 5.83 44.1 6.09 ;
      RECT 29.245 4.81 29.895 5.07 ;
      RECT 27.195 5.83 27.515 6.09 ;
      RECT 12.66 4.81 13.31 5.07 ;
      RECT 10.61 5.83 10.93 6.09 ;
    LAYER mcon ;
      RECT 85.18 6.32 85.35 6.49 ;
      RECT 85.185 6.315 85.355 6.485 ;
      RECT 68.6 6.32 68.77 6.49 ;
      RECT 68.605 6.315 68.775 6.485 ;
      RECT 52.015 6.32 52.185 6.49 ;
      RECT 52.02 6.315 52.19 6.485 ;
      RECT 35.43 6.32 35.6 6.49 ;
      RECT 35.435 6.315 35.605 6.485 ;
      RECT 18.845 6.32 19.015 6.49 ;
      RECT 18.85 6.315 19.02 6.485 ;
      RECT 85.18 7.8 85.35 7.97 ;
      RECT 84.81 2.76 84.98 2.93 ;
      RECT 84.81 5.95 84.98 6.12 ;
      RECT 84.19 0.91 84.36 1.08 ;
      RECT 84.19 2.39 84.36 2.56 ;
      RECT 84.19 6.32 84.36 6.49 ;
      RECT 84.19 7.8 84.36 7.97 ;
      RECT 83.82 2.76 83.99 2.93 ;
      RECT 83.82 5.95 83.99 6.12 ;
      RECT 82.83 2.025 83 2.195 ;
      RECT 82.83 6.685 83 6.855 ;
      RECT 82.4 0.915 82.57 1.085 ;
      RECT 82.4 1.655 82.57 1.825 ;
      RECT 82.4 7.055 82.57 7.225 ;
      RECT 82.4 7.795 82.57 7.965 ;
      RECT 82.025 2.395 82.195 2.565 ;
      RECT 82.025 6.315 82.195 6.485 ;
      RECT 79.395 2.81 79.565 2.98 ;
      RECT 79.055 4.85 79.225 5.02 ;
      RECT 78.975 3.15 79.145 3.32 ;
      RECT 78.375 5.87 78.545 6.04 ;
      RECT 78.035 2.13 78.205 2.3 ;
      RECT 77.695 5.87 77.865 6.04 ;
      RECT 77.245 2.13 77.415 2.3 ;
      RECT 77.015 3.83 77.185 4 ;
      RECT 77.015 5.87 77.185 6.04 ;
      RECT 76.335 2.47 76.505 2.64 ;
      RECT 75.815 2.47 75.985 2.64 ;
      RECT 75.315 5.87 75.485 6.04 ;
      RECT 74.975 2.47 75.145 2.64 ;
      RECT 74.805 3.83 74.975 4 ;
      RECT 73.615 4.85 73.785 5.02 ;
      RECT 72.945 2.81 73.115 2.98 ;
      RECT 71.605 6.685 71.775 6.855 ;
      RECT 71.175 7.055 71.345 7.225 ;
      RECT 71.175 7.795 71.345 7.965 ;
      RECT 68.6 7.8 68.77 7.97 ;
      RECT 68.23 2.76 68.4 2.93 ;
      RECT 68.23 5.95 68.4 6.12 ;
      RECT 67.61 0.91 67.78 1.08 ;
      RECT 67.61 2.39 67.78 2.56 ;
      RECT 67.61 6.32 67.78 6.49 ;
      RECT 67.61 7.8 67.78 7.97 ;
      RECT 67.24 2.76 67.41 2.93 ;
      RECT 67.24 5.95 67.41 6.12 ;
      RECT 66.25 2.025 66.42 2.195 ;
      RECT 66.25 6.685 66.42 6.855 ;
      RECT 65.82 0.915 65.99 1.085 ;
      RECT 65.82 1.655 65.99 1.825 ;
      RECT 65.82 7.055 65.99 7.225 ;
      RECT 65.82 7.795 65.99 7.965 ;
      RECT 65.445 2.395 65.615 2.565 ;
      RECT 65.445 6.315 65.615 6.485 ;
      RECT 62.815 2.81 62.985 2.98 ;
      RECT 62.475 4.85 62.645 5.02 ;
      RECT 62.395 3.15 62.565 3.32 ;
      RECT 61.795 5.87 61.965 6.04 ;
      RECT 61.455 2.13 61.625 2.3 ;
      RECT 61.115 5.87 61.285 6.04 ;
      RECT 60.665 2.13 60.835 2.3 ;
      RECT 60.435 3.83 60.605 4 ;
      RECT 60.435 5.87 60.605 6.04 ;
      RECT 59.755 2.47 59.925 2.64 ;
      RECT 59.235 2.47 59.405 2.64 ;
      RECT 58.735 5.87 58.905 6.04 ;
      RECT 58.395 2.47 58.565 2.64 ;
      RECT 58.225 3.83 58.395 4 ;
      RECT 57.035 4.85 57.205 5.02 ;
      RECT 56.365 2.81 56.535 2.98 ;
      RECT 55.025 6.685 55.195 6.855 ;
      RECT 54.595 7.055 54.765 7.225 ;
      RECT 54.595 7.795 54.765 7.965 ;
      RECT 52.015 7.8 52.185 7.97 ;
      RECT 51.645 2.76 51.815 2.93 ;
      RECT 51.645 5.95 51.815 6.12 ;
      RECT 51.025 0.91 51.195 1.08 ;
      RECT 51.025 2.39 51.195 2.56 ;
      RECT 51.025 6.32 51.195 6.49 ;
      RECT 51.025 7.8 51.195 7.97 ;
      RECT 50.655 2.76 50.825 2.93 ;
      RECT 50.655 5.95 50.825 6.12 ;
      RECT 49.665 2.025 49.835 2.195 ;
      RECT 49.665 6.685 49.835 6.855 ;
      RECT 49.235 0.915 49.405 1.085 ;
      RECT 49.235 1.655 49.405 1.825 ;
      RECT 49.235 7.055 49.405 7.225 ;
      RECT 49.235 7.795 49.405 7.965 ;
      RECT 48.86 2.395 49.03 2.565 ;
      RECT 48.86 6.315 49.03 6.485 ;
      RECT 46.23 2.81 46.4 2.98 ;
      RECT 45.89 4.85 46.06 5.02 ;
      RECT 45.81 3.15 45.98 3.32 ;
      RECT 45.21 5.87 45.38 6.04 ;
      RECT 44.87 2.13 45.04 2.3 ;
      RECT 44.53 5.87 44.7 6.04 ;
      RECT 44.08 2.13 44.25 2.3 ;
      RECT 43.85 3.83 44.02 4 ;
      RECT 43.85 5.87 44.02 6.04 ;
      RECT 43.17 2.47 43.34 2.64 ;
      RECT 42.65 2.47 42.82 2.64 ;
      RECT 42.15 5.87 42.32 6.04 ;
      RECT 41.81 2.47 41.98 2.64 ;
      RECT 41.64 3.83 41.81 4 ;
      RECT 40.45 4.85 40.62 5.02 ;
      RECT 39.78 2.81 39.95 2.98 ;
      RECT 38.44 6.685 38.61 6.855 ;
      RECT 38.01 7.055 38.18 7.225 ;
      RECT 38.01 7.795 38.18 7.965 ;
      RECT 35.43 7.8 35.6 7.97 ;
      RECT 35.06 2.76 35.23 2.93 ;
      RECT 35.06 5.95 35.23 6.12 ;
      RECT 34.44 0.91 34.61 1.08 ;
      RECT 34.44 2.39 34.61 2.56 ;
      RECT 34.44 6.32 34.61 6.49 ;
      RECT 34.44 7.8 34.61 7.97 ;
      RECT 34.07 2.76 34.24 2.93 ;
      RECT 34.07 5.95 34.24 6.12 ;
      RECT 33.08 2.025 33.25 2.195 ;
      RECT 33.08 6.685 33.25 6.855 ;
      RECT 32.65 0.915 32.82 1.085 ;
      RECT 32.65 1.655 32.82 1.825 ;
      RECT 32.65 7.055 32.82 7.225 ;
      RECT 32.65 7.795 32.82 7.965 ;
      RECT 32.275 2.395 32.445 2.565 ;
      RECT 32.275 6.315 32.445 6.485 ;
      RECT 29.645 2.81 29.815 2.98 ;
      RECT 29.305 4.85 29.475 5.02 ;
      RECT 29.225 3.15 29.395 3.32 ;
      RECT 28.625 5.87 28.795 6.04 ;
      RECT 28.285 2.13 28.455 2.3 ;
      RECT 27.945 5.87 28.115 6.04 ;
      RECT 27.495 2.13 27.665 2.3 ;
      RECT 27.265 3.83 27.435 4 ;
      RECT 27.265 5.87 27.435 6.04 ;
      RECT 26.585 2.47 26.755 2.64 ;
      RECT 26.065 2.47 26.235 2.64 ;
      RECT 25.565 5.87 25.735 6.04 ;
      RECT 25.225 2.47 25.395 2.64 ;
      RECT 25.055 3.83 25.225 4 ;
      RECT 23.865 4.85 24.035 5.02 ;
      RECT 23.195 2.81 23.365 2.98 ;
      RECT 21.855 6.685 22.025 6.855 ;
      RECT 21.425 7.055 21.595 7.225 ;
      RECT 21.425 7.795 21.595 7.965 ;
      RECT 18.845 7.8 19.015 7.97 ;
      RECT 18.475 2.76 18.645 2.93 ;
      RECT 18.475 5.95 18.645 6.12 ;
      RECT 17.855 0.91 18.025 1.08 ;
      RECT 17.855 2.39 18.025 2.56 ;
      RECT 17.855 6.32 18.025 6.49 ;
      RECT 17.855 7.8 18.025 7.97 ;
      RECT 17.485 2.76 17.655 2.93 ;
      RECT 17.485 5.95 17.655 6.12 ;
      RECT 16.495 2.025 16.665 2.195 ;
      RECT 16.495 6.685 16.665 6.855 ;
      RECT 16.065 0.915 16.235 1.085 ;
      RECT 16.065 1.655 16.235 1.825 ;
      RECT 16.065 7.055 16.235 7.225 ;
      RECT 16.065 7.795 16.235 7.965 ;
      RECT 15.69 2.395 15.86 2.565 ;
      RECT 15.69 6.315 15.86 6.485 ;
      RECT 13.06 2.81 13.23 2.98 ;
      RECT 12.72 4.85 12.89 5.02 ;
      RECT 12.64 3.15 12.81 3.32 ;
      RECT 12.04 5.87 12.21 6.04 ;
      RECT 11.7 2.13 11.87 2.3 ;
      RECT 11.36 5.87 11.53 6.04 ;
      RECT 10.91 2.13 11.08 2.3 ;
      RECT 10.68 3.83 10.85 4 ;
      RECT 10.68 5.87 10.85 6.04 ;
      RECT 10 2.47 10.17 2.64 ;
      RECT 9.48 2.47 9.65 2.64 ;
      RECT 8.98 5.87 9.15 6.04 ;
      RECT 8.64 2.47 8.81 2.64 ;
      RECT 8.47 3.83 8.64 4 ;
      RECT 7.28 4.85 7.45 5.02 ;
      RECT 6.61 2.81 6.78 2.98 ;
      RECT 5.27 6.685 5.44 6.855 ;
      RECT 4.84 7.055 5.01 7.225 ;
      RECT 4.84 7.795 5.01 7.965 ;
      RECT 1.61 7.055 1.78 7.225 ;
      RECT 1.61 7.795 1.78 7.965 ;
      RECT 1.235 6.315 1.405 6.485 ;
    LAYER li1 ;
      RECT 85.18 5.02 85.35 6.49 ;
      RECT 85.18 6.315 85.355 6.485 ;
      RECT 84.81 1.74 84.98 2.93 ;
      RECT 84.81 1.74 85.28 1.91 ;
      RECT 84.81 6.97 85.28 7.14 ;
      RECT 84.81 5.95 84.98 7.14 ;
      RECT 83.82 1.74 83.99 2.93 ;
      RECT 83.82 1.74 84.29 1.91 ;
      RECT 83.82 6.97 84.29 7.14 ;
      RECT 83.82 5.95 83.99 7.14 ;
      RECT 81.97 2.635 82.14 3.865 ;
      RECT 82.025 0.855 82.195 2.805 ;
      RECT 81.97 0.575 82.14 1.025 ;
      RECT 81.97 7.855 82.14 8.305 ;
      RECT 82.025 6.075 82.195 8.025 ;
      RECT 81.97 5.015 82.14 6.245 ;
      RECT 81.45 0.575 81.62 3.865 ;
      RECT 81.45 2.075 81.855 2.405 ;
      RECT 81.45 1.235 81.855 1.565 ;
      RECT 81.45 5.015 81.62 8.305 ;
      RECT 81.45 7.315 81.855 7.645 ;
      RECT 81.45 6.475 81.855 6.805 ;
      RECT 76.705 6.64 78.015 6.89 ;
      RECT 76.705 6.32 76.885 6.89 ;
      RECT 76.155 6.32 76.885 6.49 ;
      RECT 76.155 5.48 76.325 6.49 ;
      RECT 76.995 5.52 78.735 5.7 ;
      RECT 78.405 4.68 78.735 5.7 ;
      RECT 76.155 5.48 77.215 5.65 ;
      RECT 78.405 4.85 79.225 5.02 ;
      RECT 77.565 4.68 77.895 4.89 ;
      RECT 77.565 4.68 78.735 4.85 ;
      RECT 78.465 3.2 78.795 4.16 ;
      RECT 78.465 3.2 79.145 3.37 ;
      RECT 78.975 1.96 79.145 3.37 ;
      RECT 78.885 1.96 79.215 2.6 ;
      RECT 78.015 3.47 78.285 4.17 ;
      RECT 78.115 1.96 78.285 4.17 ;
      RECT 78.455 2.78 78.805 3.03 ;
      RECT 78.115 2.81 78.805 2.98 ;
      RECT 78.025 1.96 78.285 2.44 ;
      RECT 77.355 5.11 78.235 5.35 ;
      RECT 78.005 5.02 78.235 5.35 ;
      RECT 76.705 5.11 78.235 5.31 ;
      RECT 77.625 5.06 78.235 5.35 ;
      RECT 76.705 4.98 76.875 5.31 ;
      RECT 77.595 5.87 77.845 6.47 ;
      RECT 77.595 5.87 78.065 6.07 ;
      RECT 77.085 3.09 77.845 3.59 ;
      RECT 76.155 2.9 76.415 3.52 ;
      RECT 77.075 3.03 77.085 3.34 ;
      RECT 77.055 3.02 77.075 3.31 ;
      RECT 77.715 2.7 77.945 3.3 ;
      RECT 77.035 2.97 77.055 3.28 ;
      RECT 77.015 3.09 77.945 3.27 ;
      RECT 76.985 3.09 77.945 3.26 ;
      RECT 76.915 3.09 77.945 3.25 ;
      RECT 76.895 3.09 77.945 3.22 ;
      RECT 76.875 2 77.045 3.19 ;
      RECT 76.845 3.09 77.945 3.16 ;
      RECT 76.815 3.09 77.945 3.13 ;
      RECT 76.785 3.08 77.145 3.1 ;
      RECT 76.785 3.07 77.135 3.1 ;
      RECT 76.155 2.9 77.045 3.07 ;
      RECT 76.155 3.06 77.115 3.07 ;
      RECT 76.155 3.05 77.105 3.07 ;
      RECT 76.155 2.99 77.065 3.07 ;
      RECT 76.155 2 77.045 2.17 ;
      RECT 77.215 2.5 77.545 2.92 ;
      RECT 77.215 2.01 77.435 2.92 ;
      RECT 77.135 5.87 77.345 6.47 ;
      RECT 76.995 5.87 77.345 6.07 ;
      RECT 75.715 3.47 75.985 4.17 ;
      RECT 75.935 1.96 75.985 4.17 ;
      RECT 75.815 2.77 75.985 4.17 ;
      RECT 75.815 1.96 75.985 2.76 ;
      RECT 75.725 1.96 75.985 2.44 ;
      RECT 73.855 3.13 74.105 3.67 ;
      RECT 74.825 3.13 75.545 3.6 ;
      RECT 73.855 3.13 75.645 3.3 ;
      RECT 75.415 2.77 75.645 3.3 ;
      RECT 74.415 2.01 74.665 3.3 ;
      RECT 75.415 2.7 75.475 3.6 ;
      RECT 75.415 2.7 75.645 2.76 ;
      RECT 73.875 2.01 74.665 2.28 ;
      RECT 74.835 5.82 75.515 6.07 ;
      RECT 75.245 5.46 75.515 6.07 ;
      RECT 74.995 6.24 75.325 6.79 ;
      RECT 73.935 6.24 75.325 6.43 ;
      RECT 73.935 5.4 74.105 6.43 ;
      RECT 73.815 5.82 74.105 6.15 ;
      RECT 73.935 5.4 74.875 5.57 ;
      RECT 74.575 4.85 74.875 5.57 ;
      RECT 74.835 2.43 75.245 2.95 ;
      RECT 74.835 2.01 75.035 2.95 ;
      RECT 73.445 2.19 73.615 4.17 ;
      RECT 73.445 2.7 74.245 2.95 ;
      RECT 73.445 2.19 73.695 2.95 ;
      RECT 73.365 2.19 73.695 2.61 ;
      RECT 73.395 6.6 73.955 6.89 ;
      RECT 73.395 4.68 73.645 6.89 ;
      RECT 73.395 4.68 73.855 5.23 ;
      RECT 70.225 5.015 70.395 8.305 ;
      RECT 70.225 7.315 70.63 7.645 ;
      RECT 70.225 6.475 70.63 6.805 ;
      RECT 68.6 5.02 68.77 6.49 ;
      RECT 68.6 6.315 68.775 6.485 ;
      RECT 68.23 1.74 68.4 2.93 ;
      RECT 68.23 1.74 68.7 1.91 ;
      RECT 68.23 6.97 68.7 7.14 ;
      RECT 68.23 5.95 68.4 7.14 ;
      RECT 67.24 1.74 67.41 2.93 ;
      RECT 67.24 1.74 67.71 1.91 ;
      RECT 67.24 6.97 67.71 7.14 ;
      RECT 67.24 5.95 67.41 7.14 ;
      RECT 65.39 2.635 65.56 3.865 ;
      RECT 65.445 0.855 65.615 2.805 ;
      RECT 65.39 0.575 65.56 1.025 ;
      RECT 65.39 7.855 65.56 8.305 ;
      RECT 65.445 6.075 65.615 8.025 ;
      RECT 65.39 5.015 65.56 6.245 ;
      RECT 64.87 0.575 65.04 3.865 ;
      RECT 64.87 2.075 65.275 2.405 ;
      RECT 64.87 1.235 65.275 1.565 ;
      RECT 64.87 5.015 65.04 8.305 ;
      RECT 64.87 7.315 65.275 7.645 ;
      RECT 64.87 6.475 65.275 6.805 ;
      RECT 60.125 6.64 61.435 6.89 ;
      RECT 60.125 6.32 60.305 6.89 ;
      RECT 59.575 6.32 60.305 6.49 ;
      RECT 59.575 5.48 59.745 6.49 ;
      RECT 60.415 5.52 62.155 5.7 ;
      RECT 61.825 4.68 62.155 5.7 ;
      RECT 59.575 5.48 60.635 5.65 ;
      RECT 61.825 4.85 62.645 5.02 ;
      RECT 60.985 4.68 61.315 4.89 ;
      RECT 60.985 4.68 62.155 4.85 ;
      RECT 61.885 3.2 62.215 4.16 ;
      RECT 61.885 3.2 62.565 3.37 ;
      RECT 62.395 1.96 62.565 3.37 ;
      RECT 62.305 1.96 62.635 2.6 ;
      RECT 61.435 3.47 61.705 4.17 ;
      RECT 61.535 1.96 61.705 4.17 ;
      RECT 61.875 2.78 62.225 3.03 ;
      RECT 61.535 2.81 62.225 2.98 ;
      RECT 61.445 1.96 61.705 2.44 ;
      RECT 60.775 5.11 61.655 5.35 ;
      RECT 61.425 5.02 61.655 5.35 ;
      RECT 60.125 5.11 61.655 5.31 ;
      RECT 61.045 5.06 61.655 5.35 ;
      RECT 60.125 4.98 60.295 5.31 ;
      RECT 61.015 5.87 61.265 6.47 ;
      RECT 61.015 5.87 61.485 6.07 ;
      RECT 60.505 3.09 61.265 3.59 ;
      RECT 59.575 2.9 59.835 3.52 ;
      RECT 60.495 3.03 60.505 3.34 ;
      RECT 60.475 3.02 60.495 3.31 ;
      RECT 61.135 2.7 61.365 3.3 ;
      RECT 60.455 2.97 60.475 3.28 ;
      RECT 60.435 3.09 61.365 3.27 ;
      RECT 60.405 3.09 61.365 3.26 ;
      RECT 60.335 3.09 61.365 3.25 ;
      RECT 60.315 3.09 61.365 3.22 ;
      RECT 60.295 2 60.465 3.19 ;
      RECT 60.265 3.09 61.365 3.16 ;
      RECT 60.235 3.09 61.365 3.13 ;
      RECT 60.205 3.08 60.565 3.1 ;
      RECT 60.205 3.07 60.555 3.1 ;
      RECT 59.575 2.9 60.465 3.07 ;
      RECT 59.575 3.06 60.535 3.07 ;
      RECT 59.575 3.05 60.525 3.07 ;
      RECT 59.575 2.99 60.485 3.07 ;
      RECT 59.575 2 60.465 2.17 ;
      RECT 60.635 2.5 60.965 2.92 ;
      RECT 60.635 2.01 60.855 2.92 ;
      RECT 60.555 5.87 60.765 6.47 ;
      RECT 60.415 5.87 60.765 6.07 ;
      RECT 59.135 3.47 59.405 4.17 ;
      RECT 59.355 1.96 59.405 4.17 ;
      RECT 59.235 2.77 59.405 4.17 ;
      RECT 59.235 1.96 59.405 2.76 ;
      RECT 59.145 1.96 59.405 2.44 ;
      RECT 57.275 3.13 57.525 3.67 ;
      RECT 58.245 3.13 58.965 3.6 ;
      RECT 57.275 3.13 59.065 3.3 ;
      RECT 58.835 2.77 59.065 3.3 ;
      RECT 57.835 2.01 58.085 3.3 ;
      RECT 58.835 2.7 58.895 3.6 ;
      RECT 58.835 2.7 59.065 2.76 ;
      RECT 57.295 2.01 58.085 2.28 ;
      RECT 58.255 5.82 58.935 6.07 ;
      RECT 58.665 5.46 58.935 6.07 ;
      RECT 58.415 6.24 58.745 6.79 ;
      RECT 57.355 6.24 58.745 6.43 ;
      RECT 57.355 5.4 57.525 6.43 ;
      RECT 57.235 5.82 57.525 6.15 ;
      RECT 57.355 5.4 58.295 5.57 ;
      RECT 57.995 4.85 58.295 5.57 ;
      RECT 58.255 2.43 58.665 2.95 ;
      RECT 58.255 2.01 58.455 2.95 ;
      RECT 56.865 2.19 57.035 4.17 ;
      RECT 56.865 2.7 57.665 2.95 ;
      RECT 56.865 2.19 57.115 2.95 ;
      RECT 56.785 2.19 57.115 2.61 ;
      RECT 56.815 6.6 57.375 6.89 ;
      RECT 56.815 4.68 57.065 6.89 ;
      RECT 56.815 4.68 57.275 5.23 ;
      RECT 53.645 5.015 53.815 8.305 ;
      RECT 53.645 7.315 54.05 7.645 ;
      RECT 53.645 6.475 54.05 6.805 ;
      RECT 52.015 5.02 52.185 6.49 ;
      RECT 52.015 6.315 52.19 6.485 ;
      RECT 51.645 1.74 51.815 2.93 ;
      RECT 51.645 1.74 52.115 1.91 ;
      RECT 51.645 6.97 52.115 7.14 ;
      RECT 51.645 5.95 51.815 7.14 ;
      RECT 50.655 1.74 50.825 2.93 ;
      RECT 50.655 1.74 51.125 1.91 ;
      RECT 50.655 6.97 51.125 7.14 ;
      RECT 50.655 5.95 50.825 7.14 ;
      RECT 48.805 2.635 48.975 3.865 ;
      RECT 48.86 0.855 49.03 2.805 ;
      RECT 48.805 0.575 48.975 1.025 ;
      RECT 48.805 7.855 48.975 8.305 ;
      RECT 48.86 6.075 49.03 8.025 ;
      RECT 48.805 5.015 48.975 6.245 ;
      RECT 48.285 0.575 48.455 3.865 ;
      RECT 48.285 2.075 48.69 2.405 ;
      RECT 48.285 1.235 48.69 1.565 ;
      RECT 48.285 5.015 48.455 8.305 ;
      RECT 48.285 7.315 48.69 7.645 ;
      RECT 48.285 6.475 48.69 6.805 ;
      RECT 43.54 6.64 44.85 6.89 ;
      RECT 43.54 6.32 43.72 6.89 ;
      RECT 42.99 6.32 43.72 6.49 ;
      RECT 42.99 5.48 43.16 6.49 ;
      RECT 43.83 5.52 45.57 5.7 ;
      RECT 45.24 4.68 45.57 5.7 ;
      RECT 42.99 5.48 44.05 5.65 ;
      RECT 45.24 4.85 46.06 5.02 ;
      RECT 44.4 4.68 44.73 4.89 ;
      RECT 44.4 4.68 45.57 4.85 ;
      RECT 45.3 3.2 45.63 4.16 ;
      RECT 45.3 3.2 45.98 3.37 ;
      RECT 45.81 1.96 45.98 3.37 ;
      RECT 45.72 1.96 46.05 2.6 ;
      RECT 44.85 3.47 45.12 4.17 ;
      RECT 44.95 1.96 45.12 4.17 ;
      RECT 45.29 2.78 45.64 3.03 ;
      RECT 44.95 2.81 45.64 2.98 ;
      RECT 44.86 1.96 45.12 2.44 ;
      RECT 44.19 5.11 45.07 5.35 ;
      RECT 44.84 5.02 45.07 5.35 ;
      RECT 43.54 5.11 45.07 5.31 ;
      RECT 44.46 5.06 45.07 5.35 ;
      RECT 43.54 4.98 43.71 5.31 ;
      RECT 44.43 5.87 44.68 6.47 ;
      RECT 44.43 5.87 44.9 6.07 ;
      RECT 43.92 3.09 44.68 3.59 ;
      RECT 42.99 2.9 43.25 3.52 ;
      RECT 43.91 3.03 43.92 3.34 ;
      RECT 43.89 3.02 43.91 3.31 ;
      RECT 44.55 2.7 44.78 3.3 ;
      RECT 43.87 2.97 43.89 3.28 ;
      RECT 43.85 3.09 44.78 3.27 ;
      RECT 43.82 3.09 44.78 3.26 ;
      RECT 43.75 3.09 44.78 3.25 ;
      RECT 43.73 3.09 44.78 3.22 ;
      RECT 43.71 2 43.88 3.19 ;
      RECT 43.68 3.09 44.78 3.16 ;
      RECT 43.65 3.09 44.78 3.13 ;
      RECT 43.62 3.08 43.98 3.1 ;
      RECT 43.62 3.07 43.97 3.1 ;
      RECT 42.99 2.9 43.88 3.07 ;
      RECT 42.99 3.06 43.95 3.07 ;
      RECT 42.99 3.05 43.94 3.07 ;
      RECT 42.99 2.99 43.9 3.07 ;
      RECT 42.99 2 43.88 2.17 ;
      RECT 44.05 2.5 44.38 2.92 ;
      RECT 44.05 2.01 44.27 2.92 ;
      RECT 43.97 5.87 44.18 6.47 ;
      RECT 43.83 5.87 44.18 6.07 ;
      RECT 42.55 3.47 42.82 4.17 ;
      RECT 42.77 1.96 42.82 4.17 ;
      RECT 42.65 2.77 42.82 4.17 ;
      RECT 42.65 1.96 42.82 2.76 ;
      RECT 42.56 1.96 42.82 2.44 ;
      RECT 40.69 3.13 40.94 3.67 ;
      RECT 41.66 3.13 42.38 3.6 ;
      RECT 40.69 3.13 42.48 3.3 ;
      RECT 42.25 2.77 42.48 3.3 ;
      RECT 41.25 2.01 41.5 3.3 ;
      RECT 42.25 2.7 42.31 3.6 ;
      RECT 42.25 2.7 42.48 2.76 ;
      RECT 40.71 2.01 41.5 2.28 ;
      RECT 41.67 5.82 42.35 6.07 ;
      RECT 42.08 5.46 42.35 6.07 ;
      RECT 41.83 6.24 42.16 6.79 ;
      RECT 40.77 6.24 42.16 6.43 ;
      RECT 40.77 5.4 40.94 6.43 ;
      RECT 40.65 5.82 40.94 6.15 ;
      RECT 40.77 5.4 41.71 5.57 ;
      RECT 41.41 4.85 41.71 5.57 ;
      RECT 41.67 2.43 42.08 2.95 ;
      RECT 41.67 2.01 41.87 2.95 ;
      RECT 40.28 2.19 40.45 4.17 ;
      RECT 40.28 2.7 41.08 2.95 ;
      RECT 40.28 2.19 40.53 2.95 ;
      RECT 40.2 2.19 40.53 2.61 ;
      RECT 40.23 6.6 40.79 6.89 ;
      RECT 40.23 4.68 40.48 6.89 ;
      RECT 40.23 4.68 40.69 5.23 ;
      RECT 37.06 5.015 37.23 8.305 ;
      RECT 37.06 7.315 37.465 7.645 ;
      RECT 37.06 6.475 37.465 6.805 ;
      RECT 35.43 5.02 35.6 6.49 ;
      RECT 35.43 6.315 35.605 6.485 ;
      RECT 35.06 1.74 35.23 2.93 ;
      RECT 35.06 1.74 35.53 1.91 ;
      RECT 35.06 6.97 35.53 7.14 ;
      RECT 35.06 5.95 35.23 7.14 ;
      RECT 34.07 1.74 34.24 2.93 ;
      RECT 34.07 1.74 34.54 1.91 ;
      RECT 34.07 6.97 34.54 7.14 ;
      RECT 34.07 5.95 34.24 7.14 ;
      RECT 32.22 2.635 32.39 3.865 ;
      RECT 32.275 0.855 32.445 2.805 ;
      RECT 32.22 0.575 32.39 1.025 ;
      RECT 32.22 7.855 32.39 8.305 ;
      RECT 32.275 6.075 32.445 8.025 ;
      RECT 32.22 5.015 32.39 6.245 ;
      RECT 31.7 0.575 31.87 3.865 ;
      RECT 31.7 2.075 32.105 2.405 ;
      RECT 31.7 1.235 32.105 1.565 ;
      RECT 31.7 5.015 31.87 8.305 ;
      RECT 31.7 7.315 32.105 7.645 ;
      RECT 31.7 6.475 32.105 6.805 ;
      RECT 26.955 6.64 28.265 6.89 ;
      RECT 26.955 6.32 27.135 6.89 ;
      RECT 26.405 6.32 27.135 6.49 ;
      RECT 26.405 5.48 26.575 6.49 ;
      RECT 27.245 5.52 28.985 5.7 ;
      RECT 28.655 4.68 28.985 5.7 ;
      RECT 26.405 5.48 27.465 5.65 ;
      RECT 28.655 4.85 29.475 5.02 ;
      RECT 27.815 4.68 28.145 4.89 ;
      RECT 27.815 4.68 28.985 4.85 ;
      RECT 28.715 3.2 29.045 4.16 ;
      RECT 28.715 3.2 29.395 3.37 ;
      RECT 29.225 1.96 29.395 3.37 ;
      RECT 29.135 1.96 29.465 2.6 ;
      RECT 28.265 3.47 28.535 4.17 ;
      RECT 28.365 1.96 28.535 4.17 ;
      RECT 28.705 2.78 29.055 3.03 ;
      RECT 28.365 2.81 29.055 2.98 ;
      RECT 28.275 1.96 28.535 2.44 ;
      RECT 27.605 5.11 28.485 5.35 ;
      RECT 28.255 5.02 28.485 5.35 ;
      RECT 26.955 5.11 28.485 5.31 ;
      RECT 27.875 5.06 28.485 5.35 ;
      RECT 26.955 4.98 27.125 5.31 ;
      RECT 27.845 5.87 28.095 6.47 ;
      RECT 27.845 5.87 28.315 6.07 ;
      RECT 27.335 3.09 28.095 3.59 ;
      RECT 26.405 2.9 26.665 3.52 ;
      RECT 27.325 3.03 27.335 3.34 ;
      RECT 27.305 3.02 27.325 3.31 ;
      RECT 27.965 2.7 28.195 3.3 ;
      RECT 27.285 2.97 27.305 3.28 ;
      RECT 27.265 3.09 28.195 3.27 ;
      RECT 27.235 3.09 28.195 3.26 ;
      RECT 27.165 3.09 28.195 3.25 ;
      RECT 27.145 3.09 28.195 3.22 ;
      RECT 27.125 2 27.295 3.19 ;
      RECT 27.095 3.09 28.195 3.16 ;
      RECT 27.065 3.09 28.195 3.13 ;
      RECT 27.035 3.08 27.395 3.1 ;
      RECT 27.035 3.07 27.385 3.1 ;
      RECT 26.405 2.9 27.295 3.07 ;
      RECT 26.405 3.06 27.365 3.07 ;
      RECT 26.405 3.05 27.355 3.07 ;
      RECT 26.405 2.99 27.315 3.07 ;
      RECT 26.405 2 27.295 2.17 ;
      RECT 27.465 2.5 27.795 2.92 ;
      RECT 27.465 2.01 27.685 2.92 ;
      RECT 27.385 5.87 27.595 6.47 ;
      RECT 27.245 5.87 27.595 6.07 ;
      RECT 25.965 3.47 26.235 4.17 ;
      RECT 26.185 1.96 26.235 4.17 ;
      RECT 26.065 2.77 26.235 4.17 ;
      RECT 26.065 1.96 26.235 2.76 ;
      RECT 25.975 1.96 26.235 2.44 ;
      RECT 24.105 3.13 24.355 3.67 ;
      RECT 25.075 3.13 25.795 3.6 ;
      RECT 24.105 3.13 25.895 3.3 ;
      RECT 25.665 2.77 25.895 3.3 ;
      RECT 24.665 2.01 24.915 3.3 ;
      RECT 25.665 2.7 25.725 3.6 ;
      RECT 25.665 2.7 25.895 2.76 ;
      RECT 24.125 2.01 24.915 2.28 ;
      RECT 25.085 5.82 25.765 6.07 ;
      RECT 25.495 5.46 25.765 6.07 ;
      RECT 25.245 6.24 25.575 6.79 ;
      RECT 24.185 6.24 25.575 6.43 ;
      RECT 24.185 5.4 24.355 6.43 ;
      RECT 24.065 5.82 24.355 6.15 ;
      RECT 24.185 5.4 25.125 5.57 ;
      RECT 24.825 4.85 25.125 5.57 ;
      RECT 25.085 2.43 25.495 2.95 ;
      RECT 25.085 2.01 25.285 2.95 ;
      RECT 23.695 2.19 23.865 4.17 ;
      RECT 23.695 2.7 24.495 2.95 ;
      RECT 23.695 2.19 23.945 2.95 ;
      RECT 23.615 2.19 23.945 2.61 ;
      RECT 23.645 6.6 24.205 6.89 ;
      RECT 23.645 4.68 23.895 6.89 ;
      RECT 23.645 4.68 24.105 5.23 ;
      RECT 20.475 5.015 20.645 8.305 ;
      RECT 20.475 7.315 20.88 7.645 ;
      RECT 20.475 6.475 20.88 6.805 ;
      RECT 18.845 5.02 19.015 6.49 ;
      RECT 18.845 6.315 19.02 6.485 ;
      RECT 18.475 1.74 18.645 2.93 ;
      RECT 18.475 1.74 18.945 1.91 ;
      RECT 18.475 6.97 18.945 7.14 ;
      RECT 18.475 5.95 18.645 7.14 ;
      RECT 17.485 1.74 17.655 2.93 ;
      RECT 17.485 1.74 17.955 1.91 ;
      RECT 17.485 6.97 17.955 7.14 ;
      RECT 17.485 5.95 17.655 7.14 ;
      RECT 15.635 2.635 15.805 3.865 ;
      RECT 15.69 0.855 15.86 2.805 ;
      RECT 15.635 0.575 15.805 1.025 ;
      RECT 15.635 7.855 15.805 8.305 ;
      RECT 15.69 6.075 15.86 8.025 ;
      RECT 15.635 5.015 15.805 6.245 ;
      RECT 15.115 0.575 15.285 3.865 ;
      RECT 15.115 2.075 15.52 2.405 ;
      RECT 15.115 1.235 15.52 1.565 ;
      RECT 15.115 5.015 15.285 8.305 ;
      RECT 15.115 7.315 15.52 7.645 ;
      RECT 15.115 6.475 15.52 6.805 ;
      RECT 10.37 6.64 11.68 6.89 ;
      RECT 10.37 6.32 10.55 6.89 ;
      RECT 9.82 6.32 10.55 6.49 ;
      RECT 9.82 5.48 9.99 6.49 ;
      RECT 10.66 5.52 12.4 5.7 ;
      RECT 12.07 4.68 12.4 5.7 ;
      RECT 9.82 5.48 10.88 5.65 ;
      RECT 12.07 4.85 12.89 5.02 ;
      RECT 11.23 4.68 11.56 4.89 ;
      RECT 11.23 4.68 12.4 4.85 ;
      RECT 12.13 3.2 12.46 4.16 ;
      RECT 12.13 3.2 12.81 3.37 ;
      RECT 12.64 1.96 12.81 3.37 ;
      RECT 12.55 1.96 12.88 2.6 ;
      RECT 11.68 3.47 11.95 4.17 ;
      RECT 11.78 1.96 11.95 4.17 ;
      RECT 12.12 2.78 12.47 3.03 ;
      RECT 11.78 2.81 12.47 2.98 ;
      RECT 11.69 1.96 11.95 2.44 ;
      RECT 11.02 5.11 11.9 5.35 ;
      RECT 11.67 5.02 11.9 5.35 ;
      RECT 10.37 5.11 11.9 5.31 ;
      RECT 11.29 5.06 11.9 5.35 ;
      RECT 10.37 4.98 10.54 5.31 ;
      RECT 11.26 5.87 11.51 6.47 ;
      RECT 11.26 5.87 11.73 6.07 ;
      RECT 10.75 3.09 11.51 3.59 ;
      RECT 9.82 2.9 10.08 3.52 ;
      RECT 10.74 3.03 10.75 3.34 ;
      RECT 10.72 3.02 10.74 3.31 ;
      RECT 11.38 2.7 11.61 3.3 ;
      RECT 10.7 2.97 10.72 3.28 ;
      RECT 10.68 3.09 11.61 3.27 ;
      RECT 10.65 3.09 11.61 3.26 ;
      RECT 10.58 3.09 11.61 3.25 ;
      RECT 10.56 3.09 11.61 3.22 ;
      RECT 10.54 2 10.71 3.19 ;
      RECT 10.51 3.09 11.61 3.16 ;
      RECT 10.48 3.09 11.61 3.13 ;
      RECT 10.45 3.08 10.81 3.1 ;
      RECT 10.45 3.07 10.8 3.1 ;
      RECT 9.82 2.9 10.71 3.07 ;
      RECT 9.82 3.06 10.78 3.07 ;
      RECT 9.82 3.05 10.77 3.07 ;
      RECT 9.82 2.99 10.73 3.07 ;
      RECT 9.82 2 10.71 2.17 ;
      RECT 10.88 2.5 11.21 2.92 ;
      RECT 10.88 2.01 11.1 2.92 ;
      RECT 10.8 5.87 11.01 6.47 ;
      RECT 10.66 5.87 11.01 6.07 ;
      RECT 9.38 3.47 9.65 4.17 ;
      RECT 9.6 1.96 9.65 4.17 ;
      RECT 9.48 2.77 9.65 4.17 ;
      RECT 9.48 1.96 9.65 2.76 ;
      RECT 9.39 1.96 9.65 2.44 ;
      RECT 7.52 3.13 7.77 3.67 ;
      RECT 8.49 3.13 9.21 3.6 ;
      RECT 7.52 3.13 9.31 3.3 ;
      RECT 9.08 2.77 9.31 3.3 ;
      RECT 8.08 2.01 8.33 3.3 ;
      RECT 9.08 2.7 9.14 3.6 ;
      RECT 9.08 2.7 9.31 2.76 ;
      RECT 7.54 2.01 8.33 2.28 ;
      RECT 8.5 5.82 9.18 6.07 ;
      RECT 8.91 5.46 9.18 6.07 ;
      RECT 8.66 6.24 8.99 6.79 ;
      RECT 7.6 6.24 8.99 6.43 ;
      RECT 7.6 5.4 7.77 6.43 ;
      RECT 7.48 5.82 7.77 6.15 ;
      RECT 7.6 5.4 8.54 5.57 ;
      RECT 8.24 4.85 8.54 5.57 ;
      RECT 8.5 2.43 8.91 2.95 ;
      RECT 8.5 2.01 8.7 2.95 ;
      RECT 7.11 2.19 7.28 4.17 ;
      RECT 7.11 2.7 7.91 2.95 ;
      RECT 7.11 2.19 7.36 2.95 ;
      RECT 7.03 2.19 7.36 2.61 ;
      RECT 7.06 6.6 7.62 6.89 ;
      RECT 7.06 4.68 7.31 6.89 ;
      RECT 7.06 4.68 7.52 5.23 ;
      RECT 3.89 5.015 4.06 8.305 ;
      RECT 3.89 7.315 4.295 7.645 ;
      RECT 3.89 6.475 4.295 6.805 ;
      RECT 1.18 7.855 1.35 8.305 ;
      RECT 1.235 6.075 1.405 8.025 ;
      RECT 1.18 5.015 1.35 6.245 ;
      RECT 0.66 5.015 0.83 8.305 ;
      RECT 0.66 7.315 1.065 7.645 ;
      RECT 0.66 6.475 1.065 6.805 ;
      RECT 85.18 7.8 85.35 8.31 ;
      RECT 84.19 0.57 84.36 1.08 ;
      RECT 84.19 2.39 84.36 3.86 ;
      RECT 84.19 5.02 84.36 6.49 ;
      RECT 84.19 7.8 84.36 8.31 ;
      RECT 82.83 0.575 83 3.865 ;
      RECT 82.83 5.015 83 8.305 ;
      RECT 82.4 0.575 82.57 1.085 ;
      RECT 82.4 1.655 82.57 3.865 ;
      RECT 82.4 5.015 82.57 7.225 ;
      RECT 82.4 7.795 82.57 8.305 ;
      RECT 79.315 2.78 79.665 3.03 ;
      RECT 78.255 5.87 78.705 6.38 ;
      RECT 76.935 3.83 77.415 4.17 ;
      RECT 76.155 2.34 76.705 2.73 ;
      RECT 74.645 3.83 75.115 4.17 ;
      RECT 72.935 2.78 73.275 3.66 ;
      RECT 71.605 5.015 71.775 8.305 ;
      RECT 71.175 5.015 71.345 7.225 ;
      RECT 71.175 7.795 71.345 8.305 ;
      RECT 68.6 7.8 68.77 8.31 ;
      RECT 67.61 0.57 67.78 1.08 ;
      RECT 67.61 2.39 67.78 3.86 ;
      RECT 67.61 5.02 67.78 6.49 ;
      RECT 67.61 7.8 67.78 8.31 ;
      RECT 66.25 0.575 66.42 3.865 ;
      RECT 66.25 5.015 66.42 8.305 ;
      RECT 65.82 0.575 65.99 1.085 ;
      RECT 65.82 1.655 65.99 3.865 ;
      RECT 65.82 5.015 65.99 7.225 ;
      RECT 65.82 7.795 65.99 8.305 ;
      RECT 62.735 2.78 63.085 3.03 ;
      RECT 61.675 5.87 62.125 6.38 ;
      RECT 60.355 3.83 60.835 4.17 ;
      RECT 59.575 2.34 60.125 2.73 ;
      RECT 58.065 3.83 58.535 4.17 ;
      RECT 56.355 2.78 56.695 3.66 ;
      RECT 55.025 5.015 55.195 8.305 ;
      RECT 54.595 5.015 54.765 7.225 ;
      RECT 54.595 7.795 54.765 8.305 ;
      RECT 52.015 7.8 52.185 8.31 ;
      RECT 51.025 0.57 51.195 1.08 ;
      RECT 51.025 2.39 51.195 3.86 ;
      RECT 51.025 5.02 51.195 6.49 ;
      RECT 51.025 7.8 51.195 8.31 ;
      RECT 49.665 0.575 49.835 3.865 ;
      RECT 49.665 5.015 49.835 8.305 ;
      RECT 49.235 0.575 49.405 1.085 ;
      RECT 49.235 1.655 49.405 3.865 ;
      RECT 49.235 5.015 49.405 7.225 ;
      RECT 49.235 7.795 49.405 8.305 ;
      RECT 46.15 2.78 46.5 3.03 ;
      RECT 45.09 5.87 45.54 6.38 ;
      RECT 43.77 3.83 44.25 4.17 ;
      RECT 42.99 2.34 43.54 2.73 ;
      RECT 41.48 3.83 41.95 4.17 ;
      RECT 39.77 2.78 40.11 3.66 ;
      RECT 38.44 5.015 38.61 8.305 ;
      RECT 38.01 5.015 38.18 7.225 ;
      RECT 38.01 7.795 38.18 8.305 ;
      RECT 35.43 7.8 35.6 8.31 ;
      RECT 34.44 0.57 34.61 1.08 ;
      RECT 34.44 2.39 34.61 3.86 ;
      RECT 34.44 5.02 34.61 6.49 ;
      RECT 34.44 7.8 34.61 8.31 ;
      RECT 33.08 0.575 33.25 3.865 ;
      RECT 33.08 5.015 33.25 8.305 ;
      RECT 32.65 0.575 32.82 1.085 ;
      RECT 32.65 1.655 32.82 3.865 ;
      RECT 32.65 5.015 32.82 7.225 ;
      RECT 32.65 7.795 32.82 8.305 ;
      RECT 29.565 2.78 29.915 3.03 ;
      RECT 28.505 5.87 28.955 6.38 ;
      RECT 27.185 3.83 27.665 4.17 ;
      RECT 26.405 2.34 26.955 2.73 ;
      RECT 24.895 3.83 25.365 4.17 ;
      RECT 23.185 2.78 23.525 3.66 ;
      RECT 21.855 5.015 22.025 8.305 ;
      RECT 21.425 5.015 21.595 7.225 ;
      RECT 21.425 7.795 21.595 8.305 ;
      RECT 18.845 7.8 19.015 8.31 ;
      RECT 17.855 0.57 18.025 1.08 ;
      RECT 17.855 2.39 18.025 3.86 ;
      RECT 17.855 5.02 18.025 6.49 ;
      RECT 17.855 7.8 18.025 8.31 ;
      RECT 16.495 0.575 16.665 3.865 ;
      RECT 16.495 5.015 16.665 8.305 ;
      RECT 16.065 0.575 16.235 1.085 ;
      RECT 16.065 1.655 16.235 3.865 ;
      RECT 16.065 5.015 16.235 7.225 ;
      RECT 16.065 7.795 16.235 8.305 ;
      RECT 12.98 2.78 13.33 3.03 ;
      RECT 11.92 5.87 12.37 6.38 ;
      RECT 10.6 3.83 11.08 4.17 ;
      RECT 9.82 2.34 10.37 2.73 ;
      RECT 8.31 3.83 8.78 4.17 ;
      RECT 6.6 2.78 6.94 3.66 ;
      RECT 5.27 5.015 5.44 8.305 ;
      RECT 4.84 5.015 5.01 7.225 ;
      RECT 4.84 7.795 5.01 8.305 ;
      RECT 1.61 5.015 1.78 7.225 ;
      RECT 1.61 7.795 1.78 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r2 ;
  SIZE 85.88 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 19.005 2.395 19.175 2.565 ;
        RECT 19 2.39 19.17 2.56 ;
        RECT 19 0.91 19.17 1.08 ;
      LAYER li1 ;
        RECT 19 2.395 19.175 2.565 ;
        RECT 19 2.39 19.17 3.86 ;
        RECT 19 0.57 19.17 1.08 ;
      LAYER met1 ;
        RECT 18.94 2.36 19.23 2.59 ;
        RECT 18.94 0.88 19.23 1.11 ;
        RECT 19 0.88 19.17 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 35.59 2.395 35.76 2.565 ;
        RECT 35.585 2.39 35.755 2.56 ;
        RECT 35.585 0.91 35.755 1.08 ;
      LAYER li1 ;
        RECT 35.585 2.395 35.76 2.565 ;
        RECT 35.585 2.39 35.755 3.86 ;
        RECT 35.585 0.57 35.755 1.08 ;
      LAYER met1 ;
        RECT 35.525 2.36 35.815 2.59 ;
        RECT 35.525 0.88 35.815 1.11 ;
        RECT 35.585 0.88 35.755 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 52.175 2.395 52.345 2.565 ;
        RECT 52.17 2.39 52.34 2.56 ;
        RECT 52.17 0.91 52.34 1.08 ;
      LAYER li1 ;
        RECT 52.17 2.395 52.345 2.565 ;
        RECT 52.17 2.39 52.34 3.86 ;
        RECT 52.17 0.57 52.34 1.08 ;
      LAYER met1 ;
        RECT 52.11 2.36 52.4 2.59 ;
        RECT 52.11 0.88 52.4 1.11 ;
        RECT 52.17 0.88 52.34 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 68.76 2.395 68.93 2.565 ;
        RECT 68.755 2.39 68.925 2.56 ;
        RECT 68.755 0.91 68.925 1.08 ;
      LAYER li1 ;
        RECT 68.755 2.395 68.93 2.565 ;
        RECT 68.755 2.39 68.925 3.86 ;
        RECT 68.755 0.57 68.925 1.08 ;
      LAYER met1 ;
        RECT 68.695 2.36 68.985 2.59 ;
        RECT 68.695 0.88 68.985 1.11 ;
        RECT 68.755 0.88 68.925 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 85.34 2.395 85.51 2.565 ;
        RECT 85.335 2.39 85.505 2.56 ;
        RECT 85.335 0.91 85.505 1.08 ;
      LAYER li1 ;
        RECT 85.335 2.395 85.51 2.565 ;
        RECT 85.335 2.39 85.505 3.86 ;
        RECT 85.335 0.57 85.505 1.08 ;
      LAYER met1 ;
        RECT 85.275 2.36 85.565 2.59 ;
        RECT 85.275 0.88 85.565 1.11 ;
        RECT 85.335 0.88 85.505 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 14.85 1.66 15.02 2.935 ;
        RECT 14.85 5.945 15.02 7.22 ;
        RECT 3.625 5.945 3.795 7.22 ;
      LAYER met2 ;
        RECT 14.775 5.865 15.1 6.19 ;
        RECT 14.77 3.635 15.095 3.96 ;
        RECT 5.93 7.885 15.015 8.055 ;
        RECT 14.84 3.635 15.015 8.055 ;
        RECT 5.875 5.86 6.155 6.2 ;
        RECT 5.93 5.86 6.1 8.055 ;
      LAYER met1 ;
        RECT 14.79 2.765 15.25 2.935 ;
        RECT 14.77 3.635 15.095 3.96 ;
        RECT 14.79 2.735 15.08 2.965 ;
        RECT 14.845 2.735 15.025 3.96 ;
        RECT 14.775 5.945 15.25 6.115 ;
        RECT 14.775 5.865 15.1 6.19 ;
        RECT 5.845 5.89 6.185 6.17 ;
        RECT 3.565 5.945 6.185 6.115 ;
        RECT 3.565 5.915 3.855 6.145 ;
      LAYER mcon ;
        RECT 3.625 5.945 3.795 6.115 ;
        RECT 14.85 5.945 15.02 6.115 ;
        RECT 14.85 2.765 15.02 2.935 ;
      LAYER via1 ;
        RECT 5.94 5.955 6.09 6.105 ;
        RECT 14.86 3.72 15.01 3.87 ;
        RECT 14.865 5.95 15.015 6.1 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 31.435 1.66 31.605 2.935 ;
        RECT 31.435 5.945 31.605 7.22 ;
        RECT 20.21 5.945 20.38 7.22 ;
      LAYER met2 ;
        RECT 31.36 5.865 31.685 6.19 ;
        RECT 31.355 3.635 31.68 3.96 ;
        RECT 22.515 7.885 31.6 8.055 ;
        RECT 31.425 3.635 31.6 8.055 ;
        RECT 22.46 5.86 22.74 6.2 ;
        RECT 22.515 5.86 22.685 8.055 ;
      LAYER met1 ;
        RECT 31.375 2.765 31.835 2.935 ;
        RECT 31.355 3.635 31.68 3.96 ;
        RECT 31.375 2.735 31.665 2.965 ;
        RECT 31.43 2.735 31.61 3.96 ;
        RECT 31.36 5.945 31.835 6.115 ;
        RECT 31.36 5.865 31.685 6.19 ;
        RECT 22.43 5.89 22.77 6.17 ;
        RECT 20.15 5.945 22.77 6.115 ;
        RECT 20.15 5.915 20.44 6.145 ;
      LAYER mcon ;
        RECT 20.21 5.945 20.38 6.115 ;
        RECT 31.435 5.945 31.605 6.115 ;
        RECT 31.435 2.765 31.605 2.935 ;
      LAYER via1 ;
        RECT 22.525 5.955 22.675 6.105 ;
        RECT 31.445 3.72 31.595 3.87 ;
        RECT 31.45 5.95 31.6 6.1 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 48.02 1.66 48.19 2.935 ;
        RECT 48.02 5.945 48.19 7.22 ;
        RECT 36.795 5.945 36.965 7.22 ;
      LAYER met2 ;
        RECT 47.945 5.865 48.27 6.19 ;
        RECT 47.94 3.635 48.265 3.96 ;
        RECT 39.1 7.885 48.185 8.055 ;
        RECT 48.01 3.635 48.185 8.055 ;
        RECT 39.045 5.86 39.325 6.2 ;
        RECT 39.1 5.86 39.27 8.055 ;
      LAYER met1 ;
        RECT 47.96 2.765 48.42 2.935 ;
        RECT 47.94 3.635 48.265 3.96 ;
        RECT 47.96 2.735 48.25 2.965 ;
        RECT 48.015 2.735 48.195 3.96 ;
        RECT 47.945 5.945 48.42 6.115 ;
        RECT 47.945 5.865 48.27 6.19 ;
        RECT 39.015 5.89 39.355 6.17 ;
        RECT 36.735 5.945 39.355 6.115 ;
        RECT 36.735 5.915 37.025 6.145 ;
      LAYER mcon ;
        RECT 36.795 5.945 36.965 6.115 ;
        RECT 48.02 5.945 48.19 6.115 ;
        RECT 48.02 2.765 48.19 2.935 ;
      LAYER via1 ;
        RECT 39.11 5.955 39.26 6.105 ;
        RECT 48.03 3.72 48.18 3.87 ;
        RECT 48.035 5.95 48.185 6.1 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 64.605 1.66 64.775 2.935 ;
        RECT 64.605 5.945 64.775 7.22 ;
        RECT 53.38 5.945 53.55 7.22 ;
      LAYER met2 ;
        RECT 64.53 5.865 64.855 6.19 ;
        RECT 64.525 3.635 64.85 3.96 ;
        RECT 55.685 7.885 64.77 8.055 ;
        RECT 64.595 3.635 64.77 8.055 ;
        RECT 55.63 5.86 55.91 6.2 ;
        RECT 55.685 5.86 55.855 8.055 ;
      LAYER met1 ;
        RECT 64.545 2.765 65.005 2.935 ;
        RECT 64.525 3.635 64.85 3.96 ;
        RECT 64.545 2.735 64.835 2.965 ;
        RECT 64.6 2.735 64.78 3.96 ;
        RECT 64.53 5.945 65.005 6.115 ;
        RECT 64.53 5.865 64.855 6.19 ;
        RECT 55.6 5.89 55.94 6.17 ;
        RECT 53.32 5.945 55.94 6.115 ;
        RECT 53.32 5.915 53.61 6.145 ;
      LAYER mcon ;
        RECT 53.38 5.945 53.55 6.115 ;
        RECT 64.605 5.945 64.775 6.115 ;
        RECT 64.605 2.765 64.775 2.935 ;
      LAYER via1 ;
        RECT 55.695 5.955 55.845 6.105 ;
        RECT 64.615 3.72 64.765 3.87 ;
        RECT 64.62 5.95 64.77 6.1 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 81.185 1.66 81.355 2.935 ;
        RECT 81.185 5.945 81.355 7.22 ;
        RECT 69.96 5.945 70.13 7.22 ;
      LAYER met2 ;
        RECT 81.11 5.865 81.435 6.19 ;
        RECT 81.105 3.635 81.43 3.96 ;
        RECT 72.265 7.885 81.35 8.055 ;
        RECT 81.175 3.635 81.35 8.055 ;
        RECT 72.21 5.86 72.49 6.2 ;
        RECT 72.265 5.86 72.435 8.055 ;
      LAYER met1 ;
        RECT 81.125 2.765 81.585 2.935 ;
        RECT 81.105 3.635 81.43 3.96 ;
        RECT 81.125 2.735 81.415 2.965 ;
        RECT 81.18 2.735 81.36 3.96 ;
        RECT 81.11 5.945 81.585 6.115 ;
        RECT 81.11 5.865 81.435 6.19 ;
        RECT 72.18 5.89 72.52 6.17 ;
        RECT 69.9 5.945 72.52 6.115 ;
        RECT 69.9 5.915 70.19 6.145 ;
      LAYER mcon ;
        RECT 69.96 5.945 70.13 6.115 ;
        RECT 81.185 5.945 81.355 6.115 ;
        RECT 81.185 2.765 81.355 2.935 ;
      LAYER via1 ;
        RECT 72.275 5.955 72.425 6.105 ;
        RECT 81.195 3.72 81.345 3.87 ;
        RECT 81.2 5.95 81.35 6.1 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.395 5.945 0.565 7.22 ;
      LAYER met1 ;
        RECT 0.335 5.945 0.795 6.115 ;
        RECT 0.335 5.915 0.625 6.145 ;
      LAYER mcon ;
        RECT 0.395 5.945 0.565 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.34 4.23 2.145 4.61 ;
      LAYER li1 ;
        RECT 79.94 4.135 85.88 4.745 ;
        RECT 83.745 4.13 85.725 4.75 ;
        RECT 84.905 3.4 85.075 5.48 ;
        RECT 83.915 3.4 84.085 5.48 ;
        RECT 81.175 3.405 81.345 5.475 ;
        RECT 79.81 4.135 85.88 4.67 ;
        RECT 79.48 3.2 79.81 4.51 ;
        RECT 73.01 4.34 85.88 4.51 ;
        RECT 77.74 3.8 78 4.51 ;
        RECT 77.18 4.34 77.55 4.89 ;
        RECT 76.74 3.42 77.07 3.66 ;
        RECT 76.74 3.42 76.93 3.79 ;
        RECT 76.31 3.69 76.92 4.51 ;
        RECT 76.36 3.69 76.63 5.29 ;
        RECT 75.44 3.8 75.66 4.51 ;
        RECT 75.2 4.34 75.48 5.18 ;
        RECT 74.43 3.47 74.76 3.66 ;
        RECT 74.01 3.84 74.63 4.51 ;
        RECT 74.43 3.47 74.63 4.51 ;
        RECT 74.2 3.84 74.53 5.23 ;
        RECT 73.09 3.83 73.35 4.51 ;
        RECT 63.23 4.345 73.085 4.515 ;
        RECT 69.295 4.13 72.87 4.74 ;
        RECT 69.775 4.13 72.525 4.745 ;
        RECT 69.95 4.13 70.12 5.475 ;
        RECT 63.36 4.135 69.3 4.745 ;
        RECT 67.165 4.13 69.145 4.75 ;
        RECT 68.325 3.4 68.495 5.48 ;
        RECT 67.335 3.4 67.505 5.48 ;
        RECT 64.595 3.405 64.765 5.475 ;
        RECT 63.23 4.135 72.87 4.67 ;
        RECT 62.9 3.2 63.23 4.51 ;
        RECT 1.805 4.345 85.88 4.51 ;
        RECT 56.43 4.34 72.87 4.51 ;
        RECT 61.16 3.8 61.42 4.51 ;
        RECT 60.6 4.34 60.97 4.89 ;
        RECT 60.16 3.42 60.49 3.66 ;
        RECT 60.16 3.42 60.35 3.79 ;
        RECT 59.73 3.69 60.34 4.51 ;
        RECT 59.78 3.69 60.05 5.29 ;
        RECT 58.86 3.8 59.08 4.51 ;
        RECT 58.62 4.34 58.9 5.18 ;
        RECT 57.85 3.47 58.18 3.66 ;
        RECT 57.43 3.84 58.05 4.51 ;
        RECT 57.85 3.47 58.05 4.51 ;
        RECT 57.62 3.84 57.95 5.23 ;
        RECT 56.51 3.83 56.77 4.51 ;
        RECT 46.645 4.345 56.505 4.515 ;
        RECT 52.715 4.13 56.29 4.74 ;
        RECT 53.195 4.13 55.945 4.745 ;
        RECT 53.37 4.13 53.54 5.475 ;
        RECT 46.775 4.135 52.715 4.745 ;
        RECT 50.58 4.13 52.56 4.75 ;
        RECT 51.74 3.4 51.91 5.48 ;
        RECT 50.75 3.4 50.92 5.48 ;
        RECT 48.01 3.405 48.18 5.475 ;
        RECT 46.645 4.135 56.29 4.67 ;
        RECT 46.315 3.2 46.645 4.51 ;
        RECT 39.845 4.34 56.29 4.51 ;
        RECT 44.575 3.8 44.835 4.51 ;
        RECT 44.015 4.34 44.385 4.89 ;
        RECT 43.575 3.42 43.905 3.66 ;
        RECT 43.575 3.42 43.765 3.79 ;
        RECT 43.145 3.69 43.755 4.51 ;
        RECT 43.195 3.69 43.465 5.29 ;
        RECT 42.275 3.8 42.495 4.51 ;
        RECT 42.035 4.34 42.315 5.18 ;
        RECT 41.265 3.47 41.595 3.66 ;
        RECT 40.845 3.84 41.465 4.51 ;
        RECT 41.265 3.47 41.465 4.51 ;
        RECT 41.035 3.84 41.365 5.23 ;
        RECT 39.925 3.83 40.185 4.51 ;
        RECT 30.06 4.345 39.92 4.515 ;
        RECT 36.13 4.13 39.705 4.74 ;
        RECT 36.61 4.13 39.36 4.745 ;
        RECT 36.785 4.13 36.955 5.475 ;
        RECT 30.19 4.135 36.13 4.745 ;
        RECT 33.995 4.13 35.975 4.75 ;
        RECT 35.155 3.4 35.325 5.48 ;
        RECT 34.165 3.4 34.335 5.48 ;
        RECT 31.425 3.405 31.595 5.475 ;
        RECT 30.06 4.135 39.705 4.67 ;
        RECT 29.73 3.2 30.06 4.51 ;
        RECT 23.26 4.34 39.705 4.51 ;
        RECT 27.99 3.8 28.25 4.51 ;
        RECT 27.43 4.34 27.8 4.89 ;
        RECT 26.99 3.42 27.32 3.66 ;
        RECT 26.99 3.42 27.18 3.79 ;
        RECT 26.56 3.69 27.17 4.51 ;
        RECT 26.61 3.69 26.88 5.29 ;
        RECT 25.69 3.8 25.91 4.51 ;
        RECT 25.45 4.34 25.73 5.18 ;
        RECT 24.68 3.47 25.01 3.66 ;
        RECT 24.26 3.84 24.88 4.51 ;
        RECT 24.68 3.47 24.88 4.51 ;
        RECT 24.45 3.84 24.78 5.23 ;
        RECT 23.34 3.83 23.6 4.51 ;
        RECT 13.475 4.345 23.335 4.515 ;
        RECT 19.545 4.13 23.12 4.74 ;
        RECT 20.025 4.13 22.775 4.745 ;
        RECT 20.2 4.13 20.37 5.475 ;
        RECT 13.605 4.135 19.545 4.745 ;
        RECT 17.41 4.13 19.39 4.75 ;
        RECT 18.57 3.4 18.74 5.48 ;
        RECT 17.58 3.4 17.75 5.48 ;
        RECT 14.84 3.405 15.01 5.475 ;
        RECT 13.475 4.135 23.12 4.67 ;
        RECT 13.145 3.2 13.475 4.51 ;
        RECT 6.675 4.34 23.12 4.51 ;
        RECT 11.405 3.8 11.665 4.51 ;
        RECT 10.845 4.34 11.215 4.89 ;
        RECT 10.405 3.42 10.735 3.66 ;
        RECT 10.405 3.42 10.595 3.79 ;
        RECT 9.975 3.69 10.585 4.51 ;
        RECT 10.025 3.69 10.295 5.29 ;
        RECT 9.105 3.8 9.325 4.51 ;
        RECT 8.865 4.34 9.145 5.18 ;
        RECT 8.095 3.47 8.425 3.66 ;
        RECT 7.675 3.84 8.295 4.51 ;
        RECT 8.095 3.47 8.295 4.51 ;
        RECT 7.865 3.84 8.195 5.23 ;
        RECT 6.755 3.83 7.015 4.51 ;
        RECT 0 4.44 6.75 4.515 ;
        RECT 1.805 4.13 6.535 4.74 ;
        RECT 3.44 4.13 6.19 4.745 ;
        RECT 3.615 4.13 3.785 5.475 ;
        RECT 0 4.44 2.96 4.745 ;
        RECT 2.195 4.13 2.365 8.305 ;
        RECT 0 4.13 6.535 4.305 ;
        RECT 0 4.13 1.635 4.745 ;
        RECT 0.385 4.13 0.555 5.475 ;
      LAYER met2 ;
        RECT 1.53 4.23 1.91 4.61 ;
      LAYER met1 ;
        RECT 79.94 4.15 85.88 4.745 ;
        RECT 80.4 4.135 85.88 4.745 ;
        RECT 83.745 4.13 85.725 4.75 ;
        RECT 0 4.19 85.88 4.67 ;
        RECT 79.81 4.15 85.88 4.67 ;
        RECT 69.295 4.13 72.87 4.74 ;
        RECT 69.775 4.13 72.525 4.745 ;
        RECT 63.36 4.15 69.3 4.745 ;
        RECT 63.82 4.135 72.87 4.74 ;
        RECT 67.165 4.13 69.145 4.75 ;
        RECT 63.23 4.15 72.87 4.67 ;
        RECT 52.715 4.13 56.29 4.74 ;
        RECT 53.195 4.13 55.945 4.745 ;
        RECT 46.775 4.15 52.715 4.745 ;
        RECT 47.235 4.135 56.29 4.74 ;
        RECT 50.58 4.13 52.56 4.75 ;
        RECT 46.645 4.15 56.29 4.67 ;
        RECT 36.13 4.13 39.705 4.74 ;
        RECT 36.61 4.13 39.36 4.745 ;
        RECT 30.19 4.15 36.13 4.745 ;
        RECT 30.65 4.135 39.705 4.74 ;
        RECT 33.995 4.13 35.975 4.75 ;
        RECT 30.06 4.15 39.705 4.67 ;
        RECT 19.545 4.13 23.12 4.74 ;
        RECT 20.025 4.13 22.775 4.745 ;
        RECT 13.605 4.15 19.545 4.745 ;
        RECT 14.065 4.135 23.12 4.74 ;
        RECT 17.41 4.13 19.39 4.75 ;
        RECT 13.475 4.15 23.12 4.67 ;
        RECT 0 4.13 6.535 4.74 ;
        RECT 3.44 4.13 6.19 4.745 ;
        RECT 0 4.13 2.96 4.745 ;
        RECT 2.135 6.655 2.425 6.885 ;
        RECT 1.965 6.685 2.425 6.855 ;
      LAYER via2 ;
        RECT 1.62 4.32 1.82 4.52 ;
      LAYER mcon ;
        RECT 2.195 6.685 2.365 6.855 ;
        RECT 2.505 4.545 2.675 4.715 ;
        RECT 5.735 4.545 5.905 4.715 ;
        RECT 6.815 4.34 6.985 4.51 ;
        RECT 7.275 4.34 7.445 4.51 ;
        RECT 7.735 4.34 7.905 4.51 ;
        RECT 8.195 4.34 8.365 4.51 ;
        RECT 8.655 4.34 8.825 4.51 ;
        RECT 9.115 4.34 9.285 4.51 ;
        RECT 9.575 4.34 9.745 4.51 ;
        RECT 10.035 4.34 10.205 4.51 ;
        RECT 10.495 4.34 10.665 4.51 ;
        RECT 10.955 4.34 11.125 4.51 ;
        RECT 11.415 4.34 11.585 4.51 ;
        RECT 11.875 4.34 12.045 4.51 ;
        RECT 12.335 4.34 12.505 4.51 ;
        RECT 12.795 4.34 12.965 4.51 ;
        RECT 13.255 4.34 13.425 4.51 ;
        RECT 16.96 4.545 17.13 4.715 ;
        RECT 16.96 4.165 17.13 4.335 ;
        RECT 17.66 4.55 17.83 4.72 ;
        RECT 17.66 4.16 17.83 4.33 ;
        RECT 18.65 4.55 18.82 4.72 ;
        RECT 18.65 4.16 18.82 4.33 ;
        RECT 22.32 4.545 22.49 4.715 ;
        RECT 23.4 4.34 23.57 4.51 ;
        RECT 23.86 4.34 24.03 4.51 ;
        RECT 24.32 4.34 24.49 4.51 ;
        RECT 24.78 4.34 24.95 4.51 ;
        RECT 25.24 4.34 25.41 4.51 ;
        RECT 25.7 4.34 25.87 4.51 ;
        RECT 26.16 4.34 26.33 4.51 ;
        RECT 26.62 4.34 26.79 4.51 ;
        RECT 27.08 4.34 27.25 4.51 ;
        RECT 27.54 4.34 27.71 4.51 ;
        RECT 28 4.34 28.17 4.51 ;
        RECT 28.46 4.34 28.63 4.51 ;
        RECT 28.92 4.34 29.09 4.51 ;
        RECT 29.38 4.34 29.55 4.51 ;
        RECT 29.84 4.34 30.01 4.51 ;
        RECT 33.545 4.545 33.715 4.715 ;
        RECT 33.545 4.165 33.715 4.335 ;
        RECT 34.245 4.55 34.415 4.72 ;
        RECT 34.245 4.16 34.415 4.33 ;
        RECT 35.235 4.55 35.405 4.72 ;
        RECT 35.235 4.16 35.405 4.33 ;
        RECT 38.905 4.545 39.075 4.715 ;
        RECT 39.985 4.34 40.155 4.51 ;
        RECT 40.445 4.34 40.615 4.51 ;
        RECT 40.905 4.34 41.075 4.51 ;
        RECT 41.365 4.34 41.535 4.51 ;
        RECT 41.825 4.34 41.995 4.51 ;
        RECT 42.285 4.34 42.455 4.51 ;
        RECT 42.745 4.34 42.915 4.51 ;
        RECT 43.205 4.34 43.375 4.51 ;
        RECT 43.665 4.34 43.835 4.51 ;
        RECT 44.125 4.34 44.295 4.51 ;
        RECT 44.585 4.34 44.755 4.51 ;
        RECT 45.045 4.34 45.215 4.51 ;
        RECT 45.505 4.34 45.675 4.51 ;
        RECT 45.965 4.34 46.135 4.51 ;
        RECT 46.425 4.34 46.595 4.51 ;
        RECT 50.13 4.545 50.3 4.715 ;
        RECT 50.13 4.165 50.3 4.335 ;
        RECT 50.83 4.55 51 4.72 ;
        RECT 50.83 4.16 51 4.33 ;
        RECT 51.82 4.55 51.99 4.72 ;
        RECT 51.82 4.16 51.99 4.33 ;
        RECT 55.49 4.545 55.66 4.715 ;
        RECT 56.57 4.34 56.74 4.51 ;
        RECT 57.03 4.34 57.2 4.51 ;
        RECT 57.49 4.34 57.66 4.51 ;
        RECT 57.95 4.34 58.12 4.51 ;
        RECT 58.41 4.34 58.58 4.51 ;
        RECT 58.87 4.34 59.04 4.51 ;
        RECT 59.33 4.34 59.5 4.51 ;
        RECT 59.79 4.34 59.96 4.51 ;
        RECT 60.25 4.34 60.42 4.51 ;
        RECT 60.71 4.34 60.88 4.51 ;
        RECT 61.17 4.34 61.34 4.51 ;
        RECT 61.63 4.34 61.8 4.51 ;
        RECT 62.09 4.34 62.26 4.51 ;
        RECT 62.55 4.34 62.72 4.51 ;
        RECT 63.01 4.34 63.18 4.51 ;
        RECT 66.715 4.545 66.885 4.715 ;
        RECT 66.715 4.165 66.885 4.335 ;
        RECT 67.415 4.55 67.585 4.72 ;
        RECT 67.415 4.16 67.585 4.33 ;
        RECT 68.405 4.55 68.575 4.72 ;
        RECT 68.405 4.16 68.575 4.33 ;
        RECT 72.07 4.545 72.24 4.715 ;
        RECT 73.15 4.34 73.32 4.51 ;
        RECT 73.61 4.34 73.78 4.51 ;
        RECT 74.07 4.34 74.24 4.51 ;
        RECT 74.53 4.34 74.7 4.51 ;
        RECT 74.99 4.34 75.16 4.51 ;
        RECT 75.45 4.34 75.62 4.51 ;
        RECT 75.91 4.34 76.08 4.51 ;
        RECT 76.37 4.34 76.54 4.51 ;
        RECT 76.83 4.34 77 4.51 ;
        RECT 77.29 4.34 77.46 4.51 ;
        RECT 77.75 4.34 77.92 4.51 ;
        RECT 78.21 4.34 78.38 4.51 ;
        RECT 78.67 4.34 78.84 4.51 ;
        RECT 79.13 4.34 79.3 4.51 ;
        RECT 79.59 4.34 79.76 4.51 ;
        RECT 83.295 4.545 83.465 4.715 ;
        RECT 83.295 4.165 83.465 4.335 ;
        RECT 83.995 4.55 84.165 4.72 ;
        RECT 83.995 4.16 84.165 4.33 ;
        RECT 84.985 4.55 85.155 4.72 ;
        RECT 84.985 4.16 85.155 4.33 ;
      LAYER via1 ;
        RECT 1.645 4.345 1.795 4.495 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 75.38 6.47 75.71 6.8 ;
        RECT 75.35 6.49 75.65 6.9 ;
        RECT 74.91 6.49 75.71 6.79 ;
        RECT 58.8 6.47 59.13 6.8 ;
        RECT 58.77 6.49 59.07 6.9 ;
        RECT 58.33 6.49 59.13 6.79 ;
        RECT 42.215 6.47 42.545 6.8 ;
        RECT 42.185 6.49 42.485 6.9 ;
        RECT 41.745 6.49 42.545 6.79 ;
        RECT 25.63 6.47 25.96 6.8 ;
        RECT 25.6 6.49 25.9 6.9 ;
        RECT 25.16 6.49 25.96 6.79 ;
        RECT 9.045 6.47 9.375 6.8 ;
        RECT 9.015 6.49 9.315 6.9 ;
        RECT 8.575 6.49 9.375 6.79 ;
        RECT 0.17 8.5 0.975 8.88 ;
        RECT 0 0 0.805 0.38 ;
      LAYER li1 ;
        RECT 85.7 0 85.88 0.305 ;
        RECT 0.465 0 85.88 0.3 ;
        RECT 84.905 0 85.075 0.93 ;
        RECT 83.915 0 84.085 0.93 ;
        RECT 69.12 0 83.75 0.305 ;
        RECT 81.175 0 81.345 0.935 ;
        RECT 79.905 0 80.1 1.795 ;
        RECT 73.01 0 80.1 1.79 ;
        RECT 79.54 0 79.81 2.6 ;
        RECT 78.63 0 78.87 2.6 ;
        RECT 77.76 0 78.01 2.33 ;
        RECT 75.38 0 75.71 2.25 ;
        RECT 73.09 0 73.35 2.61 ;
        RECT 72.755 0 80.1 1.655 ;
        RECT 68.325 0 68.495 0.93 ;
        RECT 67.335 0 67.505 0.93 ;
        RECT 52.535 0 67.17 0.305 ;
        RECT 64.595 0 64.765 0.935 ;
        RECT 63.325 0 63.52 1.795 ;
        RECT 56.43 0 63.52 1.79 ;
        RECT 62.96 0 63.23 2.6 ;
        RECT 62.05 0 62.29 2.6 ;
        RECT 61.18 0 61.43 2.33 ;
        RECT 58.8 0 59.13 2.25 ;
        RECT 56.51 0 56.77 2.61 ;
        RECT 56.175 0 63.52 1.655 ;
        RECT 51.74 0 51.91 0.93 ;
        RECT 50.75 0 50.92 0.93 ;
        RECT 35.95 0 50.585 0.305 ;
        RECT 48.01 0 48.18 0.935 ;
        RECT 46.74 0 46.935 1.795 ;
        RECT 39.845 0 46.935 1.79 ;
        RECT 46.375 0 46.645 2.6 ;
        RECT 45.465 0 45.705 2.6 ;
        RECT 44.595 0 44.845 2.33 ;
        RECT 42.215 0 42.545 2.25 ;
        RECT 39.925 0 40.185 2.61 ;
        RECT 39.59 0 46.935 1.655 ;
        RECT 35.155 0 35.325 0.93 ;
        RECT 34.165 0 34.335 0.93 ;
        RECT 19.365 0 34 0.305 ;
        RECT 31.425 0 31.595 0.935 ;
        RECT 30.155 0 30.35 1.795 ;
        RECT 23.26 0 30.35 1.79 ;
        RECT 29.79 0 30.06 2.6 ;
        RECT 28.88 0 29.12 2.6 ;
        RECT 28.01 0 28.26 2.33 ;
        RECT 25.63 0 25.96 2.25 ;
        RECT 23.34 0 23.6 2.61 ;
        RECT 23.005 0 30.35 1.655 ;
        RECT 18.57 0 18.74 0.93 ;
        RECT 17.58 0 17.75 0.93 ;
        RECT 0 0.245 17.415 0.305 ;
        RECT 14.84 0 15.01 0.935 ;
        RECT 13.57 0 13.765 1.795 ;
        RECT 6.675 0 13.765 1.79 ;
        RECT 13.205 0 13.475 2.6 ;
        RECT 12.295 0 12.535 2.6 ;
        RECT 11.425 0 11.675 2.33 ;
        RECT 9.045 0 9.375 2.25 ;
        RECT 6.755 0 7.015 2.61 ;
        RECT 6.42 0 13.765 1.655 ;
        RECT 0 0.245 0.805 0.315 ;
        RECT 0.295 0.245 0.465 0.335 ;
        RECT 0 0 85.88 0.075 ;
        RECT 0 0 0.295 0.315 ;
        RECT 0 8.58 85.88 8.88 ;
        RECT 85.7 8.575 85.88 8.88 ;
        RECT 84.905 7.95 85.075 8.88 ;
        RECT 83.915 7.95 84.085 8.88 ;
        RECT 69.12 8.575 83.75 8.88 ;
        RECT 81.175 7.945 81.345 8.88 ;
        RECT 72.715 7.18 79.915 8.88 ;
        RECT 73.01 7.06 79.91 8.88 ;
        RECT 78.44 6.55 78.89 8.88 ;
        RECT 76.35 6.66 76.68 8.88 ;
        RECT 74.28 6.6 74.53 8.88 ;
        RECT 69.95 7.945 70.12 8.88 ;
        RECT 68.325 7.95 68.495 8.88 ;
        RECT 67.335 7.95 67.505 8.88 ;
        RECT 52.535 8.575 67.17 8.88 ;
        RECT 64.595 7.945 64.765 8.88 ;
        RECT 56.135 7.18 63.335 8.88 ;
        RECT 56.43 7.06 63.33 8.88 ;
        RECT 61.86 6.55 62.31 8.88 ;
        RECT 59.77 6.66 60.1 8.88 ;
        RECT 57.7 6.6 57.95 8.88 ;
        RECT 53.37 7.945 53.54 8.88 ;
        RECT 51.74 7.95 51.91 8.88 ;
        RECT 50.75 7.95 50.92 8.88 ;
        RECT 35.95 8.575 50.585 8.88 ;
        RECT 48.01 7.945 48.18 8.88 ;
        RECT 39.55 7.18 46.75 8.88 ;
        RECT 39.845 7.06 46.745 8.88 ;
        RECT 45.275 6.55 45.725 8.88 ;
        RECT 43.185 6.66 43.515 8.88 ;
        RECT 41.115 6.6 41.365 8.88 ;
        RECT 36.785 7.945 36.955 8.88 ;
        RECT 35.155 7.95 35.325 8.88 ;
        RECT 34.165 7.95 34.335 8.88 ;
        RECT 19.365 8.575 34 8.88 ;
        RECT 31.425 7.945 31.595 8.88 ;
        RECT 22.965 7.18 30.165 8.88 ;
        RECT 23.26 7.06 30.16 8.88 ;
        RECT 28.69 6.55 29.14 8.88 ;
        RECT 26.6 6.66 26.93 8.88 ;
        RECT 24.53 6.6 24.78 8.88 ;
        RECT 20.2 7.945 20.37 8.88 ;
        RECT 18.57 7.95 18.74 8.88 ;
        RECT 17.58 7.95 17.75 8.88 ;
        RECT 0 8.575 17.415 8.88 ;
        RECT 14.84 7.945 15.01 8.88 ;
        RECT 6.38 7.18 13.58 8.88 ;
        RECT 6.675 7.06 13.575 8.88 ;
        RECT 12.105 6.55 12.555 8.88 ;
        RECT 10.015 6.66 10.345 8.88 ;
        RECT 7.945 6.6 8.195 8.88 ;
        RECT 3.615 7.945 3.785 8.88 ;
        RECT 0.17 8.565 0.975 8.88 ;
        RECT 0.385 8.545 0.635 8.88 ;
        RECT 0.385 7.945 0.555 8.88 ;
        RECT 76.65 5.82 76.98 6.15 ;
        RECT 74.43 5.82 74.77 6.07 ;
        RECT 70.955 6.075 71.125 8.025 ;
        RECT 70.9 7.855 71.07 8.305 ;
        RECT 70.9 5.015 71.07 6.245 ;
        RECT 60.07 5.82 60.4 6.15 ;
        RECT 57.85 5.82 58.19 6.07 ;
        RECT 54.375 6.075 54.545 8.025 ;
        RECT 54.32 7.855 54.49 8.305 ;
        RECT 54.32 5.015 54.49 6.245 ;
        RECT 43.485 5.82 43.815 6.15 ;
        RECT 41.265 5.82 41.605 6.07 ;
        RECT 37.79 6.075 37.96 8.025 ;
        RECT 37.735 7.855 37.905 8.305 ;
        RECT 37.735 5.015 37.905 6.245 ;
        RECT 26.9 5.82 27.23 6.15 ;
        RECT 24.68 5.82 25.02 6.07 ;
        RECT 21.205 6.075 21.375 8.025 ;
        RECT 21.15 7.855 21.32 8.305 ;
        RECT 21.15 5.015 21.32 6.245 ;
        RECT 10.315 5.82 10.645 6.15 ;
        RECT 8.095 5.82 8.435 6.07 ;
        RECT 4.62 6.075 4.79 8.025 ;
        RECT 4.565 7.855 4.735 8.305 ;
        RECT 4.565 5.015 4.735 6.245 ;
      LAYER met2 ;
        RECT 75.41 6.45 75.69 6.82 ;
        RECT 58.83 6.45 59.11 6.82 ;
        RECT 42.245 6.45 42.525 6.82 ;
        RECT 25.66 6.45 25.94 6.82 ;
        RECT 9.075 6.45 9.355 6.82 ;
        RECT 0.36 8.5 0.74 8.88 ;
        RECT 0.19 0 0.57 0.38 ;
        RECT 0.235 0 0.405 8.82 ;
      LAYER met1 ;
        RECT 85.7 0 85.88 0.305 ;
        RECT 0 0 85.88 0.3 ;
        RECT 69.12 0 83.75 0.305 ;
        RECT 73.01 0 80.1 1.795 ;
        RECT 73.01 0 79.91 1.95 ;
        RECT 72.755 0 80.1 1.655 ;
        RECT 52.535 0 67.17 0.305 ;
        RECT 56.43 0 63.52 1.795 ;
        RECT 56.43 0 63.33 1.95 ;
        RECT 56.175 0 63.52 1.655 ;
        RECT 35.95 0 50.585 0.305 ;
        RECT 39.845 0 46.935 1.795 ;
        RECT 39.845 0 46.745 1.95 ;
        RECT 39.59 0 46.935 1.655 ;
        RECT 19.365 0 34 0.305 ;
        RECT 23.26 0 30.35 1.795 ;
        RECT 23.26 0 30.16 1.95 ;
        RECT 23.005 0 30.35 1.655 ;
        RECT 0 0 17.415 0.305 ;
        RECT 6.675 0 13.765 1.795 ;
        RECT 6.675 0 13.575 1.95 ;
        RECT 6.42 0 13.765 1.655 ;
        RECT 0 0 0.805 0.315 ;
        RECT 0.205 0 0.555 0.335 ;
        RECT 0 8.58 85.88 8.88 ;
        RECT 85.7 8.575 85.88 8.88 ;
        RECT 69.12 8.575 83.75 8.88 ;
        RECT 72.715 7.18 79.915 8.88 ;
        RECT 73.01 6.91 79.91 8.88 ;
        RECT 76.6 5.84 76.89 6.07 ;
        RECT 74.47 6.57 76.82 6.71 ;
        RECT 76.68 5.84 76.82 6.71 ;
        RECT 75.4 6.51 75.72 6.77 ;
        RECT 75.435 6.51 75.69 8.88 ;
        RECT 74.39 5.84 74.68 6.07 ;
        RECT 74.47 5.84 74.61 6.71 ;
        RECT 70.895 6.285 71.185 6.515 ;
        RECT 70.735 6.315 70.905 8.88 ;
        RECT 70.725 6.315 71.185 6.485 ;
        RECT 52.535 8.575 67.17 8.88 ;
        RECT 56.135 7.18 63.335 8.88 ;
        RECT 56.43 6.91 63.33 8.88 ;
        RECT 60.02 5.84 60.31 6.07 ;
        RECT 57.89 6.57 60.24 6.71 ;
        RECT 60.1 5.84 60.24 6.71 ;
        RECT 58.82 6.51 59.14 6.77 ;
        RECT 58.855 6.51 59.11 8.88 ;
        RECT 57.81 5.84 58.1 6.07 ;
        RECT 57.89 5.84 58.03 6.71 ;
        RECT 54.315 6.285 54.605 6.515 ;
        RECT 54.155 6.315 54.325 8.88 ;
        RECT 54.145 6.315 54.605 6.485 ;
        RECT 35.95 8.575 50.585 8.88 ;
        RECT 39.55 7.18 46.75 8.88 ;
        RECT 39.845 6.91 46.745 8.88 ;
        RECT 43.435 5.84 43.725 6.07 ;
        RECT 41.305 6.57 43.655 6.71 ;
        RECT 43.515 5.84 43.655 6.71 ;
        RECT 42.235 6.51 42.555 6.77 ;
        RECT 42.27 6.51 42.525 8.88 ;
        RECT 41.225 5.84 41.515 6.07 ;
        RECT 41.305 5.84 41.445 6.71 ;
        RECT 37.73 6.285 38.02 6.515 ;
        RECT 37.57 6.315 37.74 8.88 ;
        RECT 37.56 6.315 38.02 6.485 ;
        RECT 19.365 8.575 34 8.88 ;
        RECT 22.965 7.18 30.165 8.88 ;
        RECT 23.26 6.91 30.16 8.88 ;
        RECT 26.85 5.84 27.14 6.07 ;
        RECT 24.72 6.57 27.07 6.71 ;
        RECT 26.93 5.84 27.07 6.71 ;
        RECT 25.65 6.51 25.97 6.77 ;
        RECT 25.685 6.51 25.94 8.88 ;
        RECT 24.64 5.84 24.93 6.07 ;
        RECT 24.72 5.84 24.86 6.71 ;
        RECT 21.145 6.285 21.435 6.515 ;
        RECT 20.985 6.315 21.155 8.88 ;
        RECT 20.975 6.315 21.435 6.485 ;
        RECT 0 8.575 17.415 8.88 ;
        RECT 6.38 7.18 13.58 8.88 ;
        RECT 6.675 6.91 13.575 8.88 ;
        RECT 10.265 5.84 10.555 6.07 ;
        RECT 8.135 6.57 10.485 6.71 ;
        RECT 10.345 5.84 10.485 6.71 ;
        RECT 9.065 6.51 9.385 6.77 ;
        RECT 9.1 6.51 9.355 8.88 ;
        RECT 8.055 5.84 8.345 6.07 ;
        RECT 8.135 5.84 8.275 6.71 ;
        RECT 4.56 6.285 4.85 6.515 ;
        RECT 4.4 6.315 4.57 8.88 ;
        RECT 4.39 6.315 4.85 6.485 ;
        RECT 0.17 8.565 0.975 8.88 ;
        RECT 0.375 8.545 0.725 8.88 ;
      LAYER via2 ;
        RECT 0.28 0.09 0.48 0.29 ;
        RECT 0.45 8.59 0.65 8.79 ;
        RECT 9.115 6.54 9.315 6.74 ;
        RECT 25.7 6.54 25.9 6.74 ;
        RECT 42.285 6.54 42.485 6.74 ;
        RECT 58.87 6.54 59.07 6.74 ;
        RECT 75.45 6.54 75.65 6.74 ;
      LAYER mcon ;
        RECT 0.465 8.605 0.635 8.775 ;
        RECT 1.145 8.605 1.315 8.775 ;
        RECT 1.825 8.605 1.995 8.775 ;
        RECT 2.505 8.605 2.675 8.775 ;
        RECT 3.695 8.605 3.865 8.775 ;
        RECT 4.375 8.605 4.545 8.775 ;
        RECT 4.62 6.315 4.79 6.485 ;
        RECT 5.055 8.605 5.225 8.775 ;
        RECT 5.735 8.605 5.905 8.775 ;
        RECT 6.815 7.06 6.985 7.23 ;
        RECT 7.275 7.06 7.445 7.23 ;
        RECT 7.735 7.06 7.905 7.23 ;
        RECT 8.115 5.87 8.285 6.04 ;
        RECT 8.195 7.06 8.365 7.23 ;
        RECT 8.655 7.06 8.825 7.23 ;
        RECT 9.115 7.06 9.285 7.23 ;
        RECT 9.575 7.06 9.745 7.23 ;
        RECT 10.035 7.06 10.205 7.23 ;
        RECT 10.325 5.87 10.495 6.04 ;
        RECT 10.495 7.06 10.665 7.23 ;
        RECT 10.955 7.06 11.125 7.23 ;
        RECT 11.415 7.06 11.585 7.23 ;
        RECT 11.875 7.06 12.045 7.23 ;
        RECT 12.335 7.06 12.505 7.23 ;
        RECT 12.795 7.06 12.965 7.23 ;
        RECT 13.255 7.06 13.425 7.23 ;
        RECT 14.92 8.605 15.09 8.775 ;
        RECT 14.92 0.105 15.09 0.275 ;
        RECT 15.6 8.605 15.77 8.775 ;
        RECT 15.6 0.105 15.77 0.275 ;
        RECT 16.28 8.605 16.45 8.775 ;
        RECT 16.28 0.105 16.45 0.275 ;
        RECT 16.96 8.605 17.13 8.775 ;
        RECT 16.96 0.105 17.13 0.275 ;
        RECT 17.66 8.61 17.83 8.78 ;
        RECT 17.66 0.1 17.83 0.27 ;
        RECT 18.65 8.61 18.82 8.78 ;
        RECT 18.65 0.1 18.82 0.27 ;
        RECT 20.28 8.605 20.45 8.775 ;
        RECT 20.96 8.605 21.13 8.775 ;
        RECT 21.205 6.315 21.375 6.485 ;
        RECT 21.64 8.605 21.81 8.775 ;
        RECT 22.32 8.605 22.49 8.775 ;
        RECT 23.4 7.06 23.57 7.23 ;
        RECT 23.86 7.06 24.03 7.23 ;
        RECT 24.32 7.06 24.49 7.23 ;
        RECT 24.7 5.87 24.87 6.04 ;
        RECT 24.78 7.06 24.95 7.23 ;
        RECT 25.24 7.06 25.41 7.23 ;
        RECT 25.7 7.06 25.87 7.23 ;
        RECT 26.16 7.06 26.33 7.23 ;
        RECT 26.62 7.06 26.79 7.23 ;
        RECT 26.91 5.87 27.08 6.04 ;
        RECT 27.08 7.06 27.25 7.23 ;
        RECT 27.54 7.06 27.71 7.23 ;
        RECT 28 7.06 28.17 7.23 ;
        RECT 28.46 7.06 28.63 7.23 ;
        RECT 28.92 7.06 29.09 7.23 ;
        RECT 29.38 7.06 29.55 7.23 ;
        RECT 29.84 7.06 30.01 7.23 ;
        RECT 31.505 8.605 31.675 8.775 ;
        RECT 31.505 0.105 31.675 0.275 ;
        RECT 32.185 8.605 32.355 8.775 ;
        RECT 32.185 0.105 32.355 0.275 ;
        RECT 32.865 8.605 33.035 8.775 ;
        RECT 32.865 0.105 33.035 0.275 ;
        RECT 33.545 8.605 33.715 8.775 ;
        RECT 33.545 0.105 33.715 0.275 ;
        RECT 34.245 8.61 34.415 8.78 ;
        RECT 34.245 0.1 34.415 0.27 ;
        RECT 35.235 8.61 35.405 8.78 ;
        RECT 35.235 0.1 35.405 0.27 ;
        RECT 36.865 8.605 37.035 8.775 ;
        RECT 37.545 8.605 37.715 8.775 ;
        RECT 37.79 6.315 37.96 6.485 ;
        RECT 38.225 8.605 38.395 8.775 ;
        RECT 38.905 8.605 39.075 8.775 ;
        RECT 39.985 7.06 40.155 7.23 ;
        RECT 40.445 7.06 40.615 7.23 ;
        RECT 40.905 7.06 41.075 7.23 ;
        RECT 41.285 5.87 41.455 6.04 ;
        RECT 41.365 7.06 41.535 7.23 ;
        RECT 41.825 7.06 41.995 7.23 ;
        RECT 42.285 7.06 42.455 7.23 ;
        RECT 42.745 7.06 42.915 7.23 ;
        RECT 43.205 7.06 43.375 7.23 ;
        RECT 43.495 5.87 43.665 6.04 ;
        RECT 43.665 7.06 43.835 7.23 ;
        RECT 44.125 7.06 44.295 7.23 ;
        RECT 44.585 7.06 44.755 7.23 ;
        RECT 45.045 7.06 45.215 7.23 ;
        RECT 45.505 7.06 45.675 7.23 ;
        RECT 45.965 7.06 46.135 7.23 ;
        RECT 46.425 7.06 46.595 7.23 ;
        RECT 48.09 8.605 48.26 8.775 ;
        RECT 48.09 0.105 48.26 0.275 ;
        RECT 48.77 8.605 48.94 8.775 ;
        RECT 48.77 0.105 48.94 0.275 ;
        RECT 49.45 8.605 49.62 8.775 ;
        RECT 49.45 0.105 49.62 0.275 ;
        RECT 50.13 8.605 50.3 8.775 ;
        RECT 50.13 0.105 50.3 0.275 ;
        RECT 50.83 8.61 51 8.78 ;
        RECT 50.83 0.1 51 0.27 ;
        RECT 51.82 8.61 51.99 8.78 ;
        RECT 51.82 0.1 51.99 0.27 ;
        RECT 53.45 8.605 53.62 8.775 ;
        RECT 54.13 8.605 54.3 8.775 ;
        RECT 54.375 6.315 54.545 6.485 ;
        RECT 54.81 8.605 54.98 8.775 ;
        RECT 55.49 8.605 55.66 8.775 ;
        RECT 56.57 7.06 56.74 7.23 ;
        RECT 57.03 7.06 57.2 7.23 ;
        RECT 57.49 7.06 57.66 7.23 ;
        RECT 57.87 5.87 58.04 6.04 ;
        RECT 57.95 7.06 58.12 7.23 ;
        RECT 58.41 7.06 58.58 7.23 ;
        RECT 58.87 7.06 59.04 7.23 ;
        RECT 59.33 7.06 59.5 7.23 ;
        RECT 59.79 7.06 59.96 7.23 ;
        RECT 60.08 5.87 60.25 6.04 ;
        RECT 60.25 7.06 60.42 7.23 ;
        RECT 60.71 7.06 60.88 7.23 ;
        RECT 61.17 7.06 61.34 7.23 ;
        RECT 61.63 7.06 61.8 7.23 ;
        RECT 62.09 7.06 62.26 7.23 ;
        RECT 62.55 7.06 62.72 7.23 ;
        RECT 63.01 7.06 63.18 7.23 ;
        RECT 64.675 8.605 64.845 8.775 ;
        RECT 64.675 0.105 64.845 0.275 ;
        RECT 65.355 8.605 65.525 8.775 ;
        RECT 65.355 0.105 65.525 0.275 ;
        RECT 66.035 8.605 66.205 8.775 ;
        RECT 66.035 0.105 66.205 0.275 ;
        RECT 66.715 8.605 66.885 8.775 ;
        RECT 66.715 0.105 66.885 0.275 ;
        RECT 67.415 8.61 67.585 8.78 ;
        RECT 67.415 0.1 67.585 0.27 ;
        RECT 68.405 8.61 68.575 8.78 ;
        RECT 68.405 0.1 68.575 0.27 ;
        RECT 70.03 8.605 70.2 8.775 ;
        RECT 70.71 8.605 70.88 8.775 ;
        RECT 70.955 6.315 71.125 6.485 ;
        RECT 71.39 8.605 71.56 8.775 ;
        RECT 72.07 8.605 72.24 8.775 ;
        RECT 73.15 7.06 73.32 7.23 ;
        RECT 73.61 7.06 73.78 7.23 ;
        RECT 74.07 7.06 74.24 7.23 ;
        RECT 74.45 5.87 74.62 6.04 ;
        RECT 74.53 7.06 74.7 7.23 ;
        RECT 74.99 7.06 75.16 7.23 ;
        RECT 75.45 7.06 75.62 7.23 ;
        RECT 75.91 7.06 76.08 7.23 ;
        RECT 76.37 7.06 76.54 7.23 ;
        RECT 76.66 5.87 76.83 6.04 ;
        RECT 76.83 7.06 77 7.23 ;
        RECT 77.29 7.06 77.46 7.23 ;
        RECT 77.75 7.06 77.92 7.23 ;
        RECT 78.21 7.06 78.38 7.23 ;
        RECT 78.67 7.06 78.84 7.23 ;
        RECT 79.13 7.06 79.3 7.23 ;
        RECT 79.59 7.06 79.76 7.23 ;
        RECT 81.255 8.605 81.425 8.775 ;
        RECT 81.255 0.105 81.425 0.275 ;
        RECT 81.935 8.605 82.105 8.775 ;
        RECT 81.935 0.105 82.105 0.275 ;
        RECT 82.615 8.605 82.785 8.775 ;
        RECT 82.615 0.105 82.785 0.275 ;
        RECT 83.295 8.605 83.465 8.775 ;
        RECT 83.295 0.105 83.465 0.275 ;
        RECT 83.995 8.61 84.165 8.78 ;
        RECT 83.995 0.1 84.165 0.27 ;
        RECT 84.985 8.61 85.155 8.78 ;
        RECT 84.985 0.1 85.155 0.27 ;
      LAYER via1 ;
        RECT 0.305 0.115 0.455 0.265 ;
        RECT 0.475 8.615 0.625 8.765 ;
        RECT 9.15 6.565 9.3 6.715 ;
        RECT 25.735 6.565 25.885 6.715 ;
        RECT 42.32 6.565 42.47 6.715 ;
        RECT 58.905 6.565 59.055 6.715 ;
        RECT 75.485 6.565 75.635 6.715 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 77.805 2.73 78.105 3.065 ;
      RECT 77.78 2.73 78.11 3.06 ;
      RECT 77.78 2.75 78.58 3.05 ;
      RECT 72.105 7.97 76.385 8.27 ;
      RECT 76.08 5.79 76.38 8.27 ;
      RECT 72.105 7.03 72.405 8.27 ;
      RECT 71.23 6.995 71.6 7.365 ;
      RECT 71.23 7.03 72.405 7.33 ;
      RECT 75.455 5.795 76.39 6.125 ;
      RECT 76.06 5.79 76.39 6.125 ;
      RECT 77.1 5.79 77.43 6.12 ;
      RECT 75.455 5.81 77.9 6.11 ;
      RECT 75.455 5.795 77.43 6.11 ;
      RECT 75.455 3.765 75.785 6.125 ;
      RECT 75.455 3.765 77.75 4.095 ;
      RECT 75.455 3.765 78.105 4.085 ;
      RECT 77.78 3.75 78.11 4.08 ;
      RECT 75.455 3.77 78.58 4.07 ;
      RECT 77.79 3.7 78.09 4.085 ;
      RECT 77.08 3.07 77.41 3.4 ;
      RECT 77.11 3.06 77.41 3.4 ;
      RECT 76.61 3.09 77.41 3.39 ;
      RECT 76.425 4.77 76.46 5.105 ;
      RECT 76.42 4.77 76.75 5.1 ;
      RECT 76.42 4.79 77.22 5.09 ;
      RECT 76.42 4.785 76.755 5.09 ;
      RECT 75.74 2.39 76.07 2.72 ;
      RECT 75.27 2.41 75.63 2.71 ;
      RECT 75.63 2.4 76.07 2.7 ;
      RECT 61.225 2.73 61.525 3.065 ;
      RECT 61.2 2.73 61.53 3.06 ;
      RECT 61.2 2.75 62 3.05 ;
      RECT 55.525 7.97 59.805 8.27 ;
      RECT 59.5 5.79 59.8 8.27 ;
      RECT 55.525 7.03 55.825 8.27 ;
      RECT 54.65 6.995 55.02 7.365 ;
      RECT 54.65 7.03 55.825 7.33 ;
      RECT 58.875 5.795 59.81 6.125 ;
      RECT 59.48 5.79 59.81 6.125 ;
      RECT 60.52 5.79 60.85 6.12 ;
      RECT 58.875 5.81 61.32 6.11 ;
      RECT 58.875 5.795 60.85 6.11 ;
      RECT 58.875 3.765 59.205 6.125 ;
      RECT 58.875 3.765 61.17 4.095 ;
      RECT 58.875 3.765 61.525 4.085 ;
      RECT 61.2 3.75 61.53 4.08 ;
      RECT 58.875 3.77 62 4.07 ;
      RECT 61.21 3.7 61.51 4.085 ;
      RECT 60.5 3.07 60.83 3.4 ;
      RECT 60.53 3.06 60.83 3.4 ;
      RECT 60.03 3.09 60.83 3.39 ;
      RECT 59.845 4.77 59.88 5.105 ;
      RECT 59.84 4.77 60.17 5.1 ;
      RECT 59.84 4.79 60.64 5.09 ;
      RECT 59.84 4.785 60.175 5.09 ;
      RECT 59.16 2.39 59.49 2.72 ;
      RECT 58.69 2.41 59.05 2.71 ;
      RECT 59.05 2.4 59.49 2.7 ;
      RECT 44.64 2.73 44.94 3.065 ;
      RECT 44.615 2.73 44.945 3.06 ;
      RECT 44.615 2.75 45.415 3.05 ;
      RECT 38.94 7.97 43.22 8.27 ;
      RECT 42.915 5.79 43.215 8.27 ;
      RECT 38.94 7.03 39.24 8.27 ;
      RECT 38.065 6.995 38.435 7.365 ;
      RECT 38.065 7.03 39.24 7.33 ;
      RECT 42.29 5.795 43.225 6.125 ;
      RECT 42.895 5.79 43.225 6.125 ;
      RECT 43.935 5.79 44.265 6.12 ;
      RECT 42.29 5.81 44.735 6.11 ;
      RECT 42.29 5.795 44.265 6.11 ;
      RECT 42.29 3.765 42.62 6.125 ;
      RECT 42.29 3.765 44.585 4.095 ;
      RECT 42.29 3.765 44.94 4.085 ;
      RECT 44.615 3.75 44.945 4.08 ;
      RECT 42.29 3.77 45.415 4.07 ;
      RECT 44.625 3.7 44.925 4.085 ;
      RECT 43.915 3.07 44.245 3.4 ;
      RECT 43.945 3.06 44.245 3.4 ;
      RECT 43.445 3.09 44.245 3.39 ;
      RECT 43.26 4.77 43.295 5.105 ;
      RECT 43.255 4.77 43.585 5.1 ;
      RECT 43.255 4.79 44.055 5.09 ;
      RECT 43.255 4.785 43.59 5.09 ;
      RECT 42.575 2.39 42.905 2.72 ;
      RECT 42.105 2.41 42.465 2.71 ;
      RECT 42.465 2.4 42.905 2.7 ;
      RECT 28.055 2.73 28.355 3.065 ;
      RECT 28.03 2.73 28.36 3.06 ;
      RECT 28.03 2.75 28.83 3.05 ;
      RECT 22.355 7.97 26.635 8.27 ;
      RECT 26.33 5.79 26.63 8.27 ;
      RECT 22.355 7.03 22.655 8.27 ;
      RECT 21.48 6.995 21.85 7.365 ;
      RECT 21.48 7.03 22.655 7.33 ;
      RECT 25.705 5.795 26.64 6.125 ;
      RECT 26.31 5.79 26.64 6.125 ;
      RECT 27.35 5.79 27.68 6.12 ;
      RECT 25.705 5.81 28.15 6.11 ;
      RECT 25.705 5.795 27.68 6.11 ;
      RECT 25.705 3.765 26.035 6.125 ;
      RECT 25.705 3.765 28 4.095 ;
      RECT 25.705 3.765 28.355 4.085 ;
      RECT 28.03 3.75 28.36 4.08 ;
      RECT 25.705 3.77 28.83 4.07 ;
      RECT 28.04 3.7 28.34 4.085 ;
      RECT 27.33 3.07 27.66 3.4 ;
      RECT 27.36 3.06 27.66 3.4 ;
      RECT 26.86 3.09 27.66 3.39 ;
      RECT 26.675 4.77 26.71 5.105 ;
      RECT 26.67 4.77 27 5.1 ;
      RECT 26.67 4.79 27.47 5.09 ;
      RECT 26.67 4.785 27.005 5.09 ;
      RECT 25.99 2.39 26.32 2.72 ;
      RECT 25.52 2.41 25.88 2.71 ;
      RECT 25.88 2.4 26.32 2.7 ;
      RECT 11.47 2.73 11.77 3.065 ;
      RECT 11.445 2.73 11.775 3.06 ;
      RECT 11.445 2.75 12.245 3.05 ;
      RECT 5.77 7.97 10.05 8.27 ;
      RECT 9.745 5.79 10.045 8.27 ;
      RECT 5.77 7.03 6.07 8.27 ;
      RECT 4.895 6.995 5.265 7.365 ;
      RECT 4.895 7.03 6.07 7.33 ;
      RECT 9.12 5.795 10.055 6.125 ;
      RECT 9.725 5.79 10.055 6.125 ;
      RECT 10.765 5.79 11.095 6.12 ;
      RECT 9.12 5.81 11.565 6.11 ;
      RECT 9.12 5.795 11.095 6.11 ;
      RECT 9.12 3.765 9.45 6.125 ;
      RECT 9.12 3.765 11.415 4.095 ;
      RECT 9.12 3.765 11.77 4.085 ;
      RECT 11.445 3.75 11.775 4.08 ;
      RECT 9.12 3.77 12.245 4.07 ;
      RECT 11.455 3.7 11.755 4.085 ;
      RECT 10.745 3.07 11.075 3.4 ;
      RECT 10.775 3.06 11.075 3.4 ;
      RECT 10.275 3.09 11.075 3.39 ;
      RECT 10.09 4.77 10.125 5.105 ;
      RECT 10.085 4.77 10.415 5.1 ;
      RECT 10.085 4.79 10.885 5.09 ;
      RECT 10.085 4.785 10.42 5.09 ;
      RECT 9.405 2.39 9.735 2.72 ;
      RECT 8.935 2.41 9.295 2.71 ;
      RECT 9.295 2.4 9.735 2.7 ;
    LAYER via2 ;
      RECT 77.85 2.8 78.05 3 ;
      RECT 77.85 3.82 78.05 4.02 ;
      RECT 77.17 5.86 77.37 6.06 ;
      RECT 77.15 3.14 77.35 3.34 ;
      RECT 76.49 4.84 76.69 5.04 ;
      RECT 76.12 5.86 76.32 6.06 ;
      RECT 75.81 2.45 76.01 2.65 ;
      RECT 71.315 7.08 71.515 7.28 ;
      RECT 61.27 2.8 61.47 3 ;
      RECT 61.27 3.82 61.47 4.02 ;
      RECT 60.59 5.86 60.79 6.06 ;
      RECT 60.57 3.14 60.77 3.34 ;
      RECT 59.91 4.84 60.11 5.04 ;
      RECT 59.54 5.86 59.74 6.06 ;
      RECT 59.23 2.45 59.43 2.65 ;
      RECT 54.735 7.08 54.935 7.28 ;
      RECT 44.685 2.8 44.885 3 ;
      RECT 44.685 3.82 44.885 4.02 ;
      RECT 44.005 5.86 44.205 6.06 ;
      RECT 43.985 3.14 44.185 3.34 ;
      RECT 43.325 4.84 43.525 5.04 ;
      RECT 42.955 5.86 43.155 6.06 ;
      RECT 42.645 2.45 42.845 2.65 ;
      RECT 38.15 7.08 38.35 7.28 ;
      RECT 28.1 2.8 28.3 3 ;
      RECT 28.1 3.82 28.3 4.02 ;
      RECT 27.42 5.86 27.62 6.06 ;
      RECT 27.4 3.14 27.6 3.34 ;
      RECT 26.74 4.84 26.94 5.04 ;
      RECT 26.37 5.86 26.57 6.06 ;
      RECT 26.06 2.45 26.26 2.65 ;
      RECT 21.565 7.08 21.765 7.28 ;
      RECT 11.515 2.8 11.715 3 ;
      RECT 11.515 3.82 11.715 4.02 ;
      RECT 10.835 5.86 11.035 6.06 ;
      RECT 10.815 3.14 11.015 3.34 ;
      RECT 10.155 4.84 10.355 5.04 ;
      RECT 9.785 5.86 9.985 6.06 ;
      RECT 9.475 2.45 9.675 2.65 ;
      RECT 4.98 7.08 5.18 7.28 ;
    LAYER met2 ;
      RECT 1.37 8.6 85.51 8.77 ;
      RECT 85.34 7.3 85.51 8.77 ;
      RECT 1.37 6.255 1.54 8.77 ;
      RECT 85.305 7.3 85.63 7.625 ;
      RECT 1.33 6.255 1.61 6.595 ;
      RECT 82.15 6.28 82.47 6.605 ;
      RECT 82.18 5.695 82.35 6.605 ;
      RECT 82.18 5.695 82.355 6.045 ;
      RECT 82.18 5.695 83.155 5.87 ;
      RECT 82.98 1.965 83.155 5.87 ;
      RECT 82.925 1.965 83.275 2.315 ;
      RECT 71.815 8.29 81.995 8.46 ;
      RECT 81.835 2.395 81.995 8.46 ;
      RECT 71.815 6.6 71.985 8.46 ;
      RECT 82.95 6.655 83.275 6.98 ;
      RECT 68.76 6.655 69.085 6.98 ;
      RECT 71.76 6.6 72.04 6.94 ;
      RECT 81.835 6.745 83.275 6.915 ;
      RECT 68.76 6.685 72.04 6.855 ;
      RECT 82.15 2.365 82.47 2.685 ;
      RECT 81.835 2.395 82.47 2.565 ;
      RECT 75.77 2.37 76.05 2.74 ;
      RECT 75.815 1.605 75.985 2.74 ;
      RECT 80.48 1.995 80.805 2.32 ;
      RECT 80.555 1.605 80.725 2.32 ;
      RECT 75.815 1.605 80.725 1.775 ;
      RECT 79.51 4.78 79.77 5.1 ;
      RECT 79.57 2.74 79.71 5.1 ;
      RECT 79.51 2.74 79.77 3.06 ;
      RECT 78.49 5.8 78.75 6.12 ;
      RECT 77.87 5.89 78.75 6.03 ;
      RECT 77.87 3.73 78.01 6.03 ;
      RECT 77.81 3.73 78.09 4.1 ;
      RECT 77.13 5.77 77.41 6.14 ;
      RECT 77.19 3.85 77.33 6.14 ;
      RECT 77.19 3.85 77.67 3.99 ;
      RECT 77.53 2.06 77.67 3.99 ;
      RECT 77.47 2.06 77.73 2.38 ;
      RECT 76.45 4.75 76.73 5.12 ;
      RECT 76.51 2.4 76.65 5.12 ;
      RECT 76.45 2.4 76.71 2.72 ;
      RECT 76.08 5.77 76.36 6.14 ;
      RECT 76.08 5.8 76.37 6.12 ;
      RECT 71.23 6.995 71.6 7.365 ;
      RECT 71.23 6.995 71.605 7.005 ;
      RECT 65.57 6.28 65.89 6.605 ;
      RECT 65.6 5.695 65.77 6.605 ;
      RECT 65.6 5.695 65.775 6.045 ;
      RECT 65.6 5.695 66.575 5.87 ;
      RECT 66.4 1.965 66.575 5.87 ;
      RECT 66.345 1.965 66.695 2.315 ;
      RECT 55.235 8.29 65.415 8.46 ;
      RECT 65.255 2.395 65.415 8.46 ;
      RECT 55.235 6.6 55.405 8.46 ;
      RECT 66.37 6.655 66.695 6.98 ;
      RECT 52.175 6.655 52.5 6.98 ;
      RECT 55.18 6.6 55.46 6.94 ;
      RECT 65.255 6.745 66.695 6.915 ;
      RECT 52.175 6.685 55.46 6.855 ;
      RECT 65.57 2.365 65.89 2.685 ;
      RECT 65.255 2.395 65.89 2.565 ;
      RECT 59.19 2.37 59.47 2.74 ;
      RECT 59.235 1.605 59.405 2.74 ;
      RECT 63.9 1.995 64.225 2.32 ;
      RECT 63.975 1.605 64.145 2.32 ;
      RECT 59.235 1.605 64.145 1.775 ;
      RECT 62.93 4.78 63.19 5.1 ;
      RECT 62.99 2.74 63.13 5.1 ;
      RECT 62.93 2.74 63.19 3.06 ;
      RECT 61.91 5.8 62.17 6.12 ;
      RECT 61.29 5.89 62.17 6.03 ;
      RECT 61.29 3.73 61.43 6.03 ;
      RECT 61.23 3.73 61.51 4.1 ;
      RECT 60.55 5.77 60.83 6.14 ;
      RECT 60.61 3.85 60.75 6.14 ;
      RECT 60.61 3.85 61.09 3.99 ;
      RECT 60.95 2.06 61.09 3.99 ;
      RECT 60.89 2.06 61.15 2.38 ;
      RECT 59.87 4.75 60.15 5.12 ;
      RECT 59.93 2.4 60.07 5.12 ;
      RECT 59.87 2.4 60.13 2.72 ;
      RECT 59.5 5.77 59.78 6.14 ;
      RECT 59.5 5.8 59.79 6.12 ;
      RECT 48.985 6.28 49.305 6.605 ;
      RECT 49.015 5.695 49.185 6.605 ;
      RECT 49.015 5.695 49.19 6.045 ;
      RECT 49.015 5.695 49.99 5.87 ;
      RECT 49.815 1.965 49.99 5.87 ;
      RECT 49.76 1.965 50.11 2.315 ;
      RECT 38.65 8.29 48.83 8.46 ;
      RECT 48.67 2.395 48.83 8.46 ;
      RECT 38.65 6.6 38.82 8.46 ;
      RECT 49.785 6.655 50.11 6.98 ;
      RECT 35.59 6.655 35.915 6.98 ;
      RECT 38.595 6.6 38.875 6.94 ;
      RECT 48.67 6.745 50.11 6.915 ;
      RECT 35.59 6.685 38.875 6.855 ;
      RECT 48.985 2.365 49.305 2.685 ;
      RECT 48.67 2.395 49.305 2.565 ;
      RECT 42.605 2.37 42.885 2.74 ;
      RECT 42.65 1.605 42.82 2.74 ;
      RECT 47.315 1.995 47.64 2.32 ;
      RECT 47.39 1.605 47.56 2.32 ;
      RECT 42.65 1.605 47.56 1.775 ;
      RECT 46.345 4.78 46.605 5.1 ;
      RECT 46.405 2.74 46.545 5.1 ;
      RECT 46.345 2.74 46.605 3.06 ;
      RECT 45.325 5.8 45.585 6.12 ;
      RECT 44.705 5.89 45.585 6.03 ;
      RECT 44.705 3.73 44.845 6.03 ;
      RECT 44.645 3.73 44.925 4.1 ;
      RECT 43.965 5.77 44.245 6.14 ;
      RECT 44.025 3.85 44.165 6.14 ;
      RECT 44.025 3.85 44.505 3.99 ;
      RECT 44.365 2.06 44.505 3.99 ;
      RECT 44.305 2.06 44.565 2.38 ;
      RECT 43.285 4.75 43.565 5.12 ;
      RECT 43.345 2.4 43.485 5.12 ;
      RECT 43.285 2.4 43.545 2.72 ;
      RECT 42.915 5.77 43.195 6.14 ;
      RECT 42.915 5.8 43.205 6.12 ;
      RECT 32.4 6.28 32.72 6.605 ;
      RECT 32.43 5.695 32.6 6.605 ;
      RECT 32.43 5.695 32.605 6.045 ;
      RECT 32.43 5.695 33.405 5.87 ;
      RECT 33.23 1.965 33.405 5.87 ;
      RECT 33.175 1.965 33.525 2.315 ;
      RECT 22.065 8.29 32.245 8.46 ;
      RECT 32.085 2.395 32.245 8.46 ;
      RECT 22.065 6.6 22.235 8.46 ;
      RECT 33.2 6.655 33.525 6.98 ;
      RECT 19.005 6.655 19.33 6.98 ;
      RECT 22.01 6.6 22.29 6.94 ;
      RECT 32.085 6.745 33.525 6.915 ;
      RECT 19.005 6.685 22.29 6.855 ;
      RECT 32.4 2.365 32.72 2.685 ;
      RECT 32.085 2.395 32.72 2.565 ;
      RECT 26.02 2.37 26.3 2.74 ;
      RECT 26.065 1.605 26.235 2.74 ;
      RECT 30.73 1.995 31.055 2.32 ;
      RECT 30.805 1.605 30.975 2.32 ;
      RECT 26.065 1.605 30.975 1.775 ;
      RECT 29.76 4.78 30.02 5.1 ;
      RECT 29.82 2.74 29.96 5.1 ;
      RECT 29.76 2.74 30.02 3.06 ;
      RECT 28.74 5.8 29 6.12 ;
      RECT 28.12 5.89 29 6.03 ;
      RECT 28.12 3.73 28.26 6.03 ;
      RECT 28.06 3.73 28.34 4.1 ;
      RECT 27.38 5.77 27.66 6.14 ;
      RECT 27.44 3.85 27.58 6.14 ;
      RECT 27.44 3.85 27.92 3.99 ;
      RECT 27.78 2.06 27.92 3.99 ;
      RECT 27.72 2.06 27.98 2.38 ;
      RECT 26.7 4.75 26.98 5.12 ;
      RECT 26.76 2.4 26.9 5.12 ;
      RECT 26.7 2.4 26.96 2.72 ;
      RECT 26.33 5.77 26.61 6.14 ;
      RECT 26.33 5.8 26.62 6.12 ;
      RECT 15.815 6.28 16.135 6.605 ;
      RECT 15.845 5.695 16.015 6.605 ;
      RECT 15.845 5.695 16.02 6.045 ;
      RECT 15.845 5.695 16.82 5.87 ;
      RECT 16.645 1.965 16.82 5.87 ;
      RECT 16.59 1.965 16.94 2.315 ;
      RECT 5.48 8.29 15.66 8.46 ;
      RECT 15.5 2.395 15.66 8.46 ;
      RECT 5.48 6.6 5.65 8.46 ;
      RECT 1.715 6.995 1.995 7.335 ;
      RECT 1.715 7.06 2.905 7.23 ;
      RECT 2.735 6.685 2.905 7.23 ;
      RECT 16.615 6.655 16.94 6.98 ;
      RECT 5.425 6.6 5.705 6.94 ;
      RECT 15.5 6.745 16.94 6.915 ;
      RECT 2.735 6.685 5.705 6.855 ;
      RECT 15.815 2.365 16.135 2.685 ;
      RECT 15.5 2.395 16.135 2.565 ;
      RECT 9.435 2.37 9.715 2.74 ;
      RECT 9.48 1.605 9.65 2.74 ;
      RECT 14.145 1.995 14.47 2.32 ;
      RECT 14.22 1.605 14.39 2.32 ;
      RECT 9.48 1.605 14.39 1.775 ;
      RECT 13.175 4.78 13.435 5.1 ;
      RECT 13.235 2.74 13.375 5.1 ;
      RECT 13.175 2.74 13.435 3.06 ;
      RECT 12.155 5.8 12.415 6.12 ;
      RECT 11.535 5.89 12.415 6.03 ;
      RECT 11.535 3.73 11.675 6.03 ;
      RECT 11.475 3.73 11.755 4.1 ;
      RECT 10.795 5.77 11.075 6.14 ;
      RECT 10.855 3.85 10.995 6.14 ;
      RECT 10.855 3.85 11.335 3.99 ;
      RECT 11.195 2.06 11.335 3.99 ;
      RECT 11.135 2.06 11.395 2.38 ;
      RECT 10.115 4.75 10.395 5.12 ;
      RECT 10.175 2.4 10.315 5.12 ;
      RECT 10.115 2.4 10.375 2.72 ;
      RECT 9.745 5.77 10.025 6.14 ;
      RECT 9.745 5.8 10.035 6.12 ;
      RECT 77.81 2.71 78.09 3.08 ;
      RECT 77.11 3.05 77.39 3.42 ;
      RECT 61.23 2.71 61.51 3.08 ;
      RECT 60.53 3.05 60.81 3.42 ;
      RECT 54.65 6.995 55.02 7.365 ;
      RECT 44.645 2.71 44.925 3.08 ;
      RECT 43.945 3.05 44.225 3.42 ;
      RECT 38.065 6.995 38.435 7.365 ;
      RECT 28.06 2.71 28.34 3.08 ;
      RECT 27.36 3.05 27.64 3.42 ;
      RECT 21.48 6.995 21.85 7.365 ;
      RECT 11.475 2.71 11.755 3.08 ;
      RECT 10.775 3.05 11.055 3.42 ;
      RECT 4.895 6.995 5.265 7.365 ;
    LAYER via1 ;
      RECT 85.395 7.385 85.545 7.535 ;
      RECT 83.04 6.74 83.19 6.89 ;
      RECT 83.025 2.065 83.175 2.215 ;
      RECT 82.235 2.45 82.385 2.6 ;
      RECT 82.235 6.37 82.385 6.52 ;
      RECT 80.57 2.08 80.72 2.23 ;
      RECT 79.565 2.825 79.715 2.975 ;
      RECT 79.565 4.865 79.715 5.015 ;
      RECT 78.545 5.885 78.695 6.035 ;
      RECT 77.865 2.825 78.015 2.975 ;
      RECT 77.865 3.845 78.015 3.995 ;
      RECT 77.525 2.145 77.675 2.295 ;
      RECT 77.185 3.165 77.335 3.315 ;
      RECT 77.185 5.885 77.335 6.035 ;
      RECT 76.505 2.485 76.655 2.635 ;
      RECT 76.505 4.865 76.655 5.015 ;
      RECT 76.165 5.885 76.315 6.035 ;
      RECT 75.825 2.475 75.975 2.625 ;
      RECT 71.825 6.695 71.975 6.845 ;
      RECT 71.34 7.105 71.49 7.255 ;
      RECT 68.85 6.74 69 6.89 ;
      RECT 66.46 6.74 66.61 6.89 ;
      RECT 66.445 2.065 66.595 2.215 ;
      RECT 65.655 2.45 65.805 2.6 ;
      RECT 65.655 6.37 65.805 6.52 ;
      RECT 63.99 2.08 64.14 2.23 ;
      RECT 62.985 2.825 63.135 2.975 ;
      RECT 62.985 4.865 63.135 5.015 ;
      RECT 61.965 5.885 62.115 6.035 ;
      RECT 61.285 2.825 61.435 2.975 ;
      RECT 61.285 3.845 61.435 3.995 ;
      RECT 60.945 2.145 61.095 2.295 ;
      RECT 60.605 3.165 60.755 3.315 ;
      RECT 60.605 5.885 60.755 6.035 ;
      RECT 59.925 2.485 60.075 2.635 ;
      RECT 59.925 4.865 60.075 5.015 ;
      RECT 59.585 5.885 59.735 6.035 ;
      RECT 59.245 2.475 59.395 2.625 ;
      RECT 55.245 6.695 55.395 6.845 ;
      RECT 54.76 7.105 54.91 7.255 ;
      RECT 52.265 6.74 52.415 6.89 ;
      RECT 49.875 6.74 50.025 6.89 ;
      RECT 49.86 2.065 50.01 2.215 ;
      RECT 49.07 2.45 49.22 2.6 ;
      RECT 49.07 6.37 49.22 6.52 ;
      RECT 47.405 2.08 47.555 2.23 ;
      RECT 46.4 2.825 46.55 2.975 ;
      RECT 46.4 4.865 46.55 5.015 ;
      RECT 45.38 5.885 45.53 6.035 ;
      RECT 44.7 2.825 44.85 2.975 ;
      RECT 44.7 3.845 44.85 3.995 ;
      RECT 44.36 2.145 44.51 2.295 ;
      RECT 44.02 3.165 44.17 3.315 ;
      RECT 44.02 5.885 44.17 6.035 ;
      RECT 43.34 2.485 43.49 2.635 ;
      RECT 43.34 4.865 43.49 5.015 ;
      RECT 43 5.885 43.15 6.035 ;
      RECT 42.66 2.475 42.81 2.625 ;
      RECT 38.66 6.695 38.81 6.845 ;
      RECT 38.175 7.105 38.325 7.255 ;
      RECT 35.68 6.74 35.83 6.89 ;
      RECT 33.29 6.74 33.44 6.89 ;
      RECT 33.275 2.065 33.425 2.215 ;
      RECT 32.485 2.45 32.635 2.6 ;
      RECT 32.485 6.37 32.635 6.52 ;
      RECT 30.82 2.08 30.97 2.23 ;
      RECT 29.815 2.825 29.965 2.975 ;
      RECT 29.815 4.865 29.965 5.015 ;
      RECT 28.795 5.885 28.945 6.035 ;
      RECT 28.115 2.825 28.265 2.975 ;
      RECT 28.115 3.845 28.265 3.995 ;
      RECT 27.775 2.145 27.925 2.295 ;
      RECT 27.435 3.165 27.585 3.315 ;
      RECT 27.435 5.885 27.585 6.035 ;
      RECT 26.755 2.485 26.905 2.635 ;
      RECT 26.755 4.865 26.905 5.015 ;
      RECT 26.415 5.885 26.565 6.035 ;
      RECT 26.075 2.475 26.225 2.625 ;
      RECT 22.075 6.695 22.225 6.845 ;
      RECT 21.59 7.105 21.74 7.255 ;
      RECT 19.095 6.74 19.245 6.89 ;
      RECT 16.705 6.74 16.855 6.89 ;
      RECT 16.69 2.065 16.84 2.215 ;
      RECT 15.9 2.45 16.05 2.6 ;
      RECT 15.9 6.37 16.05 6.52 ;
      RECT 14.235 2.08 14.385 2.23 ;
      RECT 13.23 2.825 13.38 2.975 ;
      RECT 13.23 4.865 13.38 5.015 ;
      RECT 12.21 5.885 12.36 6.035 ;
      RECT 11.53 2.825 11.68 2.975 ;
      RECT 11.53 3.845 11.68 3.995 ;
      RECT 11.19 2.145 11.34 2.295 ;
      RECT 10.85 3.165 11 3.315 ;
      RECT 10.85 5.885 11 6.035 ;
      RECT 10.17 2.485 10.32 2.635 ;
      RECT 10.17 4.865 10.32 5.015 ;
      RECT 9.83 5.885 9.98 6.035 ;
      RECT 9.49 2.475 9.64 2.625 ;
      RECT 5.49 6.695 5.64 6.845 ;
      RECT 5.005 7.105 5.155 7.255 ;
      RECT 1.78 7.09 1.93 7.24 ;
      RECT 1.395 6.35 1.545 6.5 ;
    LAYER met1 ;
      RECT 85.275 7.77 85.565 8 ;
      RECT 85.335 6.29 85.505 8 ;
      RECT 85.305 7.3 85.63 7.625 ;
      RECT 85.275 6.29 85.565 6.52 ;
      RECT 84.87 2.395 84.975 2.965 ;
      RECT 84.87 2.73 85.195 2.96 ;
      RECT 84.87 2.76 85.365 2.93 ;
      RECT 84.87 2.395 85.06 2.96 ;
      RECT 84.285 2.36 84.575 2.59 ;
      RECT 84.285 2.395 85.06 2.565 ;
      RECT 84.345 0.88 84.515 2.59 ;
      RECT 84.285 0.88 84.575 1.11 ;
      RECT 84.285 7.77 84.575 8 ;
      RECT 84.345 6.29 84.515 8 ;
      RECT 84.285 6.29 84.575 6.52 ;
      RECT 84.285 6.325 85.14 6.485 ;
      RECT 84.97 5.92 85.14 6.485 ;
      RECT 84.285 6.32 84.68 6.485 ;
      RECT 84.905 5.92 85.195 6.15 ;
      RECT 84.905 5.95 85.365 6.12 ;
      RECT 83.915 2.73 84.205 2.96 ;
      RECT 83.915 2.76 84.375 2.93 ;
      RECT 83.98 1.655 84.145 2.96 ;
      RECT 82.495 1.625 82.785 1.855 ;
      RECT 82.495 1.655 84.145 1.825 ;
      RECT 82.555 0.885 82.725 1.855 ;
      RECT 82.495 0.885 82.785 1.115 ;
      RECT 82.495 7.765 82.785 7.995 ;
      RECT 82.555 7.025 82.725 7.995 ;
      RECT 82.555 7.12 84.145 7.29 ;
      RECT 83.975 5.92 84.145 7.29 ;
      RECT 82.495 7.025 82.785 7.255 ;
      RECT 83.915 5.92 84.205 6.15 ;
      RECT 83.915 5.95 84.375 6.12 ;
      RECT 80.48 1.995 80.805 2.32 ;
      RECT 82.925 1.965 83.275 2.315 ;
      RECT 80.48 2.025 83.275 2.195 ;
      RECT 82.95 6.655 83.275 6.98 ;
      RECT 82.925 6.655 83.275 6.885 ;
      RECT 82.755 6.685 83.275 6.855 ;
      RECT 82.15 2.365 82.47 2.685 ;
      RECT 82.12 2.365 82.47 2.595 ;
      RECT 81.835 2.395 82.47 2.565 ;
      RECT 82.15 6.28 82.47 6.605 ;
      RECT 82.12 6.285 82.47 6.515 ;
      RECT 81.95 6.315 82.47 6.485 ;
      RECT 79.48 2.77 79.8 3.03 ;
      RECT 79.2 2.83 79.8 2.97 ;
      RECT 77.1 3.11 77.42 3.37 ;
      RECT 79.07 3.12 79.36 3.35 ;
      RECT 77.1 3.17 79.365 3.31 ;
      RECT 78.46 5.83 78.78 6.09 ;
      RECT 78.46 5.89 79.05 6.03 ;
      RECT 77.78 2.77 78.1 3.03 ;
      RECT 73.04 2.78 73.33 3.01 ;
      RECT 73.04 2.83 78.1 2.97 ;
      RECT 77.87 2.49 78.01 3.03 ;
      RECT 77.87 2.49 78.35 2.63 ;
      RECT 78.21 2.1 78.35 2.63 ;
      RECT 78.13 2.1 78.42 2.33 ;
      RECT 77.78 3.79 78.1 4.05 ;
      RECT 77.11 3.8 77.4 4.03 ;
      RECT 74.9 3.8 75.19 4.03 ;
      RECT 74.9 3.85 78.1 3.99 ;
      RECT 76.08 5.83 76.4 6.09 ;
      RECT 77.79 5.84 78.08 6.07 ;
      RECT 75.41 5.84 75.7 6.07 ;
      RECT 75.41 5.89 76.4 6.03 ;
      RECT 77.87 5.55 78.01 6.07 ;
      RECT 76.17 5.55 76.31 6.09 ;
      RECT 76.17 5.55 78.01 5.69 ;
      RECT 75.07 2.44 75.36 2.67 ;
      RECT 75.15 2.15 75.29 2.67 ;
      RECT 77.44 2.09 77.76 2.35 ;
      RECT 77.34 2.1 77.76 2.33 ;
      RECT 75.15 2.15 77.76 2.29 ;
      RECT 76.42 2.43 76.74 2.69 ;
      RECT 76.42 2.49 77.01 2.63 ;
      RECT 76.42 4.81 76.74 5.07 ;
      RECT 73.71 4.82 74 5.05 ;
      RECT 73.71 4.87 76.74 5.01 ;
      RECT 75.74 2.39 76.07 2.72 ;
      RECT 75.74 2.44 76.2 2.67 ;
      RECT 75.74 2.49 76.22 2.63 ;
      RECT 75.62 2.49 75.63 2.63 ;
      RECT 75.63 2.48 76.2 2.62 ;
      RECT 71.73 6.63 72.07 6.91 ;
      RECT 71.7 6.655 72.07 6.885 ;
      RECT 71.53 6.685 72.07 6.855 ;
      RECT 71.27 7.765 71.56 7.995 ;
      RECT 71.33 6.995 71.5 7.995 ;
      RECT 71.23 6.995 71.6 7.365 ;
      RECT 68.695 7.77 68.985 8 ;
      RECT 68.755 6.29 68.925 8 ;
      RECT 68.755 6.655 69.085 6.98 ;
      RECT 68.695 6.29 68.985 6.52 ;
      RECT 68.29 2.395 68.395 2.965 ;
      RECT 68.29 2.73 68.615 2.96 ;
      RECT 68.29 2.76 68.785 2.93 ;
      RECT 68.29 2.395 68.48 2.96 ;
      RECT 67.705 2.36 67.995 2.59 ;
      RECT 67.705 2.395 68.48 2.565 ;
      RECT 67.765 0.88 67.935 2.59 ;
      RECT 67.705 0.88 67.995 1.11 ;
      RECT 67.705 7.77 67.995 8 ;
      RECT 67.765 6.29 67.935 8 ;
      RECT 67.705 6.29 67.995 6.52 ;
      RECT 67.705 6.325 68.56 6.485 ;
      RECT 68.39 5.92 68.56 6.485 ;
      RECT 67.705 6.32 68.1 6.485 ;
      RECT 68.325 5.92 68.615 6.15 ;
      RECT 68.325 5.95 68.785 6.12 ;
      RECT 67.335 2.73 67.625 2.96 ;
      RECT 67.335 2.76 67.795 2.93 ;
      RECT 67.4 1.655 67.565 2.96 ;
      RECT 65.915 1.625 66.205 1.855 ;
      RECT 65.915 1.655 67.565 1.825 ;
      RECT 65.975 0.885 66.145 1.855 ;
      RECT 65.915 0.885 66.205 1.115 ;
      RECT 65.915 7.765 66.205 7.995 ;
      RECT 65.975 7.025 66.145 7.995 ;
      RECT 65.975 7.12 67.565 7.29 ;
      RECT 67.395 5.92 67.565 7.29 ;
      RECT 65.915 7.025 66.205 7.255 ;
      RECT 67.335 5.92 67.625 6.15 ;
      RECT 67.335 5.95 67.795 6.12 ;
      RECT 63.9 1.995 64.225 2.32 ;
      RECT 66.345 1.965 66.695 2.315 ;
      RECT 63.9 2.025 66.695 2.195 ;
      RECT 66.37 6.655 66.695 6.98 ;
      RECT 66.345 6.655 66.695 6.885 ;
      RECT 66.175 6.685 66.695 6.855 ;
      RECT 65.57 2.365 65.89 2.685 ;
      RECT 65.54 2.365 65.89 2.595 ;
      RECT 65.255 2.395 65.89 2.565 ;
      RECT 65.57 6.28 65.89 6.605 ;
      RECT 65.54 6.285 65.89 6.515 ;
      RECT 65.37 6.315 65.89 6.485 ;
      RECT 62.9 2.77 63.22 3.03 ;
      RECT 62.62 2.83 63.22 2.97 ;
      RECT 60.52 3.11 60.84 3.37 ;
      RECT 62.49 3.12 62.78 3.35 ;
      RECT 60.52 3.17 62.785 3.31 ;
      RECT 61.88 5.83 62.2 6.09 ;
      RECT 61.88 5.89 62.47 6.03 ;
      RECT 61.2 2.77 61.52 3.03 ;
      RECT 56.46 2.78 56.75 3.01 ;
      RECT 56.46 2.83 61.52 2.97 ;
      RECT 61.29 2.49 61.43 3.03 ;
      RECT 61.29 2.49 61.77 2.63 ;
      RECT 61.63 2.1 61.77 2.63 ;
      RECT 61.55 2.1 61.84 2.33 ;
      RECT 61.2 3.79 61.52 4.05 ;
      RECT 60.53 3.8 60.82 4.03 ;
      RECT 58.32 3.8 58.61 4.03 ;
      RECT 58.32 3.85 61.52 3.99 ;
      RECT 59.5 5.83 59.82 6.09 ;
      RECT 61.21 5.84 61.5 6.07 ;
      RECT 58.83 5.84 59.12 6.07 ;
      RECT 58.83 5.89 59.82 6.03 ;
      RECT 61.29 5.55 61.43 6.07 ;
      RECT 59.59 5.55 59.73 6.09 ;
      RECT 59.59 5.55 61.43 5.69 ;
      RECT 58.49 2.44 58.78 2.67 ;
      RECT 58.57 2.15 58.71 2.67 ;
      RECT 60.86 2.09 61.18 2.35 ;
      RECT 60.76 2.1 61.18 2.33 ;
      RECT 58.57 2.15 61.18 2.29 ;
      RECT 59.84 2.43 60.16 2.69 ;
      RECT 59.84 2.49 60.43 2.63 ;
      RECT 59.84 4.81 60.16 5.07 ;
      RECT 57.13 4.82 57.42 5.05 ;
      RECT 57.13 4.87 60.16 5.01 ;
      RECT 59.16 2.39 59.49 2.72 ;
      RECT 59.16 2.44 59.62 2.67 ;
      RECT 59.16 2.49 59.64 2.63 ;
      RECT 59.04 2.49 59.05 2.63 ;
      RECT 59.05 2.48 59.62 2.62 ;
      RECT 55.15 6.63 55.49 6.91 ;
      RECT 55.12 6.655 55.49 6.885 ;
      RECT 54.95 6.685 55.49 6.855 ;
      RECT 54.69 7.765 54.98 7.995 ;
      RECT 54.75 6.995 54.92 7.995 ;
      RECT 54.65 6.995 55.02 7.365 ;
      RECT 52.11 7.77 52.4 8 ;
      RECT 52.17 6.29 52.34 8 ;
      RECT 52.17 6.655 52.5 6.98 ;
      RECT 52.11 6.29 52.4 6.52 ;
      RECT 51.705 2.395 51.81 2.965 ;
      RECT 51.705 2.73 52.03 2.96 ;
      RECT 51.705 2.76 52.2 2.93 ;
      RECT 51.705 2.395 51.895 2.96 ;
      RECT 51.12 2.36 51.41 2.59 ;
      RECT 51.12 2.395 51.895 2.565 ;
      RECT 51.18 0.88 51.35 2.59 ;
      RECT 51.12 0.88 51.41 1.11 ;
      RECT 51.12 7.77 51.41 8 ;
      RECT 51.18 6.29 51.35 8 ;
      RECT 51.12 6.29 51.41 6.52 ;
      RECT 51.12 6.325 51.975 6.485 ;
      RECT 51.805 5.92 51.975 6.485 ;
      RECT 51.12 6.32 51.515 6.485 ;
      RECT 51.74 5.92 52.03 6.15 ;
      RECT 51.74 5.95 52.2 6.12 ;
      RECT 50.75 2.73 51.04 2.96 ;
      RECT 50.75 2.76 51.21 2.93 ;
      RECT 50.815 1.655 50.98 2.96 ;
      RECT 49.33 1.625 49.62 1.855 ;
      RECT 49.33 1.655 50.98 1.825 ;
      RECT 49.39 0.885 49.56 1.855 ;
      RECT 49.33 0.885 49.62 1.115 ;
      RECT 49.33 7.765 49.62 7.995 ;
      RECT 49.39 7.025 49.56 7.995 ;
      RECT 49.39 7.12 50.98 7.29 ;
      RECT 50.81 5.92 50.98 7.29 ;
      RECT 49.33 7.025 49.62 7.255 ;
      RECT 50.75 5.92 51.04 6.15 ;
      RECT 50.75 5.95 51.21 6.12 ;
      RECT 47.315 1.995 47.64 2.32 ;
      RECT 49.76 1.965 50.11 2.315 ;
      RECT 47.315 2.025 50.11 2.195 ;
      RECT 49.785 6.655 50.11 6.98 ;
      RECT 49.76 6.655 50.11 6.885 ;
      RECT 49.59 6.685 50.11 6.855 ;
      RECT 48.985 2.365 49.305 2.685 ;
      RECT 48.955 2.365 49.305 2.595 ;
      RECT 48.67 2.395 49.305 2.565 ;
      RECT 48.985 6.28 49.305 6.605 ;
      RECT 48.955 6.285 49.305 6.515 ;
      RECT 48.785 6.315 49.305 6.485 ;
      RECT 46.315 2.77 46.635 3.03 ;
      RECT 46.035 2.83 46.635 2.97 ;
      RECT 43.935 3.11 44.255 3.37 ;
      RECT 45.905 3.12 46.195 3.35 ;
      RECT 43.935 3.17 46.2 3.31 ;
      RECT 45.295 5.83 45.615 6.09 ;
      RECT 45.295 5.89 45.885 6.03 ;
      RECT 44.615 2.77 44.935 3.03 ;
      RECT 39.875 2.78 40.165 3.01 ;
      RECT 39.875 2.83 44.935 2.97 ;
      RECT 44.705 2.49 44.845 3.03 ;
      RECT 44.705 2.49 45.185 2.63 ;
      RECT 45.045 2.1 45.185 2.63 ;
      RECT 44.965 2.1 45.255 2.33 ;
      RECT 44.615 3.79 44.935 4.05 ;
      RECT 43.945 3.8 44.235 4.03 ;
      RECT 41.735 3.8 42.025 4.03 ;
      RECT 41.735 3.85 44.935 3.99 ;
      RECT 42.915 5.83 43.235 6.09 ;
      RECT 44.625 5.84 44.915 6.07 ;
      RECT 42.245 5.84 42.535 6.07 ;
      RECT 42.245 5.89 43.235 6.03 ;
      RECT 44.705 5.55 44.845 6.07 ;
      RECT 43.005 5.55 43.145 6.09 ;
      RECT 43.005 5.55 44.845 5.69 ;
      RECT 41.905 2.44 42.195 2.67 ;
      RECT 41.985 2.15 42.125 2.67 ;
      RECT 44.275 2.09 44.595 2.35 ;
      RECT 44.175 2.1 44.595 2.33 ;
      RECT 41.985 2.15 44.595 2.29 ;
      RECT 43.255 2.43 43.575 2.69 ;
      RECT 43.255 2.49 43.845 2.63 ;
      RECT 43.255 4.81 43.575 5.07 ;
      RECT 40.545 4.82 40.835 5.05 ;
      RECT 40.545 4.87 43.575 5.01 ;
      RECT 42.575 2.39 42.905 2.72 ;
      RECT 42.575 2.44 43.035 2.67 ;
      RECT 42.575 2.49 43.055 2.63 ;
      RECT 42.455 2.49 42.465 2.63 ;
      RECT 42.465 2.48 43.035 2.62 ;
      RECT 38.565 6.63 38.905 6.91 ;
      RECT 38.535 6.655 38.905 6.885 ;
      RECT 38.365 6.685 38.905 6.855 ;
      RECT 38.105 7.765 38.395 7.995 ;
      RECT 38.165 6.995 38.335 7.995 ;
      RECT 38.065 6.995 38.435 7.365 ;
      RECT 35.525 7.77 35.815 8 ;
      RECT 35.585 6.29 35.755 8 ;
      RECT 35.585 6.655 35.915 6.98 ;
      RECT 35.525 6.29 35.815 6.52 ;
      RECT 35.12 2.395 35.225 2.965 ;
      RECT 35.12 2.73 35.445 2.96 ;
      RECT 35.12 2.76 35.615 2.93 ;
      RECT 35.12 2.395 35.31 2.96 ;
      RECT 34.535 2.36 34.825 2.59 ;
      RECT 34.535 2.395 35.31 2.565 ;
      RECT 34.595 0.88 34.765 2.59 ;
      RECT 34.535 0.88 34.825 1.11 ;
      RECT 34.535 7.77 34.825 8 ;
      RECT 34.595 6.29 34.765 8 ;
      RECT 34.535 6.29 34.825 6.52 ;
      RECT 34.535 6.325 35.39 6.485 ;
      RECT 35.22 5.92 35.39 6.485 ;
      RECT 34.535 6.32 34.93 6.485 ;
      RECT 35.155 5.92 35.445 6.15 ;
      RECT 35.155 5.95 35.615 6.12 ;
      RECT 34.165 2.73 34.455 2.96 ;
      RECT 34.165 2.76 34.625 2.93 ;
      RECT 34.23 1.655 34.395 2.96 ;
      RECT 32.745 1.625 33.035 1.855 ;
      RECT 32.745 1.655 34.395 1.825 ;
      RECT 32.805 0.885 32.975 1.855 ;
      RECT 32.745 0.885 33.035 1.115 ;
      RECT 32.745 7.765 33.035 7.995 ;
      RECT 32.805 7.025 32.975 7.995 ;
      RECT 32.805 7.12 34.395 7.29 ;
      RECT 34.225 5.92 34.395 7.29 ;
      RECT 32.745 7.025 33.035 7.255 ;
      RECT 34.165 5.92 34.455 6.15 ;
      RECT 34.165 5.95 34.625 6.12 ;
      RECT 30.73 1.995 31.055 2.32 ;
      RECT 33.175 1.965 33.525 2.315 ;
      RECT 30.73 2.025 33.525 2.195 ;
      RECT 33.2 6.655 33.525 6.98 ;
      RECT 33.175 6.655 33.525 6.885 ;
      RECT 33.005 6.685 33.525 6.855 ;
      RECT 32.4 2.365 32.72 2.685 ;
      RECT 32.37 2.365 32.72 2.595 ;
      RECT 32.085 2.395 32.72 2.565 ;
      RECT 32.4 6.28 32.72 6.605 ;
      RECT 32.37 6.285 32.72 6.515 ;
      RECT 32.2 6.315 32.72 6.485 ;
      RECT 29.73 2.77 30.05 3.03 ;
      RECT 29.45 2.83 30.05 2.97 ;
      RECT 27.35 3.11 27.67 3.37 ;
      RECT 29.32 3.12 29.61 3.35 ;
      RECT 27.35 3.17 29.615 3.31 ;
      RECT 28.71 5.83 29.03 6.09 ;
      RECT 28.71 5.89 29.3 6.03 ;
      RECT 28.03 2.77 28.35 3.03 ;
      RECT 23.29 2.78 23.58 3.01 ;
      RECT 23.29 2.83 28.35 2.97 ;
      RECT 28.12 2.49 28.26 3.03 ;
      RECT 28.12 2.49 28.6 2.63 ;
      RECT 28.46 2.1 28.6 2.63 ;
      RECT 28.38 2.1 28.67 2.33 ;
      RECT 28.03 3.79 28.35 4.05 ;
      RECT 27.36 3.8 27.65 4.03 ;
      RECT 25.15 3.8 25.44 4.03 ;
      RECT 25.15 3.85 28.35 3.99 ;
      RECT 26.33 5.83 26.65 6.09 ;
      RECT 28.04 5.84 28.33 6.07 ;
      RECT 25.66 5.84 25.95 6.07 ;
      RECT 25.66 5.89 26.65 6.03 ;
      RECT 28.12 5.55 28.26 6.07 ;
      RECT 26.42 5.55 26.56 6.09 ;
      RECT 26.42 5.55 28.26 5.69 ;
      RECT 25.32 2.44 25.61 2.67 ;
      RECT 25.4 2.15 25.54 2.67 ;
      RECT 27.69 2.09 28.01 2.35 ;
      RECT 27.59 2.1 28.01 2.33 ;
      RECT 25.4 2.15 28.01 2.29 ;
      RECT 26.67 2.43 26.99 2.69 ;
      RECT 26.67 2.49 27.26 2.63 ;
      RECT 26.67 4.81 26.99 5.07 ;
      RECT 23.96 4.82 24.25 5.05 ;
      RECT 23.96 4.87 26.99 5.01 ;
      RECT 25.99 2.39 26.32 2.72 ;
      RECT 25.99 2.44 26.45 2.67 ;
      RECT 25.99 2.49 26.47 2.63 ;
      RECT 25.87 2.49 25.88 2.63 ;
      RECT 25.88 2.48 26.45 2.62 ;
      RECT 21.98 6.63 22.32 6.91 ;
      RECT 21.95 6.655 22.32 6.885 ;
      RECT 21.78 6.685 22.32 6.855 ;
      RECT 21.52 7.765 21.81 7.995 ;
      RECT 21.58 6.995 21.75 7.995 ;
      RECT 21.48 6.995 21.85 7.365 ;
      RECT 18.94 7.77 19.23 8 ;
      RECT 19 6.29 19.17 8 ;
      RECT 19 6.655 19.33 6.98 ;
      RECT 18.94 6.29 19.23 6.52 ;
      RECT 18.535 2.395 18.64 2.965 ;
      RECT 18.535 2.73 18.86 2.96 ;
      RECT 18.535 2.76 19.03 2.93 ;
      RECT 18.535 2.395 18.725 2.96 ;
      RECT 17.95 2.36 18.24 2.59 ;
      RECT 17.95 2.395 18.725 2.565 ;
      RECT 18.01 0.88 18.18 2.59 ;
      RECT 17.95 0.88 18.24 1.11 ;
      RECT 17.95 7.77 18.24 8 ;
      RECT 18.01 6.29 18.18 8 ;
      RECT 17.95 6.29 18.24 6.52 ;
      RECT 17.95 6.325 18.805 6.485 ;
      RECT 18.635 5.92 18.805 6.485 ;
      RECT 17.95 6.32 18.345 6.485 ;
      RECT 18.57 5.92 18.86 6.15 ;
      RECT 18.57 5.95 19.03 6.12 ;
      RECT 17.58 2.73 17.87 2.96 ;
      RECT 17.58 2.76 18.04 2.93 ;
      RECT 17.645 1.655 17.81 2.96 ;
      RECT 16.16 1.625 16.45 1.855 ;
      RECT 16.16 1.655 17.81 1.825 ;
      RECT 16.22 0.885 16.39 1.855 ;
      RECT 16.16 0.885 16.45 1.115 ;
      RECT 16.16 7.765 16.45 7.995 ;
      RECT 16.22 7.025 16.39 7.995 ;
      RECT 16.22 7.12 17.81 7.29 ;
      RECT 17.64 5.92 17.81 7.29 ;
      RECT 16.16 7.025 16.45 7.255 ;
      RECT 17.58 5.92 17.87 6.15 ;
      RECT 17.58 5.95 18.04 6.12 ;
      RECT 14.145 1.995 14.47 2.32 ;
      RECT 16.59 1.965 16.94 2.315 ;
      RECT 14.145 2.025 16.94 2.195 ;
      RECT 16.615 6.655 16.94 6.98 ;
      RECT 16.59 6.655 16.94 6.885 ;
      RECT 16.42 6.685 16.94 6.855 ;
      RECT 15.815 2.365 16.135 2.685 ;
      RECT 15.785 2.365 16.135 2.595 ;
      RECT 15.5 2.395 16.135 2.565 ;
      RECT 15.815 6.28 16.135 6.605 ;
      RECT 15.785 6.285 16.135 6.515 ;
      RECT 15.615 6.315 16.135 6.485 ;
      RECT 13.145 2.77 13.465 3.03 ;
      RECT 12.865 2.83 13.465 2.97 ;
      RECT 10.765 3.11 11.085 3.37 ;
      RECT 12.735 3.12 13.025 3.35 ;
      RECT 10.765 3.17 13.03 3.31 ;
      RECT 12.125 5.83 12.445 6.09 ;
      RECT 12.125 5.89 12.715 6.03 ;
      RECT 11.445 2.77 11.765 3.03 ;
      RECT 6.705 2.78 6.995 3.01 ;
      RECT 6.705 2.83 11.765 2.97 ;
      RECT 11.535 2.49 11.675 3.03 ;
      RECT 11.535 2.49 12.015 2.63 ;
      RECT 11.875 2.1 12.015 2.63 ;
      RECT 11.795 2.1 12.085 2.33 ;
      RECT 11.445 3.79 11.765 4.05 ;
      RECT 10.775 3.8 11.065 4.03 ;
      RECT 8.565 3.8 8.855 4.03 ;
      RECT 8.565 3.85 11.765 3.99 ;
      RECT 9.745 5.83 10.065 6.09 ;
      RECT 11.455 5.84 11.745 6.07 ;
      RECT 9.075 5.84 9.365 6.07 ;
      RECT 9.075 5.89 10.065 6.03 ;
      RECT 11.535 5.55 11.675 6.07 ;
      RECT 9.835 5.55 9.975 6.09 ;
      RECT 9.835 5.55 11.675 5.69 ;
      RECT 8.735 2.44 9.025 2.67 ;
      RECT 8.815 2.15 8.955 2.67 ;
      RECT 11.105 2.09 11.425 2.35 ;
      RECT 11.005 2.1 11.425 2.33 ;
      RECT 8.815 2.15 11.425 2.29 ;
      RECT 10.085 2.43 10.405 2.69 ;
      RECT 10.085 2.49 10.675 2.63 ;
      RECT 10.085 4.81 10.405 5.07 ;
      RECT 7.375 4.82 7.665 5.05 ;
      RECT 7.375 4.87 10.405 5.01 ;
      RECT 9.405 2.39 9.735 2.72 ;
      RECT 9.405 2.44 9.865 2.67 ;
      RECT 9.405 2.49 9.885 2.63 ;
      RECT 9.285 2.49 9.295 2.63 ;
      RECT 9.295 2.48 9.865 2.62 ;
      RECT 5.395 6.63 5.735 6.91 ;
      RECT 5.365 6.655 5.735 6.885 ;
      RECT 5.195 6.685 5.735 6.855 ;
      RECT 4.935 7.765 5.225 7.995 ;
      RECT 4.995 6.995 5.165 7.995 ;
      RECT 4.895 6.995 5.265 7.365 ;
      RECT 1.705 7.765 1.995 7.995 ;
      RECT 1.765 7.025 1.935 7.995 ;
      RECT 1.685 7.025 2.025 7.305 ;
      RECT 1.3 6.285 1.64 6.565 ;
      RECT 1.16 6.315 1.64 6.485 ;
      RECT 79.15 4.81 79.8 5.07 ;
      RECT 77.1 5.83 77.42 6.09 ;
      RECT 62.57 4.81 63.22 5.07 ;
      RECT 60.52 5.83 60.84 6.09 ;
      RECT 45.985 4.81 46.635 5.07 ;
      RECT 43.935 5.83 44.255 6.09 ;
      RECT 29.4 4.81 30.05 5.07 ;
      RECT 27.35 5.83 27.67 6.09 ;
      RECT 12.815 4.81 13.465 5.07 ;
      RECT 10.765 5.83 11.085 6.09 ;
    LAYER mcon ;
      RECT 85.335 6.32 85.505 6.49 ;
      RECT 85.34 6.315 85.51 6.485 ;
      RECT 68.755 6.32 68.925 6.49 ;
      RECT 68.76 6.315 68.93 6.485 ;
      RECT 52.17 6.32 52.34 6.49 ;
      RECT 52.175 6.315 52.345 6.485 ;
      RECT 35.585 6.32 35.755 6.49 ;
      RECT 35.59 6.315 35.76 6.485 ;
      RECT 19 6.32 19.17 6.49 ;
      RECT 19.005 6.315 19.175 6.485 ;
      RECT 85.335 7.8 85.505 7.97 ;
      RECT 84.965 2.76 85.135 2.93 ;
      RECT 84.965 5.95 85.135 6.12 ;
      RECT 84.345 0.91 84.515 1.08 ;
      RECT 84.345 2.39 84.515 2.56 ;
      RECT 84.345 6.32 84.515 6.49 ;
      RECT 84.345 7.8 84.515 7.97 ;
      RECT 83.975 2.76 84.145 2.93 ;
      RECT 83.975 5.95 84.145 6.12 ;
      RECT 82.985 2.025 83.155 2.195 ;
      RECT 82.985 6.685 83.155 6.855 ;
      RECT 82.555 0.915 82.725 1.085 ;
      RECT 82.555 1.655 82.725 1.825 ;
      RECT 82.555 7.055 82.725 7.225 ;
      RECT 82.555 7.795 82.725 7.965 ;
      RECT 82.18 2.395 82.35 2.565 ;
      RECT 82.18 6.315 82.35 6.485 ;
      RECT 79.55 2.81 79.72 2.98 ;
      RECT 79.21 4.85 79.38 5.02 ;
      RECT 79.13 3.15 79.3 3.32 ;
      RECT 78.53 5.87 78.7 6.04 ;
      RECT 78.19 2.13 78.36 2.3 ;
      RECT 77.85 5.87 78.02 6.04 ;
      RECT 77.4 2.13 77.57 2.3 ;
      RECT 77.17 3.83 77.34 4 ;
      RECT 77.17 5.87 77.34 6.04 ;
      RECT 76.49 2.47 76.66 2.64 ;
      RECT 75.97 2.47 76.14 2.64 ;
      RECT 75.47 5.87 75.64 6.04 ;
      RECT 75.13 2.47 75.3 2.64 ;
      RECT 74.96 3.83 75.13 4 ;
      RECT 73.77 4.85 73.94 5.02 ;
      RECT 73.1 2.81 73.27 2.98 ;
      RECT 71.76 6.685 71.93 6.855 ;
      RECT 71.33 7.055 71.5 7.225 ;
      RECT 71.33 7.795 71.5 7.965 ;
      RECT 68.755 7.8 68.925 7.97 ;
      RECT 68.385 2.76 68.555 2.93 ;
      RECT 68.385 5.95 68.555 6.12 ;
      RECT 67.765 0.91 67.935 1.08 ;
      RECT 67.765 2.39 67.935 2.56 ;
      RECT 67.765 6.32 67.935 6.49 ;
      RECT 67.765 7.8 67.935 7.97 ;
      RECT 67.395 2.76 67.565 2.93 ;
      RECT 67.395 5.95 67.565 6.12 ;
      RECT 66.405 2.025 66.575 2.195 ;
      RECT 66.405 6.685 66.575 6.855 ;
      RECT 65.975 0.915 66.145 1.085 ;
      RECT 65.975 1.655 66.145 1.825 ;
      RECT 65.975 7.055 66.145 7.225 ;
      RECT 65.975 7.795 66.145 7.965 ;
      RECT 65.6 2.395 65.77 2.565 ;
      RECT 65.6 6.315 65.77 6.485 ;
      RECT 62.97 2.81 63.14 2.98 ;
      RECT 62.63 4.85 62.8 5.02 ;
      RECT 62.55 3.15 62.72 3.32 ;
      RECT 61.95 5.87 62.12 6.04 ;
      RECT 61.61 2.13 61.78 2.3 ;
      RECT 61.27 5.87 61.44 6.04 ;
      RECT 60.82 2.13 60.99 2.3 ;
      RECT 60.59 3.83 60.76 4 ;
      RECT 60.59 5.87 60.76 6.04 ;
      RECT 59.91 2.47 60.08 2.64 ;
      RECT 59.39 2.47 59.56 2.64 ;
      RECT 58.89 5.87 59.06 6.04 ;
      RECT 58.55 2.47 58.72 2.64 ;
      RECT 58.38 3.83 58.55 4 ;
      RECT 57.19 4.85 57.36 5.02 ;
      RECT 56.52 2.81 56.69 2.98 ;
      RECT 55.18 6.685 55.35 6.855 ;
      RECT 54.75 7.055 54.92 7.225 ;
      RECT 54.75 7.795 54.92 7.965 ;
      RECT 52.17 7.8 52.34 7.97 ;
      RECT 51.8 2.76 51.97 2.93 ;
      RECT 51.8 5.95 51.97 6.12 ;
      RECT 51.18 0.91 51.35 1.08 ;
      RECT 51.18 2.39 51.35 2.56 ;
      RECT 51.18 6.32 51.35 6.49 ;
      RECT 51.18 7.8 51.35 7.97 ;
      RECT 50.81 2.76 50.98 2.93 ;
      RECT 50.81 5.95 50.98 6.12 ;
      RECT 49.82 2.025 49.99 2.195 ;
      RECT 49.82 6.685 49.99 6.855 ;
      RECT 49.39 0.915 49.56 1.085 ;
      RECT 49.39 1.655 49.56 1.825 ;
      RECT 49.39 7.055 49.56 7.225 ;
      RECT 49.39 7.795 49.56 7.965 ;
      RECT 49.015 2.395 49.185 2.565 ;
      RECT 49.015 6.315 49.185 6.485 ;
      RECT 46.385 2.81 46.555 2.98 ;
      RECT 46.045 4.85 46.215 5.02 ;
      RECT 45.965 3.15 46.135 3.32 ;
      RECT 45.365 5.87 45.535 6.04 ;
      RECT 45.025 2.13 45.195 2.3 ;
      RECT 44.685 5.87 44.855 6.04 ;
      RECT 44.235 2.13 44.405 2.3 ;
      RECT 44.005 3.83 44.175 4 ;
      RECT 44.005 5.87 44.175 6.04 ;
      RECT 43.325 2.47 43.495 2.64 ;
      RECT 42.805 2.47 42.975 2.64 ;
      RECT 42.305 5.87 42.475 6.04 ;
      RECT 41.965 2.47 42.135 2.64 ;
      RECT 41.795 3.83 41.965 4 ;
      RECT 40.605 4.85 40.775 5.02 ;
      RECT 39.935 2.81 40.105 2.98 ;
      RECT 38.595 6.685 38.765 6.855 ;
      RECT 38.165 7.055 38.335 7.225 ;
      RECT 38.165 7.795 38.335 7.965 ;
      RECT 35.585 7.8 35.755 7.97 ;
      RECT 35.215 2.76 35.385 2.93 ;
      RECT 35.215 5.95 35.385 6.12 ;
      RECT 34.595 0.91 34.765 1.08 ;
      RECT 34.595 2.39 34.765 2.56 ;
      RECT 34.595 6.32 34.765 6.49 ;
      RECT 34.595 7.8 34.765 7.97 ;
      RECT 34.225 2.76 34.395 2.93 ;
      RECT 34.225 5.95 34.395 6.12 ;
      RECT 33.235 2.025 33.405 2.195 ;
      RECT 33.235 6.685 33.405 6.855 ;
      RECT 32.805 0.915 32.975 1.085 ;
      RECT 32.805 1.655 32.975 1.825 ;
      RECT 32.805 7.055 32.975 7.225 ;
      RECT 32.805 7.795 32.975 7.965 ;
      RECT 32.43 2.395 32.6 2.565 ;
      RECT 32.43 6.315 32.6 6.485 ;
      RECT 29.8 2.81 29.97 2.98 ;
      RECT 29.46 4.85 29.63 5.02 ;
      RECT 29.38 3.15 29.55 3.32 ;
      RECT 28.78 5.87 28.95 6.04 ;
      RECT 28.44 2.13 28.61 2.3 ;
      RECT 28.1 5.87 28.27 6.04 ;
      RECT 27.65 2.13 27.82 2.3 ;
      RECT 27.42 3.83 27.59 4 ;
      RECT 27.42 5.87 27.59 6.04 ;
      RECT 26.74 2.47 26.91 2.64 ;
      RECT 26.22 2.47 26.39 2.64 ;
      RECT 25.72 5.87 25.89 6.04 ;
      RECT 25.38 2.47 25.55 2.64 ;
      RECT 25.21 3.83 25.38 4 ;
      RECT 24.02 4.85 24.19 5.02 ;
      RECT 23.35 2.81 23.52 2.98 ;
      RECT 22.01 6.685 22.18 6.855 ;
      RECT 21.58 7.055 21.75 7.225 ;
      RECT 21.58 7.795 21.75 7.965 ;
      RECT 19 7.8 19.17 7.97 ;
      RECT 18.63 2.76 18.8 2.93 ;
      RECT 18.63 5.95 18.8 6.12 ;
      RECT 18.01 0.91 18.18 1.08 ;
      RECT 18.01 2.39 18.18 2.56 ;
      RECT 18.01 6.32 18.18 6.49 ;
      RECT 18.01 7.8 18.18 7.97 ;
      RECT 17.64 2.76 17.81 2.93 ;
      RECT 17.64 5.95 17.81 6.12 ;
      RECT 16.65 2.025 16.82 2.195 ;
      RECT 16.65 6.685 16.82 6.855 ;
      RECT 16.22 0.915 16.39 1.085 ;
      RECT 16.22 1.655 16.39 1.825 ;
      RECT 16.22 7.055 16.39 7.225 ;
      RECT 16.22 7.795 16.39 7.965 ;
      RECT 15.845 2.395 16.015 2.565 ;
      RECT 15.845 6.315 16.015 6.485 ;
      RECT 13.215 2.81 13.385 2.98 ;
      RECT 12.875 4.85 13.045 5.02 ;
      RECT 12.795 3.15 12.965 3.32 ;
      RECT 12.195 5.87 12.365 6.04 ;
      RECT 11.855 2.13 12.025 2.3 ;
      RECT 11.515 5.87 11.685 6.04 ;
      RECT 11.065 2.13 11.235 2.3 ;
      RECT 10.835 3.83 11.005 4 ;
      RECT 10.835 5.87 11.005 6.04 ;
      RECT 10.155 2.47 10.325 2.64 ;
      RECT 9.635 2.47 9.805 2.64 ;
      RECT 9.135 5.87 9.305 6.04 ;
      RECT 8.795 2.47 8.965 2.64 ;
      RECT 8.625 3.83 8.795 4 ;
      RECT 7.435 4.85 7.605 5.02 ;
      RECT 6.765 2.81 6.935 2.98 ;
      RECT 5.425 6.685 5.595 6.855 ;
      RECT 4.995 7.055 5.165 7.225 ;
      RECT 4.995 7.795 5.165 7.965 ;
      RECT 1.765 7.055 1.935 7.225 ;
      RECT 1.765 7.795 1.935 7.965 ;
      RECT 1.39 6.315 1.56 6.485 ;
    LAYER li1 ;
      RECT 85.335 5.02 85.505 6.49 ;
      RECT 85.335 6.315 85.51 6.485 ;
      RECT 84.965 1.74 85.135 2.93 ;
      RECT 84.965 1.74 85.435 1.91 ;
      RECT 84.965 6.97 85.435 7.14 ;
      RECT 84.965 5.95 85.135 7.14 ;
      RECT 83.975 1.74 84.145 2.93 ;
      RECT 83.975 1.74 84.445 1.91 ;
      RECT 83.975 6.97 84.445 7.14 ;
      RECT 83.975 5.95 84.145 7.14 ;
      RECT 82.125 2.635 82.295 3.865 ;
      RECT 82.18 0.855 82.35 2.805 ;
      RECT 82.125 0.575 82.295 1.025 ;
      RECT 82.125 7.855 82.295 8.305 ;
      RECT 82.18 6.075 82.35 8.025 ;
      RECT 82.125 5.015 82.295 6.245 ;
      RECT 81.605 0.575 81.775 3.865 ;
      RECT 81.605 2.075 82.01 2.405 ;
      RECT 81.605 1.235 82.01 1.565 ;
      RECT 81.605 5.015 81.775 8.305 ;
      RECT 81.605 7.315 82.01 7.645 ;
      RECT 81.605 6.475 82.01 6.805 ;
      RECT 76.86 6.64 78.17 6.89 ;
      RECT 76.86 6.32 77.04 6.89 ;
      RECT 76.31 6.32 77.04 6.49 ;
      RECT 76.31 5.48 76.48 6.49 ;
      RECT 77.15 5.52 78.89 5.7 ;
      RECT 78.56 4.68 78.89 5.7 ;
      RECT 76.31 5.48 77.37 5.65 ;
      RECT 78.56 4.85 79.38 5.02 ;
      RECT 77.72 4.68 78.05 4.89 ;
      RECT 77.72 4.68 78.89 4.85 ;
      RECT 78.62 3.2 78.95 4.16 ;
      RECT 78.62 3.2 79.3 3.37 ;
      RECT 79.13 1.96 79.3 3.37 ;
      RECT 79.04 1.96 79.37 2.6 ;
      RECT 78.17 3.47 78.44 4.17 ;
      RECT 78.27 1.96 78.44 4.17 ;
      RECT 78.61 2.78 78.96 3.03 ;
      RECT 78.27 2.81 78.96 2.98 ;
      RECT 78.18 1.96 78.44 2.44 ;
      RECT 77.51 5.11 78.39 5.35 ;
      RECT 78.16 5.02 78.39 5.35 ;
      RECT 76.86 5.11 78.39 5.31 ;
      RECT 77.78 5.06 78.39 5.35 ;
      RECT 76.86 4.98 77.03 5.31 ;
      RECT 77.75 5.87 78 6.47 ;
      RECT 77.75 5.87 78.22 6.07 ;
      RECT 77.24 3.09 78 3.59 ;
      RECT 76.31 2.9 76.57 3.52 ;
      RECT 77.23 3.03 77.24 3.34 ;
      RECT 77.21 3.02 77.23 3.31 ;
      RECT 77.87 2.7 78.1 3.3 ;
      RECT 77.19 2.97 77.21 3.28 ;
      RECT 77.17 3.09 78.1 3.27 ;
      RECT 77.14 3.09 78.1 3.26 ;
      RECT 77.07 3.09 78.1 3.25 ;
      RECT 77.05 3.09 78.1 3.22 ;
      RECT 77.03 2 77.2 3.19 ;
      RECT 77 3.09 78.1 3.16 ;
      RECT 76.97 3.09 78.1 3.13 ;
      RECT 76.94 3.08 77.3 3.1 ;
      RECT 76.94 3.07 77.29 3.1 ;
      RECT 76.31 2.9 77.2 3.07 ;
      RECT 76.31 3.06 77.27 3.07 ;
      RECT 76.31 3.05 77.26 3.07 ;
      RECT 76.31 2.99 77.22 3.07 ;
      RECT 76.31 2 77.2 2.17 ;
      RECT 77.37 2.5 77.7 2.92 ;
      RECT 77.37 2.01 77.59 2.92 ;
      RECT 77.29 5.87 77.5 6.47 ;
      RECT 77.15 5.87 77.5 6.07 ;
      RECT 75.87 3.47 76.14 4.17 ;
      RECT 76.09 1.96 76.14 4.17 ;
      RECT 75.97 2.77 76.14 4.17 ;
      RECT 75.97 1.96 76.14 2.76 ;
      RECT 75.88 1.96 76.14 2.44 ;
      RECT 74.01 3.13 74.26 3.67 ;
      RECT 74.98 3.13 75.7 3.6 ;
      RECT 74.01 3.13 75.8 3.3 ;
      RECT 75.57 2.77 75.8 3.3 ;
      RECT 74.57 2.01 74.82 3.3 ;
      RECT 75.57 2.7 75.63 3.6 ;
      RECT 75.57 2.7 75.8 2.76 ;
      RECT 74.03 2.01 74.82 2.28 ;
      RECT 74.99 5.82 75.67 6.07 ;
      RECT 75.4 5.46 75.67 6.07 ;
      RECT 75.15 6.24 75.48 6.79 ;
      RECT 74.09 6.24 75.48 6.43 ;
      RECT 74.09 5.4 74.26 6.43 ;
      RECT 73.97 5.82 74.26 6.15 ;
      RECT 74.09 5.4 75.03 5.57 ;
      RECT 74.73 4.85 75.03 5.57 ;
      RECT 74.99 2.43 75.4 2.95 ;
      RECT 74.99 2.01 75.19 2.95 ;
      RECT 73.6 2.19 73.77 4.17 ;
      RECT 73.6 2.7 74.4 2.95 ;
      RECT 73.6 2.19 73.85 2.95 ;
      RECT 73.52 2.19 73.85 2.61 ;
      RECT 73.55 6.6 74.11 6.89 ;
      RECT 73.55 4.68 73.8 6.89 ;
      RECT 73.55 4.68 74.01 5.23 ;
      RECT 70.38 5.015 70.55 8.305 ;
      RECT 70.38 7.315 70.785 7.645 ;
      RECT 70.38 6.475 70.785 6.805 ;
      RECT 68.755 5.02 68.925 6.49 ;
      RECT 68.755 6.315 68.93 6.485 ;
      RECT 68.385 1.74 68.555 2.93 ;
      RECT 68.385 1.74 68.855 1.91 ;
      RECT 68.385 6.97 68.855 7.14 ;
      RECT 68.385 5.95 68.555 7.14 ;
      RECT 67.395 1.74 67.565 2.93 ;
      RECT 67.395 1.74 67.865 1.91 ;
      RECT 67.395 6.97 67.865 7.14 ;
      RECT 67.395 5.95 67.565 7.14 ;
      RECT 65.545 2.635 65.715 3.865 ;
      RECT 65.6 0.855 65.77 2.805 ;
      RECT 65.545 0.575 65.715 1.025 ;
      RECT 65.545 7.855 65.715 8.305 ;
      RECT 65.6 6.075 65.77 8.025 ;
      RECT 65.545 5.015 65.715 6.245 ;
      RECT 65.025 0.575 65.195 3.865 ;
      RECT 65.025 2.075 65.43 2.405 ;
      RECT 65.025 1.235 65.43 1.565 ;
      RECT 65.025 5.015 65.195 8.305 ;
      RECT 65.025 7.315 65.43 7.645 ;
      RECT 65.025 6.475 65.43 6.805 ;
      RECT 60.28 6.64 61.59 6.89 ;
      RECT 60.28 6.32 60.46 6.89 ;
      RECT 59.73 6.32 60.46 6.49 ;
      RECT 59.73 5.48 59.9 6.49 ;
      RECT 60.57 5.52 62.31 5.7 ;
      RECT 61.98 4.68 62.31 5.7 ;
      RECT 59.73 5.48 60.79 5.65 ;
      RECT 61.98 4.85 62.8 5.02 ;
      RECT 61.14 4.68 61.47 4.89 ;
      RECT 61.14 4.68 62.31 4.85 ;
      RECT 62.04 3.2 62.37 4.16 ;
      RECT 62.04 3.2 62.72 3.37 ;
      RECT 62.55 1.96 62.72 3.37 ;
      RECT 62.46 1.96 62.79 2.6 ;
      RECT 61.59 3.47 61.86 4.17 ;
      RECT 61.69 1.96 61.86 4.17 ;
      RECT 62.03 2.78 62.38 3.03 ;
      RECT 61.69 2.81 62.38 2.98 ;
      RECT 61.6 1.96 61.86 2.44 ;
      RECT 60.93 5.11 61.81 5.35 ;
      RECT 61.58 5.02 61.81 5.35 ;
      RECT 60.28 5.11 61.81 5.31 ;
      RECT 61.2 5.06 61.81 5.35 ;
      RECT 60.28 4.98 60.45 5.31 ;
      RECT 61.17 5.87 61.42 6.47 ;
      RECT 61.17 5.87 61.64 6.07 ;
      RECT 60.66 3.09 61.42 3.59 ;
      RECT 59.73 2.9 59.99 3.52 ;
      RECT 60.65 3.03 60.66 3.34 ;
      RECT 60.63 3.02 60.65 3.31 ;
      RECT 61.29 2.7 61.52 3.3 ;
      RECT 60.61 2.97 60.63 3.28 ;
      RECT 60.59 3.09 61.52 3.27 ;
      RECT 60.56 3.09 61.52 3.26 ;
      RECT 60.49 3.09 61.52 3.25 ;
      RECT 60.47 3.09 61.52 3.22 ;
      RECT 60.45 2 60.62 3.19 ;
      RECT 60.42 3.09 61.52 3.16 ;
      RECT 60.39 3.09 61.52 3.13 ;
      RECT 60.36 3.08 60.72 3.1 ;
      RECT 60.36 3.07 60.71 3.1 ;
      RECT 59.73 2.9 60.62 3.07 ;
      RECT 59.73 3.06 60.69 3.07 ;
      RECT 59.73 3.05 60.68 3.07 ;
      RECT 59.73 2.99 60.64 3.07 ;
      RECT 59.73 2 60.62 2.17 ;
      RECT 60.79 2.5 61.12 2.92 ;
      RECT 60.79 2.01 61.01 2.92 ;
      RECT 60.71 5.87 60.92 6.47 ;
      RECT 60.57 5.87 60.92 6.07 ;
      RECT 59.29 3.47 59.56 4.17 ;
      RECT 59.51 1.96 59.56 4.17 ;
      RECT 59.39 2.77 59.56 4.17 ;
      RECT 59.39 1.96 59.56 2.76 ;
      RECT 59.3 1.96 59.56 2.44 ;
      RECT 57.43 3.13 57.68 3.67 ;
      RECT 58.4 3.13 59.12 3.6 ;
      RECT 57.43 3.13 59.22 3.3 ;
      RECT 58.99 2.77 59.22 3.3 ;
      RECT 57.99 2.01 58.24 3.3 ;
      RECT 58.99 2.7 59.05 3.6 ;
      RECT 58.99 2.7 59.22 2.76 ;
      RECT 57.45 2.01 58.24 2.28 ;
      RECT 58.41 5.82 59.09 6.07 ;
      RECT 58.82 5.46 59.09 6.07 ;
      RECT 58.57 6.24 58.9 6.79 ;
      RECT 57.51 6.24 58.9 6.43 ;
      RECT 57.51 5.4 57.68 6.43 ;
      RECT 57.39 5.82 57.68 6.15 ;
      RECT 57.51 5.4 58.45 5.57 ;
      RECT 58.15 4.85 58.45 5.57 ;
      RECT 58.41 2.43 58.82 2.95 ;
      RECT 58.41 2.01 58.61 2.95 ;
      RECT 57.02 2.19 57.19 4.17 ;
      RECT 57.02 2.7 57.82 2.95 ;
      RECT 57.02 2.19 57.27 2.95 ;
      RECT 56.94 2.19 57.27 2.61 ;
      RECT 56.97 6.6 57.53 6.89 ;
      RECT 56.97 4.68 57.22 6.89 ;
      RECT 56.97 4.68 57.43 5.23 ;
      RECT 53.8 5.015 53.97 8.305 ;
      RECT 53.8 7.315 54.205 7.645 ;
      RECT 53.8 6.475 54.205 6.805 ;
      RECT 52.17 5.02 52.34 6.49 ;
      RECT 52.17 6.315 52.345 6.485 ;
      RECT 51.8 1.74 51.97 2.93 ;
      RECT 51.8 1.74 52.27 1.91 ;
      RECT 51.8 6.97 52.27 7.14 ;
      RECT 51.8 5.95 51.97 7.14 ;
      RECT 50.81 1.74 50.98 2.93 ;
      RECT 50.81 1.74 51.28 1.91 ;
      RECT 50.81 6.97 51.28 7.14 ;
      RECT 50.81 5.95 50.98 7.14 ;
      RECT 48.96 2.635 49.13 3.865 ;
      RECT 49.015 0.855 49.185 2.805 ;
      RECT 48.96 0.575 49.13 1.025 ;
      RECT 48.96 7.855 49.13 8.305 ;
      RECT 49.015 6.075 49.185 8.025 ;
      RECT 48.96 5.015 49.13 6.245 ;
      RECT 48.44 0.575 48.61 3.865 ;
      RECT 48.44 2.075 48.845 2.405 ;
      RECT 48.44 1.235 48.845 1.565 ;
      RECT 48.44 5.015 48.61 8.305 ;
      RECT 48.44 7.315 48.845 7.645 ;
      RECT 48.44 6.475 48.845 6.805 ;
      RECT 43.695 6.64 45.005 6.89 ;
      RECT 43.695 6.32 43.875 6.89 ;
      RECT 43.145 6.32 43.875 6.49 ;
      RECT 43.145 5.48 43.315 6.49 ;
      RECT 43.985 5.52 45.725 5.7 ;
      RECT 45.395 4.68 45.725 5.7 ;
      RECT 43.145 5.48 44.205 5.65 ;
      RECT 45.395 4.85 46.215 5.02 ;
      RECT 44.555 4.68 44.885 4.89 ;
      RECT 44.555 4.68 45.725 4.85 ;
      RECT 45.455 3.2 45.785 4.16 ;
      RECT 45.455 3.2 46.135 3.37 ;
      RECT 45.965 1.96 46.135 3.37 ;
      RECT 45.875 1.96 46.205 2.6 ;
      RECT 45.005 3.47 45.275 4.17 ;
      RECT 45.105 1.96 45.275 4.17 ;
      RECT 45.445 2.78 45.795 3.03 ;
      RECT 45.105 2.81 45.795 2.98 ;
      RECT 45.015 1.96 45.275 2.44 ;
      RECT 44.345 5.11 45.225 5.35 ;
      RECT 44.995 5.02 45.225 5.35 ;
      RECT 43.695 5.11 45.225 5.31 ;
      RECT 44.615 5.06 45.225 5.35 ;
      RECT 43.695 4.98 43.865 5.31 ;
      RECT 44.585 5.87 44.835 6.47 ;
      RECT 44.585 5.87 45.055 6.07 ;
      RECT 44.075 3.09 44.835 3.59 ;
      RECT 43.145 2.9 43.405 3.52 ;
      RECT 44.065 3.03 44.075 3.34 ;
      RECT 44.045 3.02 44.065 3.31 ;
      RECT 44.705 2.7 44.935 3.3 ;
      RECT 44.025 2.97 44.045 3.28 ;
      RECT 44.005 3.09 44.935 3.27 ;
      RECT 43.975 3.09 44.935 3.26 ;
      RECT 43.905 3.09 44.935 3.25 ;
      RECT 43.885 3.09 44.935 3.22 ;
      RECT 43.865 2 44.035 3.19 ;
      RECT 43.835 3.09 44.935 3.16 ;
      RECT 43.805 3.09 44.935 3.13 ;
      RECT 43.775 3.08 44.135 3.1 ;
      RECT 43.775 3.07 44.125 3.1 ;
      RECT 43.145 2.9 44.035 3.07 ;
      RECT 43.145 3.06 44.105 3.07 ;
      RECT 43.145 3.05 44.095 3.07 ;
      RECT 43.145 2.99 44.055 3.07 ;
      RECT 43.145 2 44.035 2.17 ;
      RECT 44.205 2.5 44.535 2.92 ;
      RECT 44.205 2.01 44.425 2.92 ;
      RECT 44.125 5.87 44.335 6.47 ;
      RECT 43.985 5.87 44.335 6.07 ;
      RECT 42.705 3.47 42.975 4.17 ;
      RECT 42.925 1.96 42.975 4.17 ;
      RECT 42.805 2.77 42.975 4.17 ;
      RECT 42.805 1.96 42.975 2.76 ;
      RECT 42.715 1.96 42.975 2.44 ;
      RECT 40.845 3.13 41.095 3.67 ;
      RECT 41.815 3.13 42.535 3.6 ;
      RECT 40.845 3.13 42.635 3.3 ;
      RECT 42.405 2.77 42.635 3.3 ;
      RECT 41.405 2.01 41.655 3.3 ;
      RECT 42.405 2.7 42.465 3.6 ;
      RECT 42.405 2.7 42.635 2.76 ;
      RECT 40.865 2.01 41.655 2.28 ;
      RECT 41.825 5.82 42.505 6.07 ;
      RECT 42.235 5.46 42.505 6.07 ;
      RECT 41.985 6.24 42.315 6.79 ;
      RECT 40.925 6.24 42.315 6.43 ;
      RECT 40.925 5.4 41.095 6.43 ;
      RECT 40.805 5.82 41.095 6.15 ;
      RECT 40.925 5.4 41.865 5.57 ;
      RECT 41.565 4.85 41.865 5.57 ;
      RECT 41.825 2.43 42.235 2.95 ;
      RECT 41.825 2.01 42.025 2.95 ;
      RECT 40.435 2.19 40.605 4.17 ;
      RECT 40.435 2.7 41.235 2.95 ;
      RECT 40.435 2.19 40.685 2.95 ;
      RECT 40.355 2.19 40.685 2.61 ;
      RECT 40.385 6.6 40.945 6.89 ;
      RECT 40.385 4.68 40.635 6.89 ;
      RECT 40.385 4.68 40.845 5.23 ;
      RECT 37.215 5.015 37.385 8.305 ;
      RECT 37.215 7.315 37.62 7.645 ;
      RECT 37.215 6.475 37.62 6.805 ;
      RECT 35.585 5.02 35.755 6.49 ;
      RECT 35.585 6.315 35.76 6.485 ;
      RECT 35.215 1.74 35.385 2.93 ;
      RECT 35.215 1.74 35.685 1.91 ;
      RECT 35.215 6.97 35.685 7.14 ;
      RECT 35.215 5.95 35.385 7.14 ;
      RECT 34.225 1.74 34.395 2.93 ;
      RECT 34.225 1.74 34.695 1.91 ;
      RECT 34.225 6.97 34.695 7.14 ;
      RECT 34.225 5.95 34.395 7.14 ;
      RECT 32.375 2.635 32.545 3.865 ;
      RECT 32.43 0.855 32.6 2.805 ;
      RECT 32.375 0.575 32.545 1.025 ;
      RECT 32.375 7.855 32.545 8.305 ;
      RECT 32.43 6.075 32.6 8.025 ;
      RECT 32.375 5.015 32.545 6.245 ;
      RECT 31.855 0.575 32.025 3.865 ;
      RECT 31.855 2.075 32.26 2.405 ;
      RECT 31.855 1.235 32.26 1.565 ;
      RECT 31.855 5.015 32.025 8.305 ;
      RECT 31.855 7.315 32.26 7.645 ;
      RECT 31.855 6.475 32.26 6.805 ;
      RECT 27.11 6.64 28.42 6.89 ;
      RECT 27.11 6.32 27.29 6.89 ;
      RECT 26.56 6.32 27.29 6.49 ;
      RECT 26.56 5.48 26.73 6.49 ;
      RECT 27.4 5.52 29.14 5.7 ;
      RECT 28.81 4.68 29.14 5.7 ;
      RECT 26.56 5.48 27.62 5.65 ;
      RECT 28.81 4.85 29.63 5.02 ;
      RECT 27.97 4.68 28.3 4.89 ;
      RECT 27.97 4.68 29.14 4.85 ;
      RECT 28.87 3.2 29.2 4.16 ;
      RECT 28.87 3.2 29.55 3.37 ;
      RECT 29.38 1.96 29.55 3.37 ;
      RECT 29.29 1.96 29.62 2.6 ;
      RECT 28.42 3.47 28.69 4.17 ;
      RECT 28.52 1.96 28.69 4.17 ;
      RECT 28.86 2.78 29.21 3.03 ;
      RECT 28.52 2.81 29.21 2.98 ;
      RECT 28.43 1.96 28.69 2.44 ;
      RECT 27.76 5.11 28.64 5.35 ;
      RECT 28.41 5.02 28.64 5.35 ;
      RECT 27.11 5.11 28.64 5.31 ;
      RECT 28.03 5.06 28.64 5.35 ;
      RECT 27.11 4.98 27.28 5.31 ;
      RECT 28 5.87 28.25 6.47 ;
      RECT 28 5.87 28.47 6.07 ;
      RECT 27.49 3.09 28.25 3.59 ;
      RECT 26.56 2.9 26.82 3.52 ;
      RECT 27.48 3.03 27.49 3.34 ;
      RECT 27.46 3.02 27.48 3.31 ;
      RECT 28.12 2.7 28.35 3.3 ;
      RECT 27.44 2.97 27.46 3.28 ;
      RECT 27.42 3.09 28.35 3.27 ;
      RECT 27.39 3.09 28.35 3.26 ;
      RECT 27.32 3.09 28.35 3.25 ;
      RECT 27.3 3.09 28.35 3.22 ;
      RECT 27.28 2 27.45 3.19 ;
      RECT 27.25 3.09 28.35 3.16 ;
      RECT 27.22 3.09 28.35 3.13 ;
      RECT 27.19 3.08 27.55 3.1 ;
      RECT 27.19 3.07 27.54 3.1 ;
      RECT 26.56 2.9 27.45 3.07 ;
      RECT 26.56 3.06 27.52 3.07 ;
      RECT 26.56 3.05 27.51 3.07 ;
      RECT 26.56 2.99 27.47 3.07 ;
      RECT 26.56 2 27.45 2.17 ;
      RECT 27.62 2.5 27.95 2.92 ;
      RECT 27.62 2.01 27.84 2.92 ;
      RECT 27.54 5.87 27.75 6.47 ;
      RECT 27.4 5.87 27.75 6.07 ;
      RECT 26.12 3.47 26.39 4.17 ;
      RECT 26.34 1.96 26.39 4.17 ;
      RECT 26.22 2.77 26.39 4.17 ;
      RECT 26.22 1.96 26.39 2.76 ;
      RECT 26.13 1.96 26.39 2.44 ;
      RECT 24.26 3.13 24.51 3.67 ;
      RECT 25.23 3.13 25.95 3.6 ;
      RECT 24.26 3.13 26.05 3.3 ;
      RECT 25.82 2.77 26.05 3.3 ;
      RECT 24.82 2.01 25.07 3.3 ;
      RECT 25.82 2.7 25.88 3.6 ;
      RECT 25.82 2.7 26.05 2.76 ;
      RECT 24.28 2.01 25.07 2.28 ;
      RECT 25.24 5.82 25.92 6.07 ;
      RECT 25.65 5.46 25.92 6.07 ;
      RECT 25.4 6.24 25.73 6.79 ;
      RECT 24.34 6.24 25.73 6.43 ;
      RECT 24.34 5.4 24.51 6.43 ;
      RECT 24.22 5.82 24.51 6.15 ;
      RECT 24.34 5.4 25.28 5.57 ;
      RECT 24.98 4.85 25.28 5.57 ;
      RECT 25.24 2.43 25.65 2.95 ;
      RECT 25.24 2.01 25.44 2.95 ;
      RECT 23.85 2.19 24.02 4.17 ;
      RECT 23.85 2.7 24.65 2.95 ;
      RECT 23.85 2.19 24.1 2.95 ;
      RECT 23.77 2.19 24.1 2.61 ;
      RECT 23.8 6.6 24.36 6.89 ;
      RECT 23.8 4.68 24.05 6.89 ;
      RECT 23.8 4.68 24.26 5.23 ;
      RECT 20.63 5.015 20.8 8.305 ;
      RECT 20.63 7.315 21.035 7.645 ;
      RECT 20.63 6.475 21.035 6.805 ;
      RECT 19 5.02 19.17 6.49 ;
      RECT 19 6.315 19.175 6.485 ;
      RECT 18.63 1.74 18.8 2.93 ;
      RECT 18.63 1.74 19.1 1.91 ;
      RECT 18.63 6.97 19.1 7.14 ;
      RECT 18.63 5.95 18.8 7.14 ;
      RECT 17.64 1.74 17.81 2.93 ;
      RECT 17.64 1.74 18.11 1.91 ;
      RECT 17.64 6.97 18.11 7.14 ;
      RECT 17.64 5.95 17.81 7.14 ;
      RECT 15.79 2.635 15.96 3.865 ;
      RECT 15.845 0.855 16.015 2.805 ;
      RECT 15.79 0.575 15.96 1.025 ;
      RECT 15.79 7.855 15.96 8.305 ;
      RECT 15.845 6.075 16.015 8.025 ;
      RECT 15.79 5.015 15.96 6.245 ;
      RECT 15.27 0.575 15.44 3.865 ;
      RECT 15.27 2.075 15.675 2.405 ;
      RECT 15.27 1.235 15.675 1.565 ;
      RECT 15.27 5.015 15.44 8.305 ;
      RECT 15.27 7.315 15.675 7.645 ;
      RECT 15.27 6.475 15.675 6.805 ;
      RECT 10.525 6.64 11.835 6.89 ;
      RECT 10.525 6.32 10.705 6.89 ;
      RECT 9.975 6.32 10.705 6.49 ;
      RECT 9.975 5.48 10.145 6.49 ;
      RECT 10.815 5.52 12.555 5.7 ;
      RECT 12.225 4.68 12.555 5.7 ;
      RECT 9.975 5.48 11.035 5.65 ;
      RECT 12.225 4.85 13.045 5.02 ;
      RECT 11.385 4.68 11.715 4.89 ;
      RECT 11.385 4.68 12.555 4.85 ;
      RECT 12.285 3.2 12.615 4.16 ;
      RECT 12.285 3.2 12.965 3.37 ;
      RECT 12.795 1.96 12.965 3.37 ;
      RECT 12.705 1.96 13.035 2.6 ;
      RECT 11.835 3.47 12.105 4.17 ;
      RECT 11.935 1.96 12.105 4.17 ;
      RECT 12.275 2.78 12.625 3.03 ;
      RECT 11.935 2.81 12.625 2.98 ;
      RECT 11.845 1.96 12.105 2.44 ;
      RECT 11.175 5.11 12.055 5.35 ;
      RECT 11.825 5.02 12.055 5.35 ;
      RECT 10.525 5.11 12.055 5.31 ;
      RECT 11.445 5.06 12.055 5.35 ;
      RECT 10.525 4.98 10.695 5.31 ;
      RECT 11.415 5.87 11.665 6.47 ;
      RECT 11.415 5.87 11.885 6.07 ;
      RECT 10.905 3.09 11.665 3.59 ;
      RECT 9.975 2.9 10.235 3.52 ;
      RECT 10.895 3.03 10.905 3.34 ;
      RECT 10.875 3.02 10.895 3.31 ;
      RECT 11.535 2.7 11.765 3.3 ;
      RECT 10.855 2.97 10.875 3.28 ;
      RECT 10.835 3.09 11.765 3.27 ;
      RECT 10.805 3.09 11.765 3.26 ;
      RECT 10.735 3.09 11.765 3.25 ;
      RECT 10.715 3.09 11.765 3.22 ;
      RECT 10.695 2 10.865 3.19 ;
      RECT 10.665 3.09 11.765 3.16 ;
      RECT 10.635 3.09 11.765 3.13 ;
      RECT 10.605 3.08 10.965 3.1 ;
      RECT 10.605 3.07 10.955 3.1 ;
      RECT 9.975 2.9 10.865 3.07 ;
      RECT 9.975 3.06 10.935 3.07 ;
      RECT 9.975 3.05 10.925 3.07 ;
      RECT 9.975 2.99 10.885 3.07 ;
      RECT 9.975 2 10.865 2.17 ;
      RECT 11.035 2.5 11.365 2.92 ;
      RECT 11.035 2.01 11.255 2.92 ;
      RECT 10.955 5.87 11.165 6.47 ;
      RECT 10.815 5.87 11.165 6.07 ;
      RECT 9.535 3.47 9.805 4.17 ;
      RECT 9.755 1.96 9.805 4.17 ;
      RECT 9.635 2.77 9.805 4.17 ;
      RECT 9.635 1.96 9.805 2.76 ;
      RECT 9.545 1.96 9.805 2.44 ;
      RECT 7.675 3.13 7.925 3.67 ;
      RECT 8.645 3.13 9.365 3.6 ;
      RECT 7.675 3.13 9.465 3.3 ;
      RECT 9.235 2.77 9.465 3.3 ;
      RECT 8.235 2.01 8.485 3.3 ;
      RECT 9.235 2.7 9.295 3.6 ;
      RECT 9.235 2.7 9.465 2.76 ;
      RECT 7.695 2.01 8.485 2.28 ;
      RECT 8.655 5.82 9.335 6.07 ;
      RECT 9.065 5.46 9.335 6.07 ;
      RECT 8.815 6.24 9.145 6.79 ;
      RECT 7.755 6.24 9.145 6.43 ;
      RECT 7.755 5.4 7.925 6.43 ;
      RECT 7.635 5.82 7.925 6.15 ;
      RECT 7.755 5.4 8.695 5.57 ;
      RECT 8.395 4.85 8.695 5.57 ;
      RECT 8.655 2.43 9.065 2.95 ;
      RECT 8.655 2.01 8.855 2.95 ;
      RECT 7.265 2.19 7.435 4.17 ;
      RECT 7.265 2.7 8.065 2.95 ;
      RECT 7.265 2.19 7.515 2.95 ;
      RECT 7.185 2.19 7.515 2.61 ;
      RECT 7.215 6.6 7.775 6.89 ;
      RECT 7.215 4.68 7.465 6.89 ;
      RECT 7.215 4.68 7.675 5.23 ;
      RECT 4.045 5.015 4.215 8.305 ;
      RECT 4.045 7.315 4.45 7.645 ;
      RECT 4.045 6.475 4.45 6.805 ;
      RECT 1.335 7.855 1.505 8.305 ;
      RECT 1.39 6.075 1.56 8.025 ;
      RECT 1.335 5.015 1.505 6.245 ;
      RECT 0.815 5.015 0.985 8.305 ;
      RECT 0.815 7.315 1.22 7.645 ;
      RECT 0.815 6.475 1.22 6.805 ;
      RECT 85.335 7.8 85.505 8.31 ;
      RECT 84.345 0.57 84.515 1.08 ;
      RECT 84.345 2.39 84.515 3.86 ;
      RECT 84.345 5.02 84.515 6.49 ;
      RECT 84.345 7.8 84.515 8.31 ;
      RECT 82.985 0.575 83.155 3.865 ;
      RECT 82.985 5.015 83.155 8.305 ;
      RECT 82.555 0.575 82.725 1.085 ;
      RECT 82.555 1.655 82.725 3.865 ;
      RECT 82.555 5.015 82.725 7.225 ;
      RECT 82.555 7.795 82.725 8.305 ;
      RECT 79.47 2.78 79.82 3.03 ;
      RECT 78.41 5.87 78.86 6.38 ;
      RECT 77.09 3.83 77.57 4.17 ;
      RECT 76.31 2.34 76.86 2.73 ;
      RECT 74.8 3.83 75.27 4.17 ;
      RECT 73.09 2.78 73.43 3.66 ;
      RECT 71.76 5.015 71.93 8.305 ;
      RECT 71.33 5.015 71.5 7.225 ;
      RECT 71.33 7.795 71.5 8.305 ;
      RECT 68.755 7.8 68.925 8.31 ;
      RECT 67.765 0.57 67.935 1.08 ;
      RECT 67.765 2.39 67.935 3.86 ;
      RECT 67.765 5.02 67.935 6.49 ;
      RECT 67.765 7.8 67.935 8.31 ;
      RECT 66.405 0.575 66.575 3.865 ;
      RECT 66.405 5.015 66.575 8.305 ;
      RECT 65.975 0.575 66.145 1.085 ;
      RECT 65.975 1.655 66.145 3.865 ;
      RECT 65.975 5.015 66.145 7.225 ;
      RECT 65.975 7.795 66.145 8.305 ;
      RECT 62.89 2.78 63.24 3.03 ;
      RECT 61.83 5.87 62.28 6.38 ;
      RECT 60.51 3.83 60.99 4.17 ;
      RECT 59.73 2.34 60.28 2.73 ;
      RECT 58.22 3.83 58.69 4.17 ;
      RECT 56.51 2.78 56.85 3.66 ;
      RECT 55.18 5.015 55.35 8.305 ;
      RECT 54.75 5.015 54.92 7.225 ;
      RECT 54.75 7.795 54.92 8.305 ;
      RECT 52.17 7.8 52.34 8.31 ;
      RECT 51.18 0.57 51.35 1.08 ;
      RECT 51.18 2.39 51.35 3.86 ;
      RECT 51.18 5.02 51.35 6.49 ;
      RECT 51.18 7.8 51.35 8.31 ;
      RECT 49.82 0.575 49.99 3.865 ;
      RECT 49.82 5.015 49.99 8.305 ;
      RECT 49.39 0.575 49.56 1.085 ;
      RECT 49.39 1.655 49.56 3.865 ;
      RECT 49.39 5.015 49.56 7.225 ;
      RECT 49.39 7.795 49.56 8.305 ;
      RECT 46.305 2.78 46.655 3.03 ;
      RECT 45.245 5.87 45.695 6.38 ;
      RECT 43.925 3.83 44.405 4.17 ;
      RECT 43.145 2.34 43.695 2.73 ;
      RECT 41.635 3.83 42.105 4.17 ;
      RECT 39.925 2.78 40.265 3.66 ;
      RECT 38.595 5.015 38.765 8.305 ;
      RECT 38.165 5.015 38.335 7.225 ;
      RECT 38.165 7.795 38.335 8.305 ;
      RECT 35.585 7.8 35.755 8.31 ;
      RECT 34.595 0.57 34.765 1.08 ;
      RECT 34.595 2.39 34.765 3.86 ;
      RECT 34.595 5.02 34.765 6.49 ;
      RECT 34.595 7.8 34.765 8.31 ;
      RECT 33.235 0.575 33.405 3.865 ;
      RECT 33.235 5.015 33.405 8.305 ;
      RECT 32.805 0.575 32.975 1.085 ;
      RECT 32.805 1.655 32.975 3.865 ;
      RECT 32.805 5.015 32.975 7.225 ;
      RECT 32.805 7.795 32.975 8.305 ;
      RECT 29.72 2.78 30.07 3.03 ;
      RECT 28.66 5.87 29.11 6.38 ;
      RECT 27.34 3.83 27.82 4.17 ;
      RECT 26.56 2.34 27.11 2.73 ;
      RECT 25.05 3.83 25.52 4.17 ;
      RECT 23.34 2.78 23.68 3.66 ;
      RECT 22.01 5.015 22.18 8.305 ;
      RECT 21.58 5.015 21.75 7.225 ;
      RECT 21.58 7.795 21.75 8.305 ;
      RECT 19 7.8 19.17 8.31 ;
      RECT 18.01 0.57 18.18 1.08 ;
      RECT 18.01 2.39 18.18 3.86 ;
      RECT 18.01 5.02 18.18 6.49 ;
      RECT 18.01 7.8 18.18 8.31 ;
      RECT 16.65 0.575 16.82 3.865 ;
      RECT 16.65 5.015 16.82 8.305 ;
      RECT 16.22 0.575 16.39 1.085 ;
      RECT 16.22 1.655 16.39 3.865 ;
      RECT 16.22 5.015 16.39 7.225 ;
      RECT 16.22 7.795 16.39 8.305 ;
      RECT 13.135 2.78 13.485 3.03 ;
      RECT 12.075 5.87 12.525 6.38 ;
      RECT 10.755 3.83 11.235 4.17 ;
      RECT 9.975 2.34 10.525 2.73 ;
      RECT 8.465 3.83 8.935 4.17 ;
      RECT 6.755 2.78 7.095 3.66 ;
      RECT 5.425 5.015 5.595 8.305 ;
      RECT 4.995 5.015 5.165 7.225 ;
      RECT 4.995 7.795 5.165 8.305 ;
      RECT 1.765 5.015 1.935 7.225 ;
      RECT 1.765 7.795 1.935 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r1 ;
  SIZE 88.91 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 19.49 0.915 19.66 1.085 ;
        RECT 19.485 0.91 19.655 1.08 ;
        RECT 19.485 2.39 19.655 2.56 ;
      LAYER li1 ;
        RECT 19.49 0.915 19.66 1.085 ;
        RECT 19.485 0.57 19.655 1.08 ;
        RECT 19.485 2.39 19.655 3.86 ;
      LAYER met1 ;
        RECT 19.425 2.36 19.715 2.59 ;
        RECT 19.425 0.88 19.715 1.11 ;
        RECT 19.485 0.88 19.655 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 36.71 0.915 36.88 1.085 ;
        RECT 36.705 0.91 36.875 1.08 ;
        RECT 36.705 2.39 36.875 2.56 ;
      LAYER li1 ;
        RECT 36.71 0.915 36.88 1.085 ;
        RECT 36.705 0.57 36.875 1.08 ;
        RECT 36.705 2.39 36.875 3.86 ;
      LAYER met1 ;
        RECT 36.645 2.36 36.935 2.59 ;
        RECT 36.645 0.88 36.935 1.11 ;
        RECT 36.705 0.88 36.875 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 53.93 0.915 54.1 1.085 ;
        RECT 53.925 0.91 54.095 1.08 ;
        RECT 53.925 2.39 54.095 2.56 ;
      LAYER li1 ;
        RECT 53.93 0.915 54.1 1.085 ;
        RECT 53.925 0.57 54.095 1.08 ;
        RECT 53.925 2.39 54.095 3.86 ;
      LAYER met1 ;
        RECT 53.865 2.36 54.155 2.59 ;
        RECT 53.865 0.88 54.155 1.11 ;
        RECT 53.925 0.88 54.095 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 71.15 0.915 71.32 1.085 ;
        RECT 71.145 0.91 71.315 1.08 ;
        RECT 71.145 2.39 71.315 2.56 ;
      LAYER li1 ;
        RECT 71.15 0.915 71.32 1.085 ;
        RECT 71.145 0.57 71.315 1.08 ;
        RECT 71.145 2.39 71.315 3.86 ;
      LAYER met1 ;
        RECT 71.085 2.36 71.375 2.59 ;
        RECT 71.085 0.88 71.375 1.11 ;
        RECT 71.145 0.88 71.315 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 88.37 0.915 88.54 1.085 ;
        RECT 88.365 0.91 88.535 1.08 ;
        RECT 88.365 2.39 88.535 2.56 ;
      LAYER li1 ;
        RECT 88.37 0.915 88.54 1.085 ;
        RECT 88.365 0.57 88.535 1.08 ;
        RECT 88.365 2.39 88.535 3.86 ;
      LAYER met1 ;
        RECT 88.305 2.36 88.595 2.59 ;
        RECT 88.305 0.88 88.595 1.11 ;
        RECT 88.365 0.88 88.535 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 15.335 1.66 15.505 2.935 ;
        RECT 15.335 5.94 15.505 7.22 ;
        RECT 15.325 5.94 15.505 6.18 ;
        RECT 3.65 5.945 3.82 7.22 ;
      LAYER met2 ;
        RECT 15.255 5.855 15.58 6.18 ;
        RECT 15.255 3.495 15.58 3.82 ;
        RECT 5.955 7.55 15.505 7.72 ;
        RECT 15.335 5.855 15.505 7.72 ;
        RECT 15.325 3.495 15.495 6.18 ;
        RECT 5.9 5.86 6.18 6.2 ;
        RECT 5.955 5.86 6.125 7.72 ;
      LAYER met1 ;
        RECT 15.275 2.765 15.735 2.935 ;
        RECT 15.255 3.495 15.58 3.82 ;
        RECT 15.275 2.735 15.565 2.965 ;
        RECT 15.335 2.735 15.505 3.82 ;
        RECT 15.255 5.945 15.735 6.115 ;
        RECT 15.255 5.855 15.58 6.18 ;
        RECT 5.87 5.89 6.21 6.17 ;
        RECT 3.59 5.945 6.21 6.115 ;
        RECT 3.59 5.915 3.88 6.145 ;
      LAYER mcon ;
        RECT 3.65 5.945 3.82 6.115 ;
        RECT 15.335 5.945 15.505 6.115 ;
        RECT 15.335 2.765 15.505 2.935 ;
      LAYER via1 ;
        RECT 5.965 5.955 6.115 6.105 ;
        RECT 15.345 5.94 15.495 6.09 ;
        RECT 15.345 3.58 15.495 3.73 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 32.555 1.66 32.725 2.935 ;
        RECT 32.555 5.94 32.725 7.22 ;
        RECT 32.545 5.94 32.725 6.18 ;
        RECT 20.87 5.945 21.04 7.22 ;
      LAYER met2 ;
        RECT 32.475 5.855 32.8 6.18 ;
        RECT 32.475 3.495 32.8 3.82 ;
        RECT 23.175 7.55 32.725 7.72 ;
        RECT 32.555 5.855 32.725 7.72 ;
        RECT 32.545 3.495 32.715 6.18 ;
        RECT 23.12 5.86 23.4 6.2 ;
        RECT 23.175 5.86 23.345 7.72 ;
      LAYER met1 ;
        RECT 32.495 2.765 32.955 2.935 ;
        RECT 32.475 3.495 32.8 3.82 ;
        RECT 32.495 2.735 32.785 2.965 ;
        RECT 32.555 2.735 32.725 3.82 ;
        RECT 32.475 5.945 32.955 6.115 ;
        RECT 32.475 5.855 32.8 6.18 ;
        RECT 23.09 5.89 23.43 6.17 ;
        RECT 20.81 5.945 23.43 6.115 ;
        RECT 20.81 5.915 21.1 6.145 ;
      LAYER mcon ;
        RECT 20.87 5.945 21.04 6.115 ;
        RECT 32.555 5.945 32.725 6.115 ;
        RECT 32.555 2.765 32.725 2.935 ;
      LAYER via1 ;
        RECT 23.185 5.955 23.335 6.105 ;
        RECT 32.565 5.94 32.715 6.09 ;
        RECT 32.565 3.58 32.715 3.73 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 49.775 1.66 49.945 2.935 ;
        RECT 49.775 5.94 49.945 7.22 ;
        RECT 49.765 5.94 49.945 6.18 ;
        RECT 38.09 5.945 38.26 7.22 ;
      LAYER met2 ;
        RECT 49.695 5.855 50.02 6.18 ;
        RECT 49.695 3.495 50.02 3.82 ;
        RECT 40.395 7.55 49.945 7.72 ;
        RECT 49.775 5.855 49.945 7.72 ;
        RECT 49.765 3.495 49.935 6.18 ;
        RECT 40.34 5.86 40.62 6.2 ;
        RECT 40.395 5.86 40.565 7.72 ;
      LAYER met1 ;
        RECT 49.715 2.765 50.175 2.935 ;
        RECT 49.695 3.495 50.02 3.82 ;
        RECT 49.715 2.735 50.005 2.965 ;
        RECT 49.775 2.735 49.945 3.82 ;
        RECT 49.695 5.945 50.175 6.115 ;
        RECT 49.695 5.855 50.02 6.18 ;
        RECT 40.31 5.89 40.65 6.17 ;
        RECT 38.03 5.945 40.65 6.115 ;
        RECT 38.03 5.915 38.32 6.145 ;
      LAYER mcon ;
        RECT 38.09 5.945 38.26 6.115 ;
        RECT 49.775 5.945 49.945 6.115 ;
        RECT 49.775 2.765 49.945 2.935 ;
      LAYER via1 ;
        RECT 40.405 5.955 40.555 6.105 ;
        RECT 49.785 5.94 49.935 6.09 ;
        RECT 49.785 3.58 49.935 3.73 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 66.995 1.66 67.165 2.935 ;
        RECT 66.995 5.94 67.165 7.22 ;
        RECT 66.985 5.94 67.165 6.18 ;
        RECT 55.31 5.945 55.48 7.22 ;
      LAYER met2 ;
        RECT 66.915 5.855 67.24 6.18 ;
        RECT 66.915 3.495 67.24 3.82 ;
        RECT 57.615 7.55 67.165 7.72 ;
        RECT 66.995 5.855 67.165 7.72 ;
        RECT 66.985 3.495 67.155 6.18 ;
        RECT 57.56 5.86 57.84 6.2 ;
        RECT 57.615 5.86 57.785 7.72 ;
      LAYER met1 ;
        RECT 66.935 2.765 67.395 2.935 ;
        RECT 66.915 3.495 67.24 3.82 ;
        RECT 66.935 2.735 67.225 2.965 ;
        RECT 66.995 2.735 67.165 3.82 ;
        RECT 66.915 5.945 67.395 6.115 ;
        RECT 66.915 5.855 67.24 6.18 ;
        RECT 57.53 5.89 57.87 6.17 ;
        RECT 55.25 5.945 57.87 6.115 ;
        RECT 55.25 5.915 55.54 6.145 ;
      LAYER mcon ;
        RECT 55.31 5.945 55.48 6.115 ;
        RECT 66.995 5.945 67.165 6.115 ;
        RECT 66.995 2.765 67.165 2.935 ;
      LAYER via1 ;
        RECT 57.625 5.955 57.775 6.105 ;
        RECT 67.005 5.94 67.155 6.09 ;
        RECT 67.005 3.58 67.155 3.73 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 84.215 1.66 84.385 2.935 ;
        RECT 84.215 5.94 84.385 7.22 ;
        RECT 84.205 5.94 84.385 6.18 ;
        RECT 72.53 5.945 72.7 7.22 ;
      LAYER met2 ;
        RECT 84.135 5.855 84.46 6.18 ;
        RECT 84.135 3.495 84.46 3.82 ;
        RECT 74.835 7.55 84.385 7.72 ;
        RECT 84.215 5.855 84.385 7.72 ;
        RECT 84.205 3.495 84.375 6.18 ;
        RECT 74.78 5.86 75.06 6.2 ;
        RECT 74.835 5.86 75.005 7.72 ;
      LAYER met1 ;
        RECT 84.155 2.765 84.615 2.935 ;
        RECT 84.135 3.495 84.46 3.82 ;
        RECT 84.155 2.735 84.445 2.965 ;
        RECT 84.215 2.735 84.385 3.82 ;
        RECT 84.135 5.945 84.615 6.115 ;
        RECT 84.135 5.855 84.46 6.18 ;
        RECT 74.75 5.89 75.09 6.17 ;
        RECT 72.47 5.945 75.09 6.115 ;
        RECT 72.47 5.915 72.76 6.145 ;
      LAYER mcon ;
        RECT 72.53 5.945 72.7 6.115 ;
        RECT 84.215 5.945 84.385 6.115 ;
        RECT 84.215 2.765 84.385 2.935 ;
      LAYER via1 ;
        RECT 74.845 5.955 74.995 6.105 ;
        RECT 84.225 5.94 84.375 6.09 ;
        RECT 84.225 3.58 84.375 3.73 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.24 5.945 0.41 7.22 ;
      LAYER met1 ;
        RECT 0.18 5.945 0.64 6.115 ;
        RECT 0.18 5.915 0.47 6.145 ;
      LAYER mcon ;
        RECT 0.24 5.945 0.41 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.38 4.255 2.185 4.635 ;
      LAYER li1 ;
        RECT 82.925 4.135 88.91 4.745 ;
        RECT 86.775 4.13 88.755 4.75 ;
        RECT 87.935 3.4 88.105 5.48 ;
        RECT 86.945 3.4 87.115 5.48 ;
        RECT 84.205 3.405 84.375 5.475 ;
        RECT 82.92 4.135 88.91 4.515 ;
        RECT 1.845 4.345 88.91 4.515 ;
        RECT 82.01 4.345 82.29 5.655 ;
        RECT 81.61 3.495 81.78 4.515 ;
        RECT 81.08 4.345 81.34 5.655 ;
        RECT 80.77 3.835 80.94 4.515 ;
        RECT 80.63 4.345 80.91 5.655 ;
        RECT 79.7 4.345 79.96 5.655 ;
        RECT 79.27 4.345 79.53 5.655 ;
        RECT 79.19 3.205 79.52 4.515 ;
        RECT 78.32 4.345 78.6 5.655 ;
        RECT 76.95 3.205 77.28 4.515 ;
        RECT 76.97 3.205 77.23 5.655 ;
        RECT 76.5 3.205 76.73 4.515 ;
        RECT 76.02 4.345 76.3 5.655 ;
        RECT 65.705 4.345 75.85 4.74 ;
        RECT 65.7 4.135 75.83 4.515 ;
        RECT 75.62 3.205 75.83 4.74 ;
        RECT 71.685 4.13 75.83 4.74 ;
        RECT 72.345 4.13 75.095 4.745 ;
        RECT 72.52 4.13 72.69 5.475 ;
        RECT 65.705 4.135 71.69 4.745 ;
        RECT 69.555 4.13 71.535 4.75 ;
        RECT 70.715 3.4 70.885 5.48 ;
        RECT 69.725 3.4 69.895 5.48 ;
        RECT 66.985 3.405 67.155 5.475 ;
        RECT 64.79 4.345 65.07 5.655 ;
        RECT 64.39 3.495 64.56 4.515 ;
        RECT 63.86 4.345 64.12 5.655 ;
        RECT 63.55 3.835 63.72 4.515 ;
        RECT 63.41 4.345 63.69 5.655 ;
        RECT 62.48 4.345 62.74 5.655 ;
        RECT 62.05 4.345 62.31 5.655 ;
        RECT 61.97 3.205 62.3 4.515 ;
        RECT 61.1 4.345 61.38 5.655 ;
        RECT 59.73 3.205 60.06 4.515 ;
        RECT 59.75 3.205 60.01 5.655 ;
        RECT 59.28 3.205 59.51 4.515 ;
        RECT 58.8 4.345 59.08 5.655 ;
        RECT 48.485 4.345 58.63 4.74 ;
        RECT 48.48 4.135 58.61 4.515 ;
        RECT 58.4 3.205 58.61 4.74 ;
        RECT 54.465 4.13 58.61 4.74 ;
        RECT 55.125 4.13 57.875 4.745 ;
        RECT 55.3 4.13 55.47 5.475 ;
        RECT 48.485 4.135 54.47 4.745 ;
        RECT 52.335 4.13 54.315 4.75 ;
        RECT 53.495 3.4 53.665 5.48 ;
        RECT 52.505 3.4 52.675 5.48 ;
        RECT 49.765 3.405 49.935 5.475 ;
        RECT 47.57 4.345 47.85 5.655 ;
        RECT 47.17 3.495 47.34 4.515 ;
        RECT 46.64 4.345 46.9 5.655 ;
        RECT 46.33 3.835 46.5 4.515 ;
        RECT 46.19 4.345 46.47 5.655 ;
        RECT 45.26 4.345 45.52 5.655 ;
        RECT 44.83 4.345 45.09 5.655 ;
        RECT 44.75 3.205 45.08 4.515 ;
        RECT 43.88 4.345 44.16 5.655 ;
        RECT 42.51 3.205 42.84 4.515 ;
        RECT 42.53 3.205 42.79 5.655 ;
        RECT 42.06 3.205 42.29 4.515 ;
        RECT 41.58 4.345 41.86 5.655 ;
        RECT 31.265 4.345 41.41 4.74 ;
        RECT 31.26 4.135 41.39 4.515 ;
        RECT 41.18 3.205 41.39 4.74 ;
        RECT 37.245 4.13 41.39 4.74 ;
        RECT 37.905 4.13 40.655 4.745 ;
        RECT 38.08 4.13 38.25 5.475 ;
        RECT 31.265 4.135 37.25 4.745 ;
        RECT 35.115 4.13 37.095 4.75 ;
        RECT 36.275 3.4 36.445 5.48 ;
        RECT 35.285 3.4 35.455 5.48 ;
        RECT 32.545 3.405 32.715 5.475 ;
        RECT 30.35 4.345 30.63 5.655 ;
        RECT 29.95 3.495 30.12 4.515 ;
        RECT 29.42 4.345 29.68 5.655 ;
        RECT 29.11 3.835 29.28 4.515 ;
        RECT 28.97 4.345 29.25 5.655 ;
        RECT 28.04 4.345 28.3 5.655 ;
        RECT 27.61 4.345 27.87 5.655 ;
        RECT 27.53 3.205 27.86 4.515 ;
        RECT 26.66 4.345 26.94 5.655 ;
        RECT 25.29 3.205 25.62 4.515 ;
        RECT 25.31 3.205 25.57 5.655 ;
        RECT 24.84 3.205 25.07 4.515 ;
        RECT 24.36 4.345 24.64 5.655 ;
        RECT 14.045 4.345 24.19 4.74 ;
        RECT 14.04 4.135 24.17 4.515 ;
        RECT 23.96 3.205 24.17 4.74 ;
        RECT 20.025 4.13 24.17 4.74 ;
        RECT 20.685 4.13 23.435 4.745 ;
        RECT 20.86 4.13 21.03 5.475 ;
        RECT 14.045 4.135 20.03 4.745 ;
        RECT 17.895 4.13 19.875 4.75 ;
        RECT 19.055 3.4 19.225 5.48 ;
        RECT 18.065 3.4 18.235 5.48 ;
        RECT 15.325 3.405 15.495 5.475 ;
        RECT 13.13 4.345 13.41 5.655 ;
        RECT 12.73 3.495 12.9 4.515 ;
        RECT 12.2 4.345 12.46 5.655 ;
        RECT 11.89 3.835 12.06 4.515 ;
        RECT 11.75 4.345 12.03 5.655 ;
        RECT 10.82 4.345 11.08 5.655 ;
        RECT 10.39 4.345 10.65 5.655 ;
        RECT 10.31 3.205 10.64 4.515 ;
        RECT 9.44 4.345 9.72 5.655 ;
        RECT 8.07 3.205 8.4 4.515 ;
        RECT 8.09 3.205 8.35 5.655 ;
        RECT 7.62 3.205 7.85 4.515 ;
        RECT 7.14 4.345 7.42 5.655 ;
        RECT 0 4.44 6.97 4.74 ;
        RECT 1.845 4.13 6.95 4.74 ;
        RECT 6.74 3.205 6.95 4.74 ;
        RECT 3.465 4.13 6.215 4.745 ;
        RECT 3.64 4.13 3.81 5.475 ;
        RECT 0.055 4.44 2.805 4.745 ;
        RECT 2.04 4.13 2.21 8.305 ;
        RECT 0 4.13 6.95 4.33 ;
        RECT 0 4.13 1.675 4.74 ;
        RECT 0.23 4.13 0.4 5.475 ;
      LAYER met2 ;
        RECT 1.57 4.255 1.95 4.635 ;
      LAYER met1 ;
        RECT 82.925 4.135 88.91 4.745 ;
        RECT 86.775 4.13 88.755 4.75 ;
        RECT 0 4.19 88.91 4.67 ;
        RECT 82.92 4.135 88.91 4.67 ;
        RECT 65.705 4.19 75.85 4.74 ;
        RECT 65.7 4.135 75.83 4.67 ;
        RECT 71.685 4.13 75.83 4.74 ;
        RECT 72.345 4.13 75.095 4.745 ;
        RECT 65.705 4.135 71.69 4.745 ;
        RECT 69.555 4.13 71.535 4.75 ;
        RECT 48.485 4.19 58.63 4.74 ;
        RECT 48.48 4.135 58.61 4.67 ;
        RECT 54.465 4.13 58.61 4.74 ;
        RECT 55.125 4.13 57.875 4.745 ;
        RECT 48.485 4.135 54.47 4.745 ;
        RECT 52.335 4.13 54.315 4.75 ;
        RECT 31.265 4.19 41.41 4.74 ;
        RECT 31.26 4.135 41.39 4.67 ;
        RECT 37.245 4.13 41.39 4.74 ;
        RECT 37.905 4.13 40.655 4.745 ;
        RECT 31.265 4.135 37.25 4.745 ;
        RECT 35.115 4.13 37.095 4.75 ;
        RECT 14.045 4.19 24.19 4.74 ;
        RECT 14.04 4.135 24.17 4.67 ;
        RECT 20.025 4.13 24.17 4.74 ;
        RECT 20.685 4.13 23.435 4.745 ;
        RECT 14.045 4.135 20.03 4.745 ;
        RECT 17.895 4.13 19.875 4.75 ;
        RECT 0 4.19 6.97 4.74 ;
        RECT 0 4.13 6.95 4.74 ;
        RECT 3.465 4.13 6.215 4.745 ;
        RECT 0.055 4.13 2.805 4.745 ;
        RECT 1.98 6.655 2.27 6.885 ;
        RECT 1.81 6.685 2.27 6.855 ;
      LAYER via2 ;
        RECT 1.66 4.345 1.86 4.545 ;
      LAYER mcon ;
        RECT 2.04 6.685 2.21 6.855 ;
        RECT 2.35 4.545 2.52 4.715 ;
        RECT 5.76 4.545 5.93 4.715 ;
        RECT 6.74 4.345 6.91 4.515 ;
        RECT 7.2 4.345 7.37 4.515 ;
        RECT 7.66 4.345 7.83 4.515 ;
        RECT 8.12 4.345 8.29 4.515 ;
        RECT 8.58 4.345 8.75 4.515 ;
        RECT 9.04 4.345 9.21 4.515 ;
        RECT 9.5 4.345 9.67 4.515 ;
        RECT 9.96 4.345 10.13 4.515 ;
        RECT 10.42 4.345 10.59 4.515 ;
        RECT 10.88 4.345 11.05 4.515 ;
        RECT 11.34 4.345 11.51 4.515 ;
        RECT 11.8 4.345 11.97 4.515 ;
        RECT 12.26 4.345 12.43 4.515 ;
        RECT 12.72 4.345 12.89 4.515 ;
        RECT 13.18 4.345 13.35 4.515 ;
        RECT 13.64 4.345 13.81 4.515 ;
        RECT 17.445 4.545 17.615 4.715 ;
        RECT 17.445 4.165 17.615 4.335 ;
        RECT 18.145 4.55 18.315 4.72 ;
        RECT 18.145 4.16 18.315 4.33 ;
        RECT 19.135 4.55 19.305 4.72 ;
        RECT 19.135 4.16 19.305 4.33 ;
        RECT 22.98 4.545 23.15 4.715 ;
        RECT 23.96 4.345 24.13 4.515 ;
        RECT 24.42 4.345 24.59 4.515 ;
        RECT 24.88 4.345 25.05 4.515 ;
        RECT 25.34 4.345 25.51 4.515 ;
        RECT 25.8 4.345 25.97 4.515 ;
        RECT 26.26 4.345 26.43 4.515 ;
        RECT 26.72 4.345 26.89 4.515 ;
        RECT 27.18 4.345 27.35 4.515 ;
        RECT 27.64 4.345 27.81 4.515 ;
        RECT 28.1 4.345 28.27 4.515 ;
        RECT 28.56 4.345 28.73 4.515 ;
        RECT 29.02 4.345 29.19 4.515 ;
        RECT 29.48 4.345 29.65 4.515 ;
        RECT 29.94 4.345 30.11 4.515 ;
        RECT 30.4 4.345 30.57 4.515 ;
        RECT 30.86 4.345 31.03 4.515 ;
        RECT 34.665 4.545 34.835 4.715 ;
        RECT 34.665 4.165 34.835 4.335 ;
        RECT 35.365 4.55 35.535 4.72 ;
        RECT 35.365 4.16 35.535 4.33 ;
        RECT 36.355 4.55 36.525 4.72 ;
        RECT 36.355 4.16 36.525 4.33 ;
        RECT 40.2 4.545 40.37 4.715 ;
        RECT 41.18 4.345 41.35 4.515 ;
        RECT 41.64 4.345 41.81 4.515 ;
        RECT 42.1 4.345 42.27 4.515 ;
        RECT 42.56 4.345 42.73 4.515 ;
        RECT 43.02 4.345 43.19 4.515 ;
        RECT 43.48 4.345 43.65 4.515 ;
        RECT 43.94 4.345 44.11 4.515 ;
        RECT 44.4 4.345 44.57 4.515 ;
        RECT 44.86 4.345 45.03 4.515 ;
        RECT 45.32 4.345 45.49 4.515 ;
        RECT 45.78 4.345 45.95 4.515 ;
        RECT 46.24 4.345 46.41 4.515 ;
        RECT 46.7 4.345 46.87 4.515 ;
        RECT 47.16 4.345 47.33 4.515 ;
        RECT 47.62 4.345 47.79 4.515 ;
        RECT 48.08 4.345 48.25 4.515 ;
        RECT 51.885 4.545 52.055 4.715 ;
        RECT 51.885 4.165 52.055 4.335 ;
        RECT 52.585 4.55 52.755 4.72 ;
        RECT 52.585 4.16 52.755 4.33 ;
        RECT 53.575 4.55 53.745 4.72 ;
        RECT 53.575 4.16 53.745 4.33 ;
        RECT 57.42 4.545 57.59 4.715 ;
        RECT 58.4 4.345 58.57 4.515 ;
        RECT 58.86 4.345 59.03 4.515 ;
        RECT 59.32 4.345 59.49 4.515 ;
        RECT 59.78 4.345 59.95 4.515 ;
        RECT 60.24 4.345 60.41 4.515 ;
        RECT 60.7 4.345 60.87 4.515 ;
        RECT 61.16 4.345 61.33 4.515 ;
        RECT 61.62 4.345 61.79 4.515 ;
        RECT 62.08 4.345 62.25 4.515 ;
        RECT 62.54 4.345 62.71 4.515 ;
        RECT 63 4.345 63.17 4.515 ;
        RECT 63.46 4.345 63.63 4.515 ;
        RECT 63.92 4.345 64.09 4.515 ;
        RECT 64.38 4.345 64.55 4.515 ;
        RECT 64.84 4.345 65.01 4.515 ;
        RECT 65.3 4.345 65.47 4.515 ;
        RECT 69.105 4.545 69.275 4.715 ;
        RECT 69.105 4.165 69.275 4.335 ;
        RECT 69.805 4.55 69.975 4.72 ;
        RECT 69.805 4.16 69.975 4.33 ;
        RECT 70.795 4.55 70.965 4.72 ;
        RECT 70.795 4.16 70.965 4.33 ;
        RECT 74.64 4.545 74.81 4.715 ;
        RECT 75.62 4.345 75.79 4.515 ;
        RECT 76.08 4.345 76.25 4.515 ;
        RECT 76.54 4.345 76.71 4.515 ;
        RECT 77 4.345 77.17 4.515 ;
        RECT 77.46 4.345 77.63 4.515 ;
        RECT 77.92 4.345 78.09 4.515 ;
        RECT 78.38 4.345 78.55 4.515 ;
        RECT 78.84 4.345 79.01 4.515 ;
        RECT 79.3 4.345 79.47 4.515 ;
        RECT 79.76 4.345 79.93 4.515 ;
        RECT 80.22 4.345 80.39 4.515 ;
        RECT 80.68 4.345 80.85 4.515 ;
        RECT 81.14 4.345 81.31 4.515 ;
        RECT 81.6 4.345 81.77 4.515 ;
        RECT 82.06 4.345 82.23 4.515 ;
        RECT 82.52 4.345 82.69 4.515 ;
        RECT 86.325 4.545 86.495 4.715 ;
        RECT 86.325 4.165 86.495 4.335 ;
        RECT 87.025 4.55 87.195 4.72 ;
        RECT 87.025 4.16 87.195 4.33 ;
        RECT 88.015 4.55 88.185 4.72 ;
        RECT 88.015 4.16 88.185 4.33 ;
      LAYER via1 ;
        RECT 1.685 4.37 1.835 4.52 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 77.86 5.79 78.19 6.12 ;
        RECT 77.39 5.805 78.19 6.105 ;
        RECT 60.64 5.79 60.97 6.12 ;
        RECT 60.17 5.805 60.97 6.105 ;
        RECT 43.42 5.79 43.75 6.12 ;
        RECT 42.95 5.805 43.75 6.105 ;
        RECT 26.2 5.79 26.53 6.12 ;
        RECT 25.73 5.805 26.53 6.105 ;
        RECT 8.98 5.79 9.31 6.12 ;
        RECT 8.51 5.805 9.31 6.105 ;
        RECT 0.015 8.5 0.82 8.88 ;
        RECT 0 0 0.805 0.38 ;
      LAYER li1 ;
        RECT 88.73 0 88.91 0.305 ;
        RECT 0.465 0 88.91 0.3 ;
        RECT 87.935 0 88.105 0.93 ;
        RECT 86.945 0 87.115 0.93 ;
        RECT 71.51 0 86.78 0.305 ;
        RECT 84.205 0 84.375 0.935 ;
        RECT 75.475 0 83.13 1.795 ;
        RECT 82.37 0 82.7 2.185 ;
        RECT 81.53 0 81.86 2.185 ;
        RECT 79.7 0 79.99 2.63 ;
        RECT 79.25 0 79.52 2.605 ;
        RECT 78.34 0 78.58 2.605 ;
        RECT 77.89 0 78.13 2.605 ;
        RECT 76.95 0 77.22 2.605 ;
        RECT 76.5 0 76.73 2.615 ;
        RECT 75.62 0 75.83 2.615 ;
        RECT 75.47 0 83.13 1.635 ;
        RECT 70.715 0 70.885 0.93 ;
        RECT 69.725 0 69.895 0.93 ;
        RECT 54.29 0 69.56 0.305 ;
        RECT 66.985 0 67.155 0.935 ;
        RECT 58.255 0 65.91 1.795 ;
        RECT 65.15 0 65.48 2.185 ;
        RECT 64.31 0 64.64 2.185 ;
        RECT 62.48 0 62.77 2.63 ;
        RECT 62.03 0 62.3 2.605 ;
        RECT 61.12 0 61.36 2.605 ;
        RECT 60.67 0 60.91 2.605 ;
        RECT 59.73 0 60 2.605 ;
        RECT 59.28 0 59.51 2.615 ;
        RECT 58.4 0 58.61 2.615 ;
        RECT 58.25 0 65.91 1.635 ;
        RECT 53.495 0 53.665 0.93 ;
        RECT 52.505 0 52.675 0.93 ;
        RECT 37.07 0 52.34 0.305 ;
        RECT 49.765 0 49.935 0.935 ;
        RECT 41.035 0 48.69 1.795 ;
        RECT 47.93 0 48.26 2.185 ;
        RECT 47.09 0 47.42 2.185 ;
        RECT 45.26 0 45.55 2.63 ;
        RECT 44.81 0 45.08 2.605 ;
        RECT 43.9 0 44.14 2.605 ;
        RECT 43.45 0 43.69 2.605 ;
        RECT 42.51 0 42.78 2.605 ;
        RECT 42.06 0 42.29 2.615 ;
        RECT 41.18 0 41.39 2.615 ;
        RECT 41.03 0 48.69 1.635 ;
        RECT 36.275 0 36.445 0.93 ;
        RECT 35.285 0 35.455 0.93 ;
        RECT 19.85 0 35.12 0.305 ;
        RECT 32.545 0 32.715 0.935 ;
        RECT 23.815 0 31.47 1.795 ;
        RECT 30.71 0 31.04 2.185 ;
        RECT 29.87 0 30.2 2.185 ;
        RECT 28.04 0 28.33 2.63 ;
        RECT 27.59 0 27.86 2.605 ;
        RECT 26.68 0 26.92 2.605 ;
        RECT 26.23 0 26.47 2.605 ;
        RECT 25.29 0 25.56 2.605 ;
        RECT 24.84 0 25.07 2.615 ;
        RECT 23.96 0 24.17 2.615 ;
        RECT 23.81 0 31.47 1.635 ;
        RECT 19.055 0 19.225 0.93 ;
        RECT 18.065 0 18.235 0.93 ;
        RECT 0 0.245 17.9 0.305 ;
        RECT 15.325 0 15.495 0.935 ;
        RECT 6.595 0 14.25 1.795 ;
        RECT 13.49 0 13.82 2.185 ;
        RECT 12.65 0 12.98 2.185 ;
        RECT 10.82 0 11.11 2.63 ;
        RECT 10.37 0 10.64 2.605 ;
        RECT 9.46 0 9.7 2.605 ;
        RECT 9.01 0 9.25 2.605 ;
        RECT 8.07 0 8.34 2.605 ;
        RECT 7.62 0 7.85 2.615 ;
        RECT 6.74 0 6.95 2.615 ;
        RECT 6.59 0 14.25 1.635 ;
        RECT 0 0.245 0.805 0.315 ;
        RECT 0.295 0.245 0.465 0.335 ;
        RECT 0 0 88.91 0.075 ;
        RECT 0 0 0.295 0.315 ;
        RECT 0 8.58 88.91 8.88 ;
        RECT 88.73 8.575 88.91 8.88 ;
        RECT 87.935 7.95 88.105 8.88 ;
        RECT 86.945 7.95 87.115 8.88 ;
        RECT 71.51 8.575 86.78 8.88 ;
        RECT 84.205 7.945 84.375 8.88 ;
        RECT 75.745 7.18 82.945 8.88 ;
        RECT 75.475 7.065 82.835 7.235 ;
        RECT 81.98 6.265 82.29 8.88 ;
        RECT 80.6 6.265 80.91 8.88 ;
        RECT 78.33 5.825 78.665 6.095 ;
        RECT 78.32 6.265 78.63 8.88 ;
        RECT 77.94 5.875 78.665 6.045 ;
        RECT 77.95 5.875 78.12 8.88 ;
        RECT 76.02 6.265 76.33 8.88 ;
        RECT 72.52 7.945 72.69 8.88 ;
        RECT 70.715 7.95 70.885 8.88 ;
        RECT 69.725 7.95 69.895 8.88 ;
        RECT 54.29 8.575 69.56 8.88 ;
        RECT 66.985 7.945 67.155 8.88 ;
        RECT 58.525 7.18 65.725 8.88 ;
        RECT 58.255 7.065 65.615 7.235 ;
        RECT 64.76 6.265 65.07 8.88 ;
        RECT 63.38 6.265 63.69 8.88 ;
        RECT 61.11 5.825 61.445 6.095 ;
        RECT 61.1 6.265 61.41 8.88 ;
        RECT 60.72 5.875 61.445 6.045 ;
        RECT 60.73 5.875 60.9 8.88 ;
        RECT 58.8 6.265 59.11 8.88 ;
        RECT 55.3 7.945 55.47 8.88 ;
        RECT 53.495 7.95 53.665 8.88 ;
        RECT 52.505 7.95 52.675 8.88 ;
        RECT 37.07 8.575 52.34 8.88 ;
        RECT 49.765 7.945 49.935 8.88 ;
        RECT 41.305 7.18 48.505 8.88 ;
        RECT 41.035 7.065 48.395 7.235 ;
        RECT 47.54 6.265 47.85 8.88 ;
        RECT 46.16 6.265 46.47 8.88 ;
        RECT 43.89 5.825 44.225 6.095 ;
        RECT 43.88 6.265 44.19 8.88 ;
        RECT 43.5 5.875 44.225 6.045 ;
        RECT 43.51 5.875 43.68 8.88 ;
        RECT 41.58 6.265 41.89 8.88 ;
        RECT 38.08 7.945 38.25 8.88 ;
        RECT 36.275 7.95 36.445 8.88 ;
        RECT 35.285 7.95 35.455 8.88 ;
        RECT 19.85 8.575 35.12 8.88 ;
        RECT 32.545 7.945 32.715 8.88 ;
        RECT 24.085 7.18 31.285 8.88 ;
        RECT 23.815 7.065 31.175 7.235 ;
        RECT 30.32 6.265 30.63 8.88 ;
        RECT 28.94 6.265 29.25 8.88 ;
        RECT 26.67 5.825 27.005 6.095 ;
        RECT 26.66 6.265 26.97 8.88 ;
        RECT 26.28 5.875 27.005 6.045 ;
        RECT 26.29 5.875 26.46 8.88 ;
        RECT 24.36 6.265 24.67 8.88 ;
        RECT 20.86 7.945 21.03 8.88 ;
        RECT 19.055 7.95 19.225 8.88 ;
        RECT 18.065 7.95 18.235 8.88 ;
        RECT 0 8.575 17.9 8.88 ;
        RECT 15.325 7.945 15.495 8.88 ;
        RECT 6.865 7.18 14.065 8.88 ;
        RECT 6.595 7.065 13.955 7.235 ;
        RECT 13.1 6.265 13.41 8.88 ;
        RECT 11.72 6.265 12.03 8.88 ;
        RECT 9.45 5.825 9.785 6.095 ;
        RECT 9.44 6.265 9.75 8.88 ;
        RECT 9.06 5.875 9.785 6.045 ;
        RECT 9.07 5.875 9.24 8.88 ;
        RECT 7.14 6.265 7.45 8.88 ;
        RECT 3.64 7.945 3.81 8.88 ;
        RECT 0.015 8.565 0.82 8.88 ;
        RECT 0.23 8.545 0.48 8.88 ;
        RECT 0.23 7.945 0.4 8.88 ;
        RECT 76.03 5.825 76.365 6.095 ;
        RECT 75.56 5.875 76.365 6.045 ;
        RECT 73.525 6.075 73.695 8.025 ;
        RECT 73.47 7.855 73.64 8.305 ;
        RECT 73.47 5.015 73.64 6.245 ;
        RECT 58.81 5.825 59.145 6.095 ;
        RECT 58.34 5.875 59.145 6.045 ;
        RECT 56.305 6.075 56.475 8.025 ;
        RECT 56.25 7.855 56.42 8.305 ;
        RECT 56.25 5.015 56.42 6.245 ;
        RECT 41.59 5.825 41.925 6.095 ;
        RECT 41.12 5.875 41.925 6.045 ;
        RECT 39.085 6.075 39.255 8.025 ;
        RECT 39.03 7.855 39.2 8.305 ;
        RECT 39.03 5.015 39.2 6.245 ;
        RECT 24.37 5.825 24.705 6.095 ;
        RECT 23.9 5.875 24.705 6.045 ;
        RECT 21.865 6.075 22.035 8.025 ;
        RECT 21.81 7.855 21.98 8.305 ;
        RECT 21.81 5.015 21.98 6.245 ;
        RECT 7.15 5.825 7.485 6.095 ;
        RECT 6.68 5.875 7.485 6.045 ;
        RECT 4.645 6.075 4.815 8.025 ;
        RECT 4.59 7.855 4.76 8.305 ;
        RECT 4.59 5.015 4.76 6.245 ;
      LAYER met2 ;
        RECT 77.885 5.77 78.165 6.14 ;
        RECT 60.665 5.77 60.945 6.14 ;
        RECT 43.445 5.77 43.725 6.14 ;
        RECT 26.225 5.77 26.505 6.14 ;
        RECT 9.005 5.77 9.285 6.14 ;
        RECT 0.205 8.5 0.585 8.88 ;
        RECT 0.19 0 0.57 0.38 ;
        RECT 0.235 0 0.385 8.88 ;
      LAYER met1 ;
        RECT 88.73 0 88.91 0.305 ;
        RECT 0 0 88.91 0.3 ;
        RECT 71.51 0 86.78 0.305 ;
        RECT 75.475 0 83.13 1.795 ;
        RECT 75.475 0 82.835 1.95 ;
        RECT 75.47 0 83.13 1.635 ;
        RECT 54.29 0 69.56 0.305 ;
        RECT 58.255 0 65.91 1.795 ;
        RECT 58.255 0 65.615 1.95 ;
        RECT 58.25 0 65.91 1.635 ;
        RECT 37.07 0 52.34 0.305 ;
        RECT 41.035 0 48.69 1.795 ;
        RECT 41.035 0 48.395 1.95 ;
        RECT 41.03 0 48.69 1.635 ;
        RECT 19.85 0 35.12 0.305 ;
        RECT 23.815 0 31.47 1.795 ;
        RECT 23.815 0 31.175 1.95 ;
        RECT 23.81 0 31.47 1.635 ;
        RECT 0 0 17.9 0.305 ;
        RECT 6.595 0 14.25 1.795 ;
        RECT 6.595 0 13.955 1.95 ;
        RECT 6.59 0 14.25 1.635 ;
        RECT 0 0 0.805 0.315 ;
        RECT 0.205 0 0.555 0.335 ;
        RECT 0 8.58 88.91 8.88 ;
        RECT 88.73 8.575 88.91 8.88 ;
        RECT 71.51 8.575 86.78 8.88 ;
        RECT 75.745 7.18 82.945 8.88 ;
        RECT 75.475 6.91 82.835 7.39 ;
        RECT 73.465 6.285 73.755 6.515 ;
        RECT 73.065 6.315 73.755 6.485 ;
        RECT 73.065 6.315 73.235 8.88 ;
        RECT 54.29 8.575 69.56 8.88 ;
        RECT 58.525 7.18 65.725 8.88 ;
        RECT 58.255 6.91 65.615 7.39 ;
        RECT 56.245 6.285 56.535 6.515 ;
        RECT 55.845 6.315 56.535 6.485 ;
        RECT 55.845 6.315 56.015 8.88 ;
        RECT 37.07 8.575 52.34 8.88 ;
        RECT 41.305 7.18 48.505 8.88 ;
        RECT 41.035 6.91 48.395 7.39 ;
        RECT 39.025 6.285 39.315 6.515 ;
        RECT 38.625 6.315 39.315 6.485 ;
        RECT 38.625 6.315 38.795 8.88 ;
        RECT 19.85 8.575 35.12 8.88 ;
        RECT 24.085 7.18 31.285 8.88 ;
        RECT 23.815 6.91 31.175 7.39 ;
        RECT 21.805 6.285 22.095 6.515 ;
        RECT 21.405 6.315 22.095 6.485 ;
        RECT 21.405 6.315 21.575 8.88 ;
        RECT 0 8.575 17.9 8.88 ;
        RECT 6.865 7.18 14.065 8.88 ;
        RECT 6.595 6.91 13.955 7.39 ;
        RECT 4.585 6.285 4.875 6.515 ;
        RECT 4.185 6.315 4.875 6.485 ;
        RECT 4.185 6.315 4.355 8.88 ;
        RECT 0.015 8.565 0.82 8.88 ;
        RECT 0.22 8.545 0.57 8.88 ;
        RECT 77.865 5.83 78.185 6.09 ;
        RECT 75.5 5.89 78.185 6.03 ;
        RECT 75.5 5.845 75.79 6.075 ;
        RECT 60.645 5.83 60.965 6.09 ;
        RECT 58.28 5.89 60.965 6.03 ;
        RECT 58.28 5.845 58.57 6.075 ;
        RECT 43.425 5.83 43.745 6.09 ;
        RECT 41.06 5.89 43.745 6.03 ;
        RECT 41.06 5.845 41.35 6.075 ;
        RECT 26.205 5.83 26.525 6.09 ;
        RECT 23.84 5.89 26.525 6.03 ;
        RECT 23.84 5.845 24.13 6.075 ;
        RECT 8.985 5.83 9.305 6.09 ;
        RECT 6.62 5.89 9.305 6.03 ;
        RECT 6.62 5.845 6.91 6.075 ;
      LAYER via2 ;
        RECT 0.28 0.09 0.48 0.29 ;
        RECT 0.295 8.59 0.495 8.79 ;
        RECT 9.045 5.855 9.245 6.055 ;
        RECT 26.265 5.855 26.465 6.055 ;
        RECT 43.485 5.855 43.685 6.055 ;
        RECT 60.705 5.855 60.905 6.055 ;
        RECT 77.925 5.855 78.125 6.055 ;
      LAYER mcon ;
        RECT 0.31 8.605 0.48 8.775 ;
        RECT 0.99 8.605 1.16 8.775 ;
        RECT 1.67 8.605 1.84 8.775 ;
        RECT 2.35 8.605 2.52 8.775 ;
        RECT 3.72 8.605 3.89 8.775 ;
        RECT 4.4 8.605 4.57 8.775 ;
        RECT 4.645 6.315 4.815 6.485 ;
        RECT 5.08 8.605 5.25 8.775 ;
        RECT 5.76 8.605 5.93 8.775 ;
        RECT 6.68 5.875 6.85 6.045 ;
        RECT 6.74 7.065 6.91 7.235 ;
        RECT 6.74 1.625 6.91 1.795 ;
        RECT 7.2 7.065 7.37 7.235 ;
        RECT 7.2 1.625 7.37 1.795 ;
        RECT 7.66 7.065 7.83 7.235 ;
        RECT 7.66 1.625 7.83 1.795 ;
        RECT 8.12 7.065 8.29 7.235 ;
        RECT 8.12 1.625 8.29 1.795 ;
        RECT 8.58 7.065 8.75 7.235 ;
        RECT 8.58 1.625 8.75 1.795 ;
        RECT 9.04 7.065 9.21 7.235 ;
        RECT 9.04 1.625 9.21 1.795 ;
        RECT 9.06 5.875 9.23 6.045 ;
        RECT 9.5 7.065 9.67 7.235 ;
        RECT 9.5 1.625 9.67 1.795 ;
        RECT 9.96 7.065 10.13 7.235 ;
        RECT 9.96 1.625 10.13 1.795 ;
        RECT 10.42 7.065 10.59 7.235 ;
        RECT 10.42 1.625 10.59 1.795 ;
        RECT 10.88 7.065 11.05 7.235 ;
        RECT 10.88 1.625 11.05 1.795 ;
        RECT 11.34 7.065 11.51 7.235 ;
        RECT 11.34 1.625 11.51 1.795 ;
        RECT 11.8 7.065 11.97 7.235 ;
        RECT 11.8 1.625 11.97 1.795 ;
        RECT 12.26 7.065 12.43 7.235 ;
        RECT 12.26 1.625 12.43 1.795 ;
        RECT 12.72 7.065 12.89 7.235 ;
        RECT 12.72 1.625 12.89 1.795 ;
        RECT 13.18 7.065 13.35 7.235 ;
        RECT 13.18 1.625 13.35 1.795 ;
        RECT 13.64 7.065 13.81 7.235 ;
        RECT 13.64 1.625 13.81 1.795 ;
        RECT 15.405 8.605 15.575 8.775 ;
        RECT 15.405 0.105 15.575 0.275 ;
        RECT 16.085 8.605 16.255 8.775 ;
        RECT 16.085 0.105 16.255 0.275 ;
        RECT 16.765 8.605 16.935 8.775 ;
        RECT 16.765 0.105 16.935 0.275 ;
        RECT 17.445 8.605 17.615 8.775 ;
        RECT 17.445 0.105 17.615 0.275 ;
        RECT 18.145 8.61 18.315 8.78 ;
        RECT 18.145 0.1 18.315 0.27 ;
        RECT 19.135 8.61 19.305 8.78 ;
        RECT 19.135 0.1 19.305 0.27 ;
        RECT 20.94 8.605 21.11 8.775 ;
        RECT 21.62 8.605 21.79 8.775 ;
        RECT 21.865 6.315 22.035 6.485 ;
        RECT 22.3 8.605 22.47 8.775 ;
        RECT 22.98 8.605 23.15 8.775 ;
        RECT 23.9 5.875 24.07 6.045 ;
        RECT 23.96 7.065 24.13 7.235 ;
        RECT 23.96 1.625 24.13 1.795 ;
        RECT 24.42 7.065 24.59 7.235 ;
        RECT 24.42 1.625 24.59 1.795 ;
        RECT 24.88 7.065 25.05 7.235 ;
        RECT 24.88 1.625 25.05 1.795 ;
        RECT 25.34 7.065 25.51 7.235 ;
        RECT 25.34 1.625 25.51 1.795 ;
        RECT 25.8 7.065 25.97 7.235 ;
        RECT 25.8 1.625 25.97 1.795 ;
        RECT 26.26 7.065 26.43 7.235 ;
        RECT 26.26 1.625 26.43 1.795 ;
        RECT 26.28 5.875 26.45 6.045 ;
        RECT 26.72 7.065 26.89 7.235 ;
        RECT 26.72 1.625 26.89 1.795 ;
        RECT 27.18 7.065 27.35 7.235 ;
        RECT 27.18 1.625 27.35 1.795 ;
        RECT 27.64 7.065 27.81 7.235 ;
        RECT 27.64 1.625 27.81 1.795 ;
        RECT 28.1 7.065 28.27 7.235 ;
        RECT 28.1 1.625 28.27 1.795 ;
        RECT 28.56 7.065 28.73 7.235 ;
        RECT 28.56 1.625 28.73 1.795 ;
        RECT 29.02 7.065 29.19 7.235 ;
        RECT 29.02 1.625 29.19 1.795 ;
        RECT 29.48 7.065 29.65 7.235 ;
        RECT 29.48 1.625 29.65 1.795 ;
        RECT 29.94 7.065 30.11 7.235 ;
        RECT 29.94 1.625 30.11 1.795 ;
        RECT 30.4 7.065 30.57 7.235 ;
        RECT 30.4 1.625 30.57 1.795 ;
        RECT 30.86 7.065 31.03 7.235 ;
        RECT 30.86 1.625 31.03 1.795 ;
        RECT 32.625 8.605 32.795 8.775 ;
        RECT 32.625 0.105 32.795 0.275 ;
        RECT 33.305 8.605 33.475 8.775 ;
        RECT 33.305 0.105 33.475 0.275 ;
        RECT 33.985 8.605 34.155 8.775 ;
        RECT 33.985 0.105 34.155 0.275 ;
        RECT 34.665 8.605 34.835 8.775 ;
        RECT 34.665 0.105 34.835 0.275 ;
        RECT 35.365 8.61 35.535 8.78 ;
        RECT 35.365 0.1 35.535 0.27 ;
        RECT 36.355 8.61 36.525 8.78 ;
        RECT 36.355 0.1 36.525 0.27 ;
        RECT 38.16 8.605 38.33 8.775 ;
        RECT 38.84 8.605 39.01 8.775 ;
        RECT 39.085 6.315 39.255 6.485 ;
        RECT 39.52 8.605 39.69 8.775 ;
        RECT 40.2 8.605 40.37 8.775 ;
        RECT 41.12 5.875 41.29 6.045 ;
        RECT 41.18 7.065 41.35 7.235 ;
        RECT 41.18 1.625 41.35 1.795 ;
        RECT 41.64 7.065 41.81 7.235 ;
        RECT 41.64 1.625 41.81 1.795 ;
        RECT 42.1 7.065 42.27 7.235 ;
        RECT 42.1 1.625 42.27 1.795 ;
        RECT 42.56 7.065 42.73 7.235 ;
        RECT 42.56 1.625 42.73 1.795 ;
        RECT 43.02 7.065 43.19 7.235 ;
        RECT 43.02 1.625 43.19 1.795 ;
        RECT 43.48 7.065 43.65 7.235 ;
        RECT 43.48 1.625 43.65 1.795 ;
        RECT 43.5 5.875 43.67 6.045 ;
        RECT 43.94 7.065 44.11 7.235 ;
        RECT 43.94 1.625 44.11 1.795 ;
        RECT 44.4 7.065 44.57 7.235 ;
        RECT 44.4 1.625 44.57 1.795 ;
        RECT 44.86 7.065 45.03 7.235 ;
        RECT 44.86 1.625 45.03 1.795 ;
        RECT 45.32 7.065 45.49 7.235 ;
        RECT 45.32 1.625 45.49 1.795 ;
        RECT 45.78 7.065 45.95 7.235 ;
        RECT 45.78 1.625 45.95 1.795 ;
        RECT 46.24 7.065 46.41 7.235 ;
        RECT 46.24 1.625 46.41 1.795 ;
        RECT 46.7 7.065 46.87 7.235 ;
        RECT 46.7 1.625 46.87 1.795 ;
        RECT 47.16 7.065 47.33 7.235 ;
        RECT 47.16 1.625 47.33 1.795 ;
        RECT 47.62 7.065 47.79 7.235 ;
        RECT 47.62 1.625 47.79 1.795 ;
        RECT 48.08 7.065 48.25 7.235 ;
        RECT 48.08 1.625 48.25 1.795 ;
        RECT 49.845 8.605 50.015 8.775 ;
        RECT 49.845 0.105 50.015 0.275 ;
        RECT 50.525 8.605 50.695 8.775 ;
        RECT 50.525 0.105 50.695 0.275 ;
        RECT 51.205 8.605 51.375 8.775 ;
        RECT 51.205 0.105 51.375 0.275 ;
        RECT 51.885 8.605 52.055 8.775 ;
        RECT 51.885 0.105 52.055 0.275 ;
        RECT 52.585 8.61 52.755 8.78 ;
        RECT 52.585 0.1 52.755 0.27 ;
        RECT 53.575 8.61 53.745 8.78 ;
        RECT 53.575 0.1 53.745 0.27 ;
        RECT 55.38 8.605 55.55 8.775 ;
        RECT 56.06 8.605 56.23 8.775 ;
        RECT 56.305 6.315 56.475 6.485 ;
        RECT 56.74 8.605 56.91 8.775 ;
        RECT 57.42 8.605 57.59 8.775 ;
        RECT 58.34 5.875 58.51 6.045 ;
        RECT 58.4 7.065 58.57 7.235 ;
        RECT 58.4 1.625 58.57 1.795 ;
        RECT 58.86 7.065 59.03 7.235 ;
        RECT 58.86 1.625 59.03 1.795 ;
        RECT 59.32 7.065 59.49 7.235 ;
        RECT 59.32 1.625 59.49 1.795 ;
        RECT 59.78 7.065 59.95 7.235 ;
        RECT 59.78 1.625 59.95 1.795 ;
        RECT 60.24 7.065 60.41 7.235 ;
        RECT 60.24 1.625 60.41 1.795 ;
        RECT 60.7 7.065 60.87 7.235 ;
        RECT 60.7 1.625 60.87 1.795 ;
        RECT 60.72 5.875 60.89 6.045 ;
        RECT 61.16 7.065 61.33 7.235 ;
        RECT 61.16 1.625 61.33 1.795 ;
        RECT 61.62 7.065 61.79 7.235 ;
        RECT 61.62 1.625 61.79 1.795 ;
        RECT 62.08 7.065 62.25 7.235 ;
        RECT 62.08 1.625 62.25 1.795 ;
        RECT 62.54 7.065 62.71 7.235 ;
        RECT 62.54 1.625 62.71 1.795 ;
        RECT 63 7.065 63.17 7.235 ;
        RECT 63 1.625 63.17 1.795 ;
        RECT 63.46 7.065 63.63 7.235 ;
        RECT 63.46 1.625 63.63 1.795 ;
        RECT 63.92 7.065 64.09 7.235 ;
        RECT 63.92 1.625 64.09 1.795 ;
        RECT 64.38 7.065 64.55 7.235 ;
        RECT 64.38 1.625 64.55 1.795 ;
        RECT 64.84 7.065 65.01 7.235 ;
        RECT 64.84 1.625 65.01 1.795 ;
        RECT 65.3 7.065 65.47 7.235 ;
        RECT 65.3 1.625 65.47 1.795 ;
        RECT 67.065 8.605 67.235 8.775 ;
        RECT 67.065 0.105 67.235 0.275 ;
        RECT 67.745 8.605 67.915 8.775 ;
        RECT 67.745 0.105 67.915 0.275 ;
        RECT 68.425 8.605 68.595 8.775 ;
        RECT 68.425 0.105 68.595 0.275 ;
        RECT 69.105 8.605 69.275 8.775 ;
        RECT 69.105 0.105 69.275 0.275 ;
        RECT 69.805 8.61 69.975 8.78 ;
        RECT 69.805 0.1 69.975 0.27 ;
        RECT 70.795 8.61 70.965 8.78 ;
        RECT 70.795 0.1 70.965 0.27 ;
        RECT 72.6 8.605 72.77 8.775 ;
        RECT 73.28 8.605 73.45 8.775 ;
        RECT 73.525 6.315 73.695 6.485 ;
        RECT 73.96 8.605 74.13 8.775 ;
        RECT 74.64 8.605 74.81 8.775 ;
        RECT 75.56 5.875 75.73 6.045 ;
        RECT 75.62 7.065 75.79 7.235 ;
        RECT 75.62 1.625 75.79 1.795 ;
        RECT 76.08 7.065 76.25 7.235 ;
        RECT 76.08 1.625 76.25 1.795 ;
        RECT 76.54 7.065 76.71 7.235 ;
        RECT 76.54 1.625 76.71 1.795 ;
        RECT 77 7.065 77.17 7.235 ;
        RECT 77 1.625 77.17 1.795 ;
        RECT 77.46 7.065 77.63 7.235 ;
        RECT 77.46 1.625 77.63 1.795 ;
        RECT 77.92 7.065 78.09 7.235 ;
        RECT 77.92 1.625 78.09 1.795 ;
        RECT 77.94 5.875 78.11 6.045 ;
        RECT 78.38 7.065 78.55 7.235 ;
        RECT 78.38 1.625 78.55 1.795 ;
        RECT 78.84 7.065 79.01 7.235 ;
        RECT 78.84 1.625 79.01 1.795 ;
        RECT 79.3 7.065 79.47 7.235 ;
        RECT 79.3 1.625 79.47 1.795 ;
        RECT 79.76 7.065 79.93 7.235 ;
        RECT 79.76 1.625 79.93 1.795 ;
        RECT 80.22 7.065 80.39 7.235 ;
        RECT 80.22 1.625 80.39 1.795 ;
        RECT 80.68 7.065 80.85 7.235 ;
        RECT 80.68 1.625 80.85 1.795 ;
        RECT 81.14 7.065 81.31 7.235 ;
        RECT 81.14 1.625 81.31 1.795 ;
        RECT 81.6 7.065 81.77 7.235 ;
        RECT 81.6 1.625 81.77 1.795 ;
        RECT 82.06 7.065 82.23 7.235 ;
        RECT 82.06 1.625 82.23 1.795 ;
        RECT 82.52 7.065 82.69 7.235 ;
        RECT 82.52 1.625 82.69 1.795 ;
        RECT 84.285 8.605 84.455 8.775 ;
        RECT 84.285 0.105 84.455 0.275 ;
        RECT 84.965 8.605 85.135 8.775 ;
        RECT 84.965 0.105 85.135 0.275 ;
        RECT 85.645 8.605 85.815 8.775 ;
        RECT 85.645 0.105 85.815 0.275 ;
        RECT 86.325 8.605 86.495 8.775 ;
        RECT 86.325 0.105 86.495 0.275 ;
        RECT 87.025 8.61 87.195 8.78 ;
        RECT 87.025 0.1 87.195 0.27 ;
        RECT 88.015 8.61 88.185 8.78 ;
        RECT 88.015 0.1 88.185 0.27 ;
      LAYER via1 ;
        RECT 0.305 0.115 0.455 0.265 ;
        RECT 0.32 8.615 0.47 8.765 ;
        RECT 9.07 5.885 9.22 6.035 ;
        RECT 26.29 5.885 26.44 6.035 ;
        RECT 43.51 5.885 43.66 6.035 ;
        RECT 60.73 5.885 60.88 6.035 ;
        RECT 77.95 5.885 78.1 6.035 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 74.94 7.435 80.955 7.735 ;
      RECT 80.655 5.805 80.955 7.735 ;
      RECT 79.6 5.785 79.9 7.735 ;
      RECT 78.57 6.48 78.87 7.735 ;
      RECT 74.94 7.035 75.24 7.735 ;
      RECT 73.805 7 74.175 7.37 ;
      RECT 73.805 7.035 75.24 7.335 ;
      RECT 78.54 6.48 78.87 6.81 ;
      RECT 78.07 6.495 78.87 6.795 ;
      RECT 78.45 6.455 78.75 6.795 ;
      RECT 80.58 5.805 80.955 6.17 ;
      RECT 80.645 5.765 80.945 6.17 ;
      RECT 79.56 5.785 79.9 6.135 ;
      RECT 79.575 5.745 79.875 6.135 ;
      RECT 79.55 5.79 79.9 6.12 ;
      RECT 80.58 5.805 81.39 6.105 ;
      RECT 79.08 5.805 79.9 6.105 ;
      RECT 80.59 5.79 80.945 6.17 ;
      RECT 80.24 3.755 80.57 4.085 ;
      RECT 80.24 3.77 81.04 4.07 ;
      RECT 80.255 3.725 80.555 4.085 ;
      RECT 79.9 3.075 80.23 3.405 ;
      RECT 79.9 3.09 80.7 3.39 ;
      RECT 79.985 3.065 80.285 3.39 ;
      RECT 79.22 4.155 79.55 4.485 ;
      RECT 77.18 4.155 77.51 4.485 ;
      RECT 77.18 4.17 79.55 4.47 ;
      RECT 78.87 3.415 79.2 3.745 ;
      RECT 78.41 3.43 79.21 3.73 ;
      RECT 78.54 2.225 78.87 2.555 ;
      RECT 78.07 2.24 78.87 2.54 ;
      RECT 78.53 2.235 78.87 2.54 ;
      RECT 57.72 7.435 63.735 7.735 ;
      RECT 63.435 5.805 63.735 7.735 ;
      RECT 62.38 5.785 62.68 7.735 ;
      RECT 61.35 6.48 61.65 7.735 ;
      RECT 57.72 7.035 58.02 7.735 ;
      RECT 56.585 7 56.955 7.37 ;
      RECT 56.585 7.035 58.02 7.335 ;
      RECT 61.32 6.48 61.65 6.81 ;
      RECT 60.85 6.495 61.65 6.795 ;
      RECT 61.23 6.455 61.53 6.795 ;
      RECT 63.36 5.805 63.735 6.17 ;
      RECT 63.425 5.765 63.725 6.17 ;
      RECT 62.34 5.785 62.68 6.135 ;
      RECT 62.355 5.745 62.655 6.135 ;
      RECT 62.33 5.79 62.68 6.12 ;
      RECT 63.36 5.805 64.17 6.105 ;
      RECT 61.86 5.805 62.68 6.105 ;
      RECT 63.37 5.79 63.725 6.17 ;
      RECT 63.02 3.755 63.35 4.085 ;
      RECT 63.02 3.77 63.82 4.07 ;
      RECT 63.035 3.725 63.335 4.085 ;
      RECT 62.68 3.075 63.01 3.405 ;
      RECT 62.68 3.09 63.48 3.39 ;
      RECT 62.765 3.065 63.065 3.39 ;
      RECT 62 4.155 62.33 4.485 ;
      RECT 59.96 4.155 60.29 4.485 ;
      RECT 59.96 4.17 62.33 4.47 ;
      RECT 61.65 3.415 61.98 3.745 ;
      RECT 61.19 3.43 61.99 3.73 ;
      RECT 61.32 2.225 61.65 2.555 ;
      RECT 60.85 2.24 61.65 2.54 ;
      RECT 61.31 2.235 61.65 2.54 ;
      RECT 40.5 7.435 46.515 7.735 ;
      RECT 46.215 5.805 46.515 7.735 ;
      RECT 45.16 5.785 45.46 7.735 ;
      RECT 44.13 6.48 44.43 7.735 ;
      RECT 40.5 7.035 40.8 7.735 ;
      RECT 39.365 7 39.735 7.37 ;
      RECT 39.365 7.035 40.8 7.335 ;
      RECT 44.1 6.48 44.43 6.81 ;
      RECT 43.63 6.495 44.43 6.795 ;
      RECT 44.01 6.455 44.31 6.795 ;
      RECT 46.14 5.805 46.515 6.17 ;
      RECT 46.205 5.765 46.505 6.17 ;
      RECT 45.12 5.785 45.46 6.135 ;
      RECT 45.135 5.745 45.435 6.135 ;
      RECT 45.11 5.79 45.46 6.12 ;
      RECT 46.14 5.805 46.95 6.105 ;
      RECT 44.64 5.805 45.46 6.105 ;
      RECT 46.15 5.79 46.505 6.17 ;
      RECT 45.8 3.755 46.13 4.085 ;
      RECT 45.8 3.77 46.6 4.07 ;
      RECT 45.815 3.725 46.115 4.085 ;
      RECT 45.46 3.075 45.79 3.405 ;
      RECT 45.46 3.09 46.26 3.39 ;
      RECT 45.545 3.065 45.845 3.39 ;
      RECT 44.78 4.155 45.11 4.485 ;
      RECT 42.74 4.155 43.07 4.485 ;
      RECT 42.74 4.17 45.11 4.47 ;
      RECT 44.43 3.415 44.76 3.745 ;
      RECT 43.97 3.43 44.77 3.73 ;
      RECT 44.1 2.225 44.43 2.555 ;
      RECT 43.63 2.24 44.43 2.54 ;
      RECT 44.09 2.235 44.43 2.54 ;
      RECT 23.28 7.435 29.295 7.735 ;
      RECT 28.995 5.805 29.295 7.735 ;
      RECT 27.94 5.785 28.24 7.735 ;
      RECT 26.91 6.48 27.21 7.735 ;
      RECT 23.28 7.035 23.58 7.735 ;
      RECT 22.145 7 22.515 7.37 ;
      RECT 22.145 7.035 23.58 7.335 ;
      RECT 26.88 6.48 27.21 6.81 ;
      RECT 26.41 6.495 27.21 6.795 ;
      RECT 26.79 6.455 27.09 6.795 ;
      RECT 28.92 5.805 29.295 6.17 ;
      RECT 28.985 5.765 29.285 6.17 ;
      RECT 27.9 5.785 28.24 6.135 ;
      RECT 27.915 5.745 28.215 6.135 ;
      RECT 27.89 5.79 28.24 6.12 ;
      RECT 28.92 5.805 29.73 6.105 ;
      RECT 27.42 5.805 28.24 6.105 ;
      RECT 28.93 5.79 29.285 6.17 ;
      RECT 28.58 3.755 28.91 4.085 ;
      RECT 28.58 3.77 29.38 4.07 ;
      RECT 28.595 3.725 28.895 4.085 ;
      RECT 28.24 3.075 28.57 3.405 ;
      RECT 28.24 3.09 29.04 3.39 ;
      RECT 28.325 3.065 28.625 3.39 ;
      RECT 27.56 4.155 27.89 4.485 ;
      RECT 25.52 4.155 25.85 4.485 ;
      RECT 25.52 4.17 27.89 4.47 ;
      RECT 27.21 3.415 27.54 3.745 ;
      RECT 26.75 3.43 27.55 3.73 ;
      RECT 26.88 2.225 27.21 2.555 ;
      RECT 26.41 2.24 27.21 2.54 ;
      RECT 26.87 2.235 27.21 2.54 ;
      RECT 6.06 7.435 12.075 7.735 ;
      RECT 11.775 5.805 12.075 7.735 ;
      RECT 10.72 5.785 11.02 7.735 ;
      RECT 9.69 6.48 9.99 7.735 ;
      RECT 6.06 7.035 6.36 7.735 ;
      RECT 4.925 7 5.295 7.37 ;
      RECT 4.925 7.035 6.36 7.335 ;
      RECT 9.66 6.48 9.99 6.81 ;
      RECT 9.19 6.495 9.99 6.795 ;
      RECT 9.57 6.455 9.87 6.795 ;
      RECT 11.7 5.805 12.075 6.17 ;
      RECT 11.765 5.765 12.065 6.17 ;
      RECT 10.68 5.785 11.02 6.135 ;
      RECT 10.695 5.745 10.995 6.135 ;
      RECT 10.67 5.79 11.02 6.12 ;
      RECT 11.7 5.805 12.51 6.105 ;
      RECT 10.2 5.805 11.02 6.105 ;
      RECT 11.71 5.79 12.065 6.17 ;
      RECT 11.36 3.755 11.69 4.085 ;
      RECT 11.36 3.77 12.16 4.07 ;
      RECT 11.375 3.725 11.675 4.085 ;
      RECT 11.02 3.075 11.35 3.405 ;
      RECT 11.02 3.09 11.82 3.39 ;
      RECT 11.105 3.065 11.405 3.39 ;
      RECT 10.34 4.155 10.67 4.485 ;
      RECT 8.3 4.155 8.63 4.485 ;
      RECT 8.3 4.17 10.67 4.47 ;
      RECT 9.99 3.415 10.32 3.745 ;
      RECT 9.53 3.43 10.33 3.73 ;
      RECT 9.66 2.225 9.99 2.555 ;
      RECT 9.19 2.24 9.99 2.54 ;
      RECT 9.65 2.235 9.99 2.54 ;
    LAYER via2 ;
      RECT 80.655 5.855 80.855 6.055 ;
      RECT 80.305 3.82 80.505 4.02 ;
      RECT 79.965 3.14 80.165 3.34 ;
      RECT 79.615 5.855 79.815 6.055 ;
      RECT 79.285 4.22 79.485 4.42 ;
      RECT 78.935 3.48 79.135 3.68 ;
      RECT 78.605 2.29 78.805 2.49 ;
      RECT 78.605 6.545 78.805 6.745 ;
      RECT 77.245 4.22 77.445 4.42 ;
      RECT 73.89 7.085 74.09 7.285 ;
      RECT 63.435 5.855 63.635 6.055 ;
      RECT 63.085 3.82 63.285 4.02 ;
      RECT 62.745 3.14 62.945 3.34 ;
      RECT 62.395 5.855 62.595 6.055 ;
      RECT 62.065 4.22 62.265 4.42 ;
      RECT 61.715 3.48 61.915 3.68 ;
      RECT 61.385 2.29 61.585 2.49 ;
      RECT 61.385 6.545 61.585 6.745 ;
      RECT 60.025 4.22 60.225 4.42 ;
      RECT 56.67 7.085 56.87 7.285 ;
      RECT 46.215 5.855 46.415 6.055 ;
      RECT 45.865 3.82 46.065 4.02 ;
      RECT 45.525 3.14 45.725 3.34 ;
      RECT 45.175 5.855 45.375 6.055 ;
      RECT 44.845 4.22 45.045 4.42 ;
      RECT 44.495 3.48 44.695 3.68 ;
      RECT 44.165 2.29 44.365 2.49 ;
      RECT 44.165 6.545 44.365 6.745 ;
      RECT 42.805 4.22 43.005 4.42 ;
      RECT 39.45 7.085 39.65 7.285 ;
      RECT 28.995 5.855 29.195 6.055 ;
      RECT 28.645 3.82 28.845 4.02 ;
      RECT 28.305 3.14 28.505 3.34 ;
      RECT 27.955 5.855 28.155 6.055 ;
      RECT 27.625 4.22 27.825 4.42 ;
      RECT 27.275 3.48 27.475 3.68 ;
      RECT 26.945 2.29 27.145 2.49 ;
      RECT 26.945 6.545 27.145 6.745 ;
      RECT 25.585 4.22 25.785 4.42 ;
      RECT 22.23 7.085 22.43 7.285 ;
      RECT 11.775 5.855 11.975 6.055 ;
      RECT 11.425 3.82 11.625 4.02 ;
      RECT 11.085 3.14 11.285 3.34 ;
      RECT 10.735 5.855 10.935 6.055 ;
      RECT 10.405 4.22 10.605 4.42 ;
      RECT 10.055 3.48 10.255 3.68 ;
      RECT 9.725 2.29 9.925 2.49 ;
      RECT 9.725 6.545 9.925 6.745 ;
      RECT 8.365 4.22 8.565 4.42 ;
      RECT 5.01 7.085 5.21 7.285 ;
    LAYER met2 ;
      RECT 1.23 8.6 88.54 8.77 ;
      RECT 88.37 7.3 88.54 8.77 ;
      RECT 1.23 6.255 1.4 8.77 ;
      RECT 88.335 7.3 88.66 7.625 ;
      RECT 1.175 6.255 1.455 6.595 ;
      RECT 85.18 6.28 85.5 6.605 ;
      RECT 85.21 5.695 85.38 6.605 ;
      RECT 85.21 5.695 85.385 6.045 ;
      RECT 85.21 5.695 86.185 5.87 ;
      RECT 86.01 1.965 86.185 5.87 ;
      RECT 79.925 3.055 80.205 3.425 ;
      RECT 79.995 2.345 80.17 3.425 ;
      RECT 79.995 2.345 83.215 2.52 ;
      RECT 83.04 2.025 83.215 2.52 ;
      RECT 83.51 1.995 83.835 2.32 ;
      RECT 85.955 1.965 86.305 2.315 ;
      RECT 83.04 2.025 86.305 2.195 ;
      RECT 74.33 8.29 85.025 8.46 ;
      RECT 84.865 2.395 85.025 8.46 ;
      RECT 74.33 6.545 74.5 8.46 ;
      RECT 85.98 6.655 86.305 6.98 ;
      RECT 71.15 6.655 71.475 6.98 ;
      RECT 84.865 6.745 86.305 6.915 ;
      RECT 74.28 6.545 74.56 6.885 ;
      RECT 71.15 6.685 74.56 6.855 ;
      RECT 85.18 2.365 85.5 2.685 ;
      RECT 84.865 2.395 85.5 2.565 ;
      RECT 81.635 6.48 81.895 6.8 ;
      RECT 81.695 2.74 81.835 6.8 ;
      RECT 81.635 2.74 81.895 3.06 ;
      RECT 80.955 4.78 81.215 5.1 ;
      RECT 81.015 3.76 81.155 5.1 ;
      RECT 80.955 3.76 81.215 4.08 ;
      RECT 79.935 6.48 80.195 6.8 ;
      RECT 79.995 5.21 80.135 6.8 ;
      RECT 79.315 5.21 80.135 5.35 ;
      RECT 79.315 2.74 79.455 5.35 ;
      RECT 79.245 4.135 79.525 4.505 ;
      RECT 79.255 2.74 79.515 3.06 ;
      RECT 77.205 4.135 77.485 4.505 ;
      RECT 77.275 2.4 77.415 4.505 ;
      RECT 77.215 2.4 77.475 2.72 ;
      RECT 76.535 4.78 76.795 5.1 ;
      RECT 76.595 2.74 76.735 5.1 ;
      RECT 76.535 2.74 76.795 3.06 ;
      RECT 67.96 6.28 68.28 6.605 ;
      RECT 67.99 5.695 68.16 6.605 ;
      RECT 67.99 5.695 68.165 6.045 ;
      RECT 67.99 5.695 68.965 5.87 ;
      RECT 68.79 1.965 68.965 5.87 ;
      RECT 62.705 3.055 62.985 3.425 ;
      RECT 62.775 2.345 62.95 3.425 ;
      RECT 62.775 2.345 65.995 2.52 ;
      RECT 65.82 2.025 65.995 2.52 ;
      RECT 66.29 1.995 66.615 2.32 ;
      RECT 68.735 1.965 69.085 2.315 ;
      RECT 65.82 2.025 69.085 2.195 ;
      RECT 57.11 8.29 67.805 8.46 ;
      RECT 67.645 2.395 67.805 8.46 ;
      RECT 57.11 6.545 57.28 8.46 ;
      RECT 68.76 6.655 69.085 6.98 ;
      RECT 53.93 6.655 54.255 6.98 ;
      RECT 67.645 6.745 69.085 6.915 ;
      RECT 57.06 6.545 57.34 6.885 ;
      RECT 53.93 6.685 57.34 6.855 ;
      RECT 67.96 2.365 68.28 2.685 ;
      RECT 67.645 2.395 68.28 2.565 ;
      RECT 64.415 6.48 64.675 6.8 ;
      RECT 64.475 2.74 64.615 6.8 ;
      RECT 64.415 2.74 64.675 3.06 ;
      RECT 63.735 4.78 63.995 5.1 ;
      RECT 63.795 3.76 63.935 5.1 ;
      RECT 63.735 3.76 63.995 4.08 ;
      RECT 62.715 6.48 62.975 6.8 ;
      RECT 62.775 5.21 62.915 6.8 ;
      RECT 62.095 5.21 62.915 5.35 ;
      RECT 62.095 2.74 62.235 5.35 ;
      RECT 62.025 4.135 62.305 4.505 ;
      RECT 62.035 2.74 62.295 3.06 ;
      RECT 59.985 4.135 60.265 4.505 ;
      RECT 60.055 2.4 60.195 4.505 ;
      RECT 59.995 2.4 60.255 2.72 ;
      RECT 59.315 4.78 59.575 5.1 ;
      RECT 59.375 2.74 59.515 5.1 ;
      RECT 59.315 2.74 59.575 3.06 ;
      RECT 50.74 6.28 51.06 6.605 ;
      RECT 50.77 5.695 50.94 6.605 ;
      RECT 50.77 5.695 50.945 6.045 ;
      RECT 50.77 5.695 51.745 5.87 ;
      RECT 51.57 1.965 51.745 5.87 ;
      RECT 45.485 3.055 45.765 3.425 ;
      RECT 45.555 2.345 45.73 3.425 ;
      RECT 45.555 2.345 48.775 2.52 ;
      RECT 48.6 2.025 48.775 2.52 ;
      RECT 49.07 1.995 49.395 2.32 ;
      RECT 51.515 1.965 51.865 2.315 ;
      RECT 48.6 2.025 51.865 2.195 ;
      RECT 39.89 8.29 50.585 8.46 ;
      RECT 50.425 2.395 50.585 8.46 ;
      RECT 39.89 6.545 40.06 8.46 ;
      RECT 51.54 6.655 51.865 6.98 ;
      RECT 36.71 6.655 37.035 6.98 ;
      RECT 50.425 6.745 51.865 6.915 ;
      RECT 39.84 6.545 40.12 6.885 ;
      RECT 36.71 6.685 40.13 6.855 ;
      RECT 50.74 2.365 51.06 2.685 ;
      RECT 50.425 2.395 51.06 2.565 ;
      RECT 47.195 6.48 47.455 6.8 ;
      RECT 47.255 2.74 47.395 6.8 ;
      RECT 47.195 2.74 47.455 3.06 ;
      RECT 46.515 4.78 46.775 5.1 ;
      RECT 46.575 3.76 46.715 5.1 ;
      RECT 46.515 3.76 46.775 4.08 ;
      RECT 45.495 6.48 45.755 6.8 ;
      RECT 45.555 5.21 45.695 6.8 ;
      RECT 44.875 5.21 45.695 5.35 ;
      RECT 44.875 2.74 45.015 5.35 ;
      RECT 44.805 4.135 45.085 4.505 ;
      RECT 44.815 2.74 45.075 3.06 ;
      RECT 42.765 4.135 43.045 4.505 ;
      RECT 42.835 2.4 42.975 4.505 ;
      RECT 42.775 2.4 43.035 2.72 ;
      RECT 42.095 4.78 42.355 5.1 ;
      RECT 42.155 2.74 42.295 5.1 ;
      RECT 42.095 2.74 42.355 3.06 ;
      RECT 33.52 6.28 33.84 6.605 ;
      RECT 33.55 5.695 33.72 6.605 ;
      RECT 33.55 5.695 33.725 6.045 ;
      RECT 33.55 5.695 34.525 5.87 ;
      RECT 34.35 1.965 34.525 5.87 ;
      RECT 28.265 3.055 28.545 3.425 ;
      RECT 28.335 2.345 28.51 3.425 ;
      RECT 28.335 2.345 31.555 2.52 ;
      RECT 31.38 2.025 31.555 2.52 ;
      RECT 31.85 1.995 32.175 2.32 ;
      RECT 34.295 1.965 34.645 2.315 ;
      RECT 31.38 2.025 34.645 2.195 ;
      RECT 22.67 8.29 33.365 8.46 ;
      RECT 33.205 2.395 33.365 8.46 ;
      RECT 22.67 6.545 22.84 8.46 ;
      RECT 34.32 6.655 34.645 6.98 ;
      RECT 19.49 6.655 19.815 6.98 ;
      RECT 33.205 6.745 34.645 6.915 ;
      RECT 22.62 6.545 22.9 6.885 ;
      RECT 19.49 6.685 22.9 6.855 ;
      RECT 33.52 2.365 33.84 2.685 ;
      RECT 33.205 2.395 33.84 2.565 ;
      RECT 29.975 6.48 30.235 6.8 ;
      RECT 30.035 2.74 30.175 6.8 ;
      RECT 29.975 2.74 30.235 3.06 ;
      RECT 29.295 4.78 29.555 5.1 ;
      RECT 29.355 3.76 29.495 5.1 ;
      RECT 29.295 3.76 29.555 4.08 ;
      RECT 28.275 6.48 28.535 6.8 ;
      RECT 28.335 5.21 28.475 6.8 ;
      RECT 27.655 5.21 28.475 5.35 ;
      RECT 27.655 2.74 27.795 5.35 ;
      RECT 27.585 4.135 27.865 4.505 ;
      RECT 27.595 2.74 27.855 3.06 ;
      RECT 25.545 4.135 25.825 4.505 ;
      RECT 25.615 2.4 25.755 4.505 ;
      RECT 25.555 2.4 25.815 2.72 ;
      RECT 24.875 4.78 25.135 5.1 ;
      RECT 24.935 2.74 25.075 5.1 ;
      RECT 24.875 2.74 25.135 3.06 ;
      RECT 16.3 6.28 16.62 6.605 ;
      RECT 16.33 5.695 16.5 6.605 ;
      RECT 16.33 5.695 16.505 6.045 ;
      RECT 16.33 5.695 17.305 5.87 ;
      RECT 17.13 1.965 17.305 5.87 ;
      RECT 11.045 3.055 11.325 3.425 ;
      RECT 11.115 2.345 11.29 3.425 ;
      RECT 11.115 2.345 14.335 2.52 ;
      RECT 14.16 2.025 14.335 2.52 ;
      RECT 14.63 1.995 14.955 2.32 ;
      RECT 17.075 1.965 17.425 2.315 ;
      RECT 14.16 2.025 17.425 2.195 ;
      RECT 5.45 8.29 16.145 8.46 ;
      RECT 15.985 2.395 16.145 8.46 ;
      RECT 5.45 6.545 5.62 8.46 ;
      RECT 1.55 6.995 1.83 7.335 ;
      RECT 1.55 7.06 2.76 7.23 ;
      RECT 2.59 6.685 2.76 7.23 ;
      RECT 17.1 6.655 17.425 6.98 ;
      RECT 15.985 6.745 17.425 6.915 ;
      RECT 5.4 6.545 5.68 6.885 ;
      RECT 2.59 6.685 5.68 6.855 ;
      RECT 16.3 2.365 16.62 2.685 ;
      RECT 15.985 2.395 16.62 2.565 ;
      RECT 12.755 6.48 13.015 6.8 ;
      RECT 12.815 2.74 12.955 6.8 ;
      RECT 12.755 2.74 13.015 3.06 ;
      RECT 12.075 4.78 12.335 5.1 ;
      RECT 12.135 3.76 12.275 5.1 ;
      RECT 12.075 3.76 12.335 4.08 ;
      RECT 11.055 6.48 11.315 6.8 ;
      RECT 11.115 5.21 11.255 6.8 ;
      RECT 10.435 5.21 11.255 5.35 ;
      RECT 10.435 2.74 10.575 5.35 ;
      RECT 10.365 4.135 10.645 4.505 ;
      RECT 10.375 2.74 10.635 3.06 ;
      RECT 8.325 4.135 8.605 4.505 ;
      RECT 8.395 2.4 8.535 4.505 ;
      RECT 8.335 2.4 8.595 2.72 ;
      RECT 7.655 4.78 7.915 5.1 ;
      RECT 7.715 2.74 7.855 5.1 ;
      RECT 7.655 2.74 7.915 3.06 ;
      RECT 80.615 5.77 80.895 6.14 ;
      RECT 80.265 3.735 80.545 4.105 ;
      RECT 79.575 5.77 79.855 6.14 ;
      RECT 78.895 3.395 79.175 3.765 ;
      RECT 78.565 2.205 78.845 2.575 ;
      RECT 78.565 6.46 78.845 6.83 ;
      RECT 73.805 7 74.175 7.37 ;
      RECT 63.395 5.77 63.675 6.14 ;
      RECT 63.045 3.735 63.325 4.105 ;
      RECT 62.355 5.77 62.635 6.14 ;
      RECT 61.675 3.395 61.955 3.765 ;
      RECT 61.345 2.205 61.625 2.575 ;
      RECT 61.345 6.46 61.625 6.83 ;
      RECT 56.585 7 56.955 7.37 ;
      RECT 46.175 5.77 46.455 6.14 ;
      RECT 45.825 3.735 46.105 4.105 ;
      RECT 45.135 5.77 45.415 6.14 ;
      RECT 44.455 3.395 44.735 3.765 ;
      RECT 44.125 2.205 44.405 2.575 ;
      RECT 44.125 6.46 44.405 6.83 ;
      RECT 39.365 7 39.735 7.37 ;
      RECT 28.955 5.77 29.235 6.14 ;
      RECT 28.605 3.735 28.885 4.105 ;
      RECT 27.915 5.77 28.195 6.14 ;
      RECT 27.235 3.395 27.515 3.765 ;
      RECT 26.905 2.205 27.185 2.575 ;
      RECT 26.905 6.46 27.185 6.83 ;
      RECT 22.145 7 22.515 7.37 ;
      RECT 11.735 5.77 12.015 6.14 ;
      RECT 11.385 3.735 11.665 4.105 ;
      RECT 10.695 5.77 10.975 6.14 ;
      RECT 10.015 3.395 10.295 3.765 ;
      RECT 9.685 2.205 9.965 2.575 ;
      RECT 9.685 6.46 9.965 6.83 ;
      RECT 4.925 7 5.295 7.37 ;
    LAYER via1 ;
      RECT 88.425 7.385 88.575 7.535 ;
      RECT 86.07 6.74 86.22 6.89 ;
      RECT 86.055 2.065 86.205 2.215 ;
      RECT 85.265 2.45 85.415 2.6 ;
      RECT 85.265 6.37 85.415 6.52 ;
      RECT 83.6 2.08 83.75 2.23 ;
      RECT 81.69 2.825 81.84 2.975 ;
      RECT 81.69 6.565 81.84 6.715 ;
      RECT 81.01 3.845 81.16 3.995 ;
      RECT 81.01 4.865 81.16 5.015 ;
      RECT 80.67 5.885 80.82 6.035 ;
      RECT 80.33 3.845 80.48 3.995 ;
      RECT 79.99 3.165 80.14 3.315 ;
      RECT 79.99 6.565 80.14 6.715 ;
      RECT 79.64 5.885 79.79 6.035 ;
      RECT 79.31 2.825 79.46 2.975 ;
      RECT 78.97 3.505 79.12 3.655 ;
      RECT 78.63 2.315 78.78 2.465 ;
      RECT 78.63 6.565 78.78 6.715 ;
      RECT 77.27 2.485 77.42 2.635 ;
      RECT 76.59 2.825 76.74 2.975 ;
      RECT 76.59 4.865 76.74 5.015 ;
      RECT 74.345 6.64 74.495 6.79 ;
      RECT 73.915 7.11 74.065 7.26 ;
      RECT 71.24 6.74 71.39 6.89 ;
      RECT 68.85 6.74 69 6.89 ;
      RECT 68.835 2.065 68.985 2.215 ;
      RECT 68.045 2.45 68.195 2.6 ;
      RECT 68.045 6.37 68.195 6.52 ;
      RECT 66.38 2.08 66.53 2.23 ;
      RECT 64.47 2.825 64.62 2.975 ;
      RECT 64.47 6.565 64.62 6.715 ;
      RECT 63.79 3.845 63.94 3.995 ;
      RECT 63.79 4.865 63.94 5.015 ;
      RECT 63.45 5.885 63.6 6.035 ;
      RECT 63.11 3.845 63.26 3.995 ;
      RECT 62.77 3.165 62.92 3.315 ;
      RECT 62.77 6.565 62.92 6.715 ;
      RECT 62.42 5.885 62.57 6.035 ;
      RECT 62.09 2.825 62.24 2.975 ;
      RECT 61.75 3.505 61.9 3.655 ;
      RECT 61.41 2.315 61.56 2.465 ;
      RECT 61.41 6.565 61.56 6.715 ;
      RECT 60.05 2.485 60.2 2.635 ;
      RECT 59.37 2.825 59.52 2.975 ;
      RECT 59.37 4.865 59.52 5.015 ;
      RECT 57.125 6.64 57.275 6.79 ;
      RECT 56.695 7.11 56.845 7.26 ;
      RECT 54.02 6.74 54.17 6.89 ;
      RECT 51.63 6.74 51.78 6.89 ;
      RECT 51.615 2.065 51.765 2.215 ;
      RECT 50.825 2.45 50.975 2.6 ;
      RECT 50.825 6.37 50.975 6.52 ;
      RECT 49.16 2.08 49.31 2.23 ;
      RECT 47.25 2.825 47.4 2.975 ;
      RECT 47.25 6.565 47.4 6.715 ;
      RECT 46.57 3.845 46.72 3.995 ;
      RECT 46.57 4.865 46.72 5.015 ;
      RECT 46.23 5.885 46.38 6.035 ;
      RECT 45.89 3.845 46.04 3.995 ;
      RECT 45.55 3.165 45.7 3.315 ;
      RECT 45.55 6.565 45.7 6.715 ;
      RECT 45.2 5.885 45.35 6.035 ;
      RECT 44.87 2.825 45.02 2.975 ;
      RECT 44.53 3.505 44.68 3.655 ;
      RECT 44.19 2.315 44.34 2.465 ;
      RECT 44.19 6.565 44.34 6.715 ;
      RECT 42.83 2.485 42.98 2.635 ;
      RECT 42.15 2.825 42.3 2.975 ;
      RECT 42.15 4.865 42.3 5.015 ;
      RECT 39.905 6.64 40.055 6.79 ;
      RECT 39.475 7.11 39.625 7.26 ;
      RECT 36.8 6.74 36.95 6.89 ;
      RECT 34.41 6.74 34.56 6.89 ;
      RECT 34.395 2.065 34.545 2.215 ;
      RECT 33.605 2.45 33.755 2.6 ;
      RECT 33.605 6.37 33.755 6.52 ;
      RECT 31.94 2.08 32.09 2.23 ;
      RECT 30.03 2.825 30.18 2.975 ;
      RECT 30.03 6.565 30.18 6.715 ;
      RECT 29.35 3.845 29.5 3.995 ;
      RECT 29.35 4.865 29.5 5.015 ;
      RECT 29.01 5.885 29.16 6.035 ;
      RECT 28.67 3.845 28.82 3.995 ;
      RECT 28.33 3.165 28.48 3.315 ;
      RECT 28.33 6.565 28.48 6.715 ;
      RECT 27.98 5.885 28.13 6.035 ;
      RECT 27.65 2.825 27.8 2.975 ;
      RECT 27.31 3.505 27.46 3.655 ;
      RECT 26.97 2.315 27.12 2.465 ;
      RECT 26.97 6.565 27.12 6.715 ;
      RECT 25.61 2.485 25.76 2.635 ;
      RECT 24.93 2.825 25.08 2.975 ;
      RECT 24.93 4.865 25.08 5.015 ;
      RECT 22.685 6.64 22.835 6.79 ;
      RECT 22.255 7.11 22.405 7.26 ;
      RECT 19.58 6.74 19.73 6.89 ;
      RECT 17.19 6.74 17.34 6.89 ;
      RECT 17.175 2.065 17.325 2.215 ;
      RECT 16.385 2.45 16.535 2.6 ;
      RECT 16.385 6.37 16.535 6.52 ;
      RECT 14.72 2.08 14.87 2.23 ;
      RECT 12.81 2.825 12.96 2.975 ;
      RECT 12.81 6.565 12.96 6.715 ;
      RECT 12.13 3.845 12.28 3.995 ;
      RECT 12.13 4.865 12.28 5.015 ;
      RECT 11.79 5.885 11.94 6.035 ;
      RECT 11.45 3.845 11.6 3.995 ;
      RECT 11.11 3.165 11.26 3.315 ;
      RECT 11.11 6.565 11.26 6.715 ;
      RECT 10.76 5.885 10.91 6.035 ;
      RECT 10.43 2.825 10.58 2.975 ;
      RECT 10.09 3.505 10.24 3.655 ;
      RECT 9.75 2.315 9.9 2.465 ;
      RECT 9.75 6.565 9.9 6.715 ;
      RECT 8.39 2.485 8.54 2.635 ;
      RECT 7.71 2.825 7.86 2.975 ;
      RECT 7.71 4.865 7.86 5.015 ;
      RECT 5.465 6.64 5.615 6.79 ;
      RECT 5.035 7.11 5.185 7.26 ;
      RECT 1.615 7.09 1.765 7.24 ;
      RECT 1.24 6.35 1.39 6.5 ;
    LAYER met1 ;
      RECT 88.305 7.77 88.595 8 ;
      RECT 88.365 6.29 88.535 8 ;
      RECT 88.335 7.3 88.66 7.625 ;
      RECT 88.305 6.29 88.595 6.52 ;
      RECT 87.9 2.395 88.005 2.965 ;
      RECT 87.9 2.73 88.225 2.96 ;
      RECT 87.9 2.76 88.395 2.93 ;
      RECT 87.9 2.395 88.09 2.96 ;
      RECT 87.315 2.36 87.605 2.59 ;
      RECT 87.315 2.395 88.09 2.565 ;
      RECT 87.375 0.88 87.545 2.59 ;
      RECT 87.315 0.88 87.605 1.11 ;
      RECT 87.315 7.77 87.605 8 ;
      RECT 87.375 6.29 87.545 8 ;
      RECT 87.315 6.29 87.605 6.52 ;
      RECT 87.315 6.325 88.17 6.485 ;
      RECT 88 5.92 88.17 6.485 ;
      RECT 87.315 6.32 87.71 6.485 ;
      RECT 87.935 5.92 88.225 6.15 ;
      RECT 87.935 5.95 88.395 6.12 ;
      RECT 86.945 2.73 87.235 2.96 ;
      RECT 86.945 2.76 87.405 2.93 ;
      RECT 87.01 1.655 87.175 2.96 ;
      RECT 85.525 1.625 85.815 1.855 ;
      RECT 85.525 1.655 87.175 1.825 ;
      RECT 85.585 0.885 85.755 1.855 ;
      RECT 85.525 0.885 85.815 1.115 ;
      RECT 85.525 7.765 85.815 7.995 ;
      RECT 85.585 7.025 85.755 7.995 ;
      RECT 85.585 7.12 87.175 7.29 ;
      RECT 87.005 5.92 87.175 7.29 ;
      RECT 85.525 7.025 85.815 7.255 ;
      RECT 86.945 5.92 87.235 6.15 ;
      RECT 86.945 5.95 87.405 6.12 ;
      RECT 85.955 1.965 86.305 2.315 ;
      RECT 85.785 2.025 86.305 2.195 ;
      RECT 85.98 6.655 86.305 6.98 ;
      RECT 85.955 6.655 86.305 6.885 ;
      RECT 85.785 6.685 86.305 6.855 ;
      RECT 85.18 2.365 85.5 2.685 ;
      RECT 85.15 2.365 85.5 2.595 ;
      RECT 84.865 2.395 85.5 2.565 ;
      RECT 85.18 6.28 85.5 6.605 ;
      RECT 85.15 6.285 85.5 6.515 ;
      RECT 84.98 6.315 85.5 6.485 ;
      RECT 80.925 3.79 81.245 4.05 ;
      RECT 81.96 3.805 82.25 4.035 ;
      RECT 80.925 3.85 82.25 3.99 ;
      RECT 80.585 5.83 80.905 6.09 ;
      RECT 81.96 5.845 82.25 6.075 ;
      RECT 82.035 5.55 82.175 6.075 ;
      RECT 80.675 5.55 80.815 6.09 ;
      RECT 80.675 5.55 82.175 5.69 ;
      RECT 81.605 2.77 81.925 3.03 ;
      RECT 81.33 2.83 81.925 2.97 ;
      RECT 78.545 6.51 78.865 6.77 ;
      RECT 77.54 6.525 77.83 6.755 ;
      RECT 77.54 6.57 79.455 6.71 ;
      RECT 79.315 6.23 79.455 6.71 ;
      RECT 79.315 6.23 81.325 6.37 ;
      RECT 81.185 5.845 81.325 6.37 ;
      RECT 81.11 5.845 81.4 6.075 ;
      RECT 80.925 4.81 81.245 5.07 ;
      RECT 78.78 4.825 79.07 5.055 ;
      RECT 78.78 4.87 81.245 5.01 ;
      RECT 80.245 3.79 80.565 4.05 ;
      RECT 77.88 3.805 78.17 4.035 ;
      RECT 77.88 3.85 80.565 3.99 ;
      RECT 79.905 6.51 80.225 6.77 ;
      RECT 79.905 6.57 80.5 6.71 ;
      RECT 79.905 3.11 80.225 3.37 ;
      RECT 79.63 3.17 80.225 3.31 ;
      RECT 79.225 2.77 79.545 3.03 ;
      RECT 78.95 2.83 79.545 2.97 ;
      RECT 78.885 3.45 79.205 3.71 ;
      RECT 76.01 3.465 76.3 3.695 ;
      RECT 76.01 3.51 79.205 3.65 ;
      RECT 78.465 2.79 78.605 3.65 ;
      RECT 78.39 2.79 78.68 3.02 ;
      RECT 78.545 2.26 78.865 2.52 ;
      RECT 78.545 2.275 79.05 2.505 ;
      RECT 78.455 2.32 79.05 2.46 ;
      RECT 77.88 2.79 78.17 3.02 ;
      RECT 77.275 2.835 78.17 2.975 ;
      RECT 77.275 2.43 77.415 2.975 ;
      RECT 77.185 2.43 77.505 2.69 ;
      RECT 76.505 2.77 76.825 3.03 ;
      RECT 76.23 2.83 76.825 2.97 ;
      RECT 76.505 4.81 76.825 5.07 ;
      RECT 76.23 4.87 76.825 5.01 ;
      RECT 74.27 6.575 74.56 6.885 ;
      RECT 74.1 6.685 74.59 6.855 ;
      RECT 74.25 6.575 74.59 6.855 ;
      RECT 73.84 7.765 74.13 7.995 ;
      RECT 73.9 6.995 74.07 7.995 ;
      RECT 73.805 6.995 74.175 7.37 ;
      RECT 71.085 7.77 71.375 8 ;
      RECT 71.145 6.29 71.315 8 ;
      RECT 71.145 6.655 71.475 6.98 ;
      RECT 71.085 6.29 71.375 6.52 ;
      RECT 70.68 2.395 70.785 2.965 ;
      RECT 70.68 2.73 71.005 2.96 ;
      RECT 70.68 2.76 71.175 2.93 ;
      RECT 70.68 2.395 70.87 2.96 ;
      RECT 70.095 2.36 70.385 2.59 ;
      RECT 70.095 2.395 70.87 2.565 ;
      RECT 70.155 0.88 70.325 2.59 ;
      RECT 70.095 0.88 70.385 1.11 ;
      RECT 70.095 7.77 70.385 8 ;
      RECT 70.155 6.29 70.325 8 ;
      RECT 70.095 6.29 70.385 6.52 ;
      RECT 70.095 6.325 70.95 6.485 ;
      RECT 70.78 5.92 70.95 6.485 ;
      RECT 70.095 6.32 70.49 6.485 ;
      RECT 70.715 5.92 71.005 6.15 ;
      RECT 70.715 5.95 71.175 6.12 ;
      RECT 69.725 2.73 70.015 2.96 ;
      RECT 69.725 2.76 70.185 2.93 ;
      RECT 69.79 1.655 69.955 2.96 ;
      RECT 68.305 1.625 68.595 1.855 ;
      RECT 68.305 1.655 69.955 1.825 ;
      RECT 68.365 0.885 68.535 1.855 ;
      RECT 68.305 0.885 68.595 1.115 ;
      RECT 68.305 7.765 68.595 7.995 ;
      RECT 68.365 7.025 68.535 7.995 ;
      RECT 68.365 7.12 69.955 7.29 ;
      RECT 69.785 5.92 69.955 7.29 ;
      RECT 68.305 7.025 68.595 7.255 ;
      RECT 69.725 5.92 70.015 6.15 ;
      RECT 69.725 5.95 70.185 6.12 ;
      RECT 68.735 1.965 69.085 2.315 ;
      RECT 68.565 2.025 69.085 2.195 ;
      RECT 68.76 6.655 69.085 6.98 ;
      RECT 68.735 6.655 69.085 6.885 ;
      RECT 68.565 6.685 69.085 6.855 ;
      RECT 67.96 2.365 68.28 2.685 ;
      RECT 67.93 2.365 68.28 2.595 ;
      RECT 67.645 2.395 68.28 2.565 ;
      RECT 67.96 6.28 68.28 6.605 ;
      RECT 67.93 6.285 68.28 6.515 ;
      RECT 67.76 6.315 68.28 6.485 ;
      RECT 63.705 3.79 64.025 4.05 ;
      RECT 64.74 3.805 65.03 4.035 ;
      RECT 63.705 3.85 65.03 3.99 ;
      RECT 63.365 5.83 63.685 6.09 ;
      RECT 64.74 5.845 65.03 6.075 ;
      RECT 64.815 5.55 64.955 6.075 ;
      RECT 63.455 5.55 63.595 6.09 ;
      RECT 63.455 5.55 64.955 5.69 ;
      RECT 64.385 2.77 64.705 3.03 ;
      RECT 64.11 2.83 64.705 2.97 ;
      RECT 61.325 6.51 61.645 6.77 ;
      RECT 60.32 6.525 60.61 6.755 ;
      RECT 60.32 6.57 62.235 6.71 ;
      RECT 62.095 6.23 62.235 6.71 ;
      RECT 62.095 6.23 64.105 6.37 ;
      RECT 63.965 5.845 64.105 6.37 ;
      RECT 63.89 5.845 64.18 6.075 ;
      RECT 63.705 4.81 64.025 5.07 ;
      RECT 61.56 4.825 61.85 5.055 ;
      RECT 61.56 4.87 64.025 5.01 ;
      RECT 63.025 3.79 63.345 4.05 ;
      RECT 60.66 3.805 60.95 4.035 ;
      RECT 60.66 3.85 63.345 3.99 ;
      RECT 62.685 6.51 63.005 6.77 ;
      RECT 62.685 6.57 63.28 6.71 ;
      RECT 62.685 3.11 63.005 3.37 ;
      RECT 62.41 3.17 63.005 3.31 ;
      RECT 62.005 2.77 62.325 3.03 ;
      RECT 61.73 2.83 62.325 2.97 ;
      RECT 61.665 3.45 61.985 3.71 ;
      RECT 58.79 3.465 59.08 3.695 ;
      RECT 58.79 3.51 61.985 3.65 ;
      RECT 61.245 2.79 61.385 3.65 ;
      RECT 61.17 2.79 61.46 3.02 ;
      RECT 61.325 2.26 61.645 2.52 ;
      RECT 61.325 2.275 61.83 2.505 ;
      RECT 61.235 2.32 61.83 2.46 ;
      RECT 60.66 2.79 60.95 3.02 ;
      RECT 60.055 2.835 60.95 2.975 ;
      RECT 60.055 2.43 60.195 2.975 ;
      RECT 59.965 2.43 60.285 2.69 ;
      RECT 59.285 2.77 59.605 3.03 ;
      RECT 59.01 2.83 59.605 2.97 ;
      RECT 59.285 4.81 59.605 5.07 ;
      RECT 59.01 4.87 59.605 5.01 ;
      RECT 57.05 6.575 57.34 6.885 ;
      RECT 56.88 6.685 57.37 6.855 ;
      RECT 57.03 6.575 57.37 6.855 ;
      RECT 56.62 7.765 56.91 7.995 ;
      RECT 56.68 6.995 56.85 7.995 ;
      RECT 56.585 6.995 56.955 7.37 ;
      RECT 53.865 7.77 54.155 8 ;
      RECT 53.925 6.29 54.095 8 ;
      RECT 53.925 6.655 54.255 6.98 ;
      RECT 53.865 6.29 54.155 6.52 ;
      RECT 53.46 2.395 53.565 2.965 ;
      RECT 53.46 2.73 53.785 2.96 ;
      RECT 53.46 2.76 53.955 2.93 ;
      RECT 53.46 2.395 53.65 2.96 ;
      RECT 52.875 2.36 53.165 2.59 ;
      RECT 52.875 2.395 53.65 2.565 ;
      RECT 52.935 0.88 53.105 2.59 ;
      RECT 52.875 0.88 53.165 1.11 ;
      RECT 52.875 7.77 53.165 8 ;
      RECT 52.935 6.29 53.105 8 ;
      RECT 52.875 6.29 53.165 6.52 ;
      RECT 52.875 6.325 53.73 6.485 ;
      RECT 53.56 5.92 53.73 6.485 ;
      RECT 52.875 6.32 53.27 6.485 ;
      RECT 53.495 5.92 53.785 6.15 ;
      RECT 53.495 5.95 53.955 6.12 ;
      RECT 52.505 2.73 52.795 2.96 ;
      RECT 52.505 2.76 52.965 2.93 ;
      RECT 52.57 1.655 52.735 2.96 ;
      RECT 51.085 1.625 51.375 1.855 ;
      RECT 51.085 1.655 52.735 1.825 ;
      RECT 51.145 0.885 51.315 1.855 ;
      RECT 51.085 0.885 51.375 1.115 ;
      RECT 51.085 7.765 51.375 7.995 ;
      RECT 51.145 7.025 51.315 7.995 ;
      RECT 51.145 7.12 52.735 7.29 ;
      RECT 52.565 5.92 52.735 7.29 ;
      RECT 51.085 7.025 51.375 7.255 ;
      RECT 52.505 5.92 52.795 6.15 ;
      RECT 52.505 5.95 52.965 6.12 ;
      RECT 51.515 1.965 51.865 2.315 ;
      RECT 51.345 2.025 51.865 2.195 ;
      RECT 51.54 6.655 51.865 6.98 ;
      RECT 51.515 6.655 51.865 6.885 ;
      RECT 51.345 6.685 51.865 6.855 ;
      RECT 50.74 2.365 51.06 2.685 ;
      RECT 50.71 2.365 51.06 2.595 ;
      RECT 50.425 2.395 51.06 2.565 ;
      RECT 50.74 6.28 51.06 6.605 ;
      RECT 50.71 6.285 51.06 6.515 ;
      RECT 50.54 6.315 51.06 6.485 ;
      RECT 46.485 3.79 46.805 4.05 ;
      RECT 47.52 3.805 47.81 4.035 ;
      RECT 46.485 3.85 47.81 3.99 ;
      RECT 46.145 5.83 46.465 6.09 ;
      RECT 47.52 5.845 47.81 6.075 ;
      RECT 47.595 5.55 47.735 6.075 ;
      RECT 46.235 5.55 46.375 6.09 ;
      RECT 46.235 5.55 47.735 5.69 ;
      RECT 47.165 2.77 47.485 3.03 ;
      RECT 46.89 2.83 47.485 2.97 ;
      RECT 44.105 6.51 44.425 6.77 ;
      RECT 43.1 6.525 43.39 6.755 ;
      RECT 43.1 6.57 45.015 6.71 ;
      RECT 44.875 6.23 45.015 6.71 ;
      RECT 44.875 6.23 46.885 6.37 ;
      RECT 46.745 5.845 46.885 6.37 ;
      RECT 46.67 5.845 46.96 6.075 ;
      RECT 46.485 4.81 46.805 5.07 ;
      RECT 44.34 4.825 44.63 5.055 ;
      RECT 44.34 4.87 46.805 5.01 ;
      RECT 45.805 3.79 46.125 4.05 ;
      RECT 43.44 3.805 43.73 4.035 ;
      RECT 43.44 3.85 46.125 3.99 ;
      RECT 45.465 6.51 45.785 6.77 ;
      RECT 45.465 6.57 46.06 6.71 ;
      RECT 45.465 3.11 45.785 3.37 ;
      RECT 45.19 3.17 45.785 3.31 ;
      RECT 44.785 2.77 45.105 3.03 ;
      RECT 44.51 2.83 45.105 2.97 ;
      RECT 44.445 3.45 44.765 3.71 ;
      RECT 41.57 3.465 41.86 3.695 ;
      RECT 41.57 3.51 44.765 3.65 ;
      RECT 44.025 2.79 44.165 3.65 ;
      RECT 43.95 2.79 44.24 3.02 ;
      RECT 44.105 2.26 44.425 2.52 ;
      RECT 44.105 2.275 44.61 2.505 ;
      RECT 44.015 2.32 44.61 2.46 ;
      RECT 43.44 2.79 43.73 3.02 ;
      RECT 42.835 2.835 43.73 2.975 ;
      RECT 42.835 2.43 42.975 2.975 ;
      RECT 42.745 2.43 43.065 2.69 ;
      RECT 42.065 2.77 42.385 3.03 ;
      RECT 41.79 2.83 42.385 2.97 ;
      RECT 42.065 4.81 42.385 5.07 ;
      RECT 41.79 4.87 42.385 5.01 ;
      RECT 39.83 6.575 40.12 6.885 ;
      RECT 39.66 6.685 40.15 6.855 ;
      RECT 39.81 6.575 40.15 6.855 ;
      RECT 39.4 7.765 39.69 7.995 ;
      RECT 39.46 6.995 39.63 7.995 ;
      RECT 39.365 6.995 39.735 7.37 ;
      RECT 36.645 7.77 36.935 8 ;
      RECT 36.705 6.29 36.875 8 ;
      RECT 36.705 6.655 37.035 6.98 ;
      RECT 36.645 6.29 36.935 6.52 ;
      RECT 36.24 2.395 36.345 2.965 ;
      RECT 36.24 2.73 36.565 2.96 ;
      RECT 36.24 2.76 36.735 2.93 ;
      RECT 36.24 2.395 36.43 2.96 ;
      RECT 35.655 2.36 35.945 2.59 ;
      RECT 35.655 2.395 36.43 2.565 ;
      RECT 35.715 0.88 35.885 2.59 ;
      RECT 35.655 0.88 35.945 1.11 ;
      RECT 35.655 7.77 35.945 8 ;
      RECT 35.715 6.29 35.885 8 ;
      RECT 35.655 6.29 35.945 6.52 ;
      RECT 35.655 6.325 36.51 6.485 ;
      RECT 36.34 5.92 36.51 6.485 ;
      RECT 35.655 6.32 36.05 6.485 ;
      RECT 36.275 5.92 36.565 6.15 ;
      RECT 36.275 5.95 36.735 6.12 ;
      RECT 35.285 2.73 35.575 2.96 ;
      RECT 35.285 2.76 35.745 2.93 ;
      RECT 35.35 1.655 35.515 2.96 ;
      RECT 33.865 1.625 34.155 1.855 ;
      RECT 33.865 1.655 35.515 1.825 ;
      RECT 33.925 0.885 34.095 1.855 ;
      RECT 33.865 0.885 34.155 1.115 ;
      RECT 33.865 7.765 34.155 7.995 ;
      RECT 33.925 7.025 34.095 7.995 ;
      RECT 33.925 7.12 35.515 7.29 ;
      RECT 35.345 5.92 35.515 7.29 ;
      RECT 33.865 7.025 34.155 7.255 ;
      RECT 35.285 5.92 35.575 6.15 ;
      RECT 35.285 5.95 35.745 6.12 ;
      RECT 34.295 1.965 34.645 2.315 ;
      RECT 34.125 2.025 34.645 2.195 ;
      RECT 34.32 6.655 34.645 6.98 ;
      RECT 34.295 6.655 34.645 6.885 ;
      RECT 34.125 6.685 34.645 6.855 ;
      RECT 33.52 2.365 33.84 2.685 ;
      RECT 33.49 2.365 33.84 2.595 ;
      RECT 33.205 2.395 33.84 2.565 ;
      RECT 33.52 6.28 33.84 6.605 ;
      RECT 33.49 6.285 33.84 6.515 ;
      RECT 33.32 6.315 33.84 6.485 ;
      RECT 29.265 3.79 29.585 4.05 ;
      RECT 30.3 3.805 30.59 4.035 ;
      RECT 29.265 3.85 30.59 3.99 ;
      RECT 28.925 5.83 29.245 6.09 ;
      RECT 30.3 5.845 30.59 6.075 ;
      RECT 30.375 5.55 30.515 6.075 ;
      RECT 29.015 5.55 29.155 6.09 ;
      RECT 29.015 5.55 30.515 5.69 ;
      RECT 29.945 2.77 30.265 3.03 ;
      RECT 29.67 2.83 30.265 2.97 ;
      RECT 26.885 6.51 27.205 6.77 ;
      RECT 25.88 6.525 26.17 6.755 ;
      RECT 25.88 6.57 27.795 6.71 ;
      RECT 27.655 6.23 27.795 6.71 ;
      RECT 27.655 6.23 29.665 6.37 ;
      RECT 29.525 5.845 29.665 6.37 ;
      RECT 29.45 5.845 29.74 6.075 ;
      RECT 29.265 4.81 29.585 5.07 ;
      RECT 27.12 4.825 27.41 5.055 ;
      RECT 27.12 4.87 29.585 5.01 ;
      RECT 28.585 3.79 28.905 4.05 ;
      RECT 26.22 3.805 26.51 4.035 ;
      RECT 26.22 3.85 28.905 3.99 ;
      RECT 28.245 6.51 28.565 6.77 ;
      RECT 28.245 6.57 28.84 6.71 ;
      RECT 28.245 3.11 28.565 3.37 ;
      RECT 27.97 3.17 28.565 3.31 ;
      RECT 27.565 2.77 27.885 3.03 ;
      RECT 27.29 2.83 27.885 2.97 ;
      RECT 27.225 3.45 27.545 3.71 ;
      RECT 24.35 3.465 24.64 3.695 ;
      RECT 24.35 3.51 27.545 3.65 ;
      RECT 26.805 2.79 26.945 3.65 ;
      RECT 26.73 2.79 27.02 3.02 ;
      RECT 26.885 2.26 27.205 2.52 ;
      RECT 26.885 2.275 27.39 2.505 ;
      RECT 26.795 2.32 27.39 2.46 ;
      RECT 26.22 2.79 26.51 3.02 ;
      RECT 25.615 2.835 26.51 2.975 ;
      RECT 25.615 2.43 25.755 2.975 ;
      RECT 25.525 2.43 25.845 2.69 ;
      RECT 24.845 2.77 25.165 3.03 ;
      RECT 24.57 2.83 25.165 2.97 ;
      RECT 24.845 4.81 25.165 5.07 ;
      RECT 24.57 4.87 25.165 5.01 ;
      RECT 22.61 6.575 22.9 6.885 ;
      RECT 22.44 6.685 22.93 6.855 ;
      RECT 22.59 6.575 22.93 6.855 ;
      RECT 22.18 7.765 22.47 7.995 ;
      RECT 22.24 6.995 22.41 7.995 ;
      RECT 22.145 6.995 22.515 7.37 ;
      RECT 19.425 7.77 19.715 8 ;
      RECT 19.485 6.29 19.655 8 ;
      RECT 19.485 6.655 19.815 6.98 ;
      RECT 19.425 6.29 19.715 6.52 ;
      RECT 19.02 2.395 19.125 2.965 ;
      RECT 19.02 2.73 19.345 2.96 ;
      RECT 19.02 2.76 19.515 2.93 ;
      RECT 19.02 2.395 19.21 2.96 ;
      RECT 18.435 2.36 18.725 2.59 ;
      RECT 18.435 2.395 19.21 2.565 ;
      RECT 18.495 0.88 18.665 2.59 ;
      RECT 18.435 0.88 18.725 1.11 ;
      RECT 18.435 7.77 18.725 8 ;
      RECT 18.495 6.29 18.665 8 ;
      RECT 18.435 6.29 18.725 6.52 ;
      RECT 18.435 6.325 19.29 6.485 ;
      RECT 19.12 5.92 19.29 6.485 ;
      RECT 18.435 6.32 18.83 6.485 ;
      RECT 19.055 5.92 19.345 6.15 ;
      RECT 19.055 5.95 19.515 6.12 ;
      RECT 18.065 2.73 18.355 2.96 ;
      RECT 18.065 2.76 18.525 2.93 ;
      RECT 18.13 1.655 18.295 2.96 ;
      RECT 16.645 1.625 16.935 1.855 ;
      RECT 16.645 1.655 18.295 1.825 ;
      RECT 16.705 0.885 16.875 1.855 ;
      RECT 16.645 0.885 16.935 1.115 ;
      RECT 16.645 7.765 16.935 7.995 ;
      RECT 16.705 7.025 16.875 7.995 ;
      RECT 16.705 7.12 18.295 7.29 ;
      RECT 18.125 5.92 18.295 7.29 ;
      RECT 16.645 7.025 16.935 7.255 ;
      RECT 18.065 5.92 18.355 6.15 ;
      RECT 18.065 5.95 18.525 6.12 ;
      RECT 17.075 1.965 17.425 2.315 ;
      RECT 16.905 2.025 17.425 2.195 ;
      RECT 17.1 6.655 17.425 6.98 ;
      RECT 17.075 6.655 17.425 6.885 ;
      RECT 16.905 6.685 17.425 6.855 ;
      RECT 16.3 2.365 16.62 2.685 ;
      RECT 16.27 2.365 16.62 2.595 ;
      RECT 15.985 2.395 16.62 2.565 ;
      RECT 16.3 6.28 16.62 6.605 ;
      RECT 16.27 6.285 16.62 6.515 ;
      RECT 16.1 6.315 16.62 6.485 ;
      RECT 12.045 3.79 12.365 4.05 ;
      RECT 13.08 3.805 13.37 4.035 ;
      RECT 12.045 3.85 13.37 3.99 ;
      RECT 11.705 5.83 12.025 6.09 ;
      RECT 13.08 5.845 13.37 6.075 ;
      RECT 13.155 5.55 13.295 6.075 ;
      RECT 11.795 5.55 11.935 6.09 ;
      RECT 11.795 5.55 13.295 5.69 ;
      RECT 12.725 2.77 13.045 3.03 ;
      RECT 12.45 2.83 13.045 2.97 ;
      RECT 9.665 6.51 9.985 6.77 ;
      RECT 8.66 6.525 8.95 6.755 ;
      RECT 8.66 6.57 10.575 6.71 ;
      RECT 10.435 6.23 10.575 6.71 ;
      RECT 10.435 6.23 12.445 6.37 ;
      RECT 12.305 5.845 12.445 6.37 ;
      RECT 12.23 5.845 12.52 6.075 ;
      RECT 12.045 4.81 12.365 5.07 ;
      RECT 9.9 4.825 10.19 5.055 ;
      RECT 9.9 4.87 12.365 5.01 ;
      RECT 11.365 3.79 11.685 4.05 ;
      RECT 9 3.805 9.29 4.035 ;
      RECT 9 3.85 11.685 3.99 ;
      RECT 11.025 6.51 11.345 6.77 ;
      RECT 11.025 6.57 11.62 6.71 ;
      RECT 11.025 3.11 11.345 3.37 ;
      RECT 10.75 3.17 11.345 3.31 ;
      RECT 10.345 2.77 10.665 3.03 ;
      RECT 10.07 2.83 10.665 2.97 ;
      RECT 10.005 3.45 10.325 3.71 ;
      RECT 7.13 3.465 7.42 3.695 ;
      RECT 7.13 3.51 10.325 3.65 ;
      RECT 9.585 2.79 9.725 3.65 ;
      RECT 9.51 2.79 9.8 3.02 ;
      RECT 9.665 2.26 9.985 2.52 ;
      RECT 9.665 2.275 10.17 2.505 ;
      RECT 9.575 2.32 10.17 2.46 ;
      RECT 9 2.79 9.29 3.02 ;
      RECT 8.395 2.835 9.29 2.975 ;
      RECT 8.395 2.43 8.535 2.975 ;
      RECT 8.305 2.43 8.625 2.69 ;
      RECT 7.625 2.77 7.945 3.03 ;
      RECT 7.35 2.83 7.945 2.97 ;
      RECT 7.625 4.81 7.945 5.07 ;
      RECT 7.35 4.87 7.945 5.01 ;
      RECT 5.39 6.575 5.68 6.885 ;
      RECT 5.22 6.685 5.71 6.855 ;
      RECT 5.37 6.575 5.71 6.855 ;
      RECT 4.96 7.765 5.25 7.995 ;
      RECT 5.02 6.995 5.19 7.995 ;
      RECT 4.925 6.995 5.295 7.37 ;
      RECT 1.55 7.765 1.84 7.995 ;
      RECT 1.61 7.025 1.78 7.995 ;
      RECT 1.52 7.025 1.86 7.305 ;
      RECT 1.145 6.285 1.485 6.565 ;
      RECT 1.005 6.315 1.485 6.485 ;
      RECT 83.51 1.995 83.835 2.32 ;
      RECT 81.28 6.51 81.925 6.77 ;
      RECT 79.23 5.83 79.875 6.09 ;
      RECT 66.29 1.995 66.615 2.32 ;
      RECT 64.06 6.51 64.705 6.77 ;
      RECT 62.01 5.83 62.655 6.09 ;
      RECT 49.07 1.995 49.395 2.32 ;
      RECT 46.84 6.51 47.485 6.77 ;
      RECT 44.79 5.83 45.435 6.09 ;
      RECT 31.85 1.995 32.175 2.32 ;
      RECT 29.62 6.51 30.265 6.77 ;
      RECT 27.57 5.83 28.215 6.09 ;
      RECT 14.63 1.995 14.955 2.32 ;
      RECT 12.4 6.51 13.045 6.77 ;
      RECT 10.35 5.83 10.995 6.09 ;
    LAYER mcon ;
      RECT 88.365 6.32 88.535 6.49 ;
      RECT 88.37 6.315 88.54 6.485 ;
      RECT 71.145 6.32 71.315 6.49 ;
      RECT 71.15 6.315 71.32 6.485 ;
      RECT 53.925 6.32 54.095 6.49 ;
      RECT 53.93 6.315 54.1 6.485 ;
      RECT 36.705 6.32 36.875 6.49 ;
      RECT 36.71 6.315 36.88 6.485 ;
      RECT 19.485 6.32 19.655 6.49 ;
      RECT 19.49 6.315 19.66 6.485 ;
      RECT 88.365 7.8 88.535 7.97 ;
      RECT 87.995 2.76 88.165 2.93 ;
      RECT 87.995 5.95 88.165 6.12 ;
      RECT 87.375 0.91 87.545 1.08 ;
      RECT 87.375 2.39 87.545 2.56 ;
      RECT 87.375 6.32 87.545 6.49 ;
      RECT 87.375 7.8 87.545 7.97 ;
      RECT 87.005 2.76 87.175 2.93 ;
      RECT 87.005 5.95 87.175 6.12 ;
      RECT 86.015 2.025 86.185 2.195 ;
      RECT 86.015 6.685 86.185 6.855 ;
      RECT 85.585 0.915 85.755 1.085 ;
      RECT 85.585 1.655 85.755 1.825 ;
      RECT 85.585 7.055 85.755 7.225 ;
      RECT 85.585 7.795 85.755 7.965 ;
      RECT 85.21 2.395 85.38 2.565 ;
      RECT 85.21 6.315 85.38 6.485 ;
      RECT 82.02 3.835 82.19 4.005 ;
      RECT 82.02 5.875 82.19 6.045 ;
      RECT 81.68 2.815 81.85 2.985 ;
      RECT 81.34 6.555 81.51 6.725 ;
      RECT 81.17 5.875 81.34 6.045 ;
      RECT 80.66 5.875 80.83 6.045 ;
      RECT 79.98 3.155 80.15 3.325 ;
      RECT 79.98 6.555 80.15 6.725 ;
      RECT 79.3 2.815 79.47 2.985 ;
      RECT 79.29 5.875 79.46 6.045 ;
      RECT 78.84 4.855 79.01 5.025 ;
      RECT 78.82 2.305 78.99 2.475 ;
      RECT 78.45 2.82 78.62 2.99 ;
      RECT 77.94 2.82 78.11 2.99 ;
      RECT 77.94 3.835 78.11 4.005 ;
      RECT 77.6 6.555 77.77 6.725 ;
      RECT 76.58 2.815 76.75 2.985 ;
      RECT 76.58 4.855 76.75 5.025 ;
      RECT 76.07 3.495 76.24 3.665 ;
      RECT 74.33 6.685 74.5 6.855 ;
      RECT 73.9 7.055 74.07 7.225 ;
      RECT 73.9 7.795 74.07 7.965 ;
      RECT 71.145 7.8 71.315 7.97 ;
      RECT 70.775 2.76 70.945 2.93 ;
      RECT 70.775 5.95 70.945 6.12 ;
      RECT 70.155 0.91 70.325 1.08 ;
      RECT 70.155 2.39 70.325 2.56 ;
      RECT 70.155 6.32 70.325 6.49 ;
      RECT 70.155 7.8 70.325 7.97 ;
      RECT 69.785 2.76 69.955 2.93 ;
      RECT 69.785 5.95 69.955 6.12 ;
      RECT 68.795 2.025 68.965 2.195 ;
      RECT 68.795 6.685 68.965 6.855 ;
      RECT 68.365 0.915 68.535 1.085 ;
      RECT 68.365 1.655 68.535 1.825 ;
      RECT 68.365 7.055 68.535 7.225 ;
      RECT 68.365 7.795 68.535 7.965 ;
      RECT 67.99 2.395 68.16 2.565 ;
      RECT 67.99 6.315 68.16 6.485 ;
      RECT 64.8 3.835 64.97 4.005 ;
      RECT 64.8 5.875 64.97 6.045 ;
      RECT 64.46 2.815 64.63 2.985 ;
      RECT 64.12 6.555 64.29 6.725 ;
      RECT 63.95 5.875 64.12 6.045 ;
      RECT 63.44 5.875 63.61 6.045 ;
      RECT 62.76 3.155 62.93 3.325 ;
      RECT 62.76 6.555 62.93 6.725 ;
      RECT 62.08 2.815 62.25 2.985 ;
      RECT 62.07 5.875 62.24 6.045 ;
      RECT 61.62 4.855 61.79 5.025 ;
      RECT 61.6 2.305 61.77 2.475 ;
      RECT 61.23 2.82 61.4 2.99 ;
      RECT 60.72 2.82 60.89 2.99 ;
      RECT 60.72 3.835 60.89 4.005 ;
      RECT 60.38 6.555 60.55 6.725 ;
      RECT 59.36 2.815 59.53 2.985 ;
      RECT 59.36 4.855 59.53 5.025 ;
      RECT 58.85 3.495 59.02 3.665 ;
      RECT 57.11 6.685 57.28 6.855 ;
      RECT 56.68 7.055 56.85 7.225 ;
      RECT 56.68 7.795 56.85 7.965 ;
      RECT 53.925 7.8 54.095 7.97 ;
      RECT 53.555 2.76 53.725 2.93 ;
      RECT 53.555 5.95 53.725 6.12 ;
      RECT 52.935 0.91 53.105 1.08 ;
      RECT 52.935 2.39 53.105 2.56 ;
      RECT 52.935 6.32 53.105 6.49 ;
      RECT 52.935 7.8 53.105 7.97 ;
      RECT 52.565 2.76 52.735 2.93 ;
      RECT 52.565 5.95 52.735 6.12 ;
      RECT 51.575 2.025 51.745 2.195 ;
      RECT 51.575 6.685 51.745 6.855 ;
      RECT 51.145 0.915 51.315 1.085 ;
      RECT 51.145 1.655 51.315 1.825 ;
      RECT 51.145 7.055 51.315 7.225 ;
      RECT 51.145 7.795 51.315 7.965 ;
      RECT 50.77 2.395 50.94 2.565 ;
      RECT 50.77 6.315 50.94 6.485 ;
      RECT 47.58 3.835 47.75 4.005 ;
      RECT 47.58 5.875 47.75 6.045 ;
      RECT 47.24 2.815 47.41 2.985 ;
      RECT 46.9 6.555 47.07 6.725 ;
      RECT 46.73 5.875 46.9 6.045 ;
      RECT 46.22 5.875 46.39 6.045 ;
      RECT 45.54 3.155 45.71 3.325 ;
      RECT 45.54 6.555 45.71 6.725 ;
      RECT 44.86 2.815 45.03 2.985 ;
      RECT 44.85 5.875 45.02 6.045 ;
      RECT 44.4 4.855 44.57 5.025 ;
      RECT 44.38 2.305 44.55 2.475 ;
      RECT 44.01 2.82 44.18 2.99 ;
      RECT 43.5 2.82 43.67 2.99 ;
      RECT 43.5 3.835 43.67 4.005 ;
      RECT 43.16 6.555 43.33 6.725 ;
      RECT 42.14 2.815 42.31 2.985 ;
      RECT 42.14 4.855 42.31 5.025 ;
      RECT 41.63 3.495 41.8 3.665 ;
      RECT 39.89 6.685 40.06 6.855 ;
      RECT 39.46 7.055 39.63 7.225 ;
      RECT 39.46 7.795 39.63 7.965 ;
      RECT 36.705 7.8 36.875 7.97 ;
      RECT 36.335 2.76 36.505 2.93 ;
      RECT 36.335 5.95 36.505 6.12 ;
      RECT 35.715 0.91 35.885 1.08 ;
      RECT 35.715 2.39 35.885 2.56 ;
      RECT 35.715 6.32 35.885 6.49 ;
      RECT 35.715 7.8 35.885 7.97 ;
      RECT 35.345 2.76 35.515 2.93 ;
      RECT 35.345 5.95 35.515 6.12 ;
      RECT 34.355 2.025 34.525 2.195 ;
      RECT 34.355 6.685 34.525 6.855 ;
      RECT 33.925 0.915 34.095 1.085 ;
      RECT 33.925 1.655 34.095 1.825 ;
      RECT 33.925 7.055 34.095 7.225 ;
      RECT 33.925 7.795 34.095 7.965 ;
      RECT 33.55 2.395 33.72 2.565 ;
      RECT 33.55 6.315 33.72 6.485 ;
      RECT 30.36 3.835 30.53 4.005 ;
      RECT 30.36 5.875 30.53 6.045 ;
      RECT 30.02 2.815 30.19 2.985 ;
      RECT 29.68 6.555 29.85 6.725 ;
      RECT 29.51 5.875 29.68 6.045 ;
      RECT 29 5.875 29.17 6.045 ;
      RECT 28.32 3.155 28.49 3.325 ;
      RECT 28.32 6.555 28.49 6.725 ;
      RECT 27.64 2.815 27.81 2.985 ;
      RECT 27.63 5.875 27.8 6.045 ;
      RECT 27.18 4.855 27.35 5.025 ;
      RECT 27.16 2.305 27.33 2.475 ;
      RECT 26.79 2.82 26.96 2.99 ;
      RECT 26.28 2.82 26.45 2.99 ;
      RECT 26.28 3.835 26.45 4.005 ;
      RECT 25.94 6.555 26.11 6.725 ;
      RECT 24.92 2.815 25.09 2.985 ;
      RECT 24.92 4.855 25.09 5.025 ;
      RECT 24.41 3.495 24.58 3.665 ;
      RECT 22.67 6.685 22.84 6.855 ;
      RECT 22.24 7.055 22.41 7.225 ;
      RECT 22.24 7.795 22.41 7.965 ;
      RECT 19.485 7.8 19.655 7.97 ;
      RECT 19.115 2.76 19.285 2.93 ;
      RECT 19.115 5.95 19.285 6.12 ;
      RECT 18.495 0.91 18.665 1.08 ;
      RECT 18.495 2.39 18.665 2.56 ;
      RECT 18.495 6.32 18.665 6.49 ;
      RECT 18.495 7.8 18.665 7.97 ;
      RECT 18.125 2.76 18.295 2.93 ;
      RECT 18.125 5.95 18.295 6.12 ;
      RECT 17.135 2.025 17.305 2.195 ;
      RECT 17.135 6.685 17.305 6.855 ;
      RECT 16.705 0.915 16.875 1.085 ;
      RECT 16.705 1.655 16.875 1.825 ;
      RECT 16.705 7.055 16.875 7.225 ;
      RECT 16.705 7.795 16.875 7.965 ;
      RECT 16.33 2.395 16.5 2.565 ;
      RECT 16.33 6.315 16.5 6.485 ;
      RECT 13.14 3.835 13.31 4.005 ;
      RECT 13.14 5.875 13.31 6.045 ;
      RECT 12.8 2.815 12.97 2.985 ;
      RECT 12.46 6.555 12.63 6.725 ;
      RECT 12.29 5.875 12.46 6.045 ;
      RECT 11.78 5.875 11.95 6.045 ;
      RECT 11.1 3.155 11.27 3.325 ;
      RECT 11.1 6.555 11.27 6.725 ;
      RECT 10.42 2.815 10.59 2.985 ;
      RECT 10.41 5.875 10.58 6.045 ;
      RECT 9.96 4.855 10.13 5.025 ;
      RECT 9.94 2.305 10.11 2.475 ;
      RECT 9.57 2.82 9.74 2.99 ;
      RECT 9.06 2.82 9.23 2.99 ;
      RECT 9.06 3.835 9.23 4.005 ;
      RECT 8.72 6.555 8.89 6.725 ;
      RECT 7.7 2.815 7.87 2.985 ;
      RECT 7.7 4.855 7.87 5.025 ;
      RECT 7.19 3.495 7.36 3.665 ;
      RECT 5.45 6.685 5.62 6.855 ;
      RECT 5.02 7.055 5.19 7.225 ;
      RECT 5.02 7.795 5.19 7.965 ;
      RECT 1.61 7.055 1.78 7.225 ;
      RECT 1.61 7.795 1.78 7.965 ;
      RECT 1.235 6.315 1.405 6.485 ;
    LAYER li1 ;
      RECT 88.365 5.02 88.535 6.49 ;
      RECT 88.365 6.315 88.54 6.485 ;
      RECT 87.995 1.74 88.165 2.93 ;
      RECT 87.995 1.74 88.465 1.91 ;
      RECT 87.995 6.97 88.465 7.14 ;
      RECT 87.995 5.95 88.165 7.14 ;
      RECT 87.005 1.74 87.175 2.93 ;
      RECT 87.005 1.74 87.475 1.91 ;
      RECT 87.005 6.97 87.475 7.14 ;
      RECT 87.005 5.95 87.175 7.14 ;
      RECT 85.155 2.635 85.325 3.865 ;
      RECT 85.21 0.855 85.38 2.805 ;
      RECT 85.155 0.575 85.325 1.025 ;
      RECT 85.155 7.855 85.325 8.305 ;
      RECT 85.21 6.075 85.38 8.025 ;
      RECT 85.155 5.015 85.325 6.245 ;
      RECT 84.635 0.575 84.805 3.865 ;
      RECT 84.635 2.075 85.04 2.405 ;
      RECT 84.635 1.235 85.04 1.565 ;
      RECT 84.635 5.015 84.805 8.305 ;
      RECT 84.635 7.315 85.04 7.645 ;
      RECT 84.635 6.475 85.04 6.805 ;
      RECT 82.37 3.495 82.75 4.175 ;
      RECT 82.58 2.365 82.75 4.175 ;
      RECT 80.5 2.365 80.73 3.035 ;
      RECT 80.5 2.365 82.75 2.535 ;
      RECT 82.03 2.045 82.2 2.535 ;
      RECT 82.02 3.155 82.19 4.005 ;
      RECT 81.105 3.155 82.41 3.325 ;
      RECT 82.165 2.705 82.41 3.325 ;
      RECT 81.105 2.785 81.275 3.325 ;
      RECT 80.9 2.785 81.275 2.955 ;
      RECT 81.08 6.265 81.775 6.895 ;
      RECT 81.605 4.685 81.775 6.895 ;
      RECT 81.51 4.685 81.84 5.665 ;
      RECT 81.11 3.495 81.44 4.175 ;
      RECT 80.2 3.495 80.6 4.175 ;
      RECT 80.2 3.495 81.44 3.665 ;
      RECT 79.7 3.075 80.02 4.175 ;
      RECT 79.7 3.075 80.15 3.325 ;
      RECT 79.7 3.075 80.33 3.245 ;
      RECT 80.16 2.025 80.33 3.245 ;
      RECT 80.16 2.025 81.115 2.195 ;
      RECT 79.7 6.265 80.395 6.895 ;
      RECT 80.225 4.685 80.395 6.895 ;
      RECT 80.13 4.685 80.46 5.665 ;
      RECT 79.72 5.825 80.055 6.075 ;
      RECT 79.175 5.825 79.51 6.075 ;
      RECT 79.175 5.875 80.055 6.045 ;
      RECT 78.835 6.265 79.53 6.895 ;
      RECT 78.835 4.685 79.005 6.895 ;
      RECT 78.77 4.685 79.1 5.665 ;
      RECT 78.33 3.205 78.66 4.16 ;
      RECT 78.33 3.205 79.01 3.375 ;
      RECT 78.84 1.965 79.01 3.375 ;
      RECT 78.75 1.965 79.08 2.605 ;
      RECT 77.81 3.205 78.14 4.16 ;
      RECT 77.46 3.205 78.14 3.375 ;
      RECT 77.46 1.965 77.63 3.375 ;
      RECT 77.39 1.965 77.72 2.605 ;
      RECT 77.6 5.875 77.77 6.725 ;
      RECT 76.875 5.825 77.21 6.075 ;
      RECT 76.875 5.875 77.77 6.045 ;
      RECT 76.94 2.785 77.29 3.035 ;
      RECT 76.42 2.785 76.75 3.035 ;
      RECT 76.42 2.815 77.29 2.985 ;
      RECT 76.535 6.265 77.23 6.895 ;
      RECT 76.535 4.685 76.705 6.895 ;
      RECT 76.47 4.685 76.8 5.665 ;
      RECT 76 3.195 76.33 4.175 ;
      RECT 76 1.965 76.25 4.175 ;
      RECT 76 1.965 76.33 2.595 ;
      RECT 72.95 5.015 73.12 8.305 ;
      RECT 72.95 7.315 73.355 7.645 ;
      RECT 72.95 6.475 73.355 6.805 ;
      RECT 71.145 5.02 71.315 6.49 ;
      RECT 71.145 6.315 71.32 6.485 ;
      RECT 70.775 1.74 70.945 2.93 ;
      RECT 70.775 1.74 71.245 1.91 ;
      RECT 70.775 6.97 71.245 7.14 ;
      RECT 70.775 5.95 70.945 7.14 ;
      RECT 69.785 1.74 69.955 2.93 ;
      RECT 69.785 1.74 70.255 1.91 ;
      RECT 69.785 6.97 70.255 7.14 ;
      RECT 69.785 5.95 69.955 7.14 ;
      RECT 67.935 2.635 68.105 3.865 ;
      RECT 67.99 0.855 68.16 2.805 ;
      RECT 67.935 0.575 68.105 1.025 ;
      RECT 67.935 7.855 68.105 8.305 ;
      RECT 67.99 6.075 68.16 8.025 ;
      RECT 67.935 5.015 68.105 6.245 ;
      RECT 67.415 0.575 67.585 3.865 ;
      RECT 67.415 2.075 67.82 2.405 ;
      RECT 67.415 1.235 67.82 1.565 ;
      RECT 67.415 5.015 67.585 8.305 ;
      RECT 67.415 7.315 67.82 7.645 ;
      RECT 67.415 6.475 67.82 6.805 ;
      RECT 65.15 3.495 65.53 4.175 ;
      RECT 65.36 2.365 65.53 4.175 ;
      RECT 63.28 2.365 63.51 3.035 ;
      RECT 63.28 2.365 65.53 2.535 ;
      RECT 64.81 2.045 64.98 2.535 ;
      RECT 64.8 3.155 64.97 4.005 ;
      RECT 63.885 3.155 65.19 3.325 ;
      RECT 64.945 2.705 65.19 3.325 ;
      RECT 63.885 2.785 64.055 3.325 ;
      RECT 63.68 2.785 64.055 2.955 ;
      RECT 63.86 6.265 64.555 6.895 ;
      RECT 64.385 4.685 64.555 6.895 ;
      RECT 64.29 4.685 64.62 5.665 ;
      RECT 63.89 3.495 64.22 4.175 ;
      RECT 62.98 3.495 63.38 4.175 ;
      RECT 62.98 3.495 64.22 3.665 ;
      RECT 62.48 3.075 62.8 4.175 ;
      RECT 62.48 3.075 62.93 3.325 ;
      RECT 62.48 3.075 63.11 3.245 ;
      RECT 62.94 2.025 63.11 3.245 ;
      RECT 62.94 2.025 63.895 2.195 ;
      RECT 62.48 6.265 63.175 6.895 ;
      RECT 63.005 4.685 63.175 6.895 ;
      RECT 62.91 4.685 63.24 5.665 ;
      RECT 62.5 5.825 62.835 6.075 ;
      RECT 61.955 5.825 62.29 6.075 ;
      RECT 61.955 5.875 62.835 6.045 ;
      RECT 61.615 6.265 62.31 6.895 ;
      RECT 61.615 4.685 61.785 6.895 ;
      RECT 61.55 4.685 61.88 5.665 ;
      RECT 61.11 3.205 61.44 4.16 ;
      RECT 61.11 3.205 61.79 3.375 ;
      RECT 61.62 1.965 61.79 3.375 ;
      RECT 61.53 1.965 61.86 2.605 ;
      RECT 60.59 3.205 60.92 4.16 ;
      RECT 60.24 3.205 60.92 3.375 ;
      RECT 60.24 1.965 60.41 3.375 ;
      RECT 60.17 1.965 60.5 2.605 ;
      RECT 60.38 5.875 60.55 6.725 ;
      RECT 59.655 5.825 59.99 6.075 ;
      RECT 59.655 5.875 60.55 6.045 ;
      RECT 59.72 2.785 60.07 3.035 ;
      RECT 59.2 2.785 59.53 3.035 ;
      RECT 59.2 2.815 60.07 2.985 ;
      RECT 59.315 6.265 60.01 6.895 ;
      RECT 59.315 4.685 59.485 6.895 ;
      RECT 59.25 4.685 59.58 5.665 ;
      RECT 58.78 3.195 59.11 4.175 ;
      RECT 58.78 1.965 59.03 4.175 ;
      RECT 58.78 1.965 59.11 2.595 ;
      RECT 55.73 5.015 55.9 8.305 ;
      RECT 55.73 7.315 56.135 7.645 ;
      RECT 55.73 6.475 56.135 6.805 ;
      RECT 53.925 5.02 54.095 6.49 ;
      RECT 53.925 6.315 54.1 6.485 ;
      RECT 53.555 1.74 53.725 2.93 ;
      RECT 53.555 1.74 54.025 1.91 ;
      RECT 53.555 6.97 54.025 7.14 ;
      RECT 53.555 5.95 53.725 7.14 ;
      RECT 52.565 1.74 52.735 2.93 ;
      RECT 52.565 1.74 53.035 1.91 ;
      RECT 52.565 6.97 53.035 7.14 ;
      RECT 52.565 5.95 52.735 7.14 ;
      RECT 50.715 2.635 50.885 3.865 ;
      RECT 50.77 0.855 50.94 2.805 ;
      RECT 50.715 0.575 50.885 1.025 ;
      RECT 50.715 7.855 50.885 8.305 ;
      RECT 50.77 6.075 50.94 8.025 ;
      RECT 50.715 5.015 50.885 6.245 ;
      RECT 50.195 0.575 50.365 3.865 ;
      RECT 50.195 2.075 50.6 2.405 ;
      RECT 50.195 1.235 50.6 1.565 ;
      RECT 50.195 5.015 50.365 8.305 ;
      RECT 50.195 7.315 50.6 7.645 ;
      RECT 50.195 6.475 50.6 6.805 ;
      RECT 47.93 3.495 48.31 4.175 ;
      RECT 48.14 2.365 48.31 4.175 ;
      RECT 46.06 2.365 46.29 3.035 ;
      RECT 46.06 2.365 48.31 2.535 ;
      RECT 47.59 2.045 47.76 2.535 ;
      RECT 47.58 3.155 47.75 4.005 ;
      RECT 46.665 3.155 47.97 3.325 ;
      RECT 47.725 2.705 47.97 3.325 ;
      RECT 46.665 2.785 46.835 3.325 ;
      RECT 46.46 2.785 46.835 2.955 ;
      RECT 46.64 6.265 47.335 6.895 ;
      RECT 47.165 4.685 47.335 6.895 ;
      RECT 47.07 4.685 47.4 5.665 ;
      RECT 46.67 3.495 47 4.175 ;
      RECT 45.76 3.495 46.16 4.175 ;
      RECT 45.76 3.495 47 3.665 ;
      RECT 45.26 3.075 45.58 4.175 ;
      RECT 45.26 3.075 45.71 3.325 ;
      RECT 45.26 3.075 45.89 3.245 ;
      RECT 45.72 2.025 45.89 3.245 ;
      RECT 45.72 2.025 46.675 2.195 ;
      RECT 45.26 6.265 45.955 6.895 ;
      RECT 45.785 4.685 45.955 6.895 ;
      RECT 45.69 4.685 46.02 5.665 ;
      RECT 45.28 5.825 45.615 6.075 ;
      RECT 44.735 5.825 45.07 6.075 ;
      RECT 44.735 5.875 45.615 6.045 ;
      RECT 44.395 6.265 45.09 6.895 ;
      RECT 44.395 4.685 44.565 6.895 ;
      RECT 44.33 4.685 44.66 5.665 ;
      RECT 43.89 3.205 44.22 4.16 ;
      RECT 43.89 3.205 44.57 3.375 ;
      RECT 44.4 1.965 44.57 3.375 ;
      RECT 44.31 1.965 44.64 2.605 ;
      RECT 43.37 3.205 43.7 4.16 ;
      RECT 43.02 3.205 43.7 3.375 ;
      RECT 43.02 1.965 43.19 3.375 ;
      RECT 42.95 1.965 43.28 2.605 ;
      RECT 43.16 5.875 43.33 6.725 ;
      RECT 42.435 5.825 42.77 6.075 ;
      RECT 42.435 5.875 43.33 6.045 ;
      RECT 42.5 2.785 42.85 3.035 ;
      RECT 41.98 2.785 42.31 3.035 ;
      RECT 41.98 2.815 42.85 2.985 ;
      RECT 42.095 6.265 42.79 6.895 ;
      RECT 42.095 4.685 42.265 6.895 ;
      RECT 42.03 4.685 42.36 5.665 ;
      RECT 41.56 3.195 41.89 4.175 ;
      RECT 41.56 1.965 41.81 4.175 ;
      RECT 41.56 1.965 41.89 2.595 ;
      RECT 38.51 5.015 38.68 8.305 ;
      RECT 38.51 7.315 38.915 7.645 ;
      RECT 38.51 6.475 38.915 6.805 ;
      RECT 36.705 5.02 36.875 6.49 ;
      RECT 36.705 6.315 36.88 6.485 ;
      RECT 36.335 1.74 36.505 2.93 ;
      RECT 36.335 1.74 36.805 1.91 ;
      RECT 36.335 6.97 36.805 7.14 ;
      RECT 36.335 5.95 36.505 7.14 ;
      RECT 35.345 1.74 35.515 2.93 ;
      RECT 35.345 1.74 35.815 1.91 ;
      RECT 35.345 6.97 35.815 7.14 ;
      RECT 35.345 5.95 35.515 7.14 ;
      RECT 33.495 2.635 33.665 3.865 ;
      RECT 33.55 0.855 33.72 2.805 ;
      RECT 33.495 0.575 33.665 1.025 ;
      RECT 33.495 7.855 33.665 8.305 ;
      RECT 33.55 6.075 33.72 8.025 ;
      RECT 33.495 5.015 33.665 6.245 ;
      RECT 32.975 0.575 33.145 3.865 ;
      RECT 32.975 2.075 33.38 2.405 ;
      RECT 32.975 1.235 33.38 1.565 ;
      RECT 32.975 5.015 33.145 8.305 ;
      RECT 32.975 7.315 33.38 7.645 ;
      RECT 32.975 6.475 33.38 6.805 ;
      RECT 30.71 3.495 31.09 4.175 ;
      RECT 30.92 2.365 31.09 4.175 ;
      RECT 28.84 2.365 29.07 3.035 ;
      RECT 28.84 2.365 31.09 2.535 ;
      RECT 30.37 2.045 30.54 2.535 ;
      RECT 30.36 3.155 30.53 4.005 ;
      RECT 29.445 3.155 30.75 3.325 ;
      RECT 30.505 2.705 30.75 3.325 ;
      RECT 29.445 2.785 29.615 3.325 ;
      RECT 29.24 2.785 29.615 2.955 ;
      RECT 29.42 6.265 30.115 6.895 ;
      RECT 29.945 4.685 30.115 6.895 ;
      RECT 29.85 4.685 30.18 5.665 ;
      RECT 29.45 3.495 29.78 4.175 ;
      RECT 28.54 3.495 28.94 4.175 ;
      RECT 28.54 3.495 29.78 3.665 ;
      RECT 28.04 3.075 28.36 4.175 ;
      RECT 28.04 3.075 28.49 3.325 ;
      RECT 28.04 3.075 28.67 3.245 ;
      RECT 28.5 2.025 28.67 3.245 ;
      RECT 28.5 2.025 29.455 2.195 ;
      RECT 28.04 6.265 28.735 6.895 ;
      RECT 28.565 4.685 28.735 6.895 ;
      RECT 28.47 4.685 28.8 5.665 ;
      RECT 28.06 5.825 28.395 6.075 ;
      RECT 27.515 5.825 27.85 6.075 ;
      RECT 27.515 5.875 28.395 6.045 ;
      RECT 27.175 6.265 27.87 6.895 ;
      RECT 27.175 4.685 27.345 6.895 ;
      RECT 27.11 4.685 27.44 5.665 ;
      RECT 26.67 3.205 27 4.16 ;
      RECT 26.67 3.205 27.35 3.375 ;
      RECT 27.18 1.965 27.35 3.375 ;
      RECT 27.09 1.965 27.42 2.605 ;
      RECT 26.15 3.205 26.48 4.16 ;
      RECT 25.8 3.205 26.48 3.375 ;
      RECT 25.8 1.965 25.97 3.375 ;
      RECT 25.73 1.965 26.06 2.605 ;
      RECT 25.94 5.875 26.11 6.725 ;
      RECT 25.215 5.825 25.55 6.075 ;
      RECT 25.215 5.875 26.11 6.045 ;
      RECT 25.28 2.785 25.63 3.035 ;
      RECT 24.76 2.785 25.09 3.035 ;
      RECT 24.76 2.815 25.63 2.985 ;
      RECT 24.875 6.265 25.57 6.895 ;
      RECT 24.875 4.685 25.045 6.895 ;
      RECT 24.81 4.685 25.14 5.665 ;
      RECT 24.34 3.195 24.67 4.175 ;
      RECT 24.34 1.965 24.59 4.175 ;
      RECT 24.34 1.965 24.67 2.595 ;
      RECT 21.29 5.015 21.46 8.305 ;
      RECT 21.29 7.315 21.695 7.645 ;
      RECT 21.29 6.475 21.695 6.805 ;
      RECT 19.485 5.02 19.655 6.49 ;
      RECT 19.485 6.315 19.66 6.485 ;
      RECT 19.115 1.74 19.285 2.93 ;
      RECT 19.115 1.74 19.585 1.91 ;
      RECT 19.115 6.97 19.585 7.14 ;
      RECT 19.115 5.95 19.285 7.14 ;
      RECT 18.125 1.74 18.295 2.93 ;
      RECT 18.125 1.74 18.595 1.91 ;
      RECT 18.125 6.97 18.595 7.14 ;
      RECT 18.125 5.95 18.295 7.14 ;
      RECT 16.275 2.635 16.445 3.865 ;
      RECT 16.33 0.855 16.5 2.805 ;
      RECT 16.275 0.575 16.445 1.025 ;
      RECT 16.275 7.855 16.445 8.305 ;
      RECT 16.33 6.075 16.5 8.025 ;
      RECT 16.275 5.015 16.445 6.245 ;
      RECT 15.755 0.575 15.925 3.865 ;
      RECT 15.755 2.075 16.16 2.405 ;
      RECT 15.755 1.235 16.16 1.565 ;
      RECT 15.755 5.015 15.925 8.305 ;
      RECT 15.755 7.315 16.16 7.645 ;
      RECT 15.755 6.475 16.16 6.805 ;
      RECT 13.49 3.495 13.87 4.175 ;
      RECT 13.7 2.365 13.87 4.175 ;
      RECT 11.62 2.365 11.85 3.035 ;
      RECT 11.62 2.365 13.87 2.535 ;
      RECT 13.15 2.045 13.32 2.535 ;
      RECT 13.14 3.155 13.31 4.005 ;
      RECT 12.225 3.155 13.53 3.325 ;
      RECT 13.285 2.705 13.53 3.325 ;
      RECT 12.225 2.785 12.395 3.325 ;
      RECT 12.02 2.785 12.395 2.955 ;
      RECT 12.2 6.265 12.895 6.895 ;
      RECT 12.725 4.685 12.895 6.895 ;
      RECT 12.63 4.685 12.96 5.665 ;
      RECT 12.23 3.495 12.56 4.175 ;
      RECT 11.32 3.495 11.72 4.175 ;
      RECT 11.32 3.495 12.56 3.665 ;
      RECT 10.82 3.075 11.14 4.175 ;
      RECT 10.82 3.075 11.27 3.325 ;
      RECT 10.82 3.075 11.45 3.245 ;
      RECT 11.28 2.025 11.45 3.245 ;
      RECT 11.28 2.025 12.235 2.195 ;
      RECT 10.82 6.265 11.515 6.895 ;
      RECT 11.345 4.685 11.515 6.895 ;
      RECT 11.25 4.685 11.58 5.665 ;
      RECT 10.84 5.825 11.175 6.075 ;
      RECT 10.295 5.825 10.63 6.075 ;
      RECT 10.295 5.875 11.175 6.045 ;
      RECT 9.955 6.265 10.65 6.895 ;
      RECT 9.955 4.685 10.125 6.895 ;
      RECT 9.89 4.685 10.22 5.665 ;
      RECT 9.45 3.205 9.78 4.16 ;
      RECT 9.45 3.205 10.13 3.375 ;
      RECT 9.96 1.965 10.13 3.375 ;
      RECT 9.87 1.965 10.2 2.605 ;
      RECT 8.93 3.205 9.26 4.16 ;
      RECT 8.58 3.205 9.26 3.375 ;
      RECT 8.58 1.965 8.75 3.375 ;
      RECT 8.51 1.965 8.84 2.605 ;
      RECT 8.72 5.875 8.89 6.725 ;
      RECT 7.995 5.825 8.33 6.075 ;
      RECT 7.995 5.875 8.89 6.045 ;
      RECT 8.06 2.785 8.41 3.035 ;
      RECT 7.54 2.785 7.87 3.035 ;
      RECT 7.54 2.815 8.41 2.985 ;
      RECT 7.655 6.265 8.35 6.895 ;
      RECT 7.655 4.685 7.825 6.895 ;
      RECT 7.59 4.685 7.92 5.665 ;
      RECT 7.12 3.195 7.45 4.175 ;
      RECT 7.12 1.965 7.37 4.175 ;
      RECT 7.12 1.965 7.45 2.595 ;
      RECT 4.07 5.015 4.24 8.305 ;
      RECT 4.07 7.315 4.475 7.645 ;
      RECT 4.07 6.475 4.475 6.805 ;
      RECT 1.18 7.855 1.35 8.305 ;
      RECT 1.235 6.075 1.405 8.025 ;
      RECT 1.18 5.015 1.35 6.245 ;
      RECT 0.66 5.015 0.83 8.305 ;
      RECT 0.66 7.315 1.065 7.645 ;
      RECT 0.66 6.475 1.065 6.805 ;
      RECT 88.365 7.8 88.535 8.31 ;
      RECT 87.375 0.57 87.545 1.08 ;
      RECT 87.375 2.39 87.545 3.86 ;
      RECT 87.375 5.02 87.545 6.49 ;
      RECT 87.375 7.8 87.545 8.31 ;
      RECT 86.015 0.575 86.185 3.865 ;
      RECT 86.015 5.015 86.185 8.305 ;
      RECT 85.585 0.575 85.755 1.085 ;
      RECT 85.585 1.655 85.755 3.865 ;
      RECT 85.585 5.015 85.755 7.225 ;
      RECT 85.585 7.795 85.755 8.305 ;
      RECT 81.945 5.825 82.28 6.095 ;
      RECT 81.445 2.785 81.995 2.985 ;
      RECT 81.1 5.825 81.435 6.075 ;
      RECT 80.565 5.825 80.9 6.095 ;
      RECT 79.18 2.785 79.53 3.035 ;
      RECT 78.32 2.785 78.67 3.035 ;
      RECT 77.8 2.785 78.15 3.035 ;
      RECT 74.33 5.015 74.5 8.305 ;
      RECT 73.9 5.015 74.07 7.225 ;
      RECT 73.9 7.795 74.07 8.305 ;
      RECT 71.145 7.8 71.315 8.31 ;
      RECT 70.155 0.57 70.325 1.08 ;
      RECT 70.155 2.39 70.325 3.86 ;
      RECT 70.155 5.02 70.325 6.49 ;
      RECT 70.155 7.8 70.325 8.31 ;
      RECT 68.795 0.575 68.965 3.865 ;
      RECT 68.795 5.015 68.965 8.305 ;
      RECT 68.365 0.575 68.535 1.085 ;
      RECT 68.365 1.655 68.535 3.865 ;
      RECT 68.365 5.015 68.535 7.225 ;
      RECT 68.365 7.795 68.535 8.305 ;
      RECT 64.725 5.825 65.06 6.095 ;
      RECT 64.225 2.785 64.775 2.985 ;
      RECT 63.88 5.825 64.215 6.075 ;
      RECT 63.345 5.825 63.68 6.095 ;
      RECT 61.96 2.785 62.31 3.035 ;
      RECT 61.1 2.785 61.45 3.035 ;
      RECT 60.58 2.785 60.93 3.035 ;
      RECT 57.11 5.015 57.28 8.305 ;
      RECT 56.68 5.015 56.85 7.225 ;
      RECT 56.68 7.795 56.85 8.305 ;
      RECT 53.925 7.8 54.095 8.31 ;
      RECT 52.935 0.57 53.105 1.08 ;
      RECT 52.935 2.39 53.105 3.86 ;
      RECT 52.935 5.02 53.105 6.49 ;
      RECT 52.935 7.8 53.105 8.31 ;
      RECT 51.575 0.575 51.745 3.865 ;
      RECT 51.575 5.015 51.745 8.305 ;
      RECT 51.145 0.575 51.315 1.085 ;
      RECT 51.145 1.655 51.315 3.865 ;
      RECT 51.145 5.015 51.315 7.225 ;
      RECT 51.145 7.795 51.315 8.305 ;
      RECT 47.505 5.825 47.84 6.095 ;
      RECT 47.005 2.785 47.555 2.985 ;
      RECT 46.66 5.825 46.995 6.075 ;
      RECT 46.125 5.825 46.46 6.095 ;
      RECT 44.74 2.785 45.09 3.035 ;
      RECT 43.88 2.785 44.23 3.035 ;
      RECT 43.36 2.785 43.71 3.035 ;
      RECT 39.89 5.015 40.06 8.305 ;
      RECT 39.46 5.015 39.63 7.225 ;
      RECT 39.46 7.795 39.63 8.305 ;
      RECT 36.705 7.8 36.875 8.31 ;
      RECT 35.715 0.57 35.885 1.08 ;
      RECT 35.715 2.39 35.885 3.86 ;
      RECT 35.715 5.02 35.885 6.49 ;
      RECT 35.715 7.8 35.885 8.31 ;
      RECT 34.355 0.575 34.525 3.865 ;
      RECT 34.355 5.015 34.525 8.305 ;
      RECT 33.925 0.575 34.095 1.085 ;
      RECT 33.925 1.655 34.095 3.865 ;
      RECT 33.925 5.015 34.095 7.225 ;
      RECT 33.925 7.795 34.095 8.305 ;
      RECT 30.285 5.825 30.62 6.095 ;
      RECT 29.785 2.785 30.335 2.985 ;
      RECT 29.44 5.825 29.775 6.075 ;
      RECT 28.905 5.825 29.24 6.095 ;
      RECT 27.52 2.785 27.87 3.035 ;
      RECT 26.66 2.785 27.01 3.035 ;
      RECT 26.14 2.785 26.49 3.035 ;
      RECT 22.67 5.015 22.84 8.305 ;
      RECT 22.24 5.015 22.41 7.225 ;
      RECT 22.24 7.795 22.41 8.305 ;
      RECT 19.485 7.8 19.655 8.31 ;
      RECT 18.495 0.57 18.665 1.08 ;
      RECT 18.495 2.39 18.665 3.86 ;
      RECT 18.495 5.02 18.665 6.49 ;
      RECT 18.495 7.8 18.665 8.31 ;
      RECT 17.135 0.575 17.305 3.865 ;
      RECT 17.135 5.015 17.305 8.305 ;
      RECT 16.705 0.575 16.875 1.085 ;
      RECT 16.705 1.655 16.875 3.865 ;
      RECT 16.705 5.015 16.875 7.225 ;
      RECT 16.705 7.795 16.875 8.305 ;
      RECT 13.065 5.825 13.4 6.095 ;
      RECT 12.565 2.785 13.115 2.985 ;
      RECT 12.22 5.825 12.555 6.075 ;
      RECT 11.685 5.825 12.02 6.095 ;
      RECT 10.3 2.785 10.65 3.035 ;
      RECT 9.44 2.785 9.79 3.035 ;
      RECT 8.92 2.785 9.27 3.035 ;
      RECT 5.45 5.015 5.62 8.305 ;
      RECT 5.02 5.015 5.19 7.225 ;
      RECT 5.02 7.795 5.19 8.305 ;
      RECT 1.61 5.015 1.78 7.225 ;
      RECT 1.61 7.795 1.78 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r2 ;
  SIZE 88.9 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 19.48 0.915 19.65 1.085 ;
        RECT 19.475 0.91 19.645 1.08 ;
        RECT 19.475 2.39 19.645 2.56 ;
      LAYER li1 ;
        RECT 19.48 0.915 19.65 1.085 ;
        RECT 19.475 0.57 19.645 1.08 ;
        RECT 19.475 2.39 19.645 3.86 ;
      LAYER met1 ;
        RECT 19.415 2.36 19.705 2.59 ;
        RECT 19.415 0.88 19.705 1.11 ;
        RECT 19.475 0.88 19.645 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 36.7 0.915 36.87 1.085 ;
        RECT 36.695 0.91 36.865 1.08 ;
        RECT 36.695 2.39 36.865 2.56 ;
      LAYER li1 ;
        RECT 36.7 0.915 36.87 1.085 ;
        RECT 36.695 0.57 36.865 1.08 ;
        RECT 36.695 2.39 36.865 3.86 ;
      LAYER met1 ;
        RECT 36.635 2.36 36.925 2.59 ;
        RECT 36.635 0.88 36.925 1.11 ;
        RECT 36.695 0.88 36.865 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 53.92 0.915 54.09 1.085 ;
        RECT 53.915 0.91 54.085 1.08 ;
        RECT 53.915 2.39 54.085 2.56 ;
      LAYER li1 ;
        RECT 53.92 0.915 54.09 1.085 ;
        RECT 53.915 0.57 54.085 1.08 ;
        RECT 53.915 2.39 54.085 3.86 ;
      LAYER met1 ;
        RECT 53.855 2.36 54.145 2.59 ;
        RECT 53.855 0.88 54.145 1.11 ;
        RECT 53.915 0.88 54.085 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 71.14 0.915 71.31 1.085 ;
        RECT 71.135 0.91 71.305 1.08 ;
        RECT 71.135 2.39 71.305 2.56 ;
      LAYER li1 ;
        RECT 71.14 0.915 71.31 1.085 ;
        RECT 71.135 0.57 71.305 1.08 ;
        RECT 71.135 2.39 71.305 3.86 ;
      LAYER met1 ;
        RECT 71.075 2.36 71.365 2.59 ;
        RECT 71.075 0.88 71.365 1.11 ;
        RECT 71.135 0.88 71.305 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 88.36 0.915 88.53 1.085 ;
        RECT 88.355 0.91 88.525 1.08 ;
        RECT 88.355 2.39 88.525 2.56 ;
      LAYER li1 ;
        RECT 88.36 0.915 88.53 1.085 ;
        RECT 88.355 0.57 88.525 1.08 ;
        RECT 88.355 2.39 88.525 3.86 ;
      LAYER met1 ;
        RECT 88.295 2.36 88.585 2.59 ;
        RECT 88.295 0.88 88.585 1.11 ;
        RECT 88.355 0.88 88.525 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 15.325 1.66 15.495 2.935 ;
        RECT 15.325 5.94 15.495 7.22 ;
        RECT 15.315 5.94 15.495 6.18 ;
        RECT 3.64 5.945 3.81 7.22 ;
      LAYER met2 ;
        RECT 15.245 5.855 15.57 6.18 ;
        RECT 15.245 3.495 15.57 3.82 ;
        RECT 5.945 7.55 15.495 7.72 ;
        RECT 15.325 5.855 15.495 7.72 ;
        RECT 15.315 3.495 15.485 6.18 ;
        RECT 5.89 5.86 6.17 6.2 ;
        RECT 5.945 5.86 6.115 7.72 ;
      LAYER met1 ;
        RECT 15.265 2.765 15.725 2.935 ;
        RECT 15.245 3.495 15.57 3.82 ;
        RECT 15.265 2.735 15.555 2.965 ;
        RECT 15.325 2.735 15.495 3.82 ;
        RECT 15.245 5.945 15.725 6.115 ;
        RECT 15.245 5.855 15.57 6.18 ;
        RECT 5.86 5.89 6.2 6.17 ;
        RECT 3.58 5.945 6.2 6.115 ;
        RECT 3.58 5.915 3.87 6.145 ;
      LAYER mcon ;
        RECT 3.64 5.945 3.81 6.115 ;
        RECT 15.325 5.945 15.495 6.115 ;
        RECT 15.325 2.765 15.495 2.935 ;
      LAYER via1 ;
        RECT 5.955 5.955 6.105 6.105 ;
        RECT 15.335 5.94 15.485 6.09 ;
        RECT 15.335 3.58 15.485 3.73 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 32.545 1.66 32.715 2.935 ;
        RECT 32.545 5.94 32.715 7.22 ;
        RECT 32.535 5.94 32.715 6.18 ;
        RECT 20.86 5.945 21.03 7.22 ;
      LAYER met2 ;
        RECT 32.465 5.855 32.79 6.18 ;
        RECT 32.465 3.495 32.79 3.82 ;
        RECT 23.165 7.55 32.715 7.72 ;
        RECT 32.545 5.855 32.715 7.72 ;
        RECT 32.535 3.495 32.705 6.18 ;
        RECT 23.11 5.86 23.39 6.2 ;
        RECT 23.165 5.86 23.335 7.72 ;
      LAYER met1 ;
        RECT 32.485 2.765 32.945 2.935 ;
        RECT 32.465 3.495 32.79 3.82 ;
        RECT 32.485 2.735 32.775 2.965 ;
        RECT 32.545 2.735 32.715 3.82 ;
        RECT 32.465 5.945 32.945 6.115 ;
        RECT 32.465 5.855 32.79 6.18 ;
        RECT 23.08 5.89 23.42 6.17 ;
        RECT 20.8 5.945 23.42 6.115 ;
        RECT 20.8 5.915 21.09 6.145 ;
      LAYER mcon ;
        RECT 20.86 5.945 21.03 6.115 ;
        RECT 32.545 5.945 32.715 6.115 ;
        RECT 32.545 2.765 32.715 2.935 ;
      LAYER via1 ;
        RECT 23.175 5.955 23.325 6.105 ;
        RECT 32.555 5.94 32.705 6.09 ;
        RECT 32.555 3.58 32.705 3.73 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 49.765 1.66 49.935 2.935 ;
        RECT 49.765 5.94 49.935 7.22 ;
        RECT 49.755 5.94 49.935 6.18 ;
        RECT 38.08 5.945 38.25 7.22 ;
      LAYER met2 ;
        RECT 49.685 5.855 50.01 6.18 ;
        RECT 49.685 3.495 50.01 3.82 ;
        RECT 40.385 7.55 49.935 7.72 ;
        RECT 49.765 5.855 49.935 7.72 ;
        RECT 49.755 3.495 49.925 6.18 ;
        RECT 40.33 5.86 40.61 6.2 ;
        RECT 40.385 5.86 40.555 7.72 ;
      LAYER met1 ;
        RECT 49.705 2.765 50.165 2.935 ;
        RECT 49.685 3.495 50.01 3.82 ;
        RECT 49.705 2.735 49.995 2.965 ;
        RECT 49.765 2.735 49.935 3.82 ;
        RECT 49.685 5.945 50.165 6.115 ;
        RECT 49.685 5.855 50.01 6.18 ;
        RECT 40.3 5.89 40.64 6.17 ;
        RECT 38.02 5.945 40.64 6.115 ;
        RECT 38.02 5.915 38.31 6.145 ;
      LAYER mcon ;
        RECT 38.08 5.945 38.25 6.115 ;
        RECT 49.765 5.945 49.935 6.115 ;
        RECT 49.765 2.765 49.935 2.935 ;
      LAYER via1 ;
        RECT 40.395 5.955 40.545 6.105 ;
        RECT 49.775 5.94 49.925 6.09 ;
        RECT 49.775 3.58 49.925 3.73 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 66.985 1.66 67.155 2.935 ;
        RECT 66.985 5.94 67.155 7.22 ;
        RECT 66.975 5.94 67.155 6.18 ;
        RECT 55.3 5.945 55.47 7.22 ;
      LAYER met2 ;
        RECT 66.905 5.855 67.23 6.18 ;
        RECT 66.905 3.495 67.23 3.82 ;
        RECT 57.605 7.55 67.155 7.72 ;
        RECT 66.985 5.855 67.155 7.72 ;
        RECT 66.975 3.495 67.145 6.18 ;
        RECT 57.55 5.86 57.83 6.2 ;
        RECT 57.605 5.86 57.775 7.72 ;
      LAYER met1 ;
        RECT 66.925 2.765 67.385 2.935 ;
        RECT 66.905 3.495 67.23 3.82 ;
        RECT 66.925 2.735 67.215 2.965 ;
        RECT 66.985 2.735 67.155 3.82 ;
        RECT 66.905 5.945 67.385 6.115 ;
        RECT 66.905 5.855 67.23 6.18 ;
        RECT 57.52 5.89 57.86 6.17 ;
        RECT 55.24 5.945 57.86 6.115 ;
        RECT 55.24 5.915 55.53 6.145 ;
      LAYER mcon ;
        RECT 55.3 5.945 55.47 6.115 ;
        RECT 66.985 5.945 67.155 6.115 ;
        RECT 66.985 2.765 67.155 2.935 ;
      LAYER via1 ;
        RECT 57.615 5.955 57.765 6.105 ;
        RECT 66.995 5.94 67.145 6.09 ;
        RECT 66.995 3.58 67.145 3.73 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 84.205 1.66 84.375 2.935 ;
        RECT 84.205 5.94 84.375 7.22 ;
        RECT 84.195 5.94 84.375 6.18 ;
        RECT 72.52 5.945 72.69 7.22 ;
      LAYER met2 ;
        RECT 84.125 5.855 84.45 6.18 ;
        RECT 84.125 3.495 84.45 3.82 ;
        RECT 74.825 7.55 84.375 7.72 ;
        RECT 84.205 5.855 84.375 7.72 ;
        RECT 84.195 3.495 84.365 6.18 ;
        RECT 74.77 5.86 75.05 6.2 ;
        RECT 74.825 5.86 74.995 7.72 ;
      LAYER met1 ;
        RECT 84.145 2.765 84.605 2.935 ;
        RECT 84.125 3.495 84.45 3.82 ;
        RECT 84.145 2.735 84.435 2.965 ;
        RECT 84.205 2.735 84.375 3.82 ;
        RECT 84.125 5.945 84.605 6.115 ;
        RECT 84.125 5.855 84.45 6.18 ;
        RECT 74.74 5.89 75.08 6.17 ;
        RECT 72.46 5.945 75.08 6.115 ;
        RECT 72.46 5.915 72.75 6.145 ;
      LAYER mcon ;
        RECT 72.52 5.945 72.69 6.115 ;
        RECT 84.205 5.945 84.375 6.115 ;
        RECT 84.205 2.765 84.375 2.935 ;
      LAYER via1 ;
        RECT 74.835 5.955 74.985 6.105 ;
        RECT 84.215 5.94 84.365 6.09 ;
        RECT 84.215 3.58 84.365 3.73 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 5.945 0.4 7.22 ;
      LAYER met1 ;
        RECT 0.17 5.945 0.63 6.115 ;
        RECT 0.17 5.915 0.46 6.145 ;
      LAYER mcon ;
        RECT 0.23 5.945 0.4 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.34 4.255 2.145 4.635 ;
      LAYER li1 ;
        RECT 82.915 4.135 88.9 4.745 ;
        RECT 86.765 4.13 88.745 4.75 ;
        RECT 87.925 3.4 88.095 5.48 ;
        RECT 86.935 3.4 87.105 5.48 ;
        RECT 84.195 3.405 84.365 5.475 ;
        RECT 82.91 4.135 88.9 4.515 ;
        RECT 1.805 4.345 88.9 4.515 ;
        RECT 82 4.345 82.28 5.655 ;
        RECT 81.6 3.495 81.77 4.515 ;
        RECT 81.07 4.345 81.33 5.655 ;
        RECT 80.76 3.835 80.93 4.515 ;
        RECT 80.62 4.345 80.9 5.655 ;
        RECT 79.69 4.345 79.95 5.655 ;
        RECT 79.26 4.345 79.52 5.655 ;
        RECT 79.18 3.205 79.51 4.515 ;
        RECT 78.31 4.345 78.59 5.655 ;
        RECT 76.94 3.205 77.27 4.515 ;
        RECT 76.96 3.205 77.22 5.655 ;
        RECT 76.49 3.205 76.72 4.515 ;
        RECT 76.01 4.345 76.29 5.655 ;
        RECT 65.695 4.345 75.84 4.74 ;
        RECT 65.69 4.135 75.82 4.515 ;
        RECT 75.61 3.205 75.82 4.74 ;
        RECT 71.675 4.13 75.82 4.74 ;
        RECT 72.335 4.13 75.085 4.745 ;
        RECT 72.51 4.13 72.68 5.475 ;
        RECT 65.695 4.135 71.68 4.745 ;
        RECT 69.545 4.13 71.525 4.75 ;
        RECT 70.705 3.4 70.875 5.48 ;
        RECT 69.715 3.4 69.885 5.48 ;
        RECT 66.975 3.405 67.145 5.475 ;
        RECT 64.78 4.345 65.06 5.655 ;
        RECT 64.38 3.495 64.55 4.515 ;
        RECT 63.85 4.345 64.11 5.655 ;
        RECT 63.54 3.835 63.71 4.515 ;
        RECT 63.4 4.345 63.68 5.655 ;
        RECT 62.47 4.345 62.73 5.655 ;
        RECT 62.04 4.345 62.3 5.655 ;
        RECT 61.96 3.205 62.29 4.515 ;
        RECT 61.09 4.345 61.37 5.655 ;
        RECT 59.72 3.205 60.05 4.515 ;
        RECT 59.74 3.205 60 5.655 ;
        RECT 59.27 3.205 59.5 4.515 ;
        RECT 58.79 4.345 59.07 5.655 ;
        RECT 48.475 4.345 58.62 4.74 ;
        RECT 48.47 4.135 58.6 4.515 ;
        RECT 58.39 3.205 58.6 4.74 ;
        RECT 54.455 4.13 58.6 4.74 ;
        RECT 55.115 4.13 57.865 4.745 ;
        RECT 55.29 4.13 55.46 5.475 ;
        RECT 48.475 4.135 54.46 4.745 ;
        RECT 52.325 4.13 54.305 4.75 ;
        RECT 53.485 3.4 53.655 5.48 ;
        RECT 52.495 3.4 52.665 5.48 ;
        RECT 49.755 3.405 49.925 5.475 ;
        RECT 47.56 4.345 47.84 5.655 ;
        RECT 47.16 3.495 47.33 4.515 ;
        RECT 46.63 4.345 46.89 5.655 ;
        RECT 46.32 3.835 46.49 4.515 ;
        RECT 46.18 4.345 46.46 5.655 ;
        RECT 45.25 4.345 45.51 5.655 ;
        RECT 44.82 4.345 45.08 5.655 ;
        RECT 44.74 3.205 45.07 4.515 ;
        RECT 43.87 4.345 44.15 5.655 ;
        RECT 42.5 3.205 42.83 4.515 ;
        RECT 42.52 3.205 42.78 5.655 ;
        RECT 42.05 3.205 42.28 4.515 ;
        RECT 41.57 4.345 41.85 5.655 ;
        RECT 31.255 4.345 41.4 4.74 ;
        RECT 31.25 4.135 41.38 4.515 ;
        RECT 41.17 3.205 41.38 4.74 ;
        RECT 37.235 4.13 41.38 4.74 ;
        RECT 37.895 4.13 40.645 4.745 ;
        RECT 38.07 4.13 38.24 5.475 ;
        RECT 31.255 4.135 37.24 4.745 ;
        RECT 35.105 4.13 37.085 4.75 ;
        RECT 36.265 3.4 36.435 5.48 ;
        RECT 35.275 3.4 35.445 5.48 ;
        RECT 32.535 3.405 32.705 5.475 ;
        RECT 30.34 4.345 30.62 5.655 ;
        RECT 29.94 3.495 30.11 4.515 ;
        RECT 29.41 4.345 29.67 5.655 ;
        RECT 29.1 3.835 29.27 4.515 ;
        RECT 28.96 4.345 29.24 5.655 ;
        RECT 28.03 4.345 28.29 5.655 ;
        RECT 27.6 4.345 27.86 5.655 ;
        RECT 27.52 3.205 27.85 4.515 ;
        RECT 26.65 4.345 26.93 5.655 ;
        RECT 25.28 3.205 25.61 4.515 ;
        RECT 25.3 3.205 25.56 5.655 ;
        RECT 24.83 3.205 25.06 4.515 ;
        RECT 24.35 4.345 24.63 5.655 ;
        RECT 14.035 4.345 24.18 4.74 ;
        RECT 14.03 4.135 24.16 4.515 ;
        RECT 23.95 3.205 24.16 4.74 ;
        RECT 20.015 4.13 24.16 4.74 ;
        RECT 20.675 4.13 23.425 4.745 ;
        RECT 20.85 4.13 21.02 5.475 ;
        RECT 14.035 4.135 20.02 4.745 ;
        RECT 17.885 4.13 19.865 4.75 ;
        RECT 19.045 3.4 19.215 5.48 ;
        RECT 18.055 3.4 18.225 5.48 ;
        RECT 15.315 3.405 15.485 5.475 ;
        RECT 13.12 4.345 13.4 5.655 ;
        RECT 12.72 3.495 12.89 4.515 ;
        RECT 12.19 4.345 12.45 5.655 ;
        RECT 11.88 3.835 12.05 4.515 ;
        RECT 11.74 4.345 12.02 5.655 ;
        RECT 10.81 4.345 11.07 5.655 ;
        RECT 10.38 4.345 10.64 5.655 ;
        RECT 10.3 3.205 10.63 4.515 ;
        RECT 9.43 4.345 9.71 5.655 ;
        RECT 8.06 3.205 8.39 4.515 ;
        RECT 8.08 3.205 8.34 5.655 ;
        RECT 7.61 3.205 7.84 4.515 ;
        RECT 7.13 4.345 7.41 5.655 ;
        RECT 0 4.44 6.96 4.74 ;
        RECT 1.805 4.13 6.94 4.74 ;
        RECT 6.73 3.205 6.94 4.74 ;
        RECT 3.455 4.13 6.205 4.745 ;
        RECT 3.63 4.13 3.8 5.475 ;
        RECT 0.045 4.44 2.795 4.745 ;
        RECT 2.03 4.13 2.2 8.305 ;
        RECT 0 4.13 6.94 4.33 ;
        RECT 0 4.13 1.635 4.74 ;
        RECT 0.22 4.13 0.39 5.475 ;
      LAYER met2 ;
        RECT 1.53 4.255 1.91 4.635 ;
      LAYER met1 ;
        RECT 82.915 4.135 88.9 4.745 ;
        RECT 86.765 4.13 88.745 4.75 ;
        RECT 0 4.19 88.9 4.67 ;
        RECT 82.91 4.135 88.9 4.67 ;
        RECT 65.695 4.19 75.84 4.74 ;
        RECT 65.69 4.135 75.82 4.67 ;
        RECT 71.675 4.13 75.82 4.74 ;
        RECT 72.335 4.13 75.085 4.745 ;
        RECT 65.695 4.135 71.68 4.745 ;
        RECT 69.545 4.13 71.525 4.75 ;
        RECT 48.475 4.19 58.62 4.74 ;
        RECT 48.47 4.135 58.6 4.67 ;
        RECT 54.455 4.13 58.6 4.74 ;
        RECT 55.115 4.13 57.865 4.745 ;
        RECT 48.475 4.135 54.46 4.745 ;
        RECT 52.325 4.13 54.305 4.75 ;
        RECT 31.255 4.19 41.4 4.74 ;
        RECT 31.25 4.135 41.38 4.67 ;
        RECT 37.235 4.13 41.38 4.74 ;
        RECT 37.895 4.13 40.645 4.745 ;
        RECT 31.255 4.135 37.24 4.745 ;
        RECT 35.105 4.13 37.085 4.75 ;
        RECT 14.035 4.19 24.18 4.74 ;
        RECT 14.03 4.135 24.16 4.67 ;
        RECT 20.015 4.13 24.16 4.74 ;
        RECT 20.675 4.13 23.425 4.745 ;
        RECT 14.035 4.135 20.02 4.745 ;
        RECT 17.885 4.13 19.865 4.75 ;
        RECT 0 4.19 6.96 4.74 ;
        RECT 0 4.13 6.94 4.74 ;
        RECT 3.455 4.13 6.205 4.745 ;
        RECT 0.045 4.13 2.795 4.745 ;
        RECT 1.97 6.655 2.26 6.885 ;
        RECT 1.8 6.685 2.26 6.855 ;
      LAYER via2 ;
        RECT 1.62 4.345 1.82 4.545 ;
      LAYER mcon ;
        RECT 2.03 6.685 2.2 6.855 ;
        RECT 2.34 4.545 2.51 4.715 ;
        RECT 5.75 4.545 5.92 4.715 ;
        RECT 6.73 4.345 6.9 4.515 ;
        RECT 7.19 4.345 7.36 4.515 ;
        RECT 7.65 4.345 7.82 4.515 ;
        RECT 8.11 4.345 8.28 4.515 ;
        RECT 8.57 4.345 8.74 4.515 ;
        RECT 9.03 4.345 9.2 4.515 ;
        RECT 9.49 4.345 9.66 4.515 ;
        RECT 9.95 4.345 10.12 4.515 ;
        RECT 10.41 4.345 10.58 4.515 ;
        RECT 10.87 4.345 11.04 4.515 ;
        RECT 11.33 4.345 11.5 4.515 ;
        RECT 11.79 4.345 11.96 4.515 ;
        RECT 12.25 4.345 12.42 4.515 ;
        RECT 12.71 4.345 12.88 4.515 ;
        RECT 13.17 4.345 13.34 4.515 ;
        RECT 13.63 4.345 13.8 4.515 ;
        RECT 17.435 4.545 17.605 4.715 ;
        RECT 17.435 4.165 17.605 4.335 ;
        RECT 18.135 4.55 18.305 4.72 ;
        RECT 18.135 4.16 18.305 4.33 ;
        RECT 19.125 4.55 19.295 4.72 ;
        RECT 19.125 4.16 19.295 4.33 ;
        RECT 22.97 4.545 23.14 4.715 ;
        RECT 23.95 4.345 24.12 4.515 ;
        RECT 24.41 4.345 24.58 4.515 ;
        RECT 24.87 4.345 25.04 4.515 ;
        RECT 25.33 4.345 25.5 4.515 ;
        RECT 25.79 4.345 25.96 4.515 ;
        RECT 26.25 4.345 26.42 4.515 ;
        RECT 26.71 4.345 26.88 4.515 ;
        RECT 27.17 4.345 27.34 4.515 ;
        RECT 27.63 4.345 27.8 4.515 ;
        RECT 28.09 4.345 28.26 4.515 ;
        RECT 28.55 4.345 28.72 4.515 ;
        RECT 29.01 4.345 29.18 4.515 ;
        RECT 29.47 4.345 29.64 4.515 ;
        RECT 29.93 4.345 30.1 4.515 ;
        RECT 30.39 4.345 30.56 4.515 ;
        RECT 30.85 4.345 31.02 4.515 ;
        RECT 34.655 4.545 34.825 4.715 ;
        RECT 34.655 4.165 34.825 4.335 ;
        RECT 35.355 4.55 35.525 4.72 ;
        RECT 35.355 4.16 35.525 4.33 ;
        RECT 36.345 4.55 36.515 4.72 ;
        RECT 36.345 4.16 36.515 4.33 ;
        RECT 40.19 4.545 40.36 4.715 ;
        RECT 41.17 4.345 41.34 4.515 ;
        RECT 41.63 4.345 41.8 4.515 ;
        RECT 42.09 4.345 42.26 4.515 ;
        RECT 42.55 4.345 42.72 4.515 ;
        RECT 43.01 4.345 43.18 4.515 ;
        RECT 43.47 4.345 43.64 4.515 ;
        RECT 43.93 4.345 44.1 4.515 ;
        RECT 44.39 4.345 44.56 4.515 ;
        RECT 44.85 4.345 45.02 4.515 ;
        RECT 45.31 4.345 45.48 4.515 ;
        RECT 45.77 4.345 45.94 4.515 ;
        RECT 46.23 4.345 46.4 4.515 ;
        RECT 46.69 4.345 46.86 4.515 ;
        RECT 47.15 4.345 47.32 4.515 ;
        RECT 47.61 4.345 47.78 4.515 ;
        RECT 48.07 4.345 48.24 4.515 ;
        RECT 51.875 4.545 52.045 4.715 ;
        RECT 51.875 4.165 52.045 4.335 ;
        RECT 52.575 4.55 52.745 4.72 ;
        RECT 52.575 4.16 52.745 4.33 ;
        RECT 53.565 4.55 53.735 4.72 ;
        RECT 53.565 4.16 53.735 4.33 ;
        RECT 57.41 4.545 57.58 4.715 ;
        RECT 58.39 4.345 58.56 4.515 ;
        RECT 58.85 4.345 59.02 4.515 ;
        RECT 59.31 4.345 59.48 4.515 ;
        RECT 59.77 4.345 59.94 4.515 ;
        RECT 60.23 4.345 60.4 4.515 ;
        RECT 60.69 4.345 60.86 4.515 ;
        RECT 61.15 4.345 61.32 4.515 ;
        RECT 61.61 4.345 61.78 4.515 ;
        RECT 62.07 4.345 62.24 4.515 ;
        RECT 62.53 4.345 62.7 4.515 ;
        RECT 62.99 4.345 63.16 4.515 ;
        RECT 63.45 4.345 63.62 4.515 ;
        RECT 63.91 4.345 64.08 4.515 ;
        RECT 64.37 4.345 64.54 4.515 ;
        RECT 64.83 4.345 65 4.515 ;
        RECT 65.29 4.345 65.46 4.515 ;
        RECT 69.095 4.545 69.265 4.715 ;
        RECT 69.095 4.165 69.265 4.335 ;
        RECT 69.795 4.55 69.965 4.72 ;
        RECT 69.795 4.16 69.965 4.33 ;
        RECT 70.785 4.55 70.955 4.72 ;
        RECT 70.785 4.16 70.955 4.33 ;
        RECT 74.63 4.545 74.8 4.715 ;
        RECT 75.61 4.345 75.78 4.515 ;
        RECT 76.07 4.345 76.24 4.515 ;
        RECT 76.53 4.345 76.7 4.515 ;
        RECT 76.99 4.345 77.16 4.515 ;
        RECT 77.45 4.345 77.62 4.515 ;
        RECT 77.91 4.345 78.08 4.515 ;
        RECT 78.37 4.345 78.54 4.515 ;
        RECT 78.83 4.345 79 4.515 ;
        RECT 79.29 4.345 79.46 4.515 ;
        RECT 79.75 4.345 79.92 4.515 ;
        RECT 80.21 4.345 80.38 4.515 ;
        RECT 80.67 4.345 80.84 4.515 ;
        RECT 81.13 4.345 81.3 4.515 ;
        RECT 81.59 4.345 81.76 4.515 ;
        RECT 82.05 4.345 82.22 4.515 ;
        RECT 82.51 4.345 82.68 4.515 ;
        RECT 86.315 4.545 86.485 4.715 ;
        RECT 86.315 4.165 86.485 4.335 ;
        RECT 87.015 4.55 87.185 4.72 ;
        RECT 87.015 4.16 87.185 4.33 ;
        RECT 88.005 4.55 88.175 4.72 ;
        RECT 88.005 4.16 88.175 4.33 ;
      LAYER via1 ;
        RECT 1.645 4.37 1.795 4.52 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 77.85 5.79 78.18 6.12 ;
        RECT 77.38 5.805 78.18 6.105 ;
        RECT 60.63 5.79 60.96 6.12 ;
        RECT 60.16 5.805 60.96 6.105 ;
        RECT 43.41 5.79 43.74 6.12 ;
        RECT 42.94 5.805 43.74 6.105 ;
        RECT 26.19 5.79 26.52 6.12 ;
        RECT 25.72 5.805 26.52 6.105 ;
        RECT 8.97 5.79 9.3 6.12 ;
        RECT 8.5 5.805 9.3 6.105 ;
        RECT 0.005 8.5 0.81 8.88 ;
        RECT 0 0 0.805 0.38 ;
      LAYER li1 ;
        RECT 88.72 0 88.9 0.305 ;
        RECT 0.465 0 88.9 0.3 ;
        RECT 87.925 0 88.095 0.93 ;
        RECT 86.935 0 87.105 0.93 ;
        RECT 71.5 0 86.77 0.305 ;
        RECT 84.195 0 84.365 0.935 ;
        RECT 75.465 0 83.12 1.795 ;
        RECT 82.36 0 82.69 2.185 ;
        RECT 81.52 0 81.85 2.185 ;
        RECT 79.69 0 79.98 2.63 ;
        RECT 79.24 0 79.51 2.605 ;
        RECT 78.33 0 78.57 2.605 ;
        RECT 77.88 0 78.12 2.605 ;
        RECT 76.94 0 77.21 2.605 ;
        RECT 76.49 0 76.72 2.615 ;
        RECT 75.61 0 75.82 2.615 ;
        RECT 75.46 0 83.12 1.635 ;
        RECT 70.705 0 70.875 0.93 ;
        RECT 69.715 0 69.885 0.93 ;
        RECT 54.28 0 69.55 0.305 ;
        RECT 66.975 0 67.145 0.935 ;
        RECT 58.245 0 65.9 1.795 ;
        RECT 65.14 0 65.47 2.185 ;
        RECT 64.3 0 64.63 2.185 ;
        RECT 62.47 0 62.76 2.63 ;
        RECT 62.02 0 62.29 2.605 ;
        RECT 61.11 0 61.35 2.605 ;
        RECT 60.66 0 60.9 2.605 ;
        RECT 59.72 0 59.99 2.605 ;
        RECT 59.27 0 59.5 2.615 ;
        RECT 58.39 0 58.6 2.615 ;
        RECT 58.24 0 65.9 1.635 ;
        RECT 53.485 0 53.655 0.93 ;
        RECT 52.495 0 52.665 0.93 ;
        RECT 37.06 0 52.33 0.305 ;
        RECT 49.755 0 49.925 0.935 ;
        RECT 41.025 0 48.68 1.795 ;
        RECT 47.92 0 48.25 2.185 ;
        RECT 47.08 0 47.41 2.185 ;
        RECT 45.25 0 45.54 2.63 ;
        RECT 44.8 0 45.07 2.605 ;
        RECT 43.89 0 44.13 2.605 ;
        RECT 43.44 0 43.68 2.605 ;
        RECT 42.5 0 42.77 2.605 ;
        RECT 42.05 0 42.28 2.615 ;
        RECT 41.17 0 41.38 2.615 ;
        RECT 41.02 0 48.68 1.635 ;
        RECT 36.265 0 36.435 0.93 ;
        RECT 35.275 0 35.445 0.93 ;
        RECT 19.84 0 35.11 0.305 ;
        RECT 32.535 0 32.705 0.935 ;
        RECT 23.805 0 31.46 1.795 ;
        RECT 30.7 0 31.03 2.185 ;
        RECT 29.86 0 30.19 2.185 ;
        RECT 28.03 0 28.32 2.63 ;
        RECT 27.58 0 27.85 2.605 ;
        RECT 26.67 0 26.91 2.605 ;
        RECT 26.22 0 26.46 2.605 ;
        RECT 25.28 0 25.55 2.605 ;
        RECT 24.83 0 25.06 2.615 ;
        RECT 23.95 0 24.16 2.615 ;
        RECT 23.8 0 31.46 1.635 ;
        RECT 19.045 0 19.215 0.93 ;
        RECT 18.055 0 18.225 0.93 ;
        RECT 0 0.245 17.89 0.305 ;
        RECT 15.315 0 15.485 0.935 ;
        RECT 6.585 0 14.24 1.795 ;
        RECT 13.48 0 13.81 2.185 ;
        RECT 12.64 0 12.97 2.185 ;
        RECT 10.81 0 11.1 2.63 ;
        RECT 10.36 0 10.63 2.605 ;
        RECT 9.45 0 9.69 2.605 ;
        RECT 9 0 9.24 2.605 ;
        RECT 8.06 0 8.33 2.605 ;
        RECT 7.61 0 7.84 2.615 ;
        RECT 6.73 0 6.94 2.615 ;
        RECT 6.58 0 14.24 1.635 ;
        RECT 0 0.245 0.805 0.315 ;
        RECT 0.295 0.245 0.465 0.335 ;
        RECT 0 0 88.9 0.075 ;
        RECT 0 0 0.295 0.315 ;
        RECT 0 8.58 88.9 8.88 ;
        RECT 88.72 8.575 88.9 8.88 ;
        RECT 87.925 7.95 88.095 8.88 ;
        RECT 86.935 7.95 87.105 8.88 ;
        RECT 71.5 8.575 86.77 8.88 ;
        RECT 84.195 7.945 84.365 8.88 ;
        RECT 75.735 7.18 82.935 8.88 ;
        RECT 75.465 7.065 82.825 7.235 ;
        RECT 81.97 6.265 82.28 8.88 ;
        RECT 80.59 6.265 80.9 8.88 ;
        RECT 78.32 5.825 78.655 6.095 ;
        RECT 78.31 6.265 78.62 8.88 ;
        RECT 77.93 5.875 78.655 6.045 ;
        RECT 77.94 5.875 78.11 8.88 ;
        RECT 76.01 6.265 76.32 8.88 ;
        RECT 72.51 7.945 72.68 8.88 ;
        RECT 70.705 7.95 70.875 8.88 ;
        RECT 69.715 7.95 69.885 8.88 ;
        RECT 54.28 8.575 69.55 8.88 ;
        RECT 66.975 7.945 67.145 8.88 ;
        RECT 58.515 7.18 65.715 8.88 ;
        RECT 58.245 7.065 65.605 7.235 ;
        RECT 64.75 6.265 65.06 8.88 ;
        RECT 63.37 6.265 63.68 8.88 ;
        RECT 61.1 5.825 61.435 6.095 ;
        RECT 61.09 6.265 61.4 8.88 ;
        RECT 60.71 5.875 61.435 6.045 ;
        RECT 60.72 5.875 60.89 8.88 ;
        RECT 58.79 6.265 59.1 8.88 ;
        RECT 55.29 7.945 55.46 8.88 ;
        RECT 53.485 7.95 53.655 8.88 ;
        RECT 52.495 7.95 52.665 8.88 ;
        RECT 37.06 8.575 52.33 8.88 ;
        RECT 49.755 7.945 49.925 8.88 ;
        RECT 41.295 7.18 48.495 8.88 ;
        RECT 41.025 7.065 48.385 7.235 ;
        RECT 47.53 6.265 47.84 8.88 ;
        RECT 46.15 6.265 46.46 8.88 ;
        RECT 43.88 5.825 44.215 6.095 ;
        RECT 43.87 6.265 44.18 8.88 ;
        RECT 43.49 5.875 44.215 6.045 ;
        RECT 43.5 5.875 43.67 8.88 ;
        RECT 41.57 6.265 41.88 8.88 ;
        RECT 38.07 7.945 38.24 8.88 ;
        RECT 36.265 7.95 36.435 8.88 ;
        RECT 35.275 7.95 35.445 8.88 ;
        RECT 19.84 8.575 35.11 8.88 ;
        RECT 32.535 7.945 32.705 8.88 ;
        RECT 24.075 7.18 31.275 8.88 ;
        RECT 23.805 7.065 31.165 7.235 ;
        RECT 30.31 6.265 30.62 8.88 ;
        RECT 28.93 6.265 29.24 8.88 ;
        RECT 26.66 5.825 26.995 6.095 ;
        RECT 26.65 6.265 26.96 8.88 ;
        RECT 26.27 5.875 26.995 6.045 ;
        RECT 26.28 5.875 26.45 8.88 ;
        RECT 24.35 6.265 24.66 8.88 ;
        RECT 20.85 7.945 21.02 8.88 ;
        RECT 19.045 7.95 19.215 8.88 ;
        RECT 18.055 7.95 18.225 8.88 ;
        RECT 0 8.575 17.89 8.88 ;
        RECT 15.315 7.945 15.485 8.88 ;
        RECT 6.855 7.18 14.055 8.88 ;
        RECT 6.585 7.065 13.945 7.235 ;
        RECT 13.09 6.265 13.4 8.88 ;
        RECT 11.71 6.265 12.02 8.88 ;
        RECT 9.44 5.825 9.775 6.095 ;
        RECT 9.43 6.265 9.74 8.88 ;
        RECT 9.05 5.875 9.775 6.045 ;
        RECT 9.06 5.875 9.23 8.88 ;
        RECT 7.13 6.265 7.44 8.88 ;
        RECT 3.63 7.945 3.8 8.88 ;
        RECT 0.005 8.565 0.81 8.88 ;
        RECT 0.22 8.545 0.47 8.88 ;
        RECT 0.22 7.945 0.39 8.88 ;
        RECT 76.02 5.825 76.355 6.095 ;
        RECT 75.55 5.875 76.355 6.045 ;
        RECT 73.515 6.075 73.685 8.025 ;
        RECT 73.46 7.855 73.63 8.305 ;
        RECT 73.46 5.015 73.63 6.245 ;
        RECT 58.8 5.825 59.135 6.095 ;
        RECT 58.33 5.875 59.135 6.045 ;
        RECT 56.295 6.075 56.465 8.025 ;
        RECT 56.24 7.855 56.41 8.305 ;
        RECT 56.24 5.015 56.41 6.245 ;
        RECT 41.58 5.825 41.915 6.095 ;
        RECT 41.11 5.875 41.915 6.045 ;
        RECT 39.075 6.075 39.245 8.025 ;
        RECT 39.02 7.855 39.19 8.305 ;
        RECT 39.02 5.015 39.19 6.245 ;
        RECT 24.36 5.825 24.695 6.095 ;
        RECT 23.89 5.875 24.695 6.045 ;
        RECT 21.855 6.075 22.025 8.025 ;
        RECT 21.8 7.855 21.97 8.305 ;
        RECT 21.8 5.015 21.97 6.245 ;
        RECT 7.14 5.825 7.475 6.095 ;
        RECT 6.67 5.875 7.475 6.045 ;
        RECT 4.635 6.075 4.805 8.025 ;
        RECT 4.58 7.855 4.75 8.305 ;
        RECT 4.58 5.015 4.75 6.245 ;
      LAYER met2 ;
        RECT 77.875 5.77 78.155 6.14 ;
        RECT 60.655 5.77 60.935 6.14 ;
        RECT 43.435 5.77 43.715 6.14 ;
        RECT 26.215 5.77 26.495 6.14 ;
        RECT 8.995 5.77 9.275 6.14 ;
        RECT 0.195 8.5 0.575 8.88 ;
        RECT 0.19 0 0.57 0.38 ;
        RECT 0.235 0 0.39 8.88 ;
      LAYER met1 ;
        RECT 88.72 0 88.9 0.305 ;
        RECT 0 0 88.9 0.3 ;
        RECT 71.5 0 86.77 0.305 ;
        RECT 75.465 0 83.12 1.795 ;
        RECT 75.465 0 82.825 1.95 ;
        RECT 75.46 0 83.12 1.635 ;
        RECT 54.28 0 69.55 0.305 ;
        RECT 58.245 0 65.9 1.795 ;
        RECT 58.245 0 65.605 1.95 ;
        RECT 58.24 0 65.9 1.635 ;
        RECT 37.06 0 52.33 0.305 ;
        RECT 41.025 0 48.68 1.795 ;
        RECT 41.025 0 48.385 1.95 ;
        RECT 41.02 0 48.68 1.635 ;
        RECT 19.84 0 35.11 0.305 ;
        RECT 23.805 0 31.46 1.795 ;
        RECT 23.805 0 31.165 1.95 ;
        RECT 23.8 0 31.46 1.635 ;
        RECT 0 0 17.89 0.305 ;
        RECT 6.585 0 14.24 1.795 ;
        RECT 6.585 0 13.945 1.95 ;
        RECT 6.58 0 14.24 1.635 ;
        RECT 0 0 0.805 0.315 ;
        RECT 0.205 0 0.555 0.335 ;
        RECT 0 8.58 88.9 8.88 ;
        RECT 88.72 8.575 88.9 8.88 ;
        RECT 71.5 8.575 86.77 8.88 ;
        RECT 75.735 7.18 82.935 8.88 ;
        RECT 75.465 6.91 82.825 7.39 ;
        RECT 73.455 6.285 73.745 6.515 ;
        RECT 73.055 6.315 73.745 6.485 ;
        RECT 73.055 6.315 73.225 8.88 ;
        RECT 54.28 8.575 69.55 8.88 ;
        RECT 58.515 7.18 65.715 8.88 ;
        RECT 58.245 6.91 65.605 7.39 ;
        RECT 56.235 6.285 56.525 6.515 ;
        RECT 55.835 6.315 56.525 6.485 ;
        RECT 55.835 6.315 56.005 8.88 ;
        RECT 37.06 8.575 52.33 8.88 ;
        RECT 41.295 7.18 48.495 8.88 ;
        RECT 41.025 6.91 48.385 7.39 ;
        RECT 39.015 6.285 39.305 6.515 ;
        RECT 38.615 6.315 39.305 6.485 ;
        RECT 38.615 6.315 38.785 8.88 ;
        RECT 19.84 8.575 35.11 8.88 ;
        RECT 24.075 7.18 31.275 8.88 ;
        RECT 23.805 6.91 31.165 7.39 ;
        RECT 21.795 6.285 22.085 6.515 ;
        RECT 21.395 6.315 22.085 6.485 ;
        RECT 21.395 6.315 21.565 8.88 ;
        RECT 0 8.575 17.89 8.88 ;
        RECT 6.855 7.18 14.055 8.88 ;
        RECT 6.585 6.91 13.945 7.39 ;
        RECT 4.575 6.285 4.865 6.515 ;
        RECT 4.175 6.315 4.865 6.485 ;
        RECT 4.175 6.315 4.345 8.88 ;
        RECT 0.005 8.565 0.81 8.88 ;
        RECT 0.21 8.545 0.56 8.88 ;
        RECT 77.855 5.83 78.175 6.09 ;
        RECT 75.49 5.89 78.175 6.03 ;
        RECT 75.49 5.845 75.78 6.075 ;
        RECT 60.635 5.83 60.955 6.09 ;
        RECT 58.27 5.89 60.955 6.03 ;
        RECT 58.27 5.845 58.56 6.075 ;
        RECT 43.415 5.83 43.735 6.09 ;
        RECT 41.05 5.89 43.735 6.03 ;
        RECT 41.05 5.845 41.34 6.075 ;
        RECT 26.195 5.83 26.515 6.09 ;
        RECT 23.83 5.89 26.515 6.03 ;
        RECT 23.83 5.845 24.12 6.075 ;
        RECT 8.975 5.83 9.295 6.09 ;
        RECT 6.61 5.89 9.295 6.03 ;
        RECT 6.61 5.845 6.9 6.075 ;
      LAYER via2 ;
        RECT 0.28 0.09 0.48 0.29 ;
        RECT 0.285 8.59 0.485 8.79 ;
        RECT 9.035 5.855 9.235 6.055 ;
        RECT 26.255 5.855 26.455 6.055 ;
        RECT 43.475 5.855 43.675 6.055 ;
        RECT 60.695 5.855 60.895 6.055 ;
        RECT 77.915 5.855 78.115 6.055 ;
      LAYER mcon ;
        RECT 0.3 8.605 0.47 8.775 ;
        RECT 0.98 8.605 1.15 8.775 ;
        RECT 1.66 8.605 1.83 8.775 ;
        RECT 2.34 8.605 2.51 8.775 ;
        RECT 3.71 8.605 3.88 8.775 ;
        RECT 4.39 8.605 4.56 8.775 ;
        RECT 4.635 6.315 4.805 6.485 ;
        RECT 5.07 8.605 5.24 8.775 ;
        RECT 5.75 8.605 5.92 8.775 ;
        RECT 6.67 5.875 6.84 6.045 ;
        RECT 6.73 7.065 6.9 7.235 ;
        RECT 6.73 1.625 6.9 1.795 ;
        RECT 7.19 7.065 7.36 7.235 ;
        RECT 7.19 1.625 7.36 1.795 ;
        RECT 7.65 7.065 7.82 7.235 ;
        RECT 7.65 1.625 7.82 1.795 ;
        RECT 8.11 7.065 8.28 7.235 ;
        RECT 8.11 1.625 8.28 1.795 ;
        RECT 8.57 7.065 8.74 7.235 ;
        RECT 8.57 1.625 8.74 1.795 ;
        RECT 9.03 7.065 9.2 7.235 ;
        RECT 9.03 1.625 9.2 1.795 ;
        RECT 9.05 5.875 9.22 6.045 ;
        RECT 9.49 7.065 9.66 7.235 ;
        RECT 9.49 1.625 9.66 1.795 ;
        RECT 9.95 7.065 10.12 7.235 ;
        RECT 9.95 1.625 10.12 1.795 ;
        RECT 10.41 7.065 10.58 7.235 ;
        RECT 10.41 1.625 10.58 1.795 ;
        RECT 10.87 7.065 11.04 7.235 ;
        RECT 10.87 1.625 11.04 1.795 ;
        RECT 11.33 7.065 11.5 7.235 ;
        RECT 11.33 1.625 11.5 1.795 ;
        RECT 11.79 7.065 11.96 7.235 ;
        RECT 11.79 1.625 11.96 1.795 ;
        RECT 12.25 7.065 12.42 7.235 ;
        RECT 12.25 1.625 12.42 1.795 ;
        RECT 12.71 7.065 12.88 7.235 ;
        RECT 12.71 1.625 12.88 1.795 ;
        RECT 13.17 7.065 13.34 7.235 ;
        RECT 13.17 1.625 13.34 1.795 ;
        RECT 13.63 7.065 13.8 7.235 ;
        RECT 13.63 1.625 13.8 1.795 ;
        RECT 15.395 8.605 15.565 8.775 ;
        RECT 15.395 0.105 15.565 0.275 ;
        RECT 16.075 8.605 16.245 8.775 ;
        RECT 16.075 0.105 16.245 0.275 ;
        RECT 16.755 8.605 16.925 8.775 ;
        RECT 16.755 0.105 16.925 0.275 ;
        RECT 17.435 8.605 17.605 8.775 ;
        RECT 17.435 0.105 17.605 0.275 ;
        RECT 18.135 8.61 18.305 8.78 ;
        RECT 18.135 0.1 18.305 0.27 ;
        RECT 19.125 8.61 19.295 8.78 ;
        RECT 19.125 0.1 19.295 0.27 ;
        RECT 20.93 8.605 21.1 8.775 ;
        RECT 21.61 8.605 21.78 8.775 ;
        RECT 21.855 6.315 22.025 6.485 ;
        RECT 22.29 8.605 22.46 8.775 ;
        RECT 22.97 8.605 23.14 8.775 ;
        RECT 23.89 5.875 24.06 6.045 ;
        RECT 23.95 7.065 24.12 7.235 ;
        RECT 23.95 1.625 24.12 1.795 ;
        RECT 24.41 7.065 24.58 7.235 ;
        RECT 24.41 1.625 24.58 1.795 ;
        RECT 24.87 7.065 25.04 7.235 ;
        RECT 24.87 1.625 25.04 1.795 ;
        RECT 25.33 7.065 25.5 7.235 ;
        RECT 25.33 1.625 25.5 1.795 ;
        RECT 25.79 7.065 25.96 7.235 ;
        RECT 25.79 1.625 25.96 1.795 ;
        RECT 26.25 7.065 26.42 7.235 ;
        RECT 26.25 1.625 26.42 1.795 ;
        RECT 26.27 5.875 26.44 6.045 ;
        RECT 26.71 7.065 26.88 7.235 ;
        RECT 26.71 1.625 26.88 1.795 ;
        RECT 27.17 7.065 27.34 7.235 ;
        RECT 27.17 1.625 27.34 1.795 ;
        RECT 27.63 7.065 27.8 7.235 ;
        RECT 27.63 1.625 27.8 1.795 ;
        RECT 28.09 7.065 28.26 7.235 ;
        RECT 28.09 1.625 28.26 1.795 ;
        RECT 28.55 7.065 28.72 7.235 ;
        RECT 28.55 1.625 28.72 1.795 ;
        RECT 29.01 7.065 29.18 7.235 ;
        RECT 29.01 1.625 29.18 1.795 ;
        RECT 29.47 7.065 29.64 7.235 ;
        RECT 29.47 1.625 29.64 1.795 ;
        RECT 29.93 7.065 30.1 7.235 ;
        RECT 29.93 1.625 30.1 1.795 ;
        RECT 30.39 7.065 30.56 7.235 ;
        RECT 30.39 1.625 30.56 1.795 ;
        RECT 30.85 7.065 31.02 7.235 ;
        RECT 30.85 1.625 31.02 1.795 ;
        RECT 32.615 8.605 32.785 8.775 ;
        RECT 32.615 0.105 32.785 0.275 ;
        RECT 33.295 8.605 33.465 8.775 ;
        RECT 33.295 0.105 33.465 0.275 ;
        RECT 33.975 8.605 34.145 8.775 ;
        RECT 33.975 0.105 34.145 0.275 ;
        RECT 34.655 8.605 34.825 8.775 ;
        RECT 34.655 0.105 34.825 0.275 ;
        RECT 35.355 8.61 35.525 8.78 ;
        RECT 35.355 0.1 35.525 0.27 ;
        RECT 36.345 8.61 36.515 8.78 ;
        RECT 36.345 0.1 36.515 0.27 ;
        RECT 38.15 8.605 38.32 8.775 ;
        RECT 38.83 8.605 39 8.775 ;
        RECT 39.075 6.315 39.245 6.485 ;
        RECT 39.51 8.605 39.68 8.775 ;
        RECT 40.19 8.605 40.36 8.775 ;
        RECT 41.11 5.875 41.28 6.045 ;
        RECT 41.17 7.065 41.34 7.235 ;
        RECT 41.17 1.625 41.34 1.795 ;
        RECT 41.63 7.065 41.8 7.235 ;
        RECT 41.63 1.625 41.8 1.795 ;
        RECT 42.09 7.065 42.26 7.235 ;
        RECT 42.09 1.625 42.26 1.795 ;
        RECT 42.55 7.065 42.72 7.235 ;
        RECT 42.55 1.625 42.72 1.795 ;
        RECT 43.01 7.065 43.18 7.235 ;
        RECT 43.01 1.625 43.18 1.795 ;
        RECT 43.47 7.065 43.64 7.235 ;
        RECT 43.47 1.625 43.64 1.795 ;
        RECT 43.49 5.875 43.66 6.045 ;
        RECT 43.93 7.065 44.1 7.235 ;
        RECT 43.93 1.625 44.1 1.795 ;
        RECT 44.39 7.065 44.56 7.235 ;
        RECT 44.39 1.625 44.56 1.795 ;
        RECT 44.85 7.065 45.02 7.235 ;
        RECT 44.85 1.625 45.02 1.795 ;
        RECT 45.31 7.065 45.48 7.235 ;
        RECT 45.31 1.625 45.48 1.795 ;
        RECT 45.77 7.065 45.94 7.235 ;
        RECT 45.77 1.625 45.94 1.795 ;
        RECT 46.23 7.065 46.4 7.235 ;
        RECT 46.23 1.625 46.4 1.795 ;
        RECT 46.69 7.065 46.86 7.235 ;
        RECT 46.69 1.625 46.86 1.795 ;
        RECT 47.15 7.065 47.32 7.235 ;
        RECT 47.15 1.625 47.32 1.795 ;
        RECT 47.61 7.065 47.78 7.235 ;
        RECT 47.61 1.625 47.78 1.795 ;
        RECT 48.07 7.065 48.24 7.235 ;
        RECT 48.07 1.625 48.24 1.795 ;
        RECT 49.835 8.605 50.005 8.775 ;
        RECT 49.835 0.105 50.005 0.275 ;
        RECT 50.515 8.605 50.685 8.775 ;
        RECT 50.515 0.105 50.685 0.275 ;
        RECT 51.195 8.605 51.365 8.775 ;
        RECT 51.195 0.105 51.365 0.275 ;
        RECT 51.875 8.605 52.045 8.775 ;
        RECT 51.875 0.105 52.045 0.275 ;
        RECT 52.575 8.61 52.745 8.78 ;
        RECT 52.575 0.1 52.745 0.27 ;
        RECT 53.565 8.61 53.735 8.78 ;
        RECT 53.565 0.1 53.735 0.27 ;
        RECT 55.37 8.605 55.54 8.775 ;
        RECT 56.05 8.605 56.22 8.775 ;
        RECT 56.295 6.315 56.465 6.485 ;
        RECT 56.73 8.605 56.9 8.775 ;
        RECT 57.41 8.605 57.58 8.775 ;
        RECT 58.33 5.875 58.5 6.045 ;
        RECT 58.39 7.065 58.56 7.235 ;
        RECT 58.39 1.625 58.56 1.795 ;
        RECT 58.85 7.065 59.02 7.235 ;
        RECT 58.85 1.625 59.02 1.795 ;
        RECT 59.31 7.065 59.48 7.235 ;
        RECT 59.31 1.625 59.48 1.795 ;
        RECT 59.77 7.065 59.94 7.235 ;
        RECT 59.77 1.625 59.94 1.795 ;
        RECT 60.23 7.065 60.4 7.235 ;
        RECT 60.23 1.625 60.4 1.795 ;
        RECT 60.69 7.065 60.86 7.235 ;
        RECT 60.69 1.625 60.86 1.795 ;
        RECT 60.71 5.875 60.88 6.045 ;
        RECT 61.15 7.065 61.32 7.235 ;
        RECT 61.15 1.625 61.32 1.795 ;
        RECT 61.61 7.065 61.78 7.235 ;
        RECT 61.61 1.625 61.78 1.795 ;
        RECT 62.07 7.065 62.24 7.235 ;
        RECT 62.07 1.625 62.24 1.795 ;
        RECT 62.53 7.065 62.7 7.235 ;
        RECT 62.53 1.625 62.7 1.795 ;
        RECT 62.99 7.065 63.16 7.235 ;
        RECT 62.99 1.625 63.16 1.795 ;
        RECT 63.45 7.065 63.62 7.235 ;
        RECT 63.45 1.625 63.62 1.795 ;
        RECT 63.91 7.065 64.08 7.235 ;
        RECT 63.91 1.625 64.08 1.795 ;
        RECT 64.37 7.065 64.54 7.235 ;
        RECT 64.37 1.625 64.54 1.795 ;
        RECT 64.83 7.065 65 7.235 ;
        RECT 64.83 1.625 65 1.795 ;
        RECT 65.29 7.065 65.46 7.235 ;
        RECT 65.29 1.625 65.46 1.795 ;
        RECT 67.055 8.605 67.225 8.775 ;
        RECT 67.055 0.105 67.225 0.275 ;
        RECT 67.735 8.605 67.905 8.775 ;
        RECT 67.735 0.105 67.905 0.275 ;
        RECT 68.415 8.605 68.585 8.775 ;
        RECT 68.415 0.105 68.585 0.275 ;
        RECT 69.095 8.605 69.265 8.775 ;
        RECT 69.095 0.105 69.265 0.275 ;
        RECT 69.795 8.61 69.965 8.78 ;
        RECT 69.795 0.1 69.965 0.27 ;
        RECT 70.785 8.61 70.955 8.78 ;
        RECT 70.785 0.1 70.955 0.27 ;
        RECT 72.59 8.605 72.76 8.775 ;
        RECT 73.27 8.605 73.44 8.775 ;
        RECT 73.515 6.315 73.685 6.485 ;
        RECT 73.95 8.605 74.12 8.775 ;
        RECT 74.63 8.605 74.8 8.775 ;
        RECT 75.55 5.875 75.72 6.045 ;
        RECT 75.61 7.065 75.78 7.235 ;
        RECT 75.61 1.625 75.78 1.795 ;
        RECT 76.07 7.065 76.24 7.235 ;
        RECT 76.07 1.625 76.24 1.795 ;
        RECT 76.53 7.065 76.7 7.235 ;
        RECT 76.53 1.625 76.7 1.795 ;
        RECT 76.99 7.065 77.16 7.235 ;
        RECT 76.99 1.625 77.16 1.795 ;
        RECT 77.45 7.065 77.62 7.235 ;
        RECT 77.45 1.625 77.62 1.795 ;
        RECT 77.91 7.065 78.08 7.235 ;
        RECT 77.91 1.625 78.08 1.795 ;
        RECT 77.93 5.875 78.1 6.045 ;
        RECT 78.37 7.065 78.54 7.235 ;
        RECT 78.37 1.625 78.54 1.795 ;
        RECT 78.83 7.065 79 7.235 ;
        RECT 78.83 1.625 79 1.795 ;
        RECT 79.29 7.065 79.46 7.235 ;
        RECT 79.29 1.625 79.46 1.795 ;
        RECT 79.75 7.065 79.92 7.235 ;
        RECT 79.75 1.625 79.92 1.795 ;
        RECT 80.21 7.065 80.38 7.235 ;
        RECT 80.21 1.625 80.38 1.795 ;
        RECT 80.67 7.065 80.84 7.235 ;
        RECT 80.67 1.625 80.84 1.795 ;
        RECT 81.13 7.065 81.3 7.235 ;
        RECT 81.13 1.625 81.3 1.795 ;
        RECT 81.59 7.065 81.76 7.235 ;
        RECT 81.59 1.625 81.76 1.795 ;
        RECT 82.05 7.065 82.22 7.235 ;
        RECT 82.05 1.625 82.22 1.795 ;
        RECT 82.51 7.065 82.68 7.235 ;
        RECT 82.51 1.625 82.68 1.795 ;
        RECT 84.275 8.605 84.445 8.775 ;
        RECT 84.275 0.105 84.445 0.275 ;
        RECT 84.955 8.605 85.125 8.775 ;
        RECT 84.955 0.105 85.125 0.275 ;
        RECT 85.635 8.605 85.805 8.775 ;
        RECT 85.635 0.105 85.805 0.275 ;
        RECT 86.315 8.605 86.485 8.775 ;
        RECT 86.315 0.105 86.485 0.275 ;
        RECT 87.015 8.61 87.185 8.78 ;
        RECT 87.015 0.1 87.185 0.27 ;
        RECT 88.005 8.61 88.175 8.78 ;
        RECT 88.005 0.1 88.175 0.27 ;
      LAYER via1 ;
        RECT 0.305 0.115 0.455 0.265 ;
        RECT 0.31 8.615 0.46 8.765 ;
        RECT 9.06 5.885 9.21 6.035 ;
        RECT 26.28 5.885 26.43 6.035 ;
        RECT 43.5 5.885 43.65 6.035 ;
        RECT 60.72 5.885 60.87 6.035 ;
        RECT 77.94 5.885 78.09 6.035 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 74.93 7.435 80.945 7.735 ;
      RECT 80.645 5.805 80.945 7.735 ;
      RECT 79.59 5.785 79.89 7.735 ;
      RECT 78.56 6.48 78.86 7.735 ;
      RECT 74.93 7.035 75.23 7.735 ;
      RECT 73.795 7 74.165 7.37 ;
      RECT 73.795 7.035 75.23 7.335 ;
      RECT 78.53 6.48 78.86 6.81 ;
      RECT 78.06 6.495 78.86 6.795 ;
      RECT 78.44 6.455 78.74 6.795 ;
      RECT 80.57 5.805 80.945 6.17 ;
      RECT 80.635 5.765 80.935 6.17 ;
      RECT 79.55 5.785 79.89 6.135 ;
      RECT 79.565 5.745 79.865 6.135 ;
      RECT 79.54 5.79 79.89 6.12 ;
      RECT 80.57 5.805 81.38 6.105 ;
      RECT 79.07 5.805 79.89 6.105 ;
      RECT 80.58 5.79 80.935 6.17 ;
      RECT 80.23 3.755 80.56 4.085 ;
      RECT 80.23 3.77 81.03 4.07 ;
      RECT 80.245 3.725 80.545 4.085 ;
      RECT 79.89 3.075 80.22 3.405 ;
      RECT 79.89 3.09 80.69 3.39 ;
      RECT 79.975 3.065 80.275 3.39 ;
      RECT 79.21 4.155 79.54 4.485 ;
      RECT 77.17 4.155 77.5 4.485 ;
      RECT 77.17 4.17 79.54 4.47 ;
      RECT 78.86 3.415 79.19 3.745 ;
      RECT 78.4 3.43 79.2 3.73 ;
      RECT 78.53 2.225 78.86 2.555 ;
      RECT 78.06 2.24 78.86 2.54 ;
      RECT 78.52 2.235 78.86 2.54 ;
      RECT 57.71 7.435 63.725 7.735 ;
      RECT 63.425 5.805 63.725 7.735 ;
      RECT 62.37 5.785 62.67 7.735 ;
      RECT 61.34 6.48 61.64 7.735 ;
      RECT 57.71 7.035 58.01 7.735 ;
      RECT 56.575 7 56.945 7.37 ;
      RECT 56.575 7.035 58.01 7.335 ;
      RECT 61.31 6.48 61.64 6.81 ;
      RECT 60.84 6.495 61.64 6.795 ;
      RECT 61.22 6.455 61.52 6.795 ;
      RECT 63.35 5.805 63.725 6.17 ;
      RECT 63.415 5.765 63.715 6.17 ;
      RECT 62.33 5.785 62.67 6.135 ;
      RECT 62.345 5.745 62.645 6.135 ;
      RECT 62.32 5.79 62.67 6.12 ;
      RECT 63.35 5.805 64.16 6.105 ;
      RECT 61.85 5.805 62.67 6.105 ;
      RECT 63.36 5.79 63.715 6.17 ;
      RECT 63.01 3.755 63.34 4.085 ;
      RECT 63.01 3.77 63.81 4.07 ;
      RECT 63.025 3.725 63.325 4.085 ;
      RECT 62.67 3.075 63 3.405 ;
      RECT 62.67 3.09 63.47 3.39 ;
      RECT 62.755 3.065 63.055 3.39 ;
      RECT 61.99 4.155 62.32 4.485 ;
      RECT 59.95 4.155 60.28 4.485 ;
      RECT 59.95 4.17 62.32 4.47 ;
      RECT 61.64 3.415 61.97 3.745 ;
      RECT 61.18 3.43 61.98 3.73 ;
      RECT 61.31 2.225 61.64 2.555 ;
      RECT 60.84 2.24 61.64 2.54 ;
      RECT 61.3 2.235 61.64 2.54 ;
      RECT 40.49 7.435 46.505 7.735 ;
      RECT 46.205 5.805 46.505 7.735 ;
      RECT 45.15 5.785 45.45 7.735 ;
      RECT 44.12 6.48 44.42 7.735 ;
      RECT 40.49 7.035 40.79 7.735 ;
      RECT 39.355 7 39.725 7.37 ;
      RECT 39.355 7.035 40.79 7.335 ;
      RECT 44.09 6.48 44.42 6.81 ;
      RECT 43.62 6.495 44.42 6.795 ;
      RECT 44 6.455 44.3 6.795 ;
      RECT 46.13 5.805 46.505 6.17 ;
      RECT 46.195 5.765 46.495 6.17 ;
      RECT 45.11 5.785 45.45 6.135 ;
      RECT 45.125 5.745 45.425 6.135 ;
      RECT 45.1 5.79 45.45 6.12 ;
      RECT 46.13 5.805 46.94 6.105 ;
      RECT 44.63 5.805 45.45 6.105 ;
      RECT 46.14 5.79 46.495 6.17 ;
      RECT 45.79 3.755 46.12 4.085 ;
      RECT 45.79 3.77 46.59 4.07 ;
      RECT 45.805 3.725 46.105 4.085 ;
      RECT 45.45 3.075 45.78 3.405 ;
      RECT 45.45 3.09 46.25 3.39 ;
      RECT 45.535 3.065 45.835 3.39 ;
      RECT 44.77 4.155 45.1 4.485 ;
      RECT 42.73 4.155 43.06 4.485 ;
      RECT 42.73 4.17 45.1 4.47 ;
      RECT 44.42 3.415 44.75 3.745 ;
      RECT 43.96 3.43 44.76 3.73 ;
      RECT 44.09 2.225 44.42 2.555 ;
      RECT 43.62 2.24 44.42 2.54 ;
      RECT 44.08 2.235 44.42 2.54 ;
      RECT 23.27 7.435 29.285 7.735 ;
      RECT 28.985 5.805 29.285 7.735 ;
      RECT 27.93 5.785 28.23 7.735 ;
      RECT 26.9 6.48 27.2 7.735 ;
      RECT 23.27 7.035 23.57 7.735 ;
      RECT 22.135 7 22.505 7.37 ;
      RECT 22.135 7.035 23.57 7.335 ;
      RECT 26.87 6.48 27.2 6.81 ;
      RECT 26.4 6.495 27.2 6.795 ;
      RECT 26.78 6.455 27.08 6.795 ;
      RECT 28.91 5.805 29.285 6.17 ;
      RECT 28.975 5.765 29.275 6.17 ;
      RECT 27.89 5.785 28.23 6.135 ;
      RECT 27.905 5.745 28.205 6.135 ;
      RECT 27.88 5.79 28.23 6.12 ;
      RECT 28.91 5.805 29.72 6.105 ;
      RECT 27.41 5.805 28.23 6.105 ;
      RECT 28.92 5.79 29.275 6.17 ;
      RECT 28.57 3.755 28.9 4.085 ;
      RECT 28.57 3.77 29.37 4.07 ;
      RECT 28.585 3.725 28.885 4.085 ;
      RECT 28.23 3.075 28.56 3.405 ;
      RECT 28.23 3.09 29.03 3.39 ;
      RECT 28.315 3.065 28.615 3.39 ;
      RECT 27.55 4.155 27.88 4.485 ;
      RECT 25.51 4.155 25.84 4.485 ;
      RECT 25.51 4.17 27.88 4.47 ;
      RECT 27.2 3.415 27.53 3.745 ;
      RECT 26.74 3.43 27.54 3.73 ;
      RECT 26.87 2.225 27.2 2.555 ;
      RECT 26.4 2.24 27.2 2.54 ;
      RECT 26.86 2.235 27.2 2.54 ;
      RECT 6.05 7.435 12.065 7.735 ;
      RECT 11.765 5.805 12.065 7.735 ;
      RECT 10.71 5.785 11.01 7.735 ;
      RECT 9.68 6.48 9.98 7.735 ;
      RECT 6.05 7.035 6.35 7.735 ;
      RECT 4.915 7 5.285 7.37 ;
      RECT 4.915 7.035 6.35 7.335 ;
      RECT 9.65 6.48 9.98 6.81 ;
      RECT 9.18 6.495 9.98 6.795 ;
      RECT 9.56 6.455 9.86 6.795 ;
      RECT 11.69 5.805 12.065 6.17 ;
      RECT 11.755 5.765 12.055 6.17 ;
      RECT 10.67 5.785 11.01 6.135 ;
      RECT 10.685 5.745 10.985 6.135 ;
      RECT 10.66 5.79 11.01 6.12 ;
      RECT 11.69 5.805 12.5 6.105 ;
      RECT 10.19 5.805 11.01 6.105 ;
      RECT 11.7 5.79 12.055 6.17 ;
      RECT 11.35 3.755 11.68 4.085 ;
      RECT 11.35 3.77 12.15 4.07 ;
      RECT 11.365 3.725 11.665 4.085 ;
      RECT 11.01 3.075 11.34 3.405 ;
      RECT 11.01 3.09 11.81 3.39 ;
      RECT 11.095 3.065 11.395 3.39 ;
      RECT 10.33 4.155 10.66 4.485 ;
      RECT 8.29 4.155 8.62 4.485 ;
      RECT 8.29 4.17 10.66 4.47 ;
      RECT 9.98 3.415 10.31 3.745 ;
      RECT 9.52 3.43 10.32 3.73 ;
      RECT 9.65 2.225 9.98 2.555 ;
      RECT 9.18 2.24 9.98 2.54 ;
      RECT 9.64 2.235 9.98 2.54 ;
    LAYER via2 ;
      RECT 80.645 5.855 80.845 6.055 ;
      RECT 80.295 3.82 80.495 4.02 ;
      RECT 79.955 3.14 80.155 3.34 ;
      RECT 79.605 5.855 79.805 6.055 ;
      RECT 79.275 4.22 79.475 4.42 ;
      RECT 78.925 3.48 79.125 3.68 ;
      RECT 78.595 2.29 78.795 2.49 ;
      RECT 78.595 6.545 78.795 6.745 ;
      RECT 77.235 4.22 77.435 4.42 ;
      RECT 73.88 7.085 74.08 7.285 ;
      RECT 63.425 5.855 63.625 6.055 ;
      RECT 63.075 3.82 63.275 4.02 ;
      RECT 62.735 3.14 62.935 3.34 ;
      RECT 62.385 5.855 62.585 6.055 ;
      RECT 62.055 4.22 62.255 4.42 ;
      RECT 61.705 3.48 61.905 3.68 ;
      RECT 61.375 2.29 61.575 2.49 ;
      RECT 61.375 6.545 61.575 6.745 ;
      RECT 60.015 4.22 60.215 4.42 ;
      RECT 56.66 7.085 56.86 7.285 ;
      RECT 46.205 5.855 46.405 6.055 ;
      RECT 45.855 3.82 46.055 4.02 ;
      RECT 45.515 3.14 45.715 3.34 ;
      RECT 45.165 5.855 45.365 6.055 ;
      RECT 44.835 4.22 45.035 4.42 ;
      RECT 44.485 3.48 44.685 3.68 ;
      RECT 44.155 2.29 44.355 2.49 ;
      RECT 44.155 6.545 44.355 6.745 ;
      RECT 42.795 4.22 42.995 4.42 ;
      RECT 39.44 7.085 39.64 7.285 ;
      RECT 28.985 5.855 29.185 6.055 ;
      RECT 28.635 3.82 28.835 4.02 ;
      RECT 28.295 3.14 28.495 3.34 ;
      RECT 27.945 5.855 28.145 6.055 ;
      RECT 27.615 4.22 27.815 4.42 ;
      RECT 27.265 3.48 27.465 3.68 ;
      RECT 26.935 2.29 27.135 2.49 ;
      RECT 26.935 6.545 27.135 6.745 ;
      RECT 25.575 4.22 25.775 4.42 ;
      RECT 22.22 7.085 22.42 7.285 ;
      RECT 11.765 5.855 11.965 6.055 ;
      RECT 11.415 3.82 11.615 4.02 ;
      RECT 11.075 3.14 11.275 3.34 ;
      RECT 10.725 5.855 10.925 6.055 ;
      RECT 10.395 4.22 10.595 4.42 ;
      RECT 10.045 3.48 10.245 3.68 ;
      RECT 9.715 2.29 9.915 2.49 ;
      RECT 9.715 6.545 9.915 6.745 ;
      RECT 8.355 4.22 8.555 4.42 ;
      RECT 5 7.085 5.2 7.285 ;
    LAYER met2 ;
      RECT 1.21 8.6 88.53 8.77 ;
      RECT 88.36 7.3 88.53 8.77 ;
      RECT 1.21 6.255 1.38 8.77 ;
      RECT 88.325 7.3 88.65 7.625 ;
      RECT 1.165 6.255 1.445 6.595 ;
      RECT 85.17 6.28 85.49 6.605 ;
      RECT 85.2 5.695 85.37 6.605 ;
      RECT 85.2 5.695 85.375 6.045 ;
      RECT 85.2 5.695 86.175 5.87 ;
      RECT 86 1.965 86.175 5.87 ;
      RECT 78.555 2.205 78.835 2.575 ;
      RECT 78.555 2.345 83.205 2.52 ;
      RECT 83.03 2.025 83.205 2.52 ;
      RECT 83.5 1.995 83.825 2.32 ;
      RECT 85.945 1.965 86.295 2.315 ;
      RECT 83.03 2.025 86.295 2.195 ;
      RECT 74.32 8.29 85.015 8.46 ;
      RECT 84.855 2.395 85.015 8.46 ;
      RECT 74.32 6.545 74.49 8.46 ;
      RECT 85.97 6.655 86.295 6.98 ;
      RECT 71.14 6.655 71.465 6.98 ;
      RECT 84.855 6.745 86.295 6.915 ;
      RECT 74.27 6.545 74.55 6.885 ;
      RECT 71.14 6.685 74.55 6.855 ;
      RECT 85.17 2.365 85.49 2.685 ;
      RECT 84.855 2.395 85.49 2.565 ;
      RECT 81.625 6.48 81.885 6.8 ;
      RECT 81.685 2.74 81.825 6.8 ;
      RECT 81.625 2.74 81.885 3.06 ;
      RECT 80.945 4.78 81.205 5.1 ;
      RECT 81.005 3.76 81.145 5.1 ;
      RECT 80.945 3.76 81.205 4.08 ;
      RECT 79.925 6.48 80.185 6.8 ;
      RECT 79.985 5.21 80.125 6.8 ;
      RECT 79.305 5.21 80.125 5.35 ;
      RECT 79.305 2.74 79.445 5.35 ;
      RECT 79.235 4.135 79.515 4.505 ;
      RECT 79.245 2.74 79.505 3.06 ;
      RECT 77.195 4.135 77.475 4.505 ;
      RECT 77.265 2.4 77.405 4.505 ;
      RECT 77.205 2.4 77.465 2.72 ;
      RECT 76.525 4.78 76.785 5.1 ;
      RECT 76.585 2.74 76.725 5.1 ;
      RECT 76.525 2.74 76.785 3.06 ;
      RECT 67.95 6.28 68.27 6.605 ;
      RECT 67.98 5.695 68.15 6.605 ;
      RECT 67.98 5.695 68.155 6.045 ;
      RECT 67.98 5.695 68.955 5.87 ;
      RECT 68.78 1.965 68.955 5.87 ;
      RECT 61.335 2.205 61.615 2.575 ;
      RECT 61.335 2.345 65.985 2.52 ;
      RECT 65.81 2.025 65.985 2.52 ;
      RECT 66.28 1.995 66.605 2.32 ;
      RECT 68.725 1.965 69.075 2.315 ;
      RECT 65.81 2.025 69.075 2.195 ;
      RECT 57.1 8.29 67.795 8.46 ;
      RECT 67.635 2.395 67.795 8.46 ;
      RECT 57.1 6.545 57.27 8.46 ;
      RECT 68.75 6.655 69.075 6.98 ;
      RECT 53.92 6.655 54.245 6.98 ;
      RECT 67.635 6.745 69.075 6.915 ;
      RECT 57.05 6.545 57.33 6.885 ;
      RECT 53.92 6.685 57.33 6.855 ;
      RECT 67.95 2.365 68.27 2.685 ;
      RECT 67.635 2.395 68.27 2.565 ;
      RECT 64.405 6.48 64.665 6.8 ;
      RECT 64.465 2.74 64.605 6.8 ;
      RECT 64.405 2.74 64.665 3.06 ;
      RECT 63.725 4.78 63.985 5.1 ;
      RECT 63.785 3.76 63.925 5.1 ;
      RECT 63.725 3.76 63.985 4.08 ;
      RECT 62.705 6.48 62.965 6.8 ;
      RECT 62.765 5.21 62.905 6.8 ;
      RECT 62.085 5.21 62.905 5.35 ;
      RECT 62.085 2.74 62.225 5.35 ;
      RECT 62.015 4.135 62.295 4.505 ;
      RECT 62.025 2.74 62.285 3.06 ;
      RECT 59.975 4.135 60.255 4.505 ;
      RECT 60.045 2.4 60.185 4.505 ;
      RECT 59.985 2.4 60.245 2.72 ;
      RECT 59.305 4.78 59.565 5.1 ;
      RECT 59.365 2.74 59.505 5.1 ;
      RECT 59.305 2.74 59.565 3.06 ;
      RECT 50.73 6.28 51.05 6.605 ;
      RECT 50.76 5.695 50.93 6.605 ;
      RECT 50.76 5.695 50.935 6.045 ;
      RECT 50.76 5.695 51.735 5.87 ;
      RECT 51.56 1.965 51.735 5.87 ;
      RECT 44.115 2.205 44.395 2.575 ;
      RECT 44.115 2.345 48.765 2.52 ;
      RECT 48.59 2.025 48.765 2.52 ;
      RECT 49.06 1.995 49.385 2.32 ;
      RECT 51.505 1.965 51.855 2.315 ;
      RECT 48.59 2.025 51.855 2.195 ;
      RECT 39.88 8.29 50.575 8.46 ;
      RECT 50.415 2.395 50.575 8.46 ;
      RECT 39.88 6.545 40.05 8.46 ;
      RECT 51.53 6.655 51.855 6.98 ;
      RECT 36.7 6.655 37.025 6.98 ;
      RECT 50.415 6.745 51.855 6.915 ;
      RECT 39.83 6.545 40.11 6.885 ;
      RECT 36.7 6.685 40.12 6.855 ;
      RECT 50.73 2.365 51.05 2.685 ;
      RECT 50.415 2.395 51.05 2.565 ;
      RECT 47.185 6.48 47.445 6.8 ;
      RECT 47.245 2.74 47.385 6.8 ;
      RECT 47.185 2.74 47.445 3.06 ;
      RECT 46.505 4.78 46.765 5.1 ;
      RECT 46.565 3.76 46.705 5.1 ;
      RECT 46.505 3.76 46.765 4.08 ;
      RECT 45.485 6.48 45.745 6.8 ;
      RECT 45.545 5.21 45.685 6.8 ;
      RECT 44.865 5.21 45.685 5.35 ;
      RECT 44.865 2.74 45.005 5.35 ;
      RECT 44.795 4.135 45.075 4.505 ;
      RECT 44.805 2.74 45.065 3.06 ;
      RECT 42.755 4.135 43.035 4.505 ;
      RECT 42.825 2.4 42.965 4.505 ;
      RECT 42.765 2.4 43.025 2.72 ;
      RECT 42.085 4.78 42.345 5.1 ;
      RECT 42.145 2.74 42.285 5.1 ;
      RECT 42.085 2.74 42.345 3.06 ;
      RECT 33.51 6.28 33.83 6.605 ;
      RECT 33.54 5.695 33.71 6.605 ;
      RECT 33.54 5.695 33.715 6.045 ;
      RECT 33.54 5.695 34.515 5.87 ;
      RECT 34.34 1.965 34.515 5.87 ;
      RECT 26.895 2.205 27.175 2.575 ;
      RECT 26.895 2.345 31.545 2.52 ;
      RECT 31.37 2.025 31.545 2.52 ;
      RECT 31.84 1.995 32.165 2.32 ;
      RECT 34.285 1.965 34.635 2.315 ;
      RECT 31.37 2.025 34.635 2.195 ;
      RECT 22.66 8.29 33.355 8.46 ;
      RECT 33.195 2.395 33.355 8.46 ;
      RECT 22.66 6.545 22.83 8.46 ;
      RECT 34.31 6.655 34.635 6.98 ;
      RECT 19.48 6.655 19.805 6.98 ;
      RECT 33.195 6.745 34.635 6.915 ;
      RECT 22.61 6.545 22.89 6.885 ;
      RECT 19.48 6.685 22.89 6.855 ;
      RECT 33.51 2.365 33.83 2.685 ;
      RECT 33.195 2.395 33.83 2.565 ;
      RECT 29.965 6.48 30.225 6.8 ;
      RECT 30.025 2.74 30.165 6.8 ;
      RECT 29.965 2.74 30.225 3.06 ;
      RECT 29.285 4.78 29.545 5.1 ;
      RECT 29.345 3.76 29.485 5.1 ;
      RECT 29.285 3.76 29.545 4.08 ;
      RECT 28.265 6.48 28.525 6.8 ;
      RECT 28.325 5.21 28.465 6.8 ;
      RECT 27.645 5.21 28.465 5.35 ;
      RECT 27.645 2.74 27.785 5.35 ;
      RECT 27.575 4.135 27.855 4.505 ;
      RECT 27.585 2.74 27.845 3.06 ;
      RECT 25.535 4.135 25.815 4.505 ;
      RECT 25.605 2.4 25.745 4.505 ;
      RECT 25.545 2.4 25.805 2.72 ;
      RECT 24.865 4.78 25.125 5.1 ;
      RECT 24.925 2.74 25.065 5.1 ;
      RECT 24.865 2.74 25.125 3.06 ;
      RECT 16.29 6.28 16.61 6.605 ;
      RECT 16.32 5.695 16.49 6.605 ;
      RECT 16.32 5.695 16.495 6.045 ;
      RECT 16.32 5.695 17.295 5.87 ;
      RECT 17.12 1.965 17.295 5.87 ;
      RECT 9.675 2.205 9.955 2.575 ;
      RECT 9.675 2.345 14.325 2.52 ;
      RECT 14.15 2.025 14.325 2.52 ;
      RECT 14.62 1.995 14.945 2.32 ;
      RECT 17.065 1.965 17.415 2.315 ;
      RECT 14.15 2.025 17.415 2.195 ;
      RECT 5.44 8.29 16.135 8.46 ;
      RECT 15.975 2.395 16.135 8.46 ;
      RECT 5.44 6.545 5.61 8.46 ;
      RECT 1.54 6.995 1.82 7.335 ;
      RECT 1.54 7.06 2.745 7.23 ;
      RECT 2.575 6.685 2.745 7.23 ;
      RECT 17.09 6.655 17.415 6.98 ;
      RECT 15.975 6.745 17.415 6.915 ;
      RECT 5.39 6.545 5.67 6.885 ;
      RECT 2.575 6.685 5.67 6.855 ;
      RECT 16.29 2.365 16.61 2.685 ;
      RECT 15.975 2.395 16.61 2.565 ;
      RECT 12.745 6.48 13.005 6.8 ;
      RECT 12.805 2.74 12.945 6.8 ;
      RECT 12.745 2.74 13.005 3.06 ;
      RECT 12.065 4.78 12.325 5.1 ;
      RECT 12.125 3.76 12.265 5.1 ;
      RECT 12.065 3.76 12.325 4.08 ;
      RECT 11.045 6.48 11.305 6.8 ;
      RECT 11.105 5.21 11.245 6.8 ;
      RECT 10.425 5.21 11.245 5.35 ;
      RECT 10.425 2.74 10.565 5.35 ;
      RECT 10.355 4.135 10.635 4.505 ;
      RECT 10.365 2.74 10.625 3.06 ;
      RECT 8.315 4.135 8.595 4.505 ;
      RECT 8.385 2.4 8.525 4.505 ;
      RECT 8.325 2.4 8.585 2.72 ;
      RECT 7.645 4.78 7.905 5.1 ;
      RECT 7.705 2.74 7.845 5.1 ;
      RECT 7.645 2.74 7.905 3.06 ;
      RECT 80.605 5.77 80.885 6.14 ;
      RECT 80.255 3.735 80.535 4.105 ;
      RECT 79.915 3.055 80.195 3.425 ;
      RECT 79.565 5.77 79.845 6.14 ;
      RECT 78.885 3.395 79.165 3.765 ;
      RECT 78.555 6.46 78.835 6.83 ;
      RECT 73.795 7 74.165 7.37 ;
      RECT 63.385 5.77 63.665 6.14 ;
      RECT 63.035 3.735 63.315 4.105 ;
      RECT 62.695 3.055 62.975 3.425 ;
      RECT 62.345 5.77 62.625 6.14 ;
      RECT 61.665 3.395 61.945 3.765 ;
      RECT 61.335 6.46 61.615 6.83 ;
      RECT 56.575 7 56.945 7.37 ;
      RECT 46.165 5.77 46.445 6.14 ;
      RECT 45.815 3.735 46.095 4.105 ;
      RECT 45.475 3.055 45.755 3.425 ;
      RECT 45.125 5.77 45.405 6.14 ;
      RECT 44.445 3.395 44.725 3.765 ;
      RECT 44.115 6.46 44.395 6.83 ;
      RECT 39.355 7 39.725 7.37 ;
      RECT 28.945 5.77 29.225 6.14 ;
      RECT 28.595 3.735 28.875 4.105 ;
      RECT 28.255 3.055 28.535 3.425 ;
      RECT 27.905 5.77 28.185 6.14 ;
      RECT 27.225 3.395 27.505 3.765 ;
      RECT 26.895 6.46 27.175 6.83 ;
      RECT 22.135 7 22.505 7.37 ;
      RECT 11.725 5.77 12.005 6.14 ;
      RECT 11.375 3.735 11.655 4.105 ;
      RECT 11.035 3.055 11.315 3.425 ;
      RECT 10.685 5.77 10.965 6.14 ;
      RECT 10.005 3.395 10.285 3.765 ;
      RECT 9.675 6.46 9.955 6.83 ;
      RECT 4.915 7 5.285 7.37 ;
    LAYER via1 ;
      RECT 88.415 7.385 88.565 7.535 ;
      RECT 86.06 6.74 86.21 6.89 ;
      RECT 86.045 2.065 86.195 2.215 ;
      RECT 85.255 2.45 85.405 2.6 ;
      RECT 85.255 6.37 85.405 6.52 ;
      RECT 83.59 2.08 83.74 2.23 ;
      RECT 81.68 2.825 81.83 2.975 ;
      RECT 81.68 6.565 81.83 6.715 ;
      RECT 81 3.845 81.15 3.995 ;
      RECT 81 4.865 81.15 5.015 ;
      RECT 80.66 5.885 80.81 6.035 ;
      RECT 80.32 3.845 80.47 3.995 ;
      RECT 79.98 3.165 80.13 3.315 ;
      RECT 79.98 6.565 80.13 6.715 ;
      RECT 79.63 5.885 79.78 6.035 ;
      RECT 79.3 2.825 79.45 2.975 ;
      RECT 78.96 3.505 79.11 3.655 ;
      RECT 78.62 2.315 78.77 2.465 ;
      RECT 78.62 6.565 78.77 6.715 ;
      RECT 77.26 2.485 77.41 2.635 ;
      RECT 76.58 2.825 76.73 2.975 ;
      RECT 76.58 4.865 76.73 5.015 ;
      RECT 74.335 6.64 74.485 6.79 ;
      RECT 73.905 7.11 74.055 7.26 ;
      RECT 71.23 6.74 71.38 6.89 ;
      RECT 68.84 6.74 68.99 6.89 ;
      RECT 68.825 2.065 68.975 2.215 ;
      RECT 68.035 2.45 68.185 2.6 ;
      RECT 68.035 6.37 68.185 6.52 ;
      RECT 66.37 2.08 66.52 2.23 ;
      RECT 64.46 2.825 64.61 2.975 ;
      RECT 64.46 6.565 64.61 6.715 ;
      RECT 63.78 3.845 63.93 3.995 ;
      RECT 63.78 4.865 63.93 5.015 ;
      RECT 63.44 5.885 63.59 6.035 ;
      RECT 63.1 3.845 63.25 3.995 ;
      RECT 62.76 3.165 62.91 3.315 ;
      RECT 62.76 6.565 62.91 6.715 ;
      RECT 62.41 5.885 62.56 6.035 ;
      RECT 62.08 2.825 62.23 2.975 ;
      RECT 61.74 3.505 61.89 3.655 ;
      RECT 61.4 2.315 61.55 2.465 ;
      RECT 61.4 6.565 61.55 6.715 ;
      RECT 60.04 2.485 60.19 2.635 ;
      RECT 59.36 2.825 59.51 2.975 ;
      RECT 59.36 4.865 59.51 5.015 ;
      RECT 57.115 6.64 57.265 6.79 ;
      RECT 56.685 7.11 56.835 7.26 ;
      RECT 54.01 6.74 54.16 6.89 ;
      RECT 51.62 6.74 51.77 6.89 ;
      RECT 51.605 2.065 51.755 2.215 ;
      RECT 50.815 2.45 50.965 2.6 ;
      RECT 50.815 6.37 50.965 6.52 ;
      RECT 49.15 2.08 49.3 2.23 ;
      RECT 47.24 2.825 47.39 2.975 ;
      RECT 47.24 6.565 47.39 6.715 ;
      RECT 46.56 3.845 46.71 3.995 ;
      RECT 46.56 4.865 46.71 5.015 ;
      RECT 46.22 5.885 46.37 6.035 ;
      RECT 45.88 3.845 46.03 3.995 ;
      RECT 45.54 3.165 45.69 3.315 ;
      RECT 45.54 6.565 45.69 6.715 ;
      RECT 45.19 5.885 45.34 6.035 ;
      RECT 44.86 2.825 45.01 2.975 ;
      RECT 44.52 3.505 44.67 3.655 ;
      RECT 44.18 2.315 44.33 2.465 ;
      RECT 44.18 6.565 44.33 6.715 ;
      RECT 42.82 2.485 42.97 2.635 ;
      RECT 42.14 2.825 42.29 2.975 ;
      RECT 42.14 4.865 42.29 5.015 ;
      RECT 39.895 6.64 40.045 6.79 ;
      RECT 39.465 7.11 39.615 7.26 ;
      RECT 36.79 6.74 36.94 6.89 ;
      RECT 34.4 6.74 34.55 6.89 ;
      RECT 34.385 2.065 34.535 2.215 ;
      RECT 33.595 2.45 33.745 2.6 ;
      RECT 33.595 6.37 33.745 6.52 ;
      RECT 31.93 2.08 32.08 2.23 ;
      RECT 30.02 2.825 30.17 2.975 ;
      RECT 30.02 6.565 30.17 6.715 ;
      RECT 29.34 3.845 29.49 3.995 ;
      RECT 29.34 4.865 29.49 5.015 ;
      RECT 29 5.885 29.15 6.035 ;
      RECT 28.66 3.845 28.81 3.995 ;
      RECT 28.32 3.165 28.47 3.315 ;
      RECT 28.32 6.565 28.47 6.715 ;
      RECT 27.97 5.885 28.12 6.035 ;
      RECT 27.64 2.825 27.79 2.975 ;
      RECT 27.3 3.505 27.45 3.655 ;
      RECT 26.96 2.315 27.11 2.465 ;
      RECT 26.96 6.565 27.11 6.715 ;
      RECT 25.6 2.485 25.75 2.635 ;
      RECT 24.92 2.825 25.07 2.975 ;
      RECT 24.92 4.865 25.07 5.015 ;
      RECT 22.675 6.64 22.825 6.79 ;
      RECT 22.245 7.11 22.395 7.26 ;
      RECT 19.57 6.74 19.72 6.89 ;
      RECT 17.18 6.74 17.33 6.89 ;
      RECT 17.165 2.065 17.315 2.215 ;
      RECT 16.375 2.45 16.525 2.6 ;
      RECT 16.375 6.37 16.525 6.52 ;
      RECT 14.71 2.08 14.86 2.23 ;
      RECT 12.8 2.825 12.95 2.975 ;
      RECT 12.8 6.565 12.95 6.715 ;
      RECT 12.12 3.845 12.27 3.995 ;
      RECT 12.12 4.865 12.27 5.015 ;
      RECT 11.78 5.885 11.93 6.035 ;
      RECT 11.44 3.845 11.59 3.995 ;
      RECT 11.1 3.165 11.25 3.315 ;
      RECT 11.1 6.565 11.25 6.715 ;
      RECT 10.75 5.885 10.9 6.035 ;
      RECT 10.42 2.825 10.57 2.975 ;
      RECT 10.08 3.505 10.23 3.655 ;
      RECT 9.74 2.315 9.89 2.465 ;
      RECT 9.74 6.565 9.89 6.715 ;
      RECT 8.38 2.485 8.53 2.635 ;
      RECT 7.7 2.825 7.85 2.975 ;
      RECT 7.7 4.865 7.85 5.015 ;
      RECT 5.455 6.64 5.605 6.79 ;
      RECT 5.025 7.11 5.175 7.26 ;
      RECT 1.605 7.09 1.755 7.24 ;
      RECT 1.23 6.35 1.38 6.5 ;
    LAYER met1 ;
      RECT 88.295 7.77 88.585 8 ;
      RECT 88.355 6.29 88.525 8 ;
      RECT 88.325 7.3 88.65 7.625 ;
      RECT 88.295 6.29 88.585 6.52 ;
      RECT 87.89 2.395 87.995 2.965 ;
      RECT 87.89 2.73 88.215 2.96 ;
      RECT 87.89 2.76 88.385 2.93 ;
      RECT 87.89 2.395 88.08 2.96 ;
      RECT 87.305 2.36 87.595 2.59 ;
      RECT 87.305 2.395 88.08 2.565 ;
      RECT 87.365 0.88 87.535 2.59 ;
      RECT 87.305 0.88 87.595 1.11 ;
      RECT 87.305 7.77 87.595 8 ;
      RECT 87.365 6.29 87.535 8 ;
      RECT 87.305 6.29 87.595 6.52 ;
      RECT 87.305 6.325 88.16 6.485 ;
      RECT 87.99 5.92 88.16 6.485 ;
      RECT 87.305 6.32 87.7 6.485 ;
      RECT 87.925 5.92 88.215 6.15 ;
      RECT 87.925 5.95 88.385 6.12 ;
      RECT 86.935 2.73 87.225 2.96 ;
      RECT 86.935 2.76 87.395 2.93 ;
      RECT 87 1.655 87.165 2.96 ;
      RECT 85.515 1.625 85.805 1.855 ;
      RECT 85.515 1.655 87.165 1.825 ;
      RECT 85.575 0.885 85.745 1.855 ;
      RECT 85.515 0.885 85.805 1.115 ;
      RECT 85.515 7.765 85.805 7.995 ;
      RECT 85.575 7.025 85.745 7.995 ;
      RECT 85.575 7.12 87.165 7.29 ;
      RECT 86.995 5.92 87.165 7.29 ;
      RECT 85.515 7.025 85.805 7.255 ;
      RECT 86.935 5.92 87.225 6.15 ;
      RECT 86.935 5.95 87.395 6.12 ;
      RECT 85.945 1.965 86.295 2.315 ;
      RECT 85.775 2.025 86.295 2.195 ;
      RECT 85.97 6.655 86.295 6.98 ;
      RECT 85.945 6.655 86.295 6.885 ;
      RECT 85.775 6.685 86.295 6.855 ;
      RECT 85.17 2.365 85.49 2.685 ;
      RECT 85.14 2.365 85.49 2.595 ;
      RECT 84.855 2.395 85.49 2.565 ;
      RECT 85.17 6.28 85.49 6.605 ;
      RECT 85.14 6.285 85.49 6.515 ;
      RECT 84.97 6.315 85.49 6.485 ;
      RECT 80.915 3.79 81.235 4.05 ;
      RECT 81.95 3.805 82.24 4.035 ;
      RECT 80.915 3.85 82.24 3.99 ;
      RECT 80.575 5.83 80.895 6.09 ;
      RECT 81.95 5.845 82.24 6.075 ;
      RECT 82.025 5.55 82.165 6.075 ;
      RECT 80.665 5.55 80.805 6.09 ;
      RECT 80.665 5.55 82.165 5.69 ;
      RECT 81.595 2.77 81.915 3.03 ;
      RECT 81.32 2.83 81.915 2.97 ;
      RECT 78.535 6.51 78.855 6.77 ;
      RECT 77.53 6.525 77.82 6.755 ;
      RECT 77.53 6.57 79.445 6.71 ;
      RECT 79.305 6.23 79.445 6.71 ;
      RECT 79.305 6.23 81.315 6.37 ;
      RECT 81.175 5.845 81.315 6.37 ;
      RECT 81.1 5.845 81.39 6.075 ;
      RECT 80.915 4.81 81.235 5.07 ;
      RECT 78.77 4.825 79.06 5.055 ;
      RECT 78.77 4.87 81.235 5.01 ;
      RECT 80.235 3.79 80.555 4.05 ;
      RECT 77.87 3.805 78.16 4.035 ;
      RECT 77.87 3.85 80.555 3.99 ;
      RECT 79.895 6.51 80.215 6.77 ;
      RECT 79.895 6.57 80.49 6.71 ;
      RECT 79.895 3.11 80.215 3.37 ;
      RECT 79.62 3.17 80.215 3.31 ;
      RECT 79.215 2.77 79.535 3.03 ;
      RECT 78.94 2.83 79.535 2.97 ;
      RECT 78.875 3.45 79.195 3.71 ;
      RECT 76 3.465 76.29 3.695 ;
      RECT 76 3.51 79.195 3.65 ;
      RECT 78.455 2.79 78.595 3.65 ;
      RECT 78.38 2.79 78.67 3.02 ;
      RECT 78.535 2.26 78.855 2.52 ;
      RECT 78.535 2.275 79.04 2.505 ;
      RECT 78.445 2.32 79.04 2.46 ;
      RECT 77.87 2.79 78.16 3.02 ;
      RECT 77.265 2.835 78.16 2.975 ;
      RECT 77.265 2.43 77.405 2.975 ;
      RECT 77.175 2.43 77.495 2.69 ;
      RECT 76.495 2.77 76.815 3.03 ;
      RECT 76.22 2.83 76.815 2.97 ;
      RECT 76.495 4.81 76.815 5.07 ;
      RECT 76.22 4.87 76.815 5.01 ;
      RECT 74.26 6.575 74.55 6.885 ;
      RECT 74.09 6.685 74.58 6.855 ;
      RECT 74.24 6.575 74.58 6.855 ;
      RECT 73.83 7.765 74.12 7.995 ;
      RECT 73.89 6.995 74.06 7.995 ;
      RECT 73.795 6.995 74.165 7.37 ;
      RECT 71.075 7.77 71.365 8 ;
      RECT 71.135 6.29 71.305 8 ;
      RECT 71.135 6.655 71.465 6.98 ;
      RECT 71.075 6.29 71.365 6.52 ;
      RECT 70.67 2.395 70.775 2.965 ;
      RECT 70.67 2.73 70.995 2.96 ;
      RECT 70.67 2.76 71.165 2.93 ;
      RECT 70.67 2.395 70.86 2.96 ;
      RECT 70.085 2.36 70.375 2.59 ;
      RECT 70.085 2.395 70.86 2.565 ;
      RECT 70.145 0.88 70.315 2.59 ;
      RECT 70.085 0.88 70.375 1.11 ;
      RECT 70.085 7.77 70.375 8 ;
      RECT 70.145 6.29 70.315 8 ;
      RECT 70.085 6.29 70.375 6.52 ;
      RECT 70.085 6.325 70.94 6.485 ;
      RECT 70.77 5.92 70.94 6.485 ;
      RECT 70.085 6.32 70.48 6.485 ;
      RECT 70.705 5.92 70.995 6.15 ;
      RECT 70.705 5.95 71.165 6.12 ;
      RECT 69.715 2.73 70.005 2.96 ;
      RECT 69.715 2.76 70.175 2.93 ;
      RECT 69.78 1.655 69.945 2.96 ;
      RECT 68.295 1.625 68.585 1.855 ;
      RECT 68.295 1.655 69.945 1.825 ;
      RECT 68.355 0.885 68.525 1.855 ;
      RECT 68.295 0.885 68.585 1.115 ;
      RECT 68.295 7.765 68.585 7.995 ;
      RECT 68.355 7.025 68.525 7.995 ;
      RECT 68.355 7.12 69.945 7.29 ;
      RECT 69.775 5.92 69.945 7.29 ;
      RECT 68.295 7.025 68.585 7.255 ;
      RECT 69.715 5.92 70.005 6.15 ;
      RECT 69.715 5.95 70.175 6.12 ;
      RECT 68.725 1.965 69.075 2.315 ;
      RECT 68.555 2.025 69.075 2.195 ;
      RECT 68.75 6.655 69.075 6.98 ;
      RECT 68.725 6.655 69.075 6.885 ;
      RECT 68.555 6.685 69.075 6.855 ;
      RECT 67.95 2.365 68.27 2.685 ;
      RECT 67.92 2.365 68.27 2.595 ;
      RECT 67.635 2.395 68.27 2.565 ;
      RECT 67.95 6.28 68.27 6.605 ;
      RECT 67.92 6.285 68.27 6.515 ;
      RECT 67.75 6.315 68.27 6.485 ;
      RECT 63.695 3.79 64.015 4.05 ;
      RECT 64.73 3.805 65.02 4.035 ;
      RECT 63.695 3.85 65.02 3.99 ;
      RECT 63.355 5.83 63.675 6.09 ;
      RECT 64.73 5.845 65.02 6.075 ;
      RECT 64.805 5.55 64.945 6.075 ;
      RECT 63.445 5.55 63.585 6.09 ;
      RECT 63.445 5.55 64.945 5.69 ;
      RECT 64.375 2.77 64.695 3.03 ;
      RECT 64.1 2.83 64.695 2.97 ;
      RECT 61.315 6.51 61.635 6.77 ;
      RECT 60.31 6.525 60.6 6.755 ;
      RECT 60.31 6.57 62.225 6.71 ;
      RECT 62.085 6.23 62.225 6.71 ;
      RECT 62.085 6.23 64.095 6.37 ;
      RECT 63.955 5.845 64.095 6.37 ;
      RECT 63.88 5.845 64.17 6.075 ;
      RECT 63.695 4.81 64.015 5.07 ;
      RECT 61.55 4.825 61.84 5.055 ;
      RECT 61.55 4.87 64.015 5.01 ;
      RECT 63.015 3.79 63.335 4.05 ;
      RECT 60.65 3.805 60.94 4.035 ;
      RECT 60.65 3.85 63.335 3.99 ;
      RECT 62.675 6.51 62.995 6.77 ;
      RECT 62.675 6.57 63.27 6.71 ;
      RECT 62.675 3.11 62.995 3.37 ;
      RECT 62.4 3.17 62.995 3.31 ;
      RECT 61.995 2.77 62.315 3.03 ;
      RECT 61.72 2.83 62.315 2.97 ;
      RECT 61.655 3.45 61.975 3.71 ;
      RECT 58.78 3.465 59.07 3.695 ;
      RECT 58.78 3.51 61.975 3.65 ;
      RECT 61.235 2.79 61.375 3.65 ;
      RECT 61.16 2.79 61.45 3.02 ;
      RECT 61.315 2.26 61.635 2.52 ;
      RECT 61.315 2.275 61.82 2.505 ;
      RECT 61.225 2.32 61.82 2.46 ;
      RECT 60.65 2.79 60.94 3.02 ;
      RECT 60.045 2.835 60.94 2.975 ;
      RECT 60.045 2.43 60.185 2.975 ;
      RECT 59.955 2.43 60.275 2.69 ;
      RECT 59.275 2.77 59.595 3.03 ;
      RECT 59 2.83 59.595 2.97 ;
      RECT 59.275 4.81 59.595 5.07 ;
      RECT 59 4.87 59.595 5.01 ;
      RECT 57.04 6.575 57.33 6.885 ;
      RECT 56.87 6.685 57.36 6.855 ;
      RECT 57.02 6.575 57.36 6.855 ;
      RECT 56.61 7.765 56.9 7.995 ;
      RECT 56.67 6.995 56.84 7.995 ;
      RECT 56.575 6.995 56.945 7.37 ;
      RECT 53.855 7.77 54.145 8 ;
      RECT 53.915 6.29 54.085 8 ;
      RECT 53.915 6.655 54.245 6.98 ;
      RECT 53.855 6.29 54.145 6.52 ;
      RECT 53.45 2.395 53.555 2.965 ;
      RECT 53.45 2.73 53.775 2.96 ;
      RECT 53.45 2.76 53.945 2.93 ;
      RECT 53.45 2.395 53.64 2.96 ;
      RECT 52.865 2.36 53.155 2.59 ;
      RECT 52.865 2.395 53.64 2.565 ;
      RECT 52.925 0.88 53.095 2.59 ;
      RECT 52.865 0.88 53.155 1.11 ;
      RECT 52.865 7.77 53.155 8 ;
      RECT 52.925 6.29 53.095 8 ;
      RECT 52.865 6.29 53.155 6.52 ;
      RECT 52.865 6.325 53.72 6.485 ;
      RECT 53.55 5.92 53.72 6.485 ;
      RECT 52.865 6.32 53.26 6.485 ;
      RECT 53.485 5.92 53.775 6.15 ;
      RECT 53.485 5.95 53.945 6.12 ;
      RECT 52.495 2.73 52.785 2.96 ;
      RECT 52.495 2.76 52.955 2.93 ;
      RECT 52.56 1.655 52.725 2.96 ;
      RECT 51.075 1.625 51.365 1.855 ;
      RECT 51.075 1.655 52.725 1.825 ;
      RECT 51.135 0.885 51.305 1.855 ;
      RECT 51.075 0.885 51.365 1.115 ;
      RECT 51.075 7.765 51.365 7.995 ;
      RECT 51.135 7.025 51.305 7.995 ;
      RECT 51.135 7.12 52.725 7.29 ;
      RECT 52.555 5.92 52.725 7.29 ;
      RECT 51.075 7.025 51.365 7.255 ;
      RECT 52.495 5.92 52.785 6.15 ;
      RECT 52.495 5.95 52.955 6.12 ;
      RECT 51.505 1.965 51.855 2.315 ;
      RECT 51.335 2.025 51.855 2.195 ;
      RECT 51.53 6.655 51.855 6.98 ;
      RECT 51.505 6.655 51.855 6.885 ;
      RECT 51.335 6.685 51.855 6.855 ;
      RECT 50.73 2.365 51.05 2.685 ;
      RECT 50.7 2.365 51.05 2.595 ;
      RECT 50.415 2.395 51.05 2.565 ;
      RECT 50.73 6.28 51.05 6.605 ;
      RECT 50.7 6.285 51.05 6.515 ;
      RECT 50.53 6.315 51.05 6.485 ;
      RECT 46.475 3.79 46.795 4.05 ;
      RECT 47.51 3.805 47.8 4.035 ;
      RECT 46.475 3.85 47.8 3.99 ;
      RECT 46.135 5.83 46.455 6.09 ;
      RECT 47.51 5.845 47.8 6.075 ;
      RECT 47.585 5.55 47.725 6.075 ;
      RECT 46.225 5.55 46.365 6.09 ;
      RECT 46.225 5.55 47.725 5.69 ;
      RECT 47.155 2.77 47.475 3.03 ;
      RECT 46.88 2.83 47.475 2.97 ;
      RECT 44.095 6.51 44.415 6.77 ;
      RECT 43.09 6.525 43.38 6.755 ;
      RECT 43.09 6.57 45.005 6.71 ;
      RECT 44.865 6.23 45.005 6.71 ;
      RECT 44.865 6.23 46.875 6.37 ;
      RECT 46.735 5.845 46.875 6.37 ;
      RECT 46.66 5.845 46.95 6.075 ;
      RECT 46.475 4.81 46.795 5.07 ;
      RECT 44.33 4.825 44.62 5.055 ;
      RECT 44.33 4.87 46.795 5.01 ;
      RECT 45.795 3.79 46.115 4.05 ;
      RECT 43.43 3.805 43.72 4.035 ;
      RECT 43.43 3.85 46.115 3.99 ;
      RECT 45.455 6.51 45.775 6.77 ;
      RECT 45.455 6.57 46.05 6.71 ;
      RECT 45.455 3.11 45.775 3.37 ;
      RECT 45.18 3.17 45.775 3.31 ;
      RECT 44.775 2.77 45.095 3.03 ;
      RECT 44.5 2.83 45.095 2.97 ;
      RECT 44.435 3.45 44.755 3.71 ;
      RECT 41.56 3.465 41.85 3.695 ;
      RECT 41.56 3.51 44.755 3.65 ;
      RECT 44.015 2.79 44.155 3.65 ;
      RECT 43.94 2.79 44.23 3.02 ;
      RECT 44.095 2.26 44.415 2.52 ;
      RECT 44.095 2.275 44.6 2.505 ;
      RECT 44.005 2.32 44.6 2.46 ;
      RECT 43.43 2.79 43.72 3.02 ;
      RECT 42.825 2.835 43.72 2.975 ;
      RECT 42.825 2.43 42.965 2.975 ;
      RECT 42.735 2.43 43.055 2.69 ;
      RECT 42.055 2.77 42.375 3.03 ;
      RECT 41.78 2.83 42.375 2.97 ;
      RECT 42.055 4.81 42.375 5.07 ;
      RECT 41.78 4.87 42.375 5.01 ;
      RECT 39.82 6.575 40.11 6.885 ;
      RECT 39.65 6.685 40.14 6.855 ;
      RECT 39.8 6.575 40.14 6.855 ;
      RECT 39.39 7.765 39.68 7.995 ;
      RECT 39.45 6.995 39.62 7.995 ;
      RECT 39.355 6.995 39.725 7.37 ;
      RECT 36.635 7.77 36.925 8 ;
      RECT 36.695 6.29 36.865 8 ;
      RECT 36.695 6.655 37.025 6.98 ;
      RECT 36.635 6.29 36.925 6.52 ;
      RECT 36.23 2.395 36.335 2.965 ;
      RECT 36.23 2.73 36.555 2.96 ;
      RECT 36.23 2.76 36.725 2.93 ;
      RECT 36.23 2.395 36.42 2.96 ;
      RECT 35.645 2.36 35.935 2.59 ;
      RECT 35.645 2.395 36.42 2.565 ;
      RECT 35.705 0.88 35.875 2.59 ;
      RECT 35.645 0.88 35.935 1.11 ;
      RECT 35.645 7.77 35.935 8 ;
      RECT 35.705 6.29 35.875 8 ;
      RECT 35.645 6.29 35.935 6.52 ;
      RECT 35.645 6.325 36.5 6.485 ;
      RECT 36.33 5.92 36.5 6.485 ;
      RECT 35.645 6.32 36.04 6.485 ;
      RECT 36.265 5.92 36.555 6.15 ;
      RECT 36.265 5.95 36.725 6.12 ;
      RECT 35.275 2.73 35.565 2.96 ;
      RECT 35.275 2.76 35.735 2.93 ;
      RECT 35.34 1.655 35.505 2.96 ;
      RECT 33.855 1.625 34.145 1.855 ;
      RECT 33.855 1.655 35.505 1.825 ;
      RECT 33.915 0.885 34.085 1.855 ;
      RECT 33.855 0.885 34.145 1.115 ;
      RECT 33.855 7.765 34.145 7.995 ;
      RECT 33.915 7.025 34.085 7.995 ;
      RECT 33.915 7.12 35.505 7.29 ;
      RECT 35.335 5.92 35.505 7.29 ;
      RECT 33.855 7.025 34.145 7.255 ;
      RECT 35.275 5.92 35.565 6.15 ;
      RECT 35.275 5.95 35.735 6.12 ;
      RECT 34.285 1.965 34.635 2.315 ;
      RECT 34.115 2.025 34.635 2.195 ;
      RECT 34.31 6.655 34.635 6.98 ;
      RECT 34.285 6.655 34.635 6.885 ;
      RECT 34.115 6.685 34.635 6.855 ;
      RECT 33.51 2.365 33.83 2.685 ;
      RECT 33.48 2.365 33.83 2.595 ;
      RECT 33.195 2.395 33.83 2.565 ;
      RECT 33.51 6.28 33.83 6.605 ;
      RECT 33.48 6.285 33.83 6.515 ;
      RECT 33.31 6.315 33.83 6.485 ;
      RECT 29.255 3.79 29.575 4.05 ;
      RECT 30.29 3.805 30.58 4.035 ;
      RECT 29.255 3.85 30.58 3.99 ;
      RECT 28.915 5.83 29.235 6.09 ;
      RECT 30.29 5.845 30.58 6.075 ;
      RECT 30.365 5.55 30.505 6.075 ;
      RECT 29.005 5.55 29.145 6.09 ;
      RECT 29.005 5.55 30.505 5.69 ;
      RECT 29.935 2.77 30.255 3.03 ;
      RECT 29.66 2.83 30.255 2.97 ;
      RECT 26.875 6.51 27.195 6.77 ;
      RECT 25.87 6.525 26.16 6.755 ;
      RECT 25.87 6.57 27.785 6.71 ;
      RECT 27.645 6.23 27.785 6.71 ;
      RECT 27.645 6.23 29.655 6.37 ;
      RECT 29.515 5.845 29.655 6.37 ;
      RECT 29.44 5.845 29.73 6.075 ;
      RECT 29.255 4.81 29.575 5.07 ;
      RECT 27.11 4.825 27.4 5.055 ;
      RECT 27.11 4.87 29.575 5.01 ;
      RECT 28.575 3.79 28.895 4.05 ;
      RECT 26.21 3.805 26.5 4.035 ;
      RECT 26.21 3.85 28.895 3.99 ;
      RECT 28.235 6.51 28.555 6.77 ;
      RECT 28.235 6.57 28.83 6.71 ;
      RECT 28.235 3.11 28.555 3.37 ;
      RECT 27.96 3.17 28.555 3.31 ;
      RECT 27.555 2.77 27.875 3.03 ;
      RECT 27.28 2.83 27.875 2.97 ;
      RECT 27.215 3.45 27.535 3.71 ;
      RECT 24.34 3.465 24.63 3.695 ;
      RECT 24.34 3.51 27.535 3.65 ;
      RECT 26.795 2.79 26.935 3.65 ;
      RECT 26.72 2.79 27.01 3.02 ;
      RECT 26.875 2.26 27.195 2.52 ;
      RECT 26.875 2.275 27.38 2.505 ;
      RECT 26.785 2.32 27.38 2.46 ;
      RECT 26.21 2.79 26.5 3.02 ;
      RECT 25.605 2.835 26.5 2.975 ;
      RECT 25.605 2.43 25.745 2.975 ;
      RECT 25.515 2.43 25.835 2.69 ;
      RECT 24.835 2.77 25.155 3.03 ;
      RECT 24.56 2.83 25.155 2.97 ;
      RECT 24.835 4.81 25.155 5.07 ;
      RECT 24.56 4.87 25.155 5.01 ;
      RECT 22.6 6.575 22.89 6.885 ;
      RECT 22.43 6.685 22.92 6.855 ;
      RECT 22.58 6.575 22.92 6.855 ;
      RECT 22.17 7.765 22.46 7.995 ;
      RECT 22.23 6.995 22.4 7.995 ;
      RECT 22.135 6.995 22.505 7.37 ;
      RECT 19.415 7.77 19.705 8 ;
      RECT 19.475 6.29 19.645 8 ;
      RECT 19.475 6.655 19.805 6.98 ;
      RECT 19.415 6.29 19.705 6.52 ;
      RECT 19.01 2.395 19.115 2.965 ;
      RECT 19.01 2.73 19.335 2.96 ;
      RECT 19.01 2.76 19.505 2.93 ;
      RECT 19.01 2.395 19.2 2.96 ;
      RECT 18.425 2.36 18.715 2.59 ;
      RECT 18.425 2.395 19.2 2.565 ;
      RECT 18.485 0.88 18.655 2.59 ;
      RECT 18.425 0.88 18.715 1.11 ;
      RECT 18.425 7.77 18.715 8 ;
      RECT 18.485 6.29 18.655 8 ;
      RECT 18.425 6.29 18.715 6.52 ;
      RECT 18.425 6.325 19.28 6.485 ;
      RECT 19.11 5.92 19.28 6.485 ;
      RECT 18.425 6.32 18.82 6.485 ;
      RECT 19.045 5.92 19.335 6.15 ;
      RECT 19.045 5.95 19.505 6.12 ;
      RECT 18.055 2.73 18.345 2.96 ;
      RECT 18.055 2.76 18.515 2.93 ;
      RECT 18.12 1.655 18.285 2.96 ;
      RECT 16.635 1.625 16.925 1.855 ;
      RECT 16.635 1.655 18.285 1.825 ;
      RECT 16.695 0.885 16.865 1.855 ;
      RECT 16.635 0.885 16.925 1.115 ;
      RECT 16.635 7.765 16.925 7.995 ;
      RECT 16.695 7.025 16.865 7.995 ;
      RECT 16.695 7.12 18.285 7.29 ;
      RECT 18.115 5.92 18.285 7.29 ;
      RECT 16.635 7.025 16.925 7.255 ;
      RECT 18.055 5.92 18.345 6.15 ;
      RECT 18.055 5.95 18.515 6.12 ;
      RECT 17.065 1.965 17.415 2.315 ;
      RECT 16.895 2.025 17.415 2.195 ;
      RECT 17.09 6.655 17.415 6.98 ;
      RECT 17.065 6.655 17.415 6.885 ;
      RECT 16.895 6.685 17.415 6.855 ;
      RECT 16.29 2.365 16.61 2.685 ;
      RECT 16.26 2.365 16.61 2.595 ;
      RECT 15.975 2.395 16.61 2.565 ;
      RECT 16.29 6.28 16.61 6.605 ;
      RECT 16.26 6.285 16.61 6.515 ;
      RECT 16.09 6.315 16.61 6.485 ;
      RECT 12.035 3.79 12.355 4.05 ;
      RECT 13.07 3.805 13.36 4.035 ;
      RECT 12.035 3.85 13.36 3.99 ;
      RECT 11.695 5.83 12.015 6.09 ;
      RECT 13.07 5.845 13.36 6.075 ;
      RECT 13.145 5.55 13.285 6.075 ;
      RECT 11.785 5.55 11.925 6.09 ;
      RECT 11.785 5.55 13.285 5.69 ;
      RECT 12.715 2.77 13.035 3.03 ;
      RECT 12.44 2.83 13.035 2.97 ;
      RECT 9.655 6.51 9.975 6.77 ;
      RECT 8.65 6.525 8.94 6.755 ;
      RECT 8.65 6.57 10.565 6.71 ;
      RECT 10.425 6.23 10.565 6.71 ;
      RECT 10.425 6.23 12.435 6.37 ;
      RECT 12.295 5.845 12.435 6.37 ;
      RECT 12.22 5.845 12.51 6.075 ;
      RECT 12.035 4.81 12.355 5.07 ;
      RECT 9.89 4.825 10.18 5.055 ;
      RECT 9.89 4.87 12.355 5.01 ;
      RECT 11.355 3.79 11.675 4.05 ;
      RECT 8.99 3.805 9.28 4.035 ;
      RECT 8.99 3.85 11.675 3.99 ;
      RECT 11.015 6.51 11.335 6.77 ;
      RECT 11.015 6.57 11.61 6.71 ;
      RECT 11.015 3.11 11.335 3.37 ;
      RECT 10.74 3.17 11.335 3.31 ;
      RECT 10.335 2.77 10.655 3.03 ;
      RECT 10.06 2.83 10.655 2.97 ;
      RECT 9.995 3.45 10.315 3.71 ;
      RECT 7.12 3.465 7.41 3.695 ;
      RECT 7.12 3.51 10.315 3.65 ;
      RECT 9.575 2.79 9.715 3.65 ;
      RECT 9.5 2.79 9.79 3.02 ;
      RECT 9.655 2.26 9.975 2.52 ;
      RECT 9.655 2.275 10.16 2.505 ;
      RECT 9.565 2.32 10.16 2.46 ;
      RECT 8.99 2.79 9.28 3.02 ;
      RECT 8.385 2.835 9.28 2.975 ;
      RECT 8.385 2.43 8.525 2.975 ;
      RECT 8.295 2.43 8.615 2.69 ;
      RECT 7.615 2.77 7.935 3.03 ;
      RECT 7.34 2.83 7.935 2.97 ;
      RECT 7.615 4.81 7.935 5.07 ;
      RECT 7.34 4.87 7.935 5.01 ;
      RECT 5.38 6.575 5.67 6.885 ;
      RECT 5.21 6.685 5.7 6.855 ;
      RECT 5.36 6.575 5.7 6.855 ;
      RECT 4.95 7.765 5.24 7.995 ;
      RECT 5.01 6.995 5.18 7.995 ;
      RECT 4.915 6.995 5.285 7.37 ;
      RECT 1.54 7.765 1.83 7.995 ;
      RECT 1.6 7.025 1.77 7.995 ;
      RECT 1.51 7.025 1.85 7.305 ;
      RECT 1.135 6.285 1.475 6.565 ;
      RECT 0.995 6.315 1.475 6.485 ;
      RECT 83.5 1.995 83.825 2.32 ;
      RECT 81.27 6.51 81.915 6.77 ;
      RECT 79.22 5.83 79.865 6.09 ;
      RECT 66.28 1.995 66.605 2.32 ;
      RECT 64.05 6.51 64.695 6.77 ;
      RECT 62 5.83 62.645 6.09 ;
      RECT 49.06 1.995 49.385 2.32 ;
      RECT 46.83 6.51 47.475 6.77 ;
      RECT 44.78 5.83 45.425 6.09 ;
      RECT 31.84 1.995 32.165 2.32 ;
      RECT 29.61 6.51 30.255 6.77 ;
      RECT 27.56 5.83 28.205 6.09 ;
      RECT 14.62 1.995 14.945 2.32 ;
      RECT 12.39 6.51 13.035 6.77 ;
      RECT 10.34 5.83 10.985 6.09 ;
    LAYER mcon ;
      RECT 88.355 6.32 88.525 6.49 ;
      RECT 88.36 6.315 88.53 6.485 ;
      RECT 71.135 6.32 71.305 6.49 ;
      RECT 71.14 6.315 71.31 6.485 ;
      RECT 53.915 6.32 54.085 6.49 ;
      RECT 53.92 6.315 54.09 6.485 ;
      RECT 36.695 6.32 36.865 6.49 ;
      RECT 36.7 6.315 36.87 6.485 ;
      RECT 19.475 6.32 19.645 6.49 ;
      RECT 19.48 6.315 19.65 6.485 ;
      RECT 88.355 7.8 88.525 7.97 ;
      RECT 87.985 2.76 88.155 2.93 ;
      RECT 87.985 5.95 88.155 6.12 ;
      RECT 87.365 0.91 87.535 1.08 ;
      RECT 87.365 2.39 87.535 2.56 ;
      RECT 87.365 6.32 87.535 6.49 ;
      RECT 87.365 7.8 87.535 7.97 ;
      RECT 86.995 2.76 87.165 2.93 ;
      RECT 86.995 5.95 87.165 6.12 ;
      RECT 86.005 2.025 86.175 2.195 ;
      RECT 86.005 6.685 86.175 6.855 ;
      RECT 85.575 0.915 85.745 1.085 ;
      RECT 85.575 1.655 85.745 1.825 ;
      RECT 85.575 7.055 85.745 7.225 ;
      RECT 85.575 7.795 85.745 7.965 ;
      RECT 85.2 2.395 85.37 2.565 ;
      RECT 85.2 6.315 85.37 6.485 ;
      RECT 82.01 3.835 82.18 4.005 ;
      RECT 82.01 5.875 82.18 6.045 ;
      RECT 81.67 2.815 81.84 2.985 ;
      RECT 81.33 6.555 81.5 6.725 ;
      RECT 81.16 5.875 81.33 6.045 ;
      RECT 80.65 5.875 80.82 6.045 ;
      RECT 79.97 3.155 80.14 3.325 ;
      RECT 79.97 6.555 80.14 6.725 ;
      RECT 79.29 2.815 79.46 2.985 ;
      RECT 79.28 5.875 79.45 6.045 ;
      RECT 78.83 4.855 79 5.025 ;
      RECT 78.81 2.305 78.98 2.475 ;
      RECT 78.44 2.82 78.61 2.99 ;
      RECT 77.93 2.82 78.1 2.99 ;
      RECT 77.93 3.835 78.1 4.005 ;
      RECT 77.59 6.555 77.76 6.725 ;
      RECT 76.57 2.815 76.74 2.985 ;
      RECT 76.57 4.855 76.74 5.025 ;
      RECT 76.06 3.495 76.23 3.665 ;
      RECT 74.32 6.685 74.49 6.855 ;
      RECT 73.89 7.055 74.06 7.225 ;
      RECT 73.89 7.795 74.06 7.965 ;
      RECT 71.135 7.8 71.305 7.97 ;
      RECT 70.765 2.76 70.935 2.93 ;
      RECT 70.765 5.95 70.935 6.12 ;
      RECT 70.145 0.91 70.315 1.08 ;
      RECT 70.145 2.39 70.315 2.56 ;
      RECT 70.145 6.32 70.315 6.49 ;
      RECT 70.145 7.8 70.315 7.97 ;
      RECT 69.775 2.76 69.945 2.93 ;
      RECT 69.775 5.95 69.945 6.12 ;
      RECT 68.785 2.025 68.955 2.195 ;
      RECT 68.785 6.685 68.955 6.855 ;
      RECT 68.355 0.915 68.525 1.085 ;
      RECT 68.355 1.655 68.525 1.825 ;
      RECT 68.355 7.055 68.525 7.225 ;
      RECT 68.355 7.795 68.525 7.965 ;
      RECT 67.98 2.395 68.15 2.565 ;
      RECT 67.98 6.315 68.15 6.485 ;
      RECT 64.79 3.835 64.96 4.005 ;
      RECT 64.79 5.875 64.96 6.045 ;
      RECT 64.45 2.815 64.62 2.985 ;
      RECT 64.11 6.555 64.28 6.725 ;
      RECT 63.94 5.875 64.11 6.045 ;
      RECT 63.43 5.875 63.6 6.045 ;
      RECT 62.75 3.155 62.92 3.325 ;
      RECT 62.75 6.555 62.92 6.725 ;
      RECT 62.07 2.815 62.24 2.985 ;
      RECT 62.06 5.875 62.23 6.045 ;
      RECT 61.61 4.855 61.78 5.025 ;
      RECT 61.59 2.305 61.76 2.475 ;
      RECT 61.22 2.82 61.39 2.99 ;
      RECT 60.71 2.82 60.88 2.99 ;
      RECT 60.71 3.835 60.88 4.005 ;
      RECT 60.37 6.555 60.54 6.725 ;
      RECT 59.35 2.815 59.52 2.985 ;
      RECT 59.35 4.855 59.52 5.025 ;
      RECT 58.84 3.495 59.01 3.665 ;
      RECT 57.1 6.685 57.27 6.855 ;
      RECT 56.67 7.055 56.84 7.225 ;
      RECT 56.67 7.795 56.84 7.965 ;
      RECT 53.915 7.8 54.085 7.97 ;
      RECT 53.545 2.76 53.715 2.93 ;
      RECT 53.545 5.95 53.715 6.12 ;
      RECT 52.925 0.91 53.095 1.08 ;
      RECT 52.925 2.39 53.095 2.56 ;
      RECT 52.925 6.32 53.095 6.49 ;
      RECT 52.925 7.8 53.095 7.97 ;
      RECT 52.555 2.76 52.725 2.93 ;
      RECT 52.555 5.95 52.725 6.12 ;
      RECT 51.565 2.025 51.735 2.195 ;
      RECT 51.565 6.685 51.735 6.855 ;
      RECT 51.135 0.915 51.305 1.085 ;
      RECT 51.135 1.655 51.305 1.825 ;
      RECT 51.135 7.055 51.305 7.225 ;
      RECT 51.135 7.795 51.305 7.965 ;
      RECT 50.76 2.395 50.93 2.565 ;
      RECT 50.76 6.315 50.93 6.485 ;
      RECT 47.57 3.835 47.74 4.005 ;
      RECT 47.57 5.875 47.74 6.045 ;
      RECT 47.23 2.815 47.4 2.985 ;
      RECT 46.89 6.555 47.06 6.725 ;
      RECT 46.72 5.875 46.89 6.045 ;
      RECT 46.21 5.875 46.38 6.045 ;
      RECT 45.53 3.155 45.7 3.325 ;
      RECT 45.53 6.555 45.7 6.725 ;
      RECT 44.85 2.815 45.02 2.985 ;
      RECT 44.84 5.875 45.01 6.045 ;
      RECT 44.39 4.855 44.56 5.025 ;
      RECT 44.37 2.305 44.54 2.475 ;
      RECT 44 2.82 44.17 2.99 ;
      RECT 43.49 2.82 43.66 2.99 ;
      RECT 43.49 3.835 43.66 4.005 ;
      RECT 43.15 6.555 43.32 6.725 ;
      RECT 42.13 2.815 42.3 2.985 ;
      RECT 42.13 4.855 42.3 5.025 ;
      RECT 41.62 3.495 41.79 3.665 ;
      RECT 39.88 6.685 40.05 6.855 ;
      RECT 39.45 7.055 39.62 7.225 ;
      RECT 39.45 7.795 39.62 7.965 ;
      RECT 36.695 7.8 36.865 7.97 ;
      RECT 36.325 2.76 36.495 2.93 ;
      RECT 36.325 5.95 36.495 6.12 ;
      RECT 35.705 0.91 35.875 1.08 ;
      RECT 35.705 2.39 35.875 2.56 ;
      RECT 35.705 6.32 35.875 6.49 ;
      RECT 35.705 7.8 35.875 7.97 ;
      RECT 35.335 2.76 35.505 2.93 ;
      RECT 35.335 5.95 35.505 6.12 ;
      RECT 34.345 2.025 34.515 2.195 ;
      RECT 34.345 6.685 34.515 6.855 ;
      RECT 33.915 0.915 34.085 1.085 ;
      RECT 33.915 1.655 34.085 1.825 ;
      RECT 33.915 7.055 34.085 7.225 ;
      RECT 33.915 7.795 34.085 7.965 ;
      RECT 33.54 2.395 33.71 2.565 ;
      RECT 33.54 6.315 33.71 6.485 ;
      RECT 30.35 3.835 30.52 4.005 ;
      RECT 30.35 5.875 30.52 6.045 ;
      RECT 30.01 2.815 30.18 2.985 ;
      RECT 29.67 6.555 29.84 6.725 ;
      RECT 29.5 5.875 29.67 6.045 ;
      RECT 28.99 5.875 29.16 6.045 ;
      RECT 28.31 3.155 28.48 3.325 ;
      RECT 28.31 6.555 28.48 6.725 ;
      RECT 27.63 2.815 27.8 2.985 ;
      RECT 27.62 5.875 27.79 6.045 ;
      RECT 27.17 4.855 27.34 5.025 ;
      RECT 27.15 2.305 27.32 2.475 ;
      RECT 26.78 2.82 26.95 2.99 ;
      RECT 26.27 2.82 26.44 2.99 ;
      RECT 26.27 3.835 26.44 4.005 ;
      RECT 25.93 6.555 26.1 6.725 ;
      RECT 24.91 2.815 25.08 2.985 ;
      RECT 24.91 4.855 25.08 5.025 ;
      RECT 24.4 3.495 24.57 3.665 ;
      RECT 22.66 6.685 22.83 6.855 ;
      RECT 22.23 7.055 22.4 7.225 ;
      RECT 22.23 7.795 22.4 7.965 ;
      RECT 19.475 7.8 19.645 7.97 ;
      RECT 19.105 2.76 19.275 2.93 ;
      RECT 19.105 5.95 19.275 6.12 ;
      RECT 18.485 0.91 18.655 1.08 ;
      RECT 18.485 2.39 18.655 2.56 ;
      RECT 18.485 6.32 18.655 6.49 ;
      RECT 18.485 7.8 18.655 7.97 ;
      RECT 18.115 2.76 18.285 2.93 ;
      RECT 18.115 5.95 18.285 6.12 ;
      RECT 17.125 2.025 17.295 2.195 ;
      RECT 17.125 6.685 17.295 6.855 ;
      RECT 16.695 0.915 16.865 1.085 ;
      RECT 16.695 1.655 16.865 1.825 ;
      RECT 16.695 7.055 16.865 7.225 ;
      RECT 16.695 7.795 16.865 7.965 ;
      RECT 16.32 2.395 16.49 2.565 ;
      RECT 16.32 6.315 16.49 6.485 ;
      RECT 13.13 3.835 13.3 4.005 ;
      RECT 13.13 5.875 13.3 6.045 ;
      RECT 12.79 2.815 12.96 2.985 ;
      RECT 12.45 6.555 12.62 6.725 ;
      RECT 12.28 5.875 12.45 6.045 ;
      RECT 11.77 5.875 11.94 6.045 ;
      RECT 11.09 3.155 11.26 3.325 ;
      RECT 11.09 6.555 11.26 6.725 ;
      RECT 10.41 2.815 10.58 2.985 ;
      RECT 10.4 5.875 10.57 6.045 ;
      RECT 9.95 4.855 10.12 5.025 ;
      RECT 9.93 2.305 10.1 2.475 ;
      RECT 9.56 2.82 9.73 2.99 ;
      RECT 9.05 2.82 9.22 2.99 ;
      RECT 9.05 3.835 9.22 4.005 ;
      RECT 8.71 6.555 8.88 6.725 ;
      RECT 7.69 2.815 7.86 2.985 ;
      RECT 7.69 4.855 7.86 5.025 ;
      RECT 7.18 3.495 7.35 3.665 ;
      RECT 5.44 6.685 5.61 6.855 ;
      RECT 5.01 7.055 5.18 7.225 ;
      RECT 5.01 7.795 5.18 7.965 ;
      RECT 1.6 7.055 1.77 7.225 ;
      RECT 1.6 7.795 1.77 7.965 ;
      RECT 1.225 6.315 1.395 6.485 ;
    LAYER li1 ;
      RECT 88.355 5.02 88.525 6.49 ;
      RECT 88.355 6.315 88.53 6.485 ;
      RECT 87.985 1.74 88.155 2.93 ;
      RECT 87.985 1.74 88.455 1.91 ;
      RECT 87.985 6.97 88.455 7.14 ;
      RECT 87.985 5.95 88.155 7.14 ;
      RECT 86.995 1.74 87.165 2.93 ;
      RECT 86.995 1.74 87.465 1.91 ;
      RECT 86.995 6.97 87.465 7.14 ;
      RECT 86.995 5.95 87.165 7.14 ;
      RECT 85.145 2.635 85.315 3.865 ;
      RECT 85.2 0.855 85.37 2.805 ;
      RECT 85.145 0.575 85.315 1.025 ;
      RECT 85.145 7.855 85.315 8.305 ;
      RECT 85.2 6.075 85.37 8.025 ;
      RECT 85.145 5.015 85.315 6.245 ;
      RECT 84.625 0.575 84.795 3.865 ;
      RECT 84.625 2.075 85.03 2.405 ;
      RECT 84.625 1.235 85.03 1.565 ;
      RECT 84.625 5.015 84.795 8.305 ;
      RECT 84.625 7.315 85.03 7.645 ;
      RECT 84.625 6.475 85.03 6.805 ;
      RECT 82.36 3.495 82.74 4.175 ;
      RECT 82.57 2.365 82.74 4.175 ;
      RECT 80.49 2.365 80.72 3.035 ;
      RECT 80.49 2.365 82.74 2.535 ;
      RECT 82.02 2.045 82.19 2.535 ;
      RECT 82.01 3.155 82.18 4.005 ;
      RECT 81.095 3.155 82.4 3.325 ;
      RECT 82.155 2.705 82.4 3.325 ;
      RECT 81.095 2.785 81.265 3.325 ;
      RECT 80.89 2.785 81.265 2.955 ;
      RECT 81.07 6.265 81.765 6.895 ;
      RECT 81.595 4.685 81.765 6.895 ;
      RECT 81.5 4.685 81.83 5.665 ;
      RECT 81.1 3.495 81.43 4.175 ;
      RECT 80.19 3.495 80.59 4.175 ;
      RECT 80.19 3.495 81.43 3.665 ;
      RECT 79.69 3.075 80.01 4.175 ;
      RECT 79.69 3.075 80.14 3.325 ;
      RECT 79.69 3.075 80.32 3.245 ;
      RECT 80.15 2.025 80.32 3.245 ;
      RECT 80.15 2.025 81.105 2.195 ;
      RECT 79.69 6.265 80.385 6.895 ;
      RECT 80.215 4.685 80.385 6.895 ;
      RECT 80.12 4.685 80.45 5.665 ;
      RECT 79.71 5.825 80.045 6.075 ;
      RECT 79.165 5.825 79.5 6.075 ;
      RECT 79.165 5.875 80.045 6.045 ;
      RECT 78.825 6.265 79.52 6.895 ;
      RECT 78.825 4.685 78.995 6.895 ;
      RECT 78.76 4.685 79.09 5.665 ;
      RECT 78.32 3.205 78.65 4.16 ;
      RECT 78.32 3.205 79 3.375 ;
      RECT 78.83 1.965 79 3.375 ;
      RECT 78.74 1.965 79.07 2.605 ;
      RECT 77.8 3.205 78.13 4.16 ;
      RECT 77.45 3.205 78.13 3.375 ;
      RECT 77.45 1.965 77.62 3.375 ;
      RECT 77.38 1.965 77.71 2.605 ;
      RECT 77.59 5.875 77.76 6.725 ;
      RECT 76.865 5.825 77.2 6.075 ;
      RECT 76.865 5.875 77.76 6.045 ;
      RECT 76.93 2.785 77.28 3.035 ;
      RECT 76.41 2.785 76.74 3.035 ;
      RECT 76.41 2.815 77.28 2.985 ;
      RECT 76.525 6.265 77.22 6.895 ;
      RECT 76.525 4.685 76.695 6.895 ;
      RECT 76.46 4.685 76.79 5.665 ;
      RECT 75.99 3.195 76.32 4.175 ;
      RECT 75.99 1.965 76.24 4.175 ;
      RECT 75.99 1.965 76.32 2.595 ;
      RECT 72.94 5.015 73.11 8.305 ;
      RECT 72.94 7.315 73.345 7.645 ;
      RECT 72.94 6.475 73.345 6.805 ;
      RECT 71.135 5.02 71.305 6.49 ;
      RECT 71.135 6.315 71.31 6.485 ;
      RECT 70.765 1.74 70.935 2.93 ;
      RECT 70.765 1.74 71.235 1.91 ;
      RECT 70.765 6.97 71.235 7.14 ;
      RECT 70.765 5.95 70.935 7.14 ;
      RECT 69.775 1.74 69.945 2.93 ;
      RECT 69.775 1.74 70.245 1.91 ;
      RECT 69.775 6.97 70.245 7.14 ;
      RECT 69.775 5.95 69.945 7.14 ;
      RECT 67.925 2.635 68.095 3.865 ;
      RECT 67.98 0.855 68.15 2.805 ;
      RECT 67.925 0.575 68.095 1.025 ;
      RECT 67.925 7.855 68.095 8.305 ;
      RECT 67.98 6.075 68.15 8.025 ;
      RECT 67.925 5.015 68.095 6.245 ;
      RECT 67.405 0.575 67.575 3.865 ;
      RECT 67.405 2.075 67.81 2.405 ;
      RECT 67.405 1.235 67.81 1.565 ;
      RECT 67.405 5.015 67.575 8.305 ;
      RECT 67.405 7.315 67.81 7.645 ;
      RECT 67.405 6.475 67.81 6.805 ;
      RECT 65.14 3.495 65.52 4.175 ;
      RECT 65.35 2.365 65.52 4.175 ;
      RECT 63.27 2.365 63.5 3.035 ;
      RECT 63.27 2.365 65.52 2.535 ;
      RECT 64.8 2.045 64.97 2.535 ;
      RECT 64.79 3.155 64.96 4.005 ;
      RECT 63.875 3.155 65.18 3.325 ;
      RECT 64.935 2.705 65.18 3.325 ;
      RECT 63.875 2.785 64.045 3.325 ;
      RECT 63.67 2.785 64.045 2.955 ;
      RECT 63.85 6.265 64.545 6.895 ;
      RECT 64.375 4.685 64.545 6.895 ;
      RECT 64.28 4.685 64.61 5.665 ;
      RECT 63.88 3.495 64.21 4.175 ;
      RECT 62.97 3.495 63.37 4.175 ;
      RECT 62.97 3.495 64.21 3.665 ;
      RECT 62.47 3.075 62.79 4.175 ;
      RECT 62.47 3.075 62.92 3.325 ;
      RECT 62.47 3.075 63.1 3.245 ;
      RECT 62.93 2.025 63.1 3.245 ;
      RECT 62.93 2.025 63.885 2.195 ;
      RECT 62.47 6.265 63.165 6.895 ;
      RECT 62.995 4.685 63.165 6.895 ;
      RECT 62.9 4.685 63.23 5.665 ;
      RECT 62.49 5.825 62.825 6.075 ;
      RECT 61.945 5.825 62.28 6.075 ;
      RECT 61.945 5.875 62.825 6.045 ;
      RECT 61.605 6.265 62.3 6.895 ;
      RECT 61.605 4.685 61.775 6.895 ;
      RECT 61.54 4.685 61.87 5.665 ;
      RECT 61.1 3.205 61.43 4.16 ;
      RECT 61.1 3.205 61.78 3.375 ;
      RECT 61.61 1.965 61.78 3.375 ;
      RECT 61.52 1.965 61.85 2.605 ;
      RECT 60.58 3.205 60.91 4.16 ;
      RECT 60.23 3.205 60.91 3.375 ;
      RECT 60.23 1.965 60.4 3.375 ;
      RECT 60.16 1.965 60.49 2.605 ;
      RECT 60.37 5.875 60.54 6.725 ;
      RECT 59.645 5.825 59.98 6.075 ;
      RECT 59.645 5.875 60.54 6.045 ;
      RECT 59.71 2.785 60.06 3.035 ;
      RECT 59.19 2.785 59.52 3.035 ;
      RECT 59.19 2.815 60.06 2.985 ;
      RECT 59.305 6.265 60 6.895 ;
      RECT 59.305 4.685 59.475 6.895 ;
      RECT 59.24 4.685 59.57 5.665 ;
      RECT 58.77 3.195 59.1 4.175 ;
      RECT 58.77 1.965 59.02 4.175 ;
      RECT 58.77 1.965 59.1 2.595 ;
      RECT 55.72 5.015 55.89 8.305 ;
      RECT 55.72 7.315 56.125 7.645 ;
      RECT 55.72 6.475 56.125 6.805 ;
      RECT 53.915 5.02 54.085 6.49 ;
      RECT 53.915 6.315 54.09 6.485 ;
      RECT 53.545 1.74 53.715 2.93 ;
      RECT 53.545 1.74 54.015 1.91 ;
      RECT 53.545 6.97 54.015 7.14 ;
      RECT 53.545 5.95 53.715 7.14 ;
      RECT 52.555 1.74 52.725 2.93 ;
      RECT 52.555 1.74 53.025 1.91 ;
      RECT 52.555 6.97 53.025 7.14 ;
      RECT 52.555 5.95 52.725 7.14 ;
      RECT 50.705 2.635 50.875 3.865 ;
      RECT 50.76 0.855 50.93 2.805 ;
      RECT 50.705 0.575 50.875 1.025 ;
      RECT 50.705 7.855 50.875 8.305 ;
      RECT 50.76 6.075 50.93 8.025 ;
      RECT 50.705 5.015 50.875 6.245 ;
      RECT 50.185 0.575 50.355 3.865 ;
      RECT 50.185 2.075 50.59 2.405 ;
      RECT 50.185 1.235 50.59 1.565 ;
      RECT 50.185 5.015 50.355 8.305 ;
      RECT 50.185 7.315 50.59 7.645 ;
      RECT 50.185 6.475 50.59 6.805 ;
      RECT 47.92 3.495 48.3 4.175 ;
      RECT 48.13 2.365 48.3 4.175 ;
      RECT 46.05 2.365 46.28 3.035 ;
      RECT 46.05 2.365 48.3 2.535 ;
      RECT 47.58 2.045 47.75 2.535 ;
      RECT 47.57 3.155 47.74 4.005 ;
      RECT 46.655 3.155 47.96 3.325 ;
      RECT 47.715 2.705 47.96 3.325 ;
      RECT 46.655 2.785 46.825 3.325 ;
      RECT 46.45 2.785 46.825 2.955 ;
      RECT 46.63 6.265 47.325 6.895 ;
      RECT 47.155 4.685 47.325 6.895 ;
      RECT 47.06 4.685 47.39 5.665 ;
      RECT 46.66 3.495 46.99 4.175 ;
      RECT 45.75 3.495 46.15 4.175 ;
      RECT 45.75 3.495 46.99 3.665 ;
      RECT 45.25 3.075 45.57 4.175 ;
      RECT 45.25 3.075 45.7 3.325 ;
      RECT 45.25 3.075 45.88 3.245 ;
      RECT 45.71 2.025 45.88 3.245 ;
      RECT 45.71 2.025 46.665 2.195 ;
      RECT 45.25 6.265 45.945 6.895 ;
      RECT 45.775 4.685 45.945 6.895 ;
      RECT 45.68 4.685 46.01 5.665 ;
      RECT 45.27 5.825 45.605 6.075 ;
      RECT 44.725 5.825 45.06 6.075 ;
      RECT 44.725 5.875 45.605 6.045 ;
      RECT 44.385 6.265 45.08 6.895 ;
      RECT 44.385 4.685 44.555 6.895 ;
      RECT 44.32 4.685 44.65 5.665 ;
      RECT 43.88 3.205 44.21 4.16 ;
      RECT 43.88 3.205 44.56 3.375 ;
      RECT 44.39 1.965 44.56 3.375 ;
      RECT 44.3 1.965 44.63 2.605 ;
      RECT 43.36 3.205 43.69 4.16 ;
      RECT 43.01 3.205 43.69 3.375 ;
      RECT 43.01 1.965 43.18 3.375 ;
      RECT 42.94 1.965 43.27 2.605 ;
      RECT 43.15 5.875 43.32 6.725 ;
      RECT 42.425 5.825 42.76 6.075 ;
      RECT 42.425 5.875 43.32 6.045 ;
      RECT 42.49 2.785 42.84 3.035 ;
      RECT 41.97 2.785 42.3 3.035 ;
      RECT 41.97 2.815 42.84 2.985 ;
      RECT 42.085 6.265 42.78 6.895 ;
      RECT 42.085 4.685 42.255 6.895 ;
      RECT 42.02 4.685 42.35 5.665 ;
      RECT 41.55 3.195 41.88 4.175 ;
      RECT 41.55 1.965 41.8 4.175 ;
      RECT 41.55 1.965 41.88 2.595 ;
      RECT 38.5 5.015 38.67 8.305 ;
      RECT 38.5 7.315 38.905 7.645 ;
      RECT 38.5 6.475 38.905 6.805 ;
      RECT 36.695 5.02 36.865 6.49 ;
      RECT 36.695 6.315 36.87 6.485 ;
      RECT 36.325 1.74 36.495 2.93 ;
      RECT 36.325 1.74 36.795 1.91 ;
      RECT 36.325 6.97 36.795 7.14 ;
      RECT 36.325 5.95 36.495 7.14 ;
      RECT 35.335 1.74 35.505 2.93 ;
      RECT 35.335 1.74 35.805 1.91 ;
      RECT 35.335 6.97 35.805 7.14 ;
      RECT 35.335 5.95 35.505 7.14 ;
      RECT 33.485 2.635 33.655 3.865 ;
      RECT 33.54 0.855 33.71 2.805 ;
      RECT 33.485 0.575 33.655 1.025 ;
      RECT 33.485 7.855 33.655 8.305 ;
      RECT 33.54 6.075 33.71 8.025 ;
      RECT 33.485 5.015 33.655 6.245 ;
      RECT 32.965 0.575 33.135 3.865 ;
      RECT 32.965 2.075 33.37 2.405 ;
      RECT 32.965 1.235 33.37 1.565 ;
      RECT 32.965 5.015 33.135 8.305 ;
      RECT 32.965 7.315 33.37 7.645 ;
      RECT 32.965 6.475 33.37 6.805 ;
      RECT 30.7 3.495 31.08 4.175 ;
      RECT 30.91 2.365 31.08 4.175 ;
      RECT 28.83 2.365 29.06 3.035 ;
      RECT 28.83 2.365 31.08 2.535 ;
      RECT 30.36 2.045 30.53 2.535 ;
      RECT 30.35 3.155 30.52 4.005 ;
      RECT 29.435 3.155 30.74 3.325 ;
      RECT 30.495 2.705 30.74 3.325 ;
      RECT 29.435 2.785 29.605 3.325 ;
      RECT 29.23 2.785 29.605 2.955 ;
      RECT 29.41 6.265 30.105 6.895 ;
      RECT 29.935 4.685 30.105 6.895 ;
      RECT 29.84 4.685 30.17 5.665 ;
      RECT 29.44 3.495 29.77 4.175 ;
      RECT 28.53 3.495 28.93 4.175 ;
      RECT 28.53 3.495 29.77 3.665 ;
      RECT 28.03 3.075 28.35 4.175 ;
      RECT 28.03 3.075 28.48 3.325 ;
      RECT 28.03 3.075 28.66 3.245 ;
      RECT 28.49 2.025 28.66 3.245 ;
      RECT 28.49 2.025 29.445 2.195 ;
      RECT 28.03 6.265 28.725 6.895 ;
      RECT 28.555 4.685 28.725 6.895 ;
      RECT 28.46 4.685 28.79 5.665 ;
      RECT 28.05 5.825 28.385 6.075 ;
      RECT 27.505 5.825 27.84 6.075 ;
      RECT 27.505 5.875 28.385 6.045 ;
      RECT 27.165 6.265 27.86 6.895 ;
      RECT 27.165 4.685 27.335 6.895 ;
      RECT 27.1 4.685 27.43 5.665 ;
      RECT 26.66 3.205 26.99 4.16 ;
      RECT 26.66 3.205 27.34 3.375 ;
      RECT 27.17 1.965 27.34 3.375 ;
      RECT 27.08 1.965 27.41 2.605 ;
      RECT 26.14 3.205 26.47 4.16 ;
      RECT 25.79 3.205 26.47 3.375 ;
      RECT 25.79 1.965 25.96 3.375 ;
      RECT 25.72 1.965 26.05 2.605 ;
      RECT 25.93 5.875 26.1 6.725 ;
      RECT 25.205 5.825 25.54 6.075 ;
      RECT 25.205 5.875 26.1 6.045 ;
      RECT 25.27 2.785 25.62 3.035 ;
      RECT 24.75 2.785 25.08 3.035 ;
      RECT 24.75 2.815 25.62 2.985 ;
      RECT 24.865 6.265 25.56 6.895 ;
      RECT 24.865 4.685 25.035 6.895 ;
      RECT 24.8 4.685 25.13 5.665 ;
      RECT 24.33 3.195 24.66 4.175 ;
      RECT 24.33 1.965 24.58 4.175 ;
      RECT 24.33 1.965 24.66 2.595 ;
      RECT 21.28 5.015 21.45 8.305 ;
      RECT 21.28 7.315 21.685 7.645 ;
      RECT 21.28 6.475 21.685 6.805 ;
      RECT 19.475 5.02 19.645 6.49 ;
      RECT 19.475 6.315 19.65 6.485 ;
      RECT 19.105 1.74 19.275 2.93 ;
      RECT 19.105 1.74 19.575 1.91 ;
      RECT 19.105 6.97 19.575 7.14 ;
      RECT 19.105 5.95 19.275 7.14 ;
      RECT 18.115 1.74 18.285 2.93 ;
      RECT 18.115 1.74 18.585 1.91 ;
      RECT 18.115 6.97 18.585 7.14 ;
      RECT 18.115 5.95 18.285 7.14 ;
      RECT 16.265 2.635 16.435 3.865 ;
      RECT 16.32 0.855 16.49 2.805 ;
      RECT 16.265 0.575 16.435 1.025 ;
      RECT 16.265 7.855 16.435 8.305 ;
      RECT 16.32 6.075 16.49 8.025 ;
      RECT 16.265 5.015 16.435 6.245 ;
      RECT 15.745 0.575 15.915 3.865 ;
      RECT 15.745 2.075 16.15 2.405 ;
      RECT 15.745 1.235 16.15 1.565 ;
      RECT 15.745 5.015 15.915 8.305 ;
      RECT 15.745 7.315 16.15 7.645 ;
      RECT 15.745 6.475 16.15 6.805 ;
      RECT 13.48 3.495 13.86 4.175 ;
      RECT 13.69 2.365 13.86 4.175 ;
      RECT 11.61 2.365 11.84 3.035 ;
      RECT 11.61 2.365 13.86 2.535 ;
      RECT 13.14 2.045 13.31 2.535 ;
      RECT 13.13 3.155 13.3 4.005 ;
      RECT 12.215 3.155 13.52 3.325 ;
      RECT 13.275 2.705 13.52 3.325 ;
      RECT 12.215 2.785 12.385 3.325 ;
      RECT 12.01 2.785 12.385 2.955 ;
      RECT 12.19 6.265 12.885 6.895 ;
      RECT 12.715 4.685 12.885 6.895 ;
      RECT 12.62 4.685 12.95 5.665 ;
      RECT 12.22 3.495 12.55 4.175 ;
      RECT 11.31 3.495 11.71 4.175 ;
      RECT 11.31 3.495 12.55 3.665 ;
      RECT 10.81 3.075 11.13 4.175 ;
      RECT 10.81 3.075 11.26 3.325 ;
      RECT 10.81 3.075 11.44 3.245 ;
      RECT 11.27 2.025 11.44 3.245 ;
      RECT 11.27 2.025 12.225 2.195 ;
      RECT 10.81 6.265 11.505 6.895 ;
      RECT 11.335 4.685 11.505 6.895 ;
      RECT 11.24 4.685 11.57 5.665 ;
      RECT 10.83 5.825 11.165 6.075 ;
      RECT 10.285 5.825 10.62 6.075 ;
      RECT 10.285 5.875 11.165 6.045 ;
      RECT 9.945 6.265 10.64 6.895 ;
      RECT 9.945 4.685 10.115 6.895 ;
      RECT 9.88 4.685 10.21 5.665 ;
      RECT 9.44 3.205 9.77 4.16 ;
      RECT 9.44 3.205 10.12 3.375 ;
      RECT 9.95 1.965 10.12 3.375 ;
      RECT 9.86 1.965 10.19 2.605 ;
      RECT 8.92 3.205 9.25 4.16 ;
      RECT 8.57 3.205 9.25 3.375 ;
      RECT 8.57 1.965 8.74 3.375 ;
      RECT 8.5 1.965 8.83 2.605 ;
      RECT 8.71 5.875 8.88 6.725 ;
      RECT 7.985 5.825 8.32 6.075 ;
      RECT 7.985 5.875 8.88 6.045 ;
      RECT 8.05 2.785 8.4 3.035 ;
      RECT 7.53 2.785 7.86 3.035 ;
      RECT 7.53 2.815 8.4 2.985 ;
      RECT 7.645 6.265 8.34 6.895 ;
      RECT 7.645 4.685 7.815 6.895 ;
      RECT 7.58 4.685 7.91 5.665 ;
      RECT 7.11 3.195 7.44 4.175 ;
      RECT 7.11 1.965 7.36 4.175 ;
      RECT 7.11 1.965 7.44 2.595 ;
      RECT 4.06 5.015 4.23 8.305 ;
      RECT 4.06 7.315 4.465 7.645 ;
      RECT 4.06 6.475 4.465 6.805 ;
      RECT 1.17 7.855 1.34 8.305 ;
      RECT 1.225 6.075 1.395 8.025 ;
      RECT 1.17 5.015 1.34 6.245 ;
      RECT 0.65 5.015 0.82 8.305 ;
      RECT 0.65 7.315 1.055 7.645 ;
      RECT 0.65 6.475 1.055 6.805 ;
      RECT 88.355 7.8 88.525 8.31 ;
      RECT 87.365 0.57 87.535 1.08 ;
      RECT 87.365 2.39 87.535 3.86 ;
      RECT 87.365 5.02 87.535 6.49 ;
      RECT 87.365 7.8 87.535 8.31 ;
      RECT 86.005 0.575 86.175 3.865 ;
      RECT 86.005 5.015 86.175 8.305 ;
      RECT 85.575 0.575 85.745 1.085 ;
      RECT 85.575 1.655 85.745 3.865 ;
      RECT 85.575 5.015 85.745 7.225 ;
      RECT 85.575 7.795 85.745 8.305 ;
      RECT 81.935 5.825 82.27 6.095 ;
      RECT 81.435 2.785 81.985 2.985 ;
      RECT 81.09 5.825 81.425 6.075 ;
      RECT 80.555 5.825 80.89 6.095 ;
      RECT 79.17 2.785 79.52 3.035 ;
      RECT 78.31 2.785 78.66 3.035 ;
      RECT 77.79 2.785 78.14 3.035 ;
      RECT 74.32 5.015 74.49 8.305 ;
      RECT 73.89 5.015 74.06 7.225 ;
      RECT 73.89 7.795 74.06 8.305 ;
      RECT 71.135 7.8 71.305 8.31 ;
      RECT 70.145 0.57 70.315 1.08 ;
      RECT 70.145 2.39 70.315 3.86 ;
      RECT 70.145 5.02 70.315 6.49 ;
      RECT 70.145 7.8 70.315 8.31 ;
      RECT 68.785 0.575 68.955 3.865 ;
      RECT 68.785 5.015 68.955 8.305 ;
      RECT 68.355 0.575 68.525 1.085 ;
      RECT 68.355 1.655 68.525 3.865 ;
      RECT 68.355 5.015 68.525 7.225 ;
      RECT 68.355 7.795 68.525 8.305 ;
      RECT 64.715 5.825 65.05 6.095 ;
      RECT 64.215 2.785 64.765 2.985 ;
      RECT 63.87 5.825 64.205 6.075 ;
      RECT 63.335 5.825 63.67 6.095 ;
      RECT 61.95 2.785 62.3 3.035 ;
      RECT 61.09 2.785 61.44 3.035 ;
      RECT 60.57 2.785 60.92 3.035 ;
      RECT 57.1 5.015 57.27 8.305 ;
      RECT 56.67 5.015 56.84 7.225 ;
      RECT 56.67 7.795 56.84 8.305 ;
      RECT 53.915 7.8 54.085 8.31 ;
      RECT 52.925 0.57 53.095 1.08 ;
      RECT 52.925 2.39 53.095 3.86 ;
      RECT 52.925 5.02 53.095 6.49 ;
      RECT 52.925 7.8 53.095 8.31 ;
      RECT 51.565 0.575 51.735 3.865 ;
      RECT 51.565 5.015 51.735 8.305 ;
      RECT 51.135 0.575 51.305 1.085 ;
      RECT 51.135 1.655 51.305 3.865 ;
      RECT 51.135 5.015 51.305 7.225 ;
      RECT 51.135 7.795 51.305 8.305 ;
      RECT 47.495 5.825 47.83 6.095 ;
      RECT 46.995 2.785 47.545 2.985 ;
      RECT 46.65 5.825 46.985 6.075 ;
      RECT 46.115 5.825 46.45 6.095 ;
      RECT 44.73 2.785 45.08 3.035 ;
      RECT 43.87 2.785 44.22 3.035 ;
      RECT 43.35 2.785 43.7 3.035 ;
      RECT 39.88 5.015 40.05 8.305 ;
      RECT 39.45 5.015 39.62 7.225 ;
      RECT 39.45 7.795 39.62 8.305 ;
      RECT 36.695 7.8 36.865 8.31 ;
      RECT 35.705 0.57 35.875 1.08 ;
      RECT 35.705 2.39 35.875 3.86 ;
      RECT 35.705 5.02 35.875 6.49 ;
      RECT 35.705 7.8 35.875 8.31 ;
      RECT 34.345 0.575 34.515 3.865 ;
      RECT 34.345 5.015 34.515 8.305 ;
      RECT 33.915 0.575 34.085 1.085 ;
      RECT 33.915 1.655 34.085 3.865 ;
      RECT 33.915 5.015 34.085 7.225 ;
      RECT 33.915 7.795 34.085 8.305 ;
      RECT 30.275 5.825 30.61 6.095 ;
      RECT 29.775 2.785 30.325 2.985 ;
      RECT 29.43 5.825 29.765 6.075 ;
      RECT 28.895 5.825 29.23 6.095 ;
      RECT 27.51 2.785 27.86 3.035 ;
      RECT 26.65 2.785 27 3.035 ;
      RECT 26.13 2.785 26.48 3.035 ;
      RECT 22.66 5.015 22.83 8.305 ;
      RECT 22.23 5.015 22.4 7.225 ;
      RECT 22.23 7.795 22.4 8.305 ;
      RECT 19.475 7.8 19.645 8.31 ;
      RECT 18.485 0.57 18.655 1.08 ;
      RECT 18.485 2.39 18.655 3.86 ;
      RECT 18.485 5.02 18.655 6.49 ;
      RECT 18.485 7.8 18.655 8.31 ;
      RECT 17.125 0.575 17.295 3.865 ;
      RECT 17.125 5.015 17.295 8.305 ;
      RECT 16.695 0.575 16.865 1.085 ;
      RECT 16.695 1.655 16.865 3.865 ;
      RECT 16.695 5.015 16.865 7.225 ;
      RECT 16.695 7.795 16.865 8.305 ;
      RECT 13.055 5.825 13.39 6.095 ;
      RECT 12.555 2.785 13.105 2.985 ;
      RECT 12.21 5.825 12.545 6.075 ;
      RECT 11.675 5.825 12.01 6.095 ;
      RECT 10.29 2.785 10.64 3.035 ;
      RECT 9.43 2.785 9.78 3.035 ;
      RECT 8.91 2.785 9.26 3.035 ;
      RECT 5.44 5.015 5.61 8.305 ;
      RECT 5.01 5.015 5.18 7.225 ;
      RECT 5.01 7.795 5.18 8.305 ;
      RECT 1.6 5.015 1.77 7.225 ;
      RECT 1.6 7.795 1.77 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r1 ;
  SIZE 84.425 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 18.585 0.915 18.755 1.085 ;
        RECT 18.58 0.91 18.75 1.08 ;
        RECT 18.58 2.39 18.75 2.56 ;
      LAYER li1 ;
        RECT 18.585 0.915 18.755 1.085 ;
        RECT 18.58 0.57 18.75 1.08 ;
        RECT 18.58 2.39 18.75 3.86 ;
      LAYER met1 ;
        RECT 18.52 2.36 18.81 2.59 ;
        RECT 18.52 0.88 18.81 1.11 ;
        RECT 18.58 0.88 18.75 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 34.91 0.915 35.08 1.085 ;
        RECT 34.905 0.91 35.075 1.08 ;
        RECT 34.905 2.39 35.075 2.56 ;
      LAYER li1 ;
        RECT 34.91 0.915 35.08 1.085 ;
        RECT 34.905 0.57 35.075 1.08 ;
        RECT 34.905 2.39 35.075 3.86 ;
      LAYER met1 ;
        RECT 34.845 2.36 35.135 2.59 ;
        RECT 34.845 0.88 35.135 1.11 ;
        RECT 34.905 0.88 35.075 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 51.235 0.915 51.405 1.085 ;
        RECT 51.23 0.91 51.4 1.08 ;
        RECT 51.23 2.39 51.4 2.56 ;
      LAYER li1 ;
        RECT 51.235 0.915 51.405 1.085 ;
        RECT 51.23 0.57 51.4 1.08 ;
        RECT 51.23 2.39 51.4 3.86 ;
      LAYER met1 ;
        RECT 51.17 2.36 51.46 2.59 ;
        RECT 51.17 0.88 51.46 1.11 ;
        RECT 51.23 0.88 51.4 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 67.56 0.915 67.73 1.085 ;
        RECT 67.555 0.91 67.725 1.08 ;
        RECT 67.555 2.39 67.725 2.56 ;
      LAYER li1 ;
        RECT 67.56 0.915 67.73 1.085 ;
        RECT 67.555 0.57 67.725 1.08 ;
        RECT 67.555 2.39 67.725 3.86 ;
      LAYER met1 ;
        RECT 67.495 2.36 67.785 2.59 ;
        RECT 67.495 0.88 67.785 1.11 ;
        RECT 67.555 0.88 67.725 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 83.885 0.915 84.055 1.085 ;
        RECT 83.88 0.91 84.05 1.08 ;
        RECT 83.88 2.39 84.05 2.56 ;
      LAYER li1 ;
        RECT 83.885 0.915 84.055 1.085 ;
        RECT 83.88 0.57 84.05 1.08 ;
        RECT 83.88 2.39 84.05 3.86 ;
      LAYER met1 ;
        RECT 83.82 2.36 84.11 2.59 ;
        RECT 83.82 0.88 84.11 1.11 ;
        RECT 83.88 0.88 84.05 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 14.43 1.66 14.6 2.935 ;
        RECT 14.43 5.945 14.6 7.22 ;
        RECT 8.815 5.945 8.985 7.22 ;
      LAYER met2 ;
        RECT 14.355 2.705 14.695 3.055 ;
        RECT 14.345 5.84 14.685 6.19 ;
        RECT 14.43 2.705 14.6 6.19 ;
      LAYER met1 ;
        RECT 14.355 2.765 14.83 2.935 ;
        RECT 14.355 2.705 14.695 3.055 ;
        RECT 8.755 5.945 14.83 6.115 ;
        RECT 14.345 5.84 14.685 6.19 ;
        RECT 8.755 5.915 9.045 6.145 ;
      LAYER mcon ;
        RECT 8.815 5.945 8.985 6.115 ;
        RECT 14.43 5.945 14.6 6.115 ;
        RECT 14.43 2.765 14.6 2.935 ;
      LAYER via1 ;
        RECT 14.445 5.94 14.595 6.09 ;
        RECT 14.455 2.805 14.605 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 30.755 1.66 30.925 2.935 ;
        RECT 30.755 5.945 30.925 7.22 ;
        RECT 25.14 5.945 25.31 7.22 ;
      LAYER met2 ;
        RECT 30.68 2.705 31.02 3.055 ;
        RECT 30.67 5.84 31.01 6.19 ;
        RECT 30.755 2.705 30.925 6.19 ;
      LAYER met1 ;
        RECT 30.68 2.765 31.155 2.935 ;
        RECT 30.68 2.705 31.02 3.055 ;
        RECT 25.08 5.945 31.155 6.115 ;
        RECT 30.67 5.84 31.01 6.19 ;
        RECT 25.08 5.915 25.37 6.145 ;
      LAYER mcon ;
        RECT 25.14 5.945 25.31 6.115 ;
        RECT 30.755 5.945 30.925 6.115 ;
        RECT 30.755 2.765 30.925 2.935 ;
      LAYER via1 ;
        RECT 30.77 5.94 30.92 6.09 ;
        RECT 30.78 2.805 30.93 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 47.08 1.66 47.25 2.935 ;
        RECT 47.08 5.945 47.25 7.22 ;
        RECT 41.465 5.945 41.635 7.22 ;
      LAYER met2 ;
        RECT 47.005 2.705 47.345 3.055 ;
        RECT 46.995 5.84 47.335 6.19 ;
        RECT 47.08 2.705 47.25 6.19 ;
      LAYER met1 ;
        RECT 47.005 2.765 47.48 2.935 ;
        RECT 47.005 2.705 47.345 3.055 ;
        RECT 41.405 5.945 47.48 6.115 ;
        RECT 46.995 5.84 47.335 6.19 ;
        RECT 41.405 5.915 41.695 6.145 ;
      LAYER mcon ;
        RECT 41.465 5.945 41.635 6.115 ;
        RECT 47.08 5.945 47.25 6.115 ;
        RECT 47.08 2.765 47.25 2.935 ;
      LAYER via1 ;
        RECT 47.095 5.94 47.245 6.09 ;
        RECT 47.105 2.805 47.255 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 63.405 1.66 63.575 2.935 ;
        RECT 63.405 5.945 63.575 7.22 ;
        RECT 57.79 5.945 57.96 7.22 ;
      LAYER met2 ;
        RECT 63.33 2.705 63.67 3.055 ;
        RECT 63.32 5.84 63.66 6.19 ;
        RECT 63.405 2.705 63.575 6.19 ;
      LAYER met1 ;
        RECT 63.33 2.765 63.805 2.935 ;
        RECT 63.33 2.705 63.67 3.055 ;
        RECT 57.73 5.945 63.805 6.115 ;
        RECT 63.32 5.84 63.66 6.19 ;
        RECT 57.73 5.915 58.02 6.145 ;
      LAYER mcon ;
        RECT 57.79 5.945 57.96 6.115 ;
        RECT 63.405 5.945 63.575 6.115 ;
        RECT 63.405 2.765 63.575 2.935 ;
      LAYER via1 ;
        RECT 63.42 5.94 63.57 6.09 ;
        RECT 63.43 2.805 63.58 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 79.73 1.66 79.9 2.935 ;
        RECT 79.73 5.945 79.9 7.22 ;
        RECT 74.115 5.945 74.285 7.22 ;
      LAYER met2 ;
        RECT 79.655 2.705 79.995 3.055 ;
        RECT 79.645 5.84 79.985 6.19 ;
        RECT 79.73 2.705 79.9 6.19 ;
      LAYER met1 ;
        RECT 79.655 2.765 80.13 2.935 ;
        RECT 79.655 2.705 79.995 3.055 ;
        RECT 74.055 5.945 80.13 6.115 ;
        RECT 79.645 5.84 79.985 6.19 ;
        RECT 74.055 5.915 74.345 6.145 ;
      LAYER mcon ;
        RECT 74.115 5.945 74.285 6.115 ;
        RECT 79.73 5.945 79.9 6.115 ;
        RECT 79.73 2.765 79.9 2.935 ;
      LAYER via1 ;
        RECT 79.745 5.94 79.895 6.09 ;
        RECT 79.755 2.805 79.905 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.235 5.945 0.405 7.22 ;
      LAYER met1 ;
        RECT 0.175 5.945 0.635 6.115 ;
        RECT 0.175 5.915 0.465 6.145 ;
      LAYER mcon ;
        RECT 0.235 5.945 0.405 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.37 4.255 2.175 4.635 ;
      LAYER li1 ;
        RECT 0 4.44 84.425 4.745 ;
        RECT 1.835 4.135 84.425 4.745 ;
        RECT 82.29 4.13 84.27 4.75 ;
        RECT 83.45 3.4 83.62 5.48 ;
        RECT 82.46 3.4 82.63 5.48 ;
        RECT 79.72 3.405 79.89 5.475 ;
        RECT 77.93 3.635 78.1 4.745 ;
        RECT 76.97 3.635 77.14 4.745 ;
        RECT 74.53 3.635 74.7 4.745 ;
        RECT 74.105 4.135 74.275 5.475 ;
        RECT 73.53 3.635 73.7 4.745 ;
        RECT 72.57 3.635 72.74 4.745 ;
        RECT 70.13 3.635 70.3 4.745 ;
        RECT 65.965 4.13 67.945 4.75 ;
        RECT 67.125 3.4 67.295 5.48 ;
        RECT 66.135 3.4 66.305 5.48 ;
        RECT 63.395 3.405 63.565 5.475 ;
        RECT 61.605 3.635 61.775 4.745 ;
        RECT 60.645 3.635 60.815 4.745 ;
        RECT 58.205 3.635 58.375 4.745 ;
        RECT 57.78 4.135 57.95 5.475 ;
        RECT 57.205 3.635 57.375 4.745 ;
        RECT 56.245 3.635 56.415 4.745 ;
        RECT 53.805 3.635 53.975 4.745 ;
        RECT 49.64 4.13 51.62 4.75 ;
        RECT 50.8 3.4 50.97 5.48 ;
        RECT 49.81 3.4 49.98 5.48 ;
        RECT 47.07 3.405 47.24 5.475 ;
        RECT 45.28 3.635 45.45 4.745 ;
        RECT 44.32 3.635 44.49 4.745 ;
        RECT 41.88 3.635 42.05 4.745 ;
        RECT 41.455 4.135 41.625 5.475 ;
        RECT 40.88 3.635 41.05 4.745 ;
        RECT 39.92 3.635 40.09 4.745 ;
        RECT 37.48 3.635 37.65 4.745 ;
        RECT 33.315 4.13 35.295 4.75 ;
        RECT 34.475 3.4 34.645 5.48 ;
        RECT 33.485 3.4 33.655 5.48 ;
        RECT 30.745 3.405 30.915 5.475 ;
        RECT 28.955 3.635 29.125 4.745 ;
        RECT 27.995 3.635 28.165 4.745 ;
        RECT 25.555 3.635 25.725 4.745 ;
        RECT 25.13 4.135 25.3 5.475 ;
        RECT 24.555 3.635 24.725 4.745 ;
        RECT 23.595 3.635 23.765 4.745 ;
        RECT 21.155 3.635 21.325 4.745 ;
        RECT 16.99 4.13 18.97 4.75 ;
        RECT 18.15 3.4 18.32 5.48 ;
        RECT 17.16 3.4 17.33 5.48 ;
        RECT 14.42 3.405 14.59 5.475 ;
        RECT 12.63 3.635 12.8 4.745 ;
        RECT 11.67 3.635 11.84 4.745 ;
        RECT 9.23 3.635 9.4 4.745 ;
        RECT 8.805 4.135 8.975 5.475 ;
        RECT 8.23 3.635 8.4 4.745 ;
        RECT 7.27 3.635 7.44 4.745 ;
        RECT 4.83 3.635 5 4.745 ;
        RECT 2.035 4.135 2.205 8.305 ;
        RECT 0 4.135 84.425 4.33 ;
        RECT 0 4.135 1.665 4.745 ;
        RECT 0.225 4.135 0.395 5.475 ;
      LAYER met2 ;
        RECT 1.56 4.255 1.94 4.635 ;
      LAYER met1 ;
        RECT 0 4.135 84.425 4.745 ;
        RECT 82.29 4.13 84.27 4.75 ;
        RECT 68.84 3.98 78.5 4.745 ;
        RECT 65.965 4.13 67.945 4.75 ;
        RECT 52.515 3.98 62.175 4.745 ;
        RECT 49.64 4.13 51.62 4.75 ;
        RECT 36.19 3.98 45.85 4.745 ;
        RECT 33.315 4.13 35.295 4.75 ;
        RECT 19.865 3.98 29.525 4.745 ;
        RECT 16.99 4.13 18.97 4.75 ;
        RECT 3.54 3.98 13.2 4.745 ;
        RECT 1.975 6.655 2.265 6.885 ;
        RECT 1.805 6.685 2.265 6.855 ;
      LAYER via2 ;
        RECT 1.65 4.345 1.85 4.545 ;
      LAYER mcon ;
        RECT 2.035 6.685 2.205 6.855 ;
        RECT 2.345 4.545 2.515 4.715 ;
        RECT 3.685 4.135 3.855 4.305 ;
        RECT 4.145 4.135 4.315 4.305 ;
        RECT 4.605 4.135 4.775 4.305 ;
        RECT 5.065 4.135 5.235 4.305 ;
        RECT 5.525 4.135 5.695 4.305 ;
        RECT 5.985 4.135 6.155 4.305 ;
        RECT 6.445 4.135 6.615 4.305 ;
        RECT 6.905 4.135 7.075 4.305 ;
        RECT 7.365 4.135 7.535 4.305 ;
        RECT 7.825 4.135 7.995 4.305 ;
        RECT 8.285 4.135 8.455 4.305 ;
        RECT 8.745 4.135 8.915 4.305 ;
        RECT 9.205 4.135 9.375 4.305 ;
        RECT 9.665 4.135 9.835 4.305 ;
        RECT 10.125 4.135 10.295 4.305 ;
        RECT 10.585 4.135 10.755 4.305 ;
        RECT 10.925 4.545 11.095 4.715 ;
        RECT 11.045 4.135 11.215 4.305 ;
        RECT 11.505 4.135 11.675 4.305 ;
        RECT 11.965 4.135 12.135 4.305 ;
        RECT 12.425 4.135 12.595 4.305 ;
        RECT 12.885 4.135 13.055 4.305 ;
        RECT 16.54 4.545 16.71 4.715 ;
        RECT 16.54 4.165 16.71 4.335 ;
        RECT 17.24 4.55 17.41 4.72 ;
        RECT 17.24 4.16 17.41 4.33 ;
        RECT 18.23 4.55 18.4 4.72 ;
        RECT 18.23 4.16 18.4 4.33 ;
        RECT 20.01 4.135 20.18 4.305 ;
        RECT 20.47 4.135 20.64 4.305 ;
        RECT 20.93 4.135 21.1 4.305 ;
        RECT 21.39 4.135 21.56 4.305 ;
        RECT 21.85 4.135 22.02 4.305 ;
        RECT 22.31 4.135 22.48 4.305 ;
        RECT 22.77 4.135 22.94 4.305 ;
        RECT 23.23 4.135 23.4 4.305 ;
        RECT 23.69 4.135 23.86 4.305 ;
        RECT 24.15 4.135 24.32 4.305 ;
        RECT 24.61 4.135 24.78 4.305 ;
        RECT 25.07 4.135 25.24 4.305 ;
        RECT 25.53 4.135 25.7 4.305 ;
        RECT 25.99 4.135 26.16 4.305 ;
        RECT 26.45 4.135 26.62 4.305 ;
        RECT 26.91 4.135 27.08 4.305 ;
        RECT 27.25 4.545 27.42 4.715 ;
        RECT 27.37 4.135 27.54 4.305 ;
        RECT 27.83 4.135 28 4.305 ;
        RECT 28.29 4.135 28.46 4.305 ;
        RECT 28.75 4.135 28.92 4.305 ;
        RECT 29.21 4.135 29.38 4.305 ;
        RECT 32.865 4.545 33.035 4.715 ;
        RECT 32.865 4.165 33.035 4.335 ;
        RECT 33.565 4.55 33.735 4.72 ;
        RECT 33.565 4.16 33.735 4.33 ;
        RECT 34.555 4.55 34.725 4.72 ;
        RECT 34.555 4.16 34.725 4.33 ;
        RECT 36.335 4.135 36.505 4.305 ;
        RECT 36.795 4.135 36.965 4.305 ;
        RECT 37.255 4.135 37.425 4.305 ;
        RECT 37.715 4.135 37.885 4.305 ;
        RECT 38.175 4.135 38.345 4.305 ;
        RECT 38.635 4.135 38.805 4.305 ;
        RECT 39.095 4.135 39.265 4.305 ;
        RECT 39.555 4.135 39.725 4.305 ;
        RECT 40.015 4.135 40.185 4.305 ;
        RECT 40.475 4.135 40.645 4.305 ;
        RECT 40.935 4.135 41.105 4.305 ;
        RECT 41.395 4.135 41.565 4.305 ;
        RECT 41.855 4.135 42.025 4.305 ;
        RECT 42.315 4.135 42.485 4.305 ;
        RECT 42.775 4.135 42.945 4.305 ;
        RECT 43.235 4.135 43.405 4.305 ;
        RECT 43.575 4.545 43.745 4.715 ;
        RECT 43.695 4.135 43.865 4.305 ;
        RECT 44.155 4.135 44.325 4.305 ;
        RECT 44.615 4.135 44.785 4.305 ;
        RECT 45.075 4.135 45.245 4.305 ;
        RECT 45.535 4.135 45.705 4.305 ;
        RECT 49.19 4.545 49.36 4.715 ;
        RECT 49.19 4.165 49.36 4.335 ;
        RECT 49.89 4.55 50.06 4.72 ;
        RECT 49.89 4.16 50.06 4.33 ;
        RECT 50.88 4.55 51.05 4.72 ;
        RECT 50.88 4.16 51.05 4.33 ;
        RECT 52.66 4.135 52.83 4.305 ;
        RECT 53.12 4.135 53.29 4.305 ;
        RECT 53.58 4.135 53.75 4.305 ;
        RECT 54.04 4.135 54.21 4.305 ;
        RECT 54.5 4.135 54.67 4.305 ;
        RECT 54.96 4.135 55.13 4.305 ;
        RECT 55.42 4.135 55.59 4.305 ;
        RECT 55.88 4.135 56.05 4.305 ;
        RECT 56.34 4.135 56.51 4.305 ;
        RECT 56.8 4.135 56.97 4.305 ;
        RECT 57.26 4.135 57.43 4.305 ;
        RECT 57.72 4.135 57.89 4.305 ;
        RECT 58.18 4.135 58.35 4.305 ;
        RECT 58.64 4.135 58.81 4.305 ;
        RECT 59.1 4.135 59.27 4.305 ;
        RECT 59.56 4.135 59.73 4.305 ;
        RECT 59.9 4.545 60.07 4.715 ;
        RECT 60.02 4.135 60.19 4.305 ;
        RECT 60.48 4.135 60.65 4.305 ;
        RECT 60.94 4.135 61.11 4.305 ;
        RECT 61.4 4.135 61.57 4.305 ;
        RECT 61.86 4.135 62.03 4.305 ;
        RECT 65.515 4.545 65.685 4.715 ;
        RECT 65.515 4.165 65.685 4.335 ;
        RECT 66.215 4.55 66.385 4.72 ;
        RECT 66.215 4.16 66.385 4.33 ;
        RECT 67.205 4.55 67.375 4.72 ;
        RECT 67.205 4.16 67.375 4.33 ;
        RECT 68.985 4.135 69.155 4.305 ;
        RECT 69.445 4.135 69.615 4.305 ;
        RECT 69.905 4.135 70.075 4.305 ;
        RECT 70.365 4.135 70.535 4.305 ;
        RECT 70.825 4.135 70.995 4.305 ;
        RECT 71.285 4.135 71.455 4.305 ;
        RECT 71.745 4.135 71.915 4.305 ;
        RECT 72.205 4.135 72.375 4.305 ;
        RECT 72.665 4.135 72.835 4.305 ;
        RECT 73.125 4.135 73.295 4.305 ;
        RECT 73.585 4.135 73.755 4.305 ;
        RECT 74.045 4.135 74.215 4.305 ;
        RECT 74.505 4.135 74.675 4.305 ;
        RECT 74.965 4.135 75.135 4.305 ;
        RECT 75.425 4.135 75.595 4.305 ;
        RECT 75.885 4.135 76.055 4.305 ;
        RECT 76.225 4.545 76.395 4.715 ;
        RECT 76.345 4.135 76.515 4.305 ;
        RECT 76.805 4.135 76.975 4.305 ;
        RECT 77.265 4.135 77.435 4.305 ;
        RECT 77.725 4.135 77.895 4.305 ;
        RECT 78.185 4.135 78.355 4.305 ;
        RECT 81.84 4.545 82.01 4.715 ;
        RECT 81.84 4.165 82.01 4.335 ;
        RECT 82.54 4.55 82.71 4.72 ;
        RECT 82.54 4.16 82.71 4.33 ;
        RECT 83.53 4.55 83.7 4.72 ;
        RECT 83.53 4.16 83.7 4.33 ;
      LAYER via1 ;
        RECT 1.675 4.37 1.825 4.52 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 77.73 2.975 78.06 3.705 ;
        RECT 61.405 2.975 61.735 3.705 ;
        RECT 45.08 2.975 45.41 3.705 ;
        RECT 28.755 2.975 29.085 3.705 ;
        RECT 12.43 2.975 12.76 3.705 ;
        RECT 0.01 8.5 0.815 8.88 ;
        RECT 0 0 0.805 0.38 ;
      LAYER li1 ;
        RECT 84.245 0 84.425 0.305 ;
        RECT 0.465 0 84.425 0.3 ;
        RECT 83.45 0 83.62 0.93 ;
        RECT 82.46 0 82.63 0.93 ;
        RECT 67.92 0 82.295 0.305 ;
        RECT 79.72 0 79.89 0.935 ;
        RECT 68.84 0 78.655 1.585 ;
        RECT 76.97 0 77.14 2.085 ;
        RECT 75.01 0 75.18 2.085 ;
        RECT 74.94 0 75.18 1.595 ;
        RECT 73.39 0 73.585 1.595 ;
        RECT 72.57 0 72.74 2.085 ;
        RECT 71.61 0 71.78 2.085 ;
        RECT 71.265 0 71.46 1.595 ;
        RECT 71.09 0 71.26 2.085 ;
        RECT 70.13 0 70.3 2.085 ;
        RECT 69.17 0 69.34 2.085 ;
        RECT 68.965 0 69.16 1.595 ;
        RECT 67.125 0 67.295 0.93 ;
        RECT 66.135 0 66.305 0.93 ;
        RECT 51.595 0 65.97 0.305 ;
        RECT 63.395 0 63.565 0.935 ;
        RECT 52.515 0 62.33 1.585 ;
        RECT 60.645 0 60.815 2.085 ;
        RECT 58.685 0 58.855 2.085 ;
        RECT 58.615 0 58.855 1.595 ;
        RECT 57.065 0 57.26 1.595 ;
        RECT 56.245 0 56.415 2.085 ;
        RECT 55.285 0 55.455 2.085 ;
        RECT 54.94 0 55.135 1.595 ;
        RECT 54.765 0 54.935 2.085 ;
        RECT 53.805 0 53.975 2.085 ;
        RECT 52.845 0 53.015 2.085 ;
        RECT 52.64 0 52.835 1.595 ;
        RECT 50.8 0 50.97 0.93 ;
        RECT 49.81 0 49.98 0.93 ;
        RECT 35.27 0 49.645 0.305 ;
        RECT 47.07 0 47.24 0.935 ;
        RECT 36.19 0 46.005 1.585 ;
        RECT 44.32 0 44.49 2.085 ;
        RECT 42.36 0 42.53 2.085 ;
        RECT 42.29 0 42.53 1.595 ;
        RECT 40.74 0 40.935 1.595 ;
        RECT 39.92 0 40.09 2.085 ;
        RECT 38.96 0 39.13 2.085 ;
        RECT 38.615 0 38.81 1.595 ;
        RECT 38.44 0 38.61 2.085 ;
        RECT 37.48 0 37.65 2.085 ;
        RECT 36.52 0 36.69 2.085 ;
        RECT 36.315 0 36.51 1.595 ;
        RECT 34.475 0 34.645 0.93 ;
        RECT 33.485 0 33.655 0.93 ;
        RECT 18.945 0 33.32 0.305 ;
        RECT 30.745 0 30.915 0.935 ;
        RECT 19.865 0 29.68 1.585 ;
        RECT 27.995 0 28.165 2.085 ;
        RECT 26.035 0 26.205 2.085 ;
        RECT 25.965 0 26.205 1.595 ;
        RECT 24.415 0 24.61 1.595 ;
        RECT 23.595 0 23.765 2.085 ;
        RECT 22.635 0 22.805 2.085 ;
        RECT 22.29 0 22.485 1.595 ;
        RECT 22.115 0 22.285 2.085 ;
        RECT 21.155 0 21.325 2.085 ;
        RECT 20.195 0 20.365 2.085 ;
        RECT 19.99 0 20.185 1.595 ;
        RECT 18.15 0 18.32 0.93 ;
        RECT 17.16 0 17.33 0.93 ;
        RECT 0 0.245 16.995 0.305 ;
        RECT 14.42 0 14.59 0.935 ;
        RECT 3.54 0 13.355 1.585 ;
        RECT 11.67 0 11.84 2.085 ;
        RECT 9.71 0 9.88 2.085 ;
        RECT 9.64 0 9.88 1.595 ;
        RECT 8.09 0 8.285 1.595 ;
        RECT 7.27 0 7.44 2.085 ;
        RECT 6.31 0 6.48 2.085 ;
        RECT 5.965 0 6.16 1.595 ;
        RECT 5.79 0 5.96 2.085 ;
        RECT 4.83 0 5 2.085 ;
        RECT 3.87 0 4.04 2.085 ;
        RECT 3.665 0 3.86 1.595 ;
        RECT 0 0.245 0.805 0.315 ;
        RECT 0.295 0.245 0.465 0.335 ;
        RECT 0 0 84.425 0.075 ;
        RECT 0 0 0.295 0.315 ;
        RECT 0 8.58 84.425 8.88 ;
        RECT 84.245 8.575 84.425 8.88 ;
        RECT 83.45 7.95 83.62 8.88 ;
        RECT 82.46 7.95 82.63 8.88 ;
        RECT 67.92 8.575 82.295 8.88 ;
        RECT 79.72 7.945 79.89 8.88 ;
        RECT 74.105 7.945 74.275 8.88 ;
        RECT 67.125 7.95 67.295 8.88 ;
        RECT 66.135 7.95 66.305 8.88 ;
        RECT 51.595 8.575 65.97 8.88 ;
        RECT 63.395 7.945 63.565 8.88 ;
        RECT 57.78 7.945 57.95 8.88 ;
        RECT 50.8 7.95 50.97 8.88 ;
        RECT 49.81 7.95 49.98 8.88 ;
        RECT 35.27 8.575 49.645 8.88 ;
        RECT 47.07 7.945 47.24 8.88 ;
        RECT 41.455 7.945 41.625 8.88 ;
        RECT 34.475 7.95 34.645 8.88 ;
        RECT 33.485 7.95 33.655 8.88 ;
        RECT 18.945 8.575 33.32 8.88 ;
        RECT 30.745 7.945 30.915 8.88 ;
        RECT 25.13 7.945 25.3 8.88 ;
        RECT 18.15 7.95 18.32 8.88 ;
        RECT 17.16 7.95 17.33 8.88 ;
        RECT 0 8.575 16.995 8.88 ;
        RECT 14.42 7.945 14.59 8.88 ;
        RECT 8.805 7.945 8.975 8.88 ;
        RECT 0.01 8.565 0.815 8.88 ;
        RECT 0.225 8.545 0.475 8.88 ;
        RECT 0.225 7.945 0.395 8.88 ;
        RECT 77.93 2.575 78.1 2.945 ;
        RECT 77.61 2.575 78.1 2.745 ;
        RECT 75.97 2.575 76.14 2.945 ;
        RECT 75.65 2.575 76.14 2.745 ;
        RECT 75.11 6.075 75.28 8.025 ;
        RECT 75.055 7.855 75.225 8.305 ;
        RECT 75.055 5.015 75.225 6.245 ;
        RECT 61.605 2.575 61.775 2.945 ;
        RECT 61.285 2.575 61.775 2.745 ;
        RECT 59.645 2.575 59.815 2.945 ;
        RECT 59.325 2.575 59.815 2.745 ;
        RECT 58.785 6.075 58.955 8.025 ;
        RECT 58.73 7.855 58.9 8.305 ;
        RECT 58.73 5.015 58.9 6.245 ;
        RECT 45.28 2.575 45.45 2.945 ;
        RECT 44.96 2.575 45.45 2.745 ;
        RECT 43.32 2.575 43.49 2.945 ;
        RECT 43 2.575 43.49 2.745 ;
        RECT 42.46 6.075 42.63 8.025 ;
        RECT 42.405 7.855 42.575 8.305 ;
        RECT 42.405 5.015 42.575 6.245 ;
        RECT 28.955 2.575 29.125 2.945 ;
        RECT 28.635 2.575 29.125 2.745 ;
        RECT 26.995 2.575 27.165 2.945 ;
        RECT 26.675 2.575 27.165 2.745 ;
        RECT 26.135 6.075 26.305 8.025 ;
        RECT 26.08 7.855 26.25 8.305 ;
        RECT 26.08 5.015 26.25 6.245 ;
        RECT 12.63 2.575 12.8 2.945 ;
        RECT 12.31 2.575 12.8 2.745 ;
        RECT 10.67 2.575 10.84 2.945 ;
        RECT 10.35 2.575 10.84 2.745 ;
        RECT 9.81 6.075 9.98 8.025 ;
        RECT 9.755 7.855 9.925 8.305 ;
        RECT 9.755 5.015 9.925 6.245 ;
      LAYER met2 ;
        RECT 77.755 2.955 78.035 3.325 ;
        RECT 77.765 2.7 78.025 3.325 ;
        RECT 61.43 2.955 61.71 3.325 ;
        RECT 61.44 2.7 61.7 3.325 ;
        RECT 45.105 2.955 45.385 3.325 ;
        RECT 45.115 2.7 45.375 3.325 ;
        RECT 28.78 2.955 29.06 3.325 ;
        RECT 28.79 2.7 29.05 3.325 ;
        RECT 12.455 2.955 12.735 3.325 ;
        RECT 12.465 2.7 12.725 3.325 ;
        RECT 0.2 8.5 0.58 8.88 ;
        RECT 0.19 0 0.57 0.38 ;
        RECT 0.235 0 0.41 8.88 ;
      LAYER met1 ;
        RECT 84.245 0 84.425 0.305 ;
        RECT 0 0 84.425 0.3 ;
        RECT 67.92 0 82.295 0.305 ;
        RECT 78.47 0 78.655 2.945 ;
        RECT 77.705 2.79 78.655 2.945 ;
        RECT 77.735 2.76 78.655 2.945 ;
        RECT 68.84 0 78.655 1.74 ;
        RECT 77.735 2.745 78.16 2.975 ;
        RECT 77.735 2.73 78.055 2.99 ;
        RECT 76.245 2.93 78.01 3.055 ;
        RECT 76.245 2.93 77.845 3.07 ;
        RECT 75.91 2.79 76.385 2.975 ;
        RECT 75.91 2.745 76.2 2.975 ;
        RECT 51.595 0 65.97 0.305 ;
        RECT 62.145 0 62.33 2.945 ;
        RECT 61.38 2.79 62.33 2.945 ;
        RECT 61.41 2.76 62.33 2.945 ;
        RECT 52.515 0 62.33 1.74 ;
        RECT 61.41 2.745 61.835 2.975 ;
        RECT 61.41 2.73 61.73 2.99 ;
        RECT 59.92 2.93 61.685 3.055 ;
        RECT 59.92 2.93 61.52 3.07 ;
        RECT 59.585 2.79 60.06 2.975 ;
        RECT 59.585 2.745 59.875 2.975 ;
        RECT 35.27 0 49.645 0.305 ;
        RECT 45.82 0 46.005 2.945 ;
        RECT 45.055 2.79 46.005 2.945 ;
        RECT 45.085 2.76 46.005 2.945 ;
        RECT 36.19 0 46.005 1.74 ;
        RECT 45.085 2.745 45.51 2.975 ;
        RECT 45.085 2.73 45.405 2.99 ;
        RECT 43.595 2.93 45.36 3.055 ;
        RECT 43.595 2.93 45.195 3.07 ;
        RECT 43.26 2.79 43.735 2.975 ;
        RECT 43.26 2.745 43.55 2.975 ;
        RECT 18.945 0 33.32 0.305 ;
        RECT 29.495 0 29.68 2.945 ;
        RECT 28.73 2.79 29.68 2.945 ;
        RECT 28.76 2.76 29.68 2.945 ;
        RECT 19.865 0 29.68 1.74 ;
        RECT 28.76 2.745 29.185 2.975 ;
        RECT 28.76 2.73 29.08 2.99 ;
        RECT 27.27 2.93 29.035 3.055 ;
        RECT 27.27 2.93 28.87 3.07 ;
        RECT 26.935 2.79 27.41 2.975 ;
        RECT 26.935 2.745 27.225 2.975 ;
        RECT 0 0 16.995 0.305 ;
        RECT 13.17 0 13.355 2.945 ;
        RECT 12.405 2.79 13.355 2.945 ;
        RECT 12.435 2.76 13.355 2.945 ;
        RECT 3.54 0 13.355 1.74 ;
        RECT 12.435 2.745 12.86 2.975 ;
        RECT 12.435 2.73 12.755 2.99 ;
        RECT 10.945 2.93 12.71 3.055 ;
        RECT 10.945 2.93 12.545 3.07 ;
        RECT 10.61 2.79 11.085 2.975 ;
        RECT 10.61 2.745 10.9 2.975 ;
        RECT 0 0 0.805 0.315 ;
        RECT 0.205 0 0.555 0.335 ;
        RECT 0 8.58 84.425 8.88 ;
        RECT 84.245 8.575 84.425 8.88 ;
        RECT 67.92 8.575 82.295 8.88 ;
        RECT 75.05 6.285 75.34 6.515 ;
        RECT 74.675 6.315 75.34 6.485 ;
        RECT 74.675 6.315 74.85 8.88 ;
        RECT 51.595 8.575 65.97 8.88 ;
        RECT 58.725 6.285 59.015 6.515 ;
        RECT 58.35 6.315 59.015 6.485 ;
        RECT 58.35 6.315 58.525 8.88 ;
        RECT 35.27 8.575 49.645 8.88 ;
        RECT 42.4 6.285 42.69 6.515 ;
        RECT 42.025 6.315 42.69 6.485 ;
        RECT 42.025 6.315 42.2 8.88 ;
        RECT 18.945 8.575 33.32 8.88 ;
        RECT 26.075 6.285 26.365 6.515 ;
        RECT 25.7 6.315 26.365 6.485 ;
        RECT 25.7 6.315 25.875 8.88 ;
        RECT 0 8.575 16.995 8.88 ;
        RECT 9.75 6.285 10.04 6.515 ;
        RECT 9.375 6.315 10.04 6.485 ;
        RECT 9.375 6.315 9.55 8.88 ;
        RECT 0.01 8.565 0.815 8.88 ;
        RECT 0.215 8.545 0.565 8.88 ;
      LAYER via2 ;
        RECT 0.28 0.09 0.48 0.29 ;
        RECT 0.29 8.59 0.49 8.79 ;
        RECT 12.495 3.04 12.695 3.24 ;
        RECT 28.82 3.04 29.02 3.24 ;
        RECT 45.145 3.04 45.345 3.24 ;
        RECT 61.47 3.04 61.67 3.24 ;
        RECT 77.795 3.04 77.995 3.24 ;
      LAYER mcon ;
        RECT 0.305 8.605 0.475 8.775 ;
        RECT 0.985 8.605 1.155 8.775 ;
        RECT 1.665 8.605 1.835 8.775 ;
        RECT 2.345 8.605 2.515 8.775 ;
        RECT 3.685 1.415 3.855 1.585 ;
        RECT 4.145 1.415 4.315 1.585 ;
        RECT 4.605 1.415 4.775 1.585 ;
        RECT 5.065 1.415 5.235 1.585 ;
        RECT 5.525 1.415 5.695 1.585 ;
        RECT 5.985 1.415 6.155 1.585 ;
        RECT 6.445 1.415 6.615 1.585 ;
        RECT 6.905 1.415 7.075 1.585 ;
        RECT 7.365 1.415 7.535 1.585 ;
        RECT 7.825 1.415 7.995 1.585 ;
        RECT 8.285 1.415 8.455 1.585 ;
        RECT 8.745 1.415 8.915 1.585 ;
        RECT 8.885 8.605 9.055 8.775 ;
        RECT 9.205 1.415 9.375 1.585 ;
        RECT 9.565 8.605 9.735 8.775 ;
        RECT 9.665 1.415 9.835 1.585 ;
        RECT 9.81 6.315 9.98 6.485 ;
        RECT 10.125 1.415 10.295 1.585 ;
        RECT 10.245 8.605 10.415 8.775 ;
        RECT 10.585 1.415 10.755 1.585 ;
        RECT 10.67 2.775 10.84 2.945 ;
        RECT 10.925 8.605 11.095 8.775 ;
        RECT 11.045 1.415 11.215 1.585 ;
        RECT 11.505 1.415 11.675 1.585 ;
        RECT 11.965 1.415 12.135 1.585 ;
        RECT 12.425 1.415 12.595 1.585 ;
        RECT 12.63 2.775 12.8 2.945 ;
        RECT 12.885 1.415 13.055 1.585 ;
        RECT 14.5 8.605 14.67 8.775 ;
        RECT 14.5 0.105 14.67 0.275 ;
        RECT 15.18 8.605 15.35 8.775 ;
        RECT 15.18 0.105 15.35 0.275 ;
        RECT 15.86 8.605 16.03 8.775 ;
        RECT 15.86 0.105 16.03 0.275 ;
        RECT 16.54 8.605 16.71 8.775 ;
        RECT 16.54 0.105 16.71 0.275 ;
        RECT 17.24 8.61 17.41 8.78 ;
        RECT 17.24 0.1 17.41 0.27 ;
        RECT 18.23 8.61 18.4 8.78 ;
        RECT 18.23 0.1 18.4 0.27 ;
        RECT 20.01 1.415 20.18 1.585 ;
        RECT 20.47 1.415 20.64 1.585 ;
        RECT 20.93 1.415 21.1 1.585 ;
        RECT 21.39 1.415 21.56 1.585 ;
        RECT 21.85 1.415 22.02 1.585 ;
        RECT 22.31 1.415 22.48 1.585 ;
        RECT 22.77 1.415 22.94 1.585 ;
        RECT 23.23 1.415 23.4 1.585 ;
        RECT 23.69 1.415 23.86 1.585 ;
        RECT 24.15 1.415 24.32 1.585 ;
        RECT 24.61 1.415 24.78 1.585 ;
        RECT 25.07 1.415 25.24 1.585 ;
        RECT 25.21 8.605 25.38 8.775 ;
        RECT 25.53 1.415 25.7 1.585 ;
        RECT 25.89 8.605 26.06 8.775 ;
        RECT 25.99 1.415 26.16 1.585 ;
        RECT 26.135 6.315 26.305 6.485 ;
        RECT 26.45 1.415 26.62 1.585 ;
        RECT 26.57 8.605 26.74 8.775 ;
        RECT 26.91 1.415 27.08 1.585 ;
        RECT 26.995 2.775 27.165 2.945 ;
        RECT 27.25 8.605 27.42 8.775 ;
        RECT 27.37 1.415 27.54 1.585 ;
        RECT 27.83 1.415 28 1.585 ;
        RECT 28.29 1.415 28.46 1.585 ;
        RECT 28.75 1.415 28.92 1.585 ;
        RECT 28.955 2.775 29.125 2.945 ;
        RECT 29.21 1.415 29.38 1.585 ;
        RECT 30.825 8.605 30.995 8.775 ;
        RECT 30.825 0.105 30.995 0.275 ;
        RECT 31.505 8.605 31.675 8.775 ;
        RECT 31.505 0.105 31.675 0.275 ;
        RECT 32.185 8.605 32.355 8.775 ;
        RECT 32.185 0.105 32.355 0.275 ;
        RECT 32.865 8.605 33.035 8.775 ;
        RECT 32.865 0.105 33.035 0.275 ;
        RECT 33.565 8.61 33.735 8.78 ;
        RECT 33.565 0.1 33.735 0.27 ;
        RECT 34.555 8.61 34.725 8.78 ;
        RECT 34.555 0.1 34.725 0.27 ;
        RECT 36.335 1.415 36.505 1.585 ;
        RECT 36.795 1.415 36.965 1.585 ;
        RECT 37.255 1.415 37.425 1.585 ;
        RECT 37.715 1.415 37.885 1.585 ;
        RECT 38.175 1.415 38.345 1.585 ;
        RECT 38.635 1.415 38.805 1.585 ;
        RECT 39.095 1.415 39.265 1.585 ;
        RECT 39.555 1.415 39.725 1.585 ;
        RECT 40.015 1.415 40.185 1.585 ;
        RECT 40.475 1.415 40.645 1.585 ;
        RECT 40.935 1.415 41.105 1.585 ;
        RECT 41.395 1.415 41.565 1.585 ;
        RECT 41.535 8.605 41.705 8.775 ;
        RECT 41.855 1.415 42.025 1.585 ;
        RECT 42.215 8.605 42.385 8.775 ;
        RECT 42.315 1.415 42.485 1.585 ;
        RECT 42.46 6.315 42.63 6.485 ;
        RECT 42.775 1.415 42.945 1.585 ;
        RECT 42.895 8.605 43.065 8.775 ;
        RECT 43.235 1.415 43.405 1.585 ;
        RECT 43.32 2.775 43.49 2.945 ;
        RECT 43.575 8.605 43.745 8.775 ;
        RECT 43.695 1.415 43.865 1.585 ;
        RECT 44.155 1.415 44.325 1.585 ;
        RECT 44.615 1.415 44.785 1.585 ;
        RECT 45.075 1.415 45.245 1.585 ;
        RECT 45.28 2.775 45.45 2.945 ;
        RECT 45.535 1.415 45.705 1.585 ;
        RECT 47.15 8.605 47.32 8.775 ;
        RECT 47.15 0.105 47.32 0.275 ;
        RECT 47.83 8.605 48 8.775 ;
        RECT 47.83 0.105 48 0.275 ;
        RECT 48.51 8.605 48.68 8.775 ;
        RECT 48.51 0.105 48.68 0.275 ;
        RECT 49.19 8.605 49.36 8.775 ;
        RECT 49.19 0.105 49.36 0.275 ;
        RECT 49.89 8.61 50.06 8.78 ;
        RECT 49.89 0.1 50.06 0.27 ;
        RECT 50.88 8.61 51.05 8.78 ;
        RECT 50.88 0.1 51.05 0.27 ;
        RECT 52.66 1.415 52.83 1.585 ;
        RECT 53.12 1.415 53.29 1.585 ;
        RECT 53.58 1.415 53.75 1.585 ;
        RECT 54.04 1.415 54.21 1.585 ;
        RECT 54.5 1.415 54.67 1.585 ;
        RECT 54.96 1.415 55.13 1.585 ;
        RECT 55.42 1.415 55.59 1.585 ;
        RECT 55.88 1.415 56.05 1.585 ;
        RECT 56.34 1.415 56.51 1.585 ;
        RECT 56.8 1.415 56.97 1.585 ;
        RECT 57.26 1.415 57.43 1.585 ;
        RECT 57.72 1.415 57.89 1.585 ;
        RECT 57.86 8.605 58.03 8.775 ;
        RECT 58.18 1.415 58.35 1.585 ;
        RECT 58.54 8.605 58.71 8.775 ;
        RECT 58.64 1.415 58.81 1.585 ;
        RECT 58.785 6.315 58.955 6.485 ;
        RECT 59.1 1.415 59.27 1.585 ;
        RECT 59.22 8.605 59.39 8.775 ;
        RECT 59.56 1.415 59.73 1.585 ;
        RECT 59.645 2.775 59.815 2.945 ;
        RECT 59.9 8.605 60.07 8.775 ;
        RECT 60.02 1.415 60.19 1.585 ;
        RECT 60.48 1.415 60.65 1.585 ;
        RECT 60.94 1.415 61.11 1.585 ;
        RECT 61.4 1.415 61.57 1.585 ;
        RECT 61.605 2.775 61.775 2.945 ;
        RECT 61.86 1.415 62.03 1.585 ;
        RECT 63.475 8.605 63.645 8.775 ;
        RECT 63.475 0.105 63.645 0.275 ;
        RECT 64.155 8.605 64.325 8.775 ;
        RECT 64.155 0.105 64.325 0.275 ;
        RECT 64.835 8.605 65.005 8.775 ;
        RECT 64.835 0.105 65.005 0.275 ;
        RECT 65.515 8.605 65.685 8.775 ;
        RECT 65.515 0.105 65.685 0.275 ;
        RECT 66.215 8.61 66.385 8.78 ;
        RECT 66.215 0.1 66.385 0.27 ;
        RECT 67.205 8.61 67.375 8.78 ;
        RECT 67.205 0.1 67.375 0.27 ;
        RECT 68.985 1.415 69.155 1.585 ;
        RECT 69.445 1.415 69.615 1.585 ;
        RECT 69.905 1.415 70.075 1.585 ;
        RECT 70.365 1.415 70.535 1.585 ;
        RECT 70.825 1.415 70.995 1.585 ;
        RECT 71.285 1.415 71.455 1.585 ;
        RECT 71.745 1.415 71.915 1.585 ;
        RECT 72.205 1.415 72.375 1.585 ;
        RECT 72.665 1.415 72.835 1.585 ;
        RECT 73.125 1.415 73.295 1.585 ;
        RECT 73.585 1.415 73.755 1.585 ;
        RECT 74.045 1.415 74.215 1.585 ;
        RECT 74.185 8.605 74.355 8.775 ;
        RECT 74.505 1.415 74.675 1.585 ;
        RECT 74.865 8.605 75.035 8.775 ;
        RECT 74.965 1.415 75.135 1.585 ;
        RECT 75.11 6.315 75.28 6.485 ;
        RECT 75.425 1.415 75.595 1.585 ;
        RECT 75.545 8.605 75.715 8.775 ;
        RECT 75.885 1.415 76.055 1.585 ;
        RECT 75.97 2.775 76.14 2.945 ;
        RECT 76.225 8.605 76.395 8.775 ;
        RECT 76.345 1.415 76.515 1.585 ;
        RECT 76.805 1.415 76.975 1.585 ;
        RECT 77.265 1.415 77.435 1.585 ;
        RECT 77.725 1.415 77.895 1.585 ;
        RECT 77.93 2.775 78.1 2.945 ;
        RECT 78.185 1.415 78.355 1.585 ;
        RECT 79.8 8.605 79.97 8.775 ;
        RECT 79.8 0.105 79.97 0.275 ;
        RECT 80.48 8.605 80.65 8.775 ;
        RECT 80.48 0.105 80.65 0.275 ;
        RECT 81.16 8.605 81.33 8.775 ;
        RECT 81.16 0.105 81.33 0.275 ;
        RECT 81.84 8.605 82.01 8.775 ;
        RECT 81.84 0.105 82.01 0.275 ;
        RECT 82.54 8.61 82.71 8.78 ;
        RECT 82.54 0.1 82.71 0.27 ;
        RECT 83.53 8.61 83.7 8.78 ;
        RECT 83.53 0.1 83.7 0.27 ;
      LAYER via1 ;
        RECT 0.305 0.115 0.455 0.265 ;
        RECT 0.315 8.615 0.465 8.765 ;
        RECT 12.52 2.785 12.67 2.935 ;
        RECT 28.845 2.785 28.995 2.935 ;
        RECT 45.17 2.785 45.32 2.935 ;
        RECT 61.495 2.785 61.645 2.935 ;
        RECT 77.82 2.785 77.97 2.935 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 75.405 7.055 75.775 7.425 ;
      RECT 75.405 7.09 77.39 7.39 ;
      RECT 77.09 2.28 77.39 7.39 ;
      RECT 74.09 2.015 74.42 2.745 ;
      RECT 73.21 2.015 73.54 2.745 ;
      RECT 76.29 2.28 77.58 2.58 ;
      RECT 77.25 1.85 77.58 2.58 ;
      RECT 73.21 2.28 75.35 2.58 ;
      RECT 75.05 1.965 75.35 2.58 ;
      RECT 76.29 1.98 76.595 2.58 ;
      RECT 75.05 1.965 76.41 2.275 ;
      RECT 73.71 3.535 74.04 3.865 ;
      RECT 72.505 3.55 74.04 3.85 ;
      RECT 72.505 2.43 72.805 3.85 ;
      RECT 72.25 2.415 72.58 2.745 ;
      RECT 59.08 7.055 59.45 7.425 ;
      RECT 59.08 7.09 61.065 7.39 ;
      RECT 60.765 2.28 61.065 7.39 ;
      RECT 57.765 2.015 58.095 2.745 ;
      RECT 56.885 2.015 57.215 2.745 ;
      RECT 59.965 2.28 61.255 2.58 ;
      RECT 60.925 1.85 61.255 2.58 ;
      RECT 56.885 2.28 59.025 2.58 ;
      RECT 58.725 1.965 59.025 2.58 ;
      RECT 59.965 1.98 60.27 2.58 ;
      RECT 58.725 1.965 60.085 2.275 ;
      RECT 57.385 3.535 57.715 3.865 ;
      RECT 56.18 3.55 57.715 3.85 ;
      RECT 56.18 2.43 56.48 3.85 ;
      RECT 55.925 2.415 56.255 2.745 ;
      RECT 42.755 7.055 43.125 7.425 ;
      RECT 42.755 7.09 44.74 7.39 ;
      RECT 44.44 2.28 44.74 7.39 ;
      RECT 41.44 2.015 41.77 2.745 ;
      RECT 40.56 2.015 40.89 2.745 ;
      RECT 43.64 2.28 44.93 2.58 ;
      RECT 44.6 1.85 44.93 2.58 ;
      RECT 40.56 2.28 42.7 2.58 ;
      RECT 42.4 1.965 42.7 2.58 ;
      RECT 43.64 1.98 43.945 2.58 ;
      RECT 42.4 1.965 43.76 2.275 ;
      RECT 41.06 3.535 41.39 3.865 ;
      RECT 39.855 3.55 41.39 3.85 ;
      RECT 39.855 2.43 40.155 3.85 ;
      RECT 39.6 2.415 39.93 2.745 ;
      RECT 26.43 7.055 26.8 7.425 ;
      RECT 26.43 7.09 28.415 7.39 ;
      RECT 28.115 2.28 28.415 7.39 ;
      RECT 25.115 2.015 25.445 2.745 ;
      RECT 24.235 2.015 24.565 2.745 ;
      RECT 27.315 2.28 28.605 2.58 ;
      RECT 28.275 1.85 28.605 2.58 ;
      RECT 24.235 2.28 26.375 2.58 ;
      RECT 26.075 1.965 26.375 2.58 ;
      RECT 27.315 1.98 27.62 2.58 ;
      RECT 26.075 1.965 27.435 2.275 ;
      RECT 24.735 3.535 25.065 3.865 ;
      RECT 23.53 3.55 25.065 3.85 ;
      RECT 23.53 2.43 23.83 3.85 ;
      RECT 23.275 2.415 23.605 2.745 ;
      RECT 10.105 7.055 10.475 7.425 ;
      RECT 10.105 7.09 12.09 7.39 ;
      RECT 11.79 2.28 12.09 7.39 ;
      RECT 8.79 2.015 9.12 2.745 ;
      RECT 7.91 2.015 8.24 2.745 ;
      RECT 10.99 2.28 12.28 2.58 ;
      RECT 11.95 1.85 12.28 2.58 ;
      RECT 7.91 2.28 10.05 2.58 ;
      RECT 9.75 1.965 10.05 2.58 ;
      RECT 10.99 1.98 11.295 2.58 ;
      RECT 9.75 1.965 11.11 2.275 ;
      RECT 8.41 3.535 8.74 3.865 ;
      RECT 7.205 3.55 8.74 3.85 ;
      RECT 7.205 2.43 7.505 3.85 ;
      RECT 6.95 2.415 7.28 2.745 ;
      RECT 75.65 2.575 75.98 3.305 ;
      RECT 71.53 2.415 71.86 3.145 ;
      RECT 70.53 1.855 70.86 2.585 ;
      RECT 69.09 2.575 69.42 3.305 ;
      RECT 59.325 2.575 59.655 3.305 ;
      RECT 55.205 2.415 55.535 3.145 ;
      RECT 54.205 1.855 54.535 2.585 ;
      RECT 52.765 2.575 53.095 3.305 ;
      RECT 43 2.575 43.33 3.305 ;
      RECT 38.88 2.415 39.21 3.145 ;
      RECT 37.88 1.855 38.21 2.585 ;
      RECT 36.44 2.575 36.77 3.305 ;
      RECT 26.675 2.575 27.005 3.305 ;
      RECT 22.555 2.415 22.885 3.145 ;
      RECT 21.555 1.855 21.885 2.585 ;
      RECT 20.115 2.575 20.445 3.305 ;
      RECT 10.35 2.575 10.68 3.305 ;
      RECT 6.23 2.415 6.56 3.145 ;
      RECT 5.23 1.855 5.56 2.585 ;
      RECT 3.79 2.575 4.12 3.305 ;
    LAYER via2 ;
      RECT 77.315 2.315 77.515 2.515 ;
      RECT 75.715 3.04 75.915 3.24 ;
      RECT 75.49 7.14 75.69 7.34 ;
      RECT 74.155 2.48 74.355 2.68 ;
      RECT 73.775 3.6 73.975 3.8 ;
      RECT 73.275 2.48 73.475 2.68 ;
      RECT 72.315 2.48 72.515 2.68 ;
      RECT 71.595 2.48 71.795 2.68 ;
      RECT 70.595 1.92 70.795 2.12 ;
      RECT 69.155 3.04 69.355 3.24 ;
      RECT 60.99 2.315 61.19 2.515 ;
      RECT 59.39 3.04 59.59 3.24 ;
      RECT 59.165 7.14 59.365 7.34 ;
      RECT 57.83 2.48 58.03 2.68 ;
      RECT 57.45 3.6 57.65 3.8 ;
      RECT 56.95 2.48 57.15 2.68 ;
      RECT 55.99 2.48 56.19 2.68 ;
      RECT 55.27 2.48 55.47 2.68 ;
      RECT 54.27 1.92 54.47 2.12 ;
      RECT 52.83 3.04 53.03 3.24 ;
      RECT 44.665 2.315 44.865 2.515 ;
      RECT 43.065 3.04 43.265 3.24 ;
      RECT 42.84 7.14 43.04 7.34 ;
      RECT 41.505 2.48 41.705 2.68 ;
      RECT 41.125 3.6 41.325 3.8 ;
      RECT 40.625 2.48 40.825 2.68 ;
      RECT 39.665 2.48 39.865 2.68 ;
      RECT 38.945 2.48 39.145 2.68 ;
      RECT 37.945 1.92 38.145 2.12 ;
      RECT 36.505 3.04 36.705 3.24 ;
      RECT 28.34 2.315 28.54 2.515 ;
      RECT 26.74 3.04 26.94 3.24 ;
      RECT 26.515 7.14 26.715 7.34 ;
      RECT 25.18 2.48 25.38 2.68 ;
      RECT 24.8 3.6 25 3.8 ;
      RECT 24.3 2.48 24.5 2.68 ;
      RECT 23.34 2.48 23.54 2.68 ;
      RECT 22.62 2.48 22.82 2.68 ;
      RECT 21.62 1.92 21.82 2.12 ;
      RECT 20.18 3.04 20.38 3.24 ;
      RECT 12.015 2.315 12.215 2.515 ;
      RECT 10.415 3.04 10.615 3.24 ;
      RECT 10.19 7.14 10.39 7.34 ;
      RECT 8.855 2.48 9.055 2.68 ;
      RECT 8.475 3.6 8.675 3.8 ;
      RECT 7.975 2.48 8.175 2.68 ;
      RECT 7.015 2.48 7.215 2.68 ;
      RECT 6.295 2.48 6.495 2.68 ;
      RECT 5.295 1.92 5.495 2.12 ;
      RECT 3.855 3.04 4.055 3.24 ;
    LAYER met2 ;
      RECT 1.23 8.4 84.055 8.57 ;
      RECT 83.885 7.275 84.055 8.57 ;
      RECT 1.23 6.255 1.4 8.57 ;
      RECT 83.855 7.275 84.205 7.625 ;
      RECT 1.17 6.255 1.46 6.605 ;
      RECT 80.695 6.22 81.015 6.545 ;
      RECT 80.725 5.695 80.895 6.545 ;
      RECT 80.725 5.695 80.9 6.045 ;
      RECT 80.725 5.695 81.7 5.87 ;
      RECT 81.525 1.965 81.7 5.87 ;
      RECT 81.47 1.965 81.82 2.315 ;
      RECT 81.495 6.655 81.82 6.98 ;
      RECT 80.38 6.745 81.82 6.915 ;
      RECT 80.38 2.395 80.54 6.915 ;
      RECT 80.695 2.365 81.015 2.685 ;
      RECT 80.38 2.395 81.015 2.565 ;
      RECT 70.555 1.835 70.835 2.205 ;
      RECT 70.59 1.29 70.76 2.205 ;
      RECT 79.165 1.29 79.335 1.815 ;
      RECT 79.075 1.46 79.415 1.81 ;
      RECT 70.59 1.29 79.335 1.46 ;
      RECT 75.795 2.395 76.075 2.765 ;
      RECT 74.725 2.42 74.985 2.74 ;
      RECT 77.275 2.23 77.555 2.6 ;
      RECT 77.885 2.14 78.145 2.46 ;
      RECT 74.785 1.58 74.925 2.74 ;
      RECT 75.865 1.58 76.005 2.765 ;
      RECT 76.985 2.23 78.145 2.37 ;
      RECT 76.985 1.58 77.125 2.37 ;
      RECT 74.785 1.58 77.125 1.72 ;
      RECT 74.815 3.72 76.99 3.885 ;
      RECT 76.845 2.6 76.99 3.885 ;
      RECT 73.735 3.515 74.015 3.885 ;
      RECT 73.735 3.63 74.955 3.77 ;
      RECT 76.565 2.6 76.99 2.74 ;
      RECT 76.565 2.42 76.825 2.74 ;
      RECT 69.905 4 73.565 4.14 ;
      RECT 73.425 3.185 73.565 4.14 ;
      RECT 69.905 3.07 70.045 4.14 ;
      RECT 76.445 3.26 76.705 3.58 ;
      RECT 73.425 3.185 75.955 3.325 ;
      RECT 75.675 2.955 75.955 3.325 ;
      RECT 69.905 3.07 70.355 3.325 ;
      RECT 70.075 2.955 70.355 3.325 ;
      RECT 76.445 3.07 76.645 3.58 ;
      RECT 75.675 3.07 76.645 3.21 ;
      RECT 76.245 1.86 76.385 3.21 ;
      RECT 76.185 1.86 76.445 2.18 ;
      RECT 67.505 6.655 67.855 7.005 ;
      RECT 76.06 6.61 76.41 6.96 ;
      RECT 67.505 6.685 76.41 6.885 ;
      RECT 70.085 2.42 70.345 2.74 ;
      RECT 70.085 2.51 71.125 2.65 ;
      RECT 70.985 1.72 71.125 2.65 ;
      RECT 73.745 1.86 74.005 2.18 ;
      RECT 70.985 1.72 73.945 1.86 ;
      RECT 73.125 2.7 73.385 3.02 ;
      RECT 73.125 2.7 73.445 2.93 ;
      RECT 73.235 2.395 73.515 2.765 ;
      RECT 72.825 3.26 73.145 3.58 ;
      RECT 72.825 2.14 72.965 3.58 ;
      RECT 72.765 2.14 73.025 2.46 ;
      RECT 70.325 3.54 70.585 3.86 ;
      RECT 70.325 3.63 72.005 3.77 ;
      RECT 71.865 3.35 72.005 3.77 ;
      RECT 71.865 3.35 72.305 3.58 ;
      RECT 72.045 3.26 72.305 3.58 ;
      RECT 71.365 2.42 71.765 2.93 ;
      RECT 71.555 2.395 71.835 2.765 ;
      RECT 71.305 2.42 71.835 2.74 ;
      RECT 64.37 6.22 64.69 6.545 ;
      RECT 64.4 5.695 64.57 6.545 ;
      RECT 64.4 5.695 64.575 6.045 ;
      RECT 64.4 5.695 65.375 5.87 ;
      RECT 65.2 1.965 65.375 5.87 ;
      RECT 65.145 1.965 65.495 2.315 ;
      RECT 65.17 6.655 65.495 6.98 ;
      RECT 64.055 6.745 65.495 6.915 ;
      RECT 64.055 2.395 64.215 6.915 ;
      RECT 64.37 2.365 64.69 2.685 ;
      RECT 64.055 2.395 64.69 2.565 ;
      RECT 54.23 1.835 54.51 2.205 ;
      RECT 54.265 1.29 54.435 2.205 ;
      RECT 62.84 1.29 63.01 1.815 ;
      RECT 62.75 1.46 63.09 1.81 ;
      RECT 54.265 1.29 63.01 1.46 ;
      RECT 59.47 2.395 59.75 2.765 ;
      RECT 58.4 2.42 58.66 2.74 ;
      RECT 60.95 2.23 61.23 2.6 ;
      RECT 61.56 2.14 61.82 2.46 ;
      RECT 58.46 1.58 58.6 2.74 ;
      RECT 59.54 1.58 59.68 2.765 ;
      RECT 60.66 2.23 61.82 2.37 ;
      RECT 60.66 1.58 60.8 2.37 ;
      RECT 58.46 1.58 60.8 1.72 ;
      RECT 58.49 3.72 60.665 3.885 ;
      RECT 60.52 2.6 60.665 3.885 ;
      RECT 57.41 3.515 57.69 3.885 ;
      RECT 57.41 3.63 58.63 3.77 ;
      RECT 60.24 2.6 60.665 2.74 ;
      RECT 60.24 2.42 60.5 2.74 ;
      RECT 53.58 4 57.24 4.14 ;
      RECT 57.1 3.185 57.24 4.14 ;
      RECT 53.58 3.07 53.72 4.14 ;
      RECT 60.12 3.26 60.38 3.58 ;
      RECT 57.1 3.185 59.63 3.325 ;
      RECT 59.35 2.955 59.63 3.325 ;
      RECT 53.58 3.07 54.03 3.325 ;
      RECT 53.75 2.955 54.03 3.325 ;
      RECT 60.12 3.07 60.32 3.58 ;
      RECT 59.35 3.07 60.32 3.21 ;
      RECT 59.92 1.86 60.06 3.21 ;
      RECT 59.86 1.86 60.12 2.18 ;
      RECT 51.18 6.655 51.53 7.005 ;
      RECT 59.73 6.61 60.08 6.96 ;
      RECT 51.18 6.685 60.08 6.885 ;
      RECT 53.76 2.42 54.02 2.74 ;
      RECT 53.76 2.51 54.8 2.65 ;
      RECT 54.66 1.72 54.8 2.65 ;
      RECT 57.42 1.86 57.68 2.18 ;
      RECT 54.66 1.72 57.62 1.86 ;
      RECT 56.8 2.7 57.06 3.02 ;
      RECT 56.8 2.7 57.12 2.93 ;
      RECT 56.91 2.395 57.19 2.765 ;
      RECT 56.5 3.26 56.82 3.58 ;
      RECT 56.5 2.14 56.64 3.58 ;
      RECT 56.44 2.14 56.7 2.46 ;
      RECT 54 3.54 54.26 3.86 ;
      RECT 54 3.63 55.68 3.77 ;
      RECT 55.54 3.35 55.68 3.77 ;
      RECT 55.54 3.35 55.98 3.58 ;
      RECT 55.72 3.26 55.98 3.58 ;
      RECT 55.04 2.42 55.44 2.93 ;
      RECT 55.23 2.395 55.51 2.765 ;
      RECT 54.98 2.42 55.51 2.74 ;
      RECT 48.045 6.22 48.365 6.545 ;
      RECT 48.075 5.695 48.245 6.545 ;
      RECT 48.075 5.695 48.25 6.045 ;
      RECT 48.075 5.695 49.05 5.87 ;
      RECT 48.875 1.965 49.05 5.87 ;
      RECT 48.82 1.965 49.17 2.315 ;
      RECT 48.845 6.655 49.17 6.98 ;
      RECT 47.73 6.745 49.17 6.915 ;
      RECT 47.73 2.395 47.89 6.915 ;
      RECT 48.045 2.365 48.365 2.685 ;
      RECT 47.73 2.395 48.365 2.565 ;
      RECT 37.905 1.835 38.185 2.205 ;
      RECT 37.94 1.29 38.11 2.205 ;
      RECT 46.515 1.29 46.685 1.815 ;
      RECT 46.425 1.46 46.765 1.81 ;
      RECT 37.94 1.29 46.685 1.46 ;
      RECT 43.145 2.395 43.425 2.765 ;
      RECT 42.075 2.42 42.335 2.74 ;
      RECT 44.625 2.23 44.905 2.6 ;
      RECT 45.235 2.14 45.495 2.46 ;
      RECT 42.135 1.58 42.275 2.74 ;
      RECT 43.215 1.58 43.355 2.765 ;
      RECT 44.335 2.23 45.495 2.37 ;
      RECT 44.335 1.58 44.475 2.37 ;
      RECT 42.135 1.58 44.475 1.72 ;
      RECT 42.165 3.72 44.34 3.885 ;
      RECT 44.195 2.6 44.34 3.885 ;
      RECT 41.085 3.515 41.365 3.885 ;
      RECT 41.085 3.63 42.305 3.77 ;
      RECT 43.915 2.6 44.34 2.74 ;
      RECT 43.915 2.42 44.175 2.74 ;
      RECT 37.255 4 40.915 4.14 ;
      RECT 40.775 3.185 40.915 4.14 ;
      RECT 37.255 3.07 37.395 4.14 ;
      RECT 43.795 3.26 44.055 3.58 ;
      RECT 40.775 3.185 43.305 3.325 ;
      RECT 43.025 2.955 43.305 3.325 ;
      RECT 37.255 3.07 37.705 3.325 ;
      RECT 37.425 2.955 37.705 3.325 ;
      RECT 43.795 3.07 43.995 3.58 ;
      RECT 43.025 3.07 43.995 3.21 ;
      RECT 43.595 1.86 43.735 3.21 ;
      RECT 43.535 1.86 43.795 2.18 ;
      RECT 34.9 6.66 35.25 7.01 ;
      RECT 43.405 6.615 43.755 6.965 ;
      RECT 34.9 6.69 43.755 6.89 ;
      RECT 37.435 2.42 37.695 2.74 ;
      RECT 37.435 2.51 38.475 2.65 ;
      RECT 38.335 1.72 38.475 2.65 ;
      RECT 41.095 1.86 41.355 2.18 ;
      RECT 38.335 1.72 41.295 1.86 ;
      RECT 40.475 2.7 40.735 3.02 ;
      RECT 40.475 2.7 40.795 2.93 ;
      RECT 40.585 2.395 40.865 2.765 ;
      RECT 40.175 3.26 40.495 3.58 ;
      RECT 40.175 2.14 40.315 3.58 ;
      RECT 40.115 2.14 40.375 2.46 ;
      RECT 37.675 3.54 37.935 3.86 ;
      RECT 37.675 3.63 39.355 3.77 ;
      RECT 39.215 3.35 39.355 3.77 ;
      RECT 39.215 3.35 39.655 3.58 ;
      RECT 39.395 3.26 39.655 3.58 ;
      RECT 38.715 2.42 39.115 2.93 ;
      RECT 38.905 2.395 39.185 2.765 ;
      RECT 38.655 2.42 39.185 2.74 ;
      RECT 31.72 6.22 32.04 6.545 ;
      RECT 31.75 5.695 31.92 6.545 ;
      RECT 31.75 5.695 31.925 6.045 ;
      RECT 31.75 5.695 32.725 5.87 ;
      RECT 32.55 1.965 32.725 5.87 ;
      RECT 32.495 1.965 32.845 2.315 ;
      RECT 32.52 6.655 32.845 6.98 ;
      RECT 31.405 6.745 32.845 6.915 ;
      RECT 31.405 2.395 31.565 6.915 ;
      RECT 31.72 2.365 32.04 2.685 ;
      RECT 31.405 2.395 32.04 2.565 ;
      RECT 21.58 1.835 21.86 2.205 ;
      RECT 21.615 1.29 21.785 2.205 ;
      RECT 30.19 1.29 30.36 1.815 ;
      RECT 30.1 1.46 30.44 1.81 ;
      RECT 21.615 1.29 30.36 1.46 ;
      RECT 26.82 2.395 27.1 2.765 ;
      RECT 25.75 2.42 26.01 2.74 ;
      RECT 28.3 2.23 28.58 2.6 ;
      RECT 28.91 2.14 29.17 2.46 ;
      RECT 25.81 1.58 25.95 2.74 ;
      RECT 26.89 1.58 27.03 2.765 ;
      RECT 28.01 2.23 29.17 2.37 ;
      RECT 28.01 1.58 28.15 2.37 ;
      RECT 25.81 1.58 28.15 1.72 ;
      RECT 25.84 3.72 28.015 3.885 ;
      RECT 27.87 2.6 28.015 3.885 ;
      RECT 24.76 3.515 25.04 3.885 ;
      RECT 24.76 3.63 25.98 3.77 ;
      RECT 27.59 2.6 28.015 2.74 ;
      RECT 27.59 2.42 27.85 2.74 ;
      RECT 20.93 4 24.59 4.14 ;
      RECT 24.45 3.185 24.59 4.14 ;
      RECT 20.93 3.07 21.07 4.14 ;
      RECT 27.47 3.26 27.73 3.58 ;
      RECT 24.45 3.185 26.98 3.325 ;
      RECT 26.7 2.955 26.98 3.325 ;
      RECT 20.93 3.07 21.38 3.325 ;
      RECT 21.1 2.955 21.38 3.325 ;
      RECT 27.47 3.07 27.67 3.58 ;
      RECT 26.7 3.07 27.67 3.21 ;
      RECT 27.27 1.86 27.41 3.21 ;
      RECT 27.21 1.86 27.47 2.18 ;
      RECT 18.575 6.655 18.925 7.005 ;
      RECT 27.08 6.61 27.43 6.96 ;
      RECT 18.575 6.685 27.43 6.885 ;
      RECT 21.11 2.42 21.37 2.74 ;
      RECT 21.11 2.51 22.15 2.65 ;
      RECT 22.01 1.72 22.15 2.65 ;
      RECT 24.77 1.86 25.03 2.18 ;
      RECT 22.01 1.72 24.97 1.86 ;
      RECT 24.15 2.7 24.41 3.02 ;
      RECT 24.15 2.7 24.47 2.93 ;
      RECT 24.26 2.395 24.54 2.765 ;
      RECT 23.85 3.26 24.17 3.58 ;
      RECT 23.85 2.14 23.99 3.58 ;
      RECT 23.79 2.14 24.05 2.46 ;
      RECT 21.35 3.54 21.61 3.86 ;
      RECT 21.35 3.63 23.03 3.77 ;
      RECT 22.89 3.35 23.03 3.77 ;
      RECT 22.89 3.35 23.33 3.58 ;
      RECT 23.07 3.26 23.33 3.58 ;
      RECT 22.39 2.42 22.79 2.93 ;
      RECT 22.58 2.395 22.86 2.765 ;
      RECT 22.33 2.42 22.86 2.74 ;
      RECT 15.395 6.22 15.715 6.545 ;
      RECT 15.425 5.695 15.595 6.545 ;
      RECT 15.425 5.695 15.6 6.045 ;
      RECT 15.425 5.695 16.4 5.87 ;
      RECT 16.225 1.965 16.4 5.87 ;
      RECT 16.17 1.965 16.52 2.315 ;
      RECT 16.195 6.655 16.52 6.98 ;
      RECT 15.08 6.745 16.52 6.915 ;
      RECT 15.08 2.395 15.24 6.915 ;
      RECT 15.395 2.365 15.715 2.685 ;
      RECT 15.08 2.395 15.715 2.565 ;
      RECT 5.255 1.835 5.535 2.205 ;
      RECT 5.29 1.29 5.46 2.205 ;
      RECT 13.865 1.29 14.035 1.815 ;
      RECT 13.775 1.46 14.115 1.81 ;
      RECT 5.29 1.29 14.035 1.46 ;
      RECT 10.495 2.395 10.775 2.765 ;
      RECT 9.425 2.42 9.685 2.74 ;
      RECT 11.975 2.23 12.255 2.6 ;
      RECT 12.585 2.14 12.845 2.46 ;
      RECT 9.485 1.58 9.625 2.74 ;
      RECT 10.565 1.58 10.705 2.765 ;
      RECT 11.685 2.23 12.845 2.37 ;
      RECT 11.685 1.58 11.825 2.37 ;
      RECT 9.485 1.58 11.825 1.72 ;
      RECT 1.545 6.995 1.835 7.345 ;
      RECT 1.545 7.05 2.83 7.225 ;
      RECT 2.655 6.685 2.83 7.225 ;
      RECT 11.59 6.605 11.94 6.955 ;
      RECT 2.655 6.685 11.94 6.86 ;
      RECT 9.515 3.72 11.69 3.885 ;
      RECT 11.545 2.6 11.69 3.885 ;
      RECT 8.435 3.515 8.715 3.885 ;
      RECT 8.435 3.63 9.655 3.77 ;
      RECT 11.265 2.6 11.69 2.74 ;
      RECT 11.265 2.42 11.525 2.74 ;
      RECT 4.605 4 8.265 4.14 ;
      RECT 8.125 3.185 8.265 4.14 ;
      RECT 4.605 3.07 4.745 4.14 ;
      RECT 11.145 3.26 11.405 3.58 ;
      RECT 8.125 3.185 10.655 3.325 ;
      RECT 10.375 2.955 10.655 3.325 ;
      RECT 4.605 3.07 5.055 3.325 ;
      RECT 4.775 2.955 5.055 3.325 ;
      RECT 11.145 3.07 11.345 3.58 ;
      RECT 10.375 3.07 11.345 3.21 ;
      RECT 10.945 1.86 11.085 3.21 ;
      RECT 10.885 1.86 11.145 2.18 ;
      RECT 4.785 2.42 5.045 2.74 ;
      RECT 4.785 2.51 5.825 2.65 ;
      RECT 5.685 1.72 5.825 2.65 ;
      RECT 8.445 1.86 8.705 2.18 ;
      RECT 5.685 1.72 8.645 1.86 ;
      RECT 7.825 2.7 8.085 3.02 ;
      RECT 7.825 2.7 8.145 2.93 ;
      RECT 7.935 2.395 8.215 2.765 ;
      RECT 7.525 3.26 7.845 3.58 ;
      RECT 7.525 2.14 7.665 3.58 ;
      RECT 7.465 2.14 7.725 2.46 ;
      RECT 5.025 3.54 5.285 3.86 ;
      RECT 5.025 3.63 6.705 3.77 ;
      RECT 6.565 3.35 6.705 3.77 ;
      RECT 6.565 3.35 7.005 3.58 ;
      RECT 6.745 3.26 7.005 3.58 ;
      RECT 6.065 2.42 6.465 2.93 ;
      RECT 6.255 2.395 6.535 2.765 ;
      RECT 6.005 2.42 6.535 2.74 ;
      RECT 75.405 7.055 75.775 7.425 ;
      RECT 74.115 2.395 74.395 2.765 ;
      RECT 72.275 2.395 72.555 2.765 ;
      RECT 69.115 2.955 69.395 3.325 ;
      RECT 59.08 7.055 59.45 7.425 ;
      RECT 57.79 2.395 58.07 2.765 ;
      RECT 55.95 2.395 56.23 2.765 ;
      RECT 52.79 2.955 53.07 3.325 ;
      RECT 42.755 7.055 43.125 7.425 ;
      RECT 41.465 2.395 41.745 2.765 ;
      RECT 39.625 2.395 39.905 2.765 ;
      RECT 36.465 2.955 36.745 3.325 ;
      RECT 26.43 7.055 26.8 7.425 ;
      RECT 25.14 2.395 25.42 2.765 ;
      RECT 23.3 2.395 23.58 2.765 ;
      RECT 20.14 2.955 20.42 3.325 ;
      RECT 10.105 7.055 10.475 7.425 ;
      RECT 8.815 2.395 9.095 2.765 ;
      RECT 6.975 2.395 7.255 2.765 ;
      RECT 3.815 2.955 4.095 3.325 ;
    LAYER via1 ;
      RECT 83.955 7.375 84.105 7.525 ;
      RECT 81.585 6.74 81.735 6.89 ;
      RECT 81.57 2.065 81.72 2.215 ;
      RECT 80.78 2.45 80.93 2.6 ;
      RECT 80.78 6.325 80.93 6.475 ;
      RECT 79.175 1.56 79.325 1.71 ;
      RECT 77.94 2.225 78.09 2.375 ;
      RECT 76.62 2.505 76.77 2.655 ;
      RECT 76.5 3.345 76.65 3.495 ;
      RECT 76.24 1.945 76.39 2.095 ;
      RECT 76.16 6.71 76.31 6.86 ;
      RECT 75.515 7.165 75.665 7.315 ;
      RECT 74.78 2.505 74.93 2.655 ;
      RECT 74.18 2.505 74.33 2.655 ;
      RECT 73.8 1.945 73.95 2.095 ;
      RECT 73.18 2.785 73.33 2.935 ;
      RECT 72.94 3.345 73.09 3.495 ;
      RECT 72.82 2.225 72.97 2.375 ;
      RECT 72.34 2.505 72.49 2.655 ;
      RECT 72.1 3.345 72.25 3.495 ;
      RECT 71.36 2.505 71.51 2.655 ;
      RECT 70.62 1.945 70.77 2.095 ;
      RECT 70.38 3.625 70.53 3.775 ;
      RECT 70.14 2.505 70.29 2.655 ;
      RECT 70.14 3.065 70.29 3.215 ;
      RECT 69.18 3.065 69.33 3.215 ;
      RECT 67.605 6.755 67.755 6.905 ;
      RECT 65.26 6.74 65.41 6.89 ;
      RECT 65.245 2.065 65.395 2.215 ;
      RECT 64.455 2.45 64.605 2.6 ;
      RECT 64.455 6.325 64.605 6.475 ;
      RECT 62.85 1.56 63 1.71 ;
      RECT 61.615 2.225 61.765 2.375 ;
      RECT 60.295 2.505 60.445 2.655 ;
      RECT 60.175 3.345 60.325 3.495 ;
      RECT 59.915 1.945 60.065 2.095 ;
      RECT 59.83 6.71 59.98 6.86 ;
      RECT 59.19 7.165 59.34 7.315 ;
      RECT 58.455 2.505 58.605 2.655 ;
      RECT 57.855 2.505 58.005 2.655 ;
      RECT 57.475 1.945 57.625 2.095 ;
      RECT 56.855 2.785 57.005 2.935 ;
      RECT 56.615 3.345 56.765 3.495 ;
      RECT 56.495 2.225 56.645 2.375 ;
      RECT 56.015 2.505 56.165 2.655 ;
      RECT 55.775 3.345 55.925 3.495 ;
      RECT 55.035 2.505 55.185 2.655 ;
      RECT 54.295 1.945 54.445 2.095 ;
      RECT 54.055 3.625 54.205 3.775 ;
      RECT 53.815 2.505 53.965 2.655 ;
      RECT 53.815 3.065 53.965 3.215 ;
      RECT 52.855 3.065 53.005 3.215 ;
      RECT 51.28 6.755 51.43 6.905 ;
      RECT 48.935 6.74 49.085 6.89 ;
      RECT 48.92 2.065 49.07 2.215 ;
      RECT 48.13 2.45 48.28 2.6 ;
      RECT 48.13 6.325 48.28 6.475 ;
      RECT 46.525 1.56 46.675 1.71 ;
      RECT 45.29 2.225 45.44 2.375 ;
      RECT 43.97 2.505 44.12 2.655 ;
      RECT 43.85 3.345 44 3.495 ;
      RECT 43.59 1.945 43.74 2.095 ;
      RECT 43.505 6.715 43.655 6.865 ;
      RECT 42.865 7.165 43.015 7.315 ;
      RECT 42.13 2.505 42.28 2.655 ;
      RECT 41.53 2.505 41.68 2.655 ;
      RECT 41.15 1.945 41.3 2.095 ;
      RECT 40.53 2.785 40.68 2.935 ;
      RECT 40.29 3.345 40.44 3.495 ;
      RECT 40.17 2.225 40.32 2.375 ;
      RECT 39.69 2.505 39.84 2.655 ;
      RECT 39.45 3.345 39.6 3.495 ;
      RECT 38.71 2.505 38.86 2.655 ;
      RECT 37.97 1.945 38.12 2.095 ;
      RECT 37.73 3.625 37.88 3.775 ;
      RECT 37.49 2.505 37.64 2.655 ;
      RECT 37.49 3.065 37.64 3.215 ;
      RECT 36.53 3.065 36.68 3.215 ;
      RECT 35 6.76 35.15 6.91 ;
      RECT 32.61 6.74 32.76 6.89 ;
      RECT 32.595 2.065 32.745 2.215 ;
      RECT 31.805 2.45 31.955 2.6 ;
      RECT 31.805 6.325 31.955 6.475 ;
      RECT 30.2 1.56 30.35 1.71 ;
      RECT 28.965 2.225 29.115 2.375 ;
      RECT 27.645 2.505 27.795 2.655 ;
      RECT 27.525 3.345 27.675 3.495 ;
      RECT 27.265 1.945 27.415 2.095 ;
      RECT 27.18 6.71 27.33 6.86 ;
      RECT 26.54 7.165 26.69 7.315 ;
      RECT 25.805 2.505 25.955 2.655 ;
      RECT 25.205 2.505 25.355 2.655 ;
      RECT 24.825 1.945 24.975 2.095 ;
      RECT 24.205 2.785 24.355 2.935 ;
      RECT 23.965 3.345 24.115 3.495 ;
      RECT 23.845 2.225 23.995 2.375 ;
      RECT 23.365 2.505 23.515 2.655 ;
      RECT 23.125 3.345 23.275 3.495 ;
      RECT 22.385 2.505 22.535 2.655 ;
      RECT 21.645 1.945 21.795 2.095 ;
      RECT 21.405 3.625 21.555 3.775 ;
      RECT 21.165 2.505 21.315 2.655 ;
      RECT 21.165 3.065 21.315 3.215 ;
      RECT 20.205 3.065 20.355 3.215 ;
      RECT 18.675 6.755 18.825 6.905 ;
      RECT 16.285 6.74 16.435 6.89 ;
      RECT 16.27 2.065 16.42 2.215 ;
      RECT 15.48 2.45 15.63 2.6 ;
      RECT 15.48 6.325 15.63 6.475 ;
      RECT 13.875 1.56 14.025 1.71 ;
      RECT 12.64 2.225 12.79 2.375 ;
      RECT 11.69 6.705 11.84 6.855 ;
      RECT 11.32 2.505 11.47 2.655 ;
      RECT 11.2 3.345 11.35 3.495 ;
      RECT 10.94 1.945 11.09 2.095 ;
      RECT 10.215 7.165 10.365 7.315 ;
      RECT 9.48 2.505 9.63 2.655 ;
      RECT 8.88 2.505 9.03 2.655 ;
      RECT 8.5 1.945 8.65 2.095 ;
      RECT 7.88 2.785 8.03 2.935 ;
      RECT 7.64 3.345 7.79 3.495 ;
      RECT 7.52 2.225 7.67 2.375 ;
      RECT 7.04 2.505 7.19 2.655 ;
      RECT 6.8 3.345 6.95 3.495 ;
      RECT 6.06 2.505 6.21 2.655 ;
      RECT 5.32 1.945 5.47 2.095 ;
      RECT 5.08 3.625 5.23 3.775 ;
      RECT 4.84 2.505 4.99 2.655 ;
      RECT 4.84 3.065 4.99 3.215 ;
      RECT 3.88 3.065 4.03 3.215 ;
      RECT 1.615 7.095 1.765 7.245 ;
      RECT 1.24 6.355 1.39 6.505 ;
    LAYER met1 ;
      RECT 83.82 7.77 84.11 8 ;
      RECT 83.88 6.29 84.05 8 ;
      RECT 83.855 7.275 84.205 7.625 ;
      RECT 83.82 6.29 84.11 6.52 ;
      RECT 83.415 2.395 83.52 2.965 ;
      RECT 83.415 2.73 83.74 2.96 ;
      RECT 83.415 2.76 83.91 2.93 ;
      RECT 83.415 2.395 83.605 2.96 ;
      RECT 82.83 2.36 83.12 2.59 ;
      RECT 82.83 2.395 83.605 2.565 ;
      RECT 82.89 0.88 83.06 2.59 ;
      RECT 82.83 0.88 83.12 1.11 ;
      RECT 82.83 7.77 83.12 8 ;
      RECT 82.89 6.29 83.06 8 ;
      RECT 82.83 6.29 83.12 6.52 ;
      RECT 82.83 6.325 83.685 6.485 ;
      RECT 83.515 5.92 83.685 6.485 ;
      RECT 82.83 6.32 83.225 6.485 ;
      RECT 83.45 5.92 83.74 6.15 ;
      RECT 83.45 5.95 83.91 6.12 ;
      RECT 82.46 2.73 82.75 2.96 ;
      RECT 82.46 2.76 82.92 2.93 ;
      RECT 82.525 1.655 82.69 2.96 ;
      RECT 81.04 1.625 81.33 1.855 ;
      RECT 81.04 1.655 82.69 1.825 ;
      RECT 81.1 0.885 81.27 1.855 ;
      RECT 81.04 0.885 81.33 1.115 ;
      RECT 81.04 7.765 81.33 7.995 ;
      RECT 81.1 7.025 81.27 7.995 ;
      RECT 81.1 7.12 82.69 7.29 ;
      RECT 82.52 5.92 82.69 7.29 ;
      RECT 81.04 7.025 81.33 7.255 ;
      RECT 82.46 5.92 82.75 6.15 ;
      RECT 82.46 5.95 82.92 6.12 ;
      RECT 81.47 1.965 81.82 2.315 ;
      RECT 79.165 2.025 81.82 2.195 ;
      RECT 79.165 1.46 79.335 2.195 ;
      RECT 79.075 1.46 79.415 1.81 ;
      RECT 81.495 6.655 81.82 6.98 ;
      RECT 76.06 6.61 76.41 6.96 ;
      RECT 81.47 6.655 81.82 6.885 ;
      RECT 75.855 6.655 76.41 6.885 ;
      RECT 75.685 6.685 81.82 6.855 ;
      RECT 80.695 2.365 81.015 2.685 ;
      RECT 80.665 2.365 81.015 2.595 ;
      RECT 80.495 2.395 81.015 2.565 ;
      RECT 80.695 6.255 81.015 6.545 ;
      RECT 80.665 6.285 81.015 6.515 ;
      RECT 80.495 6.315 81.015 6.485 ;
      RECT 77.15 2.465 77.44 2.695 ;
      RECT 77.15 2.465 77.605 2.65 ;
      RECT 77.465 2.37 78.085 2.51 ;
      RECT 77.855 2.17 78.175 2.43 ;
      RECT 76.535 2.45 76.855 2.71 ;
      RECT 76.535 2.45 77 2.695 ;
      RECT 76.86 2.07 77 2.695 ;
      RECT 76.86 2.07 77.125 2.21 ;
      RECT 77.39 1.905 77.68 2.135 ;
      RECT 76.985 1.95 77.68 2.09 ;
      RECT 76.43 3.29 76.72 3.815 ;
      RECT 76.415 3.29 76.735 3.55 ;
      RECT 76.155 1.89 76.475 2.15 ;
      RECT 76.155 1.905 76.72 2.135 ;
      RECT 75.43 3.585 75.72 3.815 ;
      RECT 75.625 2.23 75.765 3.77 ;
      RECT 75.67 2.185 75.96 2.415 ;
      RECT 75.265 2.23 75.96 2.37 ;
      RECT 75.265 2.07 75.405 2.37 ;
      RECT 73.805 2.07 75.405 2.21 ;
      RECT 73.715 1.89 74.035 2.15 ;
      RECT 73.715 1.905 74.28 2.15 ;
      RECT 75.425 7.765 75.715 7.995 ;
      RECT 75.485 7.025 75.655 7.995 ;
      RECT 75.405 7.075 75.775 7.425 ;
      RECT 75.405 7.055 75.715 7.425 ;
      RECT 75.425 7.025 75.715 7.425 ;
      RECT 72.825 2.93 75.405 3.07 ;
      RECT 75.19 2.745 75.48 2.975 ;
      RECT 72.75 2.745 73.415 2.975 ;
      RECT 73.095 2.73 73.415 3.07 ;
      RECT 74.095 2.45 74.415 2.71 ;
      RECT 74.095 2.465 74.52 2.695 ;
      RECT 72.735 2.17 73.055 2.43 ;
      RECT 73.23 2.185 73.52 2.415 ;
      RECT 72.735 2.23 73.52 2.37 ;
      RECT 72.855 3.29 73.175 3.55 ;
      RECT 72.015 3.29 72.335 3.55 ;
      RECT 72.855 3.305 73.28 3.535 ;
      RECT 72.015 3.35 73.28 3.49 ;
      RECT 71.55 3.025 71.84 3.255 ;
      RECT 71.625 1.95 71.765 3.255 ;
      RECT 71.275 2.45 71.765 2.71 ;
      RECT 71.03 2.465 71.765 2.695 ;
      RECT 72.03 1.905 72.32 2.135 ;
      RECT 71.625 1.95 72.32 2.09 ;
      RECT 70.79 3.305 71.08 3.535 ;
      RECT 70.79 3.305 71.245 3.49 ;
      RECT 71.105 2.93 71.245 3.49 ;
      RECT 70.745 2.93 71.245 3.07 ;
      RECT 70.745 1.95 70.885 3.07 ;
      RECT 70.535 1.89 70.855 2.15 ;
      RECT 70.295 3.57 70.615 3.83 ;
      RECT 69.59 3.585 69.88 3.815 ;
      RECT 69.59 3.63 70.615 3.77 ;
      RECT 69.665 3.58 69.925 3.77 ;
      RECT 70.055 2.45 70.375 2.71 ;
      RECT 70.055 2.465 70.6 2.695 ;
      RECT 70.055 3.01 70.375 3.27 ;
      RECT 70.055 3.025 70.6 3.255 ;
      RECT 69.095 3.01 69.415 3.27 ;
      RECT 69.185 1.95 69.325 3.27 ;
      RECT 69.59 1.905 69.88 2.135 ;
      RECT 69.185 1.95 69.88 2.09 ;
      RECT 67.495 7.77 67.785 8 ;
      RECT 67.555 6.29 67.725 8 ;
      RECT 67.505 6.655 67.855 7.005 ;
      RECT 67.495 6.29 67.785 6.52 ;
      RECT 67.09 2.395 67.195 2.965 ;
      RECT 67.09 2.73 67.415 2.96 ;
      RECT 67.09 2.76 67.585 2.93 ;
      RECT 67.09 2.395 67.28 2.96 ;
      RECT 66.505 2.36 66.795 2.59 ;
      RECT 66.505 2.395 67.28 2.565 ;
      RECT 66.565 0.88 66.735 2.59 ;
      RECT 66.505 0.88 66.795 1.11 ;
      RECT 66.505 7.77 66.795 8 ;
      RECT 66.565 6.29 66.735 8 ;
      RECT 66.505 6.29 66.795 6.52 ;
      RECT 66.505 6.325 67.36 6.485 ;
      RECT 67.19 5.92 67.36 6.485 ;
      RECT 66.505 6.32 66.9 6.485 ;
      RECT 67.125 5.92 67.415 6.15 ;
      RECT 67.125 5.95 67.585 6.12 ;
      RECT 66.135 2.73 66.425 2.96 ;
      RECT 66.135 2.76 66.595 2.93 ;
      RECT 66.2 1.655 66.365 2.96 ;
      RECT 64.715 1.625 65.005 1.855 ;
      RECT 64.715 1.655 66.365 1.825 ;
      RECT 64.775 0.885 64.945 1.855 ;
      RECT 64.715 0.885 65.005 1.115 ;
      RECT 64.715 7.765 65.005 7.995 ;
      RECT 64.775 7.025 64.945 7.995 ;
      RECT 64.775 7.12 66.365 7.29 ;
      RECT 66.195 5.92 66.365 7.29 ;
      RECT 64.715 7.025 65.005 7.255 ;
      RECT 66.135 5.92 66.425 6.15 ;
      RECT 66.135 5.95 66.595 6.12 ;
      RECT 65.145 1.965 65.495 2.315 ;
      RECT 62.84 2.025 65.495 2.195 ;
      RECT 62.84 1.46 63.01 2.195 ;
      RECT 62.75 1.46 63.09 1.81 ;
      RECT 65.17 6.655 65.495 6.98 ;
      RECT 59.73 6.61 60.08 6.96 ;
      RECT 65.145 6.655 65.495 6.885 ;
      RECT 59.53 6.655 60.08 6.885 ;
      RECT 59.36 6.685 65.495 6.855 ;
      RECT 64.37 2.365 64.69 2.685 ;
      RECT 64.34 2.365 64.69 2.595 ;
      RECT 64.17 2.395 64.69 2.565 ;
      RECT 64.37 6.255 64.69 6.545 ;
      RECT 64.34 6.285 64.69 6.515 ;
      RECT 64.17 6.315 64.69 6.485 ;
      RECT 60.825 2.465 61.115 2.695 ;
      RECT 60.825 2.465 61.28 2.65 ;
      RECT 61.14 2.37 61.76 2.51 ;
      RECT 61.53 2.17 61.85 2.43 ;
      RECT 60.21 2.45 60.53 2.71 ;
      RECT 60.21 2.45 60.675 2.695 ;
      RECT 60.535 2.07 60.675 2.695 ;
      RECT 60.535 2.07 60.8 2.21 ;
      RECT 61.065 1.905 61.355 2.135 ;
      RECT 60.66 1.95 61.355 2.09 ;
      RECT 60.105 3.29 60.395 3.815 ;
      RECT 60.09 3.29 60.41 3.55 ;
      RECT 59.83 1.89 60.15 2.15 ;
      RECT 59.83 1.905 60.395 2.135 ;
      RECT 59.105 3.585 59.395 3.815 ;
      RECT 59.3 2.23 59.44 3.77 ;
      RECT 59.345 2.185 59.635 2.415 ;
      RECT 58.94 2.23 59.635 2.37 ;
      RECT 58.94 2.07 59.08 2.37 ;
      RECT 57.48 2.07 59.08 2.21 ;
      RECT 57.39 1.89 57.71 2.15 ;
      RECT 57.39 1.905 57.955 2.15 ;
      RECT 59.1 7.765 59.39 7.995 ;
      RECT 59.16 7.025 59.33 7.995 ;
      RECT 59.08 7.075 59.45 7.425 ;
      RECT 59.08 7.055 59.39 7.425 ;
      RECT 59.1 7.025 59.39 7.425 ;
      RECT 56.5 2.93 59.08 3.07 ;
      RECT 58.865 2.745 59.155 2.975 ;
      RECT 56.425 2.745 57.09 2.975 ;
      RECT 56.77 2.73 57.09 3.07 ;
      RECT 57.77 2.45 58.09 2.71 ;
      RECT 57.77 2.465 58.195 2.695 ;
      RECT 56.41 2.17 56.73 2.43 ;
      RECT 56.905 2.185 57.195 2.415 ;
      RECT 56.41 2.23 57.195 2.37 ;
      RECT 56.53 3.29 56.85 3.55 ;
      RECT 55.69 3.29 56.01 3.55 ;
      RECT 56.53 3.305 56.955 3.535 ;
      RECT 55.69 3.35 56.955 3.49 ;
      RECT 55.225 3.025 55.515 3.255 ;
      RECT 55.3 1.95 55.44 3.255 ;
      RECT 54.95 2.45 55.44 2.71 ;
      RECT 54.705 2.465 55.44 2.695 ;
      RECT 55.705 1.905 55.995 2.135 ;
      RECT 55.3 1.95 55.995 2.09 ;
      RECT 54.465 3.305 54.755 3.535 ;
      RECT 54.465 3.305 54.92 3.49 ;
      RECT 54.78 2.93 54.92 3.49 ;
      RECT 54.42 2.93 54.92 3.07 ;
      RECT 54.42 1.95 54.56 3.07 ;
      RECT 54.21 1.89 54.53 2.15 ;
      RECT 53.97 3.57 54.29 3.83 ;
      RECT 53.265 3.585 53.555 3.815 ;
      RECT 53.265 3.63 54.29 3.77 ;
      RECT 53.34 3.58 53.6 3.77 ;
      RECT 53.73 2.45 54.05 2.71 ;
      RECT 53.73 2.465 54.275 2.695 ;
      RECT 53.73 3.01 54.05 3.27 ;
      RECT 53.73 3.025 54.275 3.255 ;
      RECT 52.77 3.01 53.09 3.27 ;
      RECT 52.86 1.95 53 3.27 ;
      RECT 53.265 1.905 53.555 2.135 ;
      RECT 52.86 1.95 53.555 2.09 ;
      RECT 51.17 7.77 51.46 8 ;
      RECT 51.23 6.29 51.4 8 ;
      RECT 51.18 6.655 51.53 7.005 ;
      RECT 51.17 6.29 51.46 6.52 ;
      RECT 50.765 2.395 50.87 2.965 ;
      RECT 50.765 2.73 51.09 2.96 ;
      RECT 50.765 2.76 51.26 2.93 ;
      RECT 50.765 2.395 50.955 2.96 ;
      RECT 50.18 2.36 50.47 2.59 ;
      RECT 50.18 2.395 50.955 2.565 ;
      RECT 50.24 0.88 50.41 2.59 ;
      RECT 50.18 0.88 50.47 1.11 ;
      RECT 50.18 7.77 50.47 8 ;
      RECT 50.24 6.29 50.41 8 ;
      RECT 50.18 6.29 50.47 6.52 ;
      RECT 50.18 6.325 51.035 6.485 ;
      RECT 50.865 5.92 51.035 6.485 ;
      RECT 50.18 6.32 50.575 6.485 ;
      RECT 50.8 5.92 51.09 6.15 ;
      RECT 50.8 5.95 51.26 6.12 ;
      RECT 49.81 2.73 50.1 2.96 ;
      RECT 49.81 2.76 50.27 2.93 ;
      RECT 49.875 1.655 50.04 2.96 ;
      RECT 48.39 1.625 48.68 1.855 ;
      RECT 48.39 1.655 50.04 1.825 ;
      RECT 48.45 0.885 48.62 1.855 ;
      RECT 48.39 0.885 48.68 1.115 ;
      RECT 48.39 7.765 48.68 7.995 ;
      RECT 48.45 7.025 48.62 7.995 ;
      RECT 48.45 7.12 50.04 7.29 ;
      RECT 49.87 5.92 50.04 7.29 ;
      RECT 48.39 7.025 48.68 7.255 ;
      RECT 49.81 5.92 50.1 6.15 ;
      RECT 49.81 5.95 50.27 6.12 ;
      RECT 48.82 1.965 49.17 2.315 ;
      RECT 46.515 2.025 49.17 2.195 ;
      RECT 46.515 1.46 46.685 2.195 ;
      RECT 46.425 1.46 46.765 1.81 ;
      RECT 48.845 6.655 49.17 6.98 ;
      RECT 43.405 6.615 43.755 6.965 ;
      RECT 48.82 6.655 49.17 6.885 ;
      RECT 43.205 6.655 43.755 6.885 ;
      RECT 43.035 6.685 49.17 6.855 ;
      RECT 48.045 2.365 48.365 2.685 ;
      RECT 48.015 2.365 48.365 2.595 ;
      RECT 47.845 2.395 48.365 2.565 ;
      RECT 48.045 6.255 48.365 6.545 ;
      RECT 48.015 6.285 48.365 6.515 ;
      RECT 47.845 6.315 48.365 6.485 ;
      RECT 44.5 2.465 44.79 2.695 ;
      RECT 44.5 2.465 44.955 2.65 ;
      RECT 44.815 2.37 45.435 2.51 ;
      RECT 45.205 2.17 45.525 2.43 ;
      RECT 43.885 2.45 44.205 2.71 ;
      RECT 43.885 2.45 44.35 2.695 ;
      RECT 44.21 2.07 44.35 2.695 ;
      RECT 44.21 2.07 44.475 2.21 ;
      RECT 44.74 1.905 45.03 2.135 ;
      RECT 44.335 1.95 45.03 2.09 ;
      RECT 43.78 3.29 44.07 3.815 ;
      RECT 43.765 3.29 44.085 3.55 ;
      RECT 43.505 1.89 43.825 2.15 ;
      RECT 43.505 1.905 44.07 2.135 ;
      RECT 42.78 3.585 43.07 3.815 ;
      RECT 42.975 2.23 43.115 3.77 ;
      RECT 43.02 2.185 43.31 2.415 ;
      RECT 42.615 2.23 43.31 2.37 ;
      RECT 42.615 2.07 42.755 2.37 ;
      RECT 41.155 2.07 42.755 2.21 ;
      RECT 41.065 1.89 41.385 2.15 ;
      RECT 41.065 1.905 41.63 2.15 ;
      RECT 42.775 7.765 43.065 7.995 ;
      RECT 42.835 7.025 43.005 7.995 ;
      RECT 42.755 7.075 43.125 7.425 ;
      RECT 42.755 7.055 43.065 7.425 ;
      RECT 42.775 7.025 43.065 7.425 ;
      RECT 40.175 2.93 42.755 3.07 ;
      RECT 42.54 2.745 42.83 2.975 ;
      RECT 40.1 2.745 40.765 2.975 ;
      RECT 40.445 2.73 40.765 3.07 ;
      RECT 41.445 2.45 41.765 2.71 ;
      RECT 41.445 2.465 41.87 2.695 ;
      RECT 40.085 2.17 40.405 2.43 ;
      RECT 40.58 2.185 40.87 2.415 ;
      RECT 40.085 2.23 40.87 2.37 ;
      RECT 40.205 3.29 40.525 3.55 ;
      RECT 39.365 3.29 39.685 3.55 ;
      RECT 40.205 3.305 40.63 3.535 ;
      RECT 39.365 3.35 40.63 3.49 ;
      RECT 38.9 3.025 39.19 3.255 ;
      RECT 38.975 1.95 39.115 3.255 ;
      RECT 38.625 2.45 39.115 2.71 ;
      RECT 38.38 2.465 39.115 2.695 ;
      RECT 39.38 1.905 39.67 2.135 ;
      RECT 38.975 1.95 39.67 2.09 ;
      RECT 38.14 3.305 38.43 3.535 ;
      RECT 38.14 3.305 38.595 3.49 ;
      RECT 38.455 2.93 38.595 3.49 ;
      RECT 38.095 2.93 38.595 3.07 ;
      RECT 38.095 1.95 38.235 3.07 ;
      RECT 37.885 1.89 38.205 2.15 ;
      RECT 37.645 3.57 37.965 3.83 ;
      RECT 36.94 3.585 37.23 3.815 ;
      RECT 36.94 3.63 37.965 3.77 ;
      RECT 37.015 3.58 37.275 3.77 ;
      RECT 37.405 2.45 37.725 2.71 ;
      RECT 37.405 2.465 37.95 2.695 ;
      RECT 37.405 3.01 37.725 3.27 ;
      RECT 37.405 3.025 37.95 3.255 ;
      RECT 36.445 3.01 36.765 3.27 ;
      RECT 36.535 1.95 36.675 3.27 ;
      RECT 36.94 1.905 37.23 2.135 ;
      RECT 36.535 1.95 37.23 2.09 ;
      RECT 34.845 7.77 35.135 8 ;
      RECT 34.905 6.29 35.075 8 ;
      RECT 34.895 6.66 35.25 7.015 ;
      RECT 34.845 6.29 35.135 6.52 ;
      RECT 34.44 2.395 34.545 2.965 ;
      RECT 34.44 2.73 34.765 2.96 ;
      RECT 34.44 2.76 34.935 2.93 ;
      RECT 34.44 2.395 34.63 2.96 ;
      RECT 33.855 2.36 34.145 2.59 ;
      RECT 33.855 2.395 34.63 2.565 ;
      RECT 33.915 0.88 34.085 2.59 ;
      RECT 33.855 0.88 34.145 1.11 ;
      RECT 33.855 7.77 34.145 8 ;
      RECT 33.915 6.29 34.085 8 ;
      RECT 33.855 6.29 34.145 6.52 ;
      RECT 33.855 6.325 34.71 6.485 ;
      RECT 34.54 5.92 34.71 6.485 ;
      RECT 33.855 6.32 34.25 6.485 ;
      RECT 34.475 5.92 34.765 6.15 ;
      RECT 34.475 5.95 34.935 6.12 ;
      RECT 33.485 2.73 33.775 2.96 ;
      RECT 33.485 2.76 33.945 2.93 ;
      RECT 33.55 1.655 33.715 2.96 ;
      RECT 32.065 1.625 32.355 1.855 ;
      RECT 32.065 1.655 33.715 1.825 ;
      RECT 32.125 0.885 32.295 1.855 ;
      RECT 32.065 0.885 32.355 1.115 ;
      RECT 32.065 7.765 32.355 7.995 ;
      RECT 32.125 7.025 32.295 7.995 ;
      RECT 32.125 7.12 33.715 7.29 ;
      RECT 33.545 5.92 33.715 7.29 ;
      RECT 32.065 7.025 32.355 7.255 ;
      RECT 33.485 5.92 33.775 6.15 ;
      RECT 33.485 5.95 33.945 6.12 ;
      RECT 32.495 1.965 32.845 2.315 ;
      RECT 30.19 2.025 32.845 2.195 ;
      RECT 30.19 1.46 30.36 2.195 ;
      RECT 30.1 1.46 30.44 1.81 ;
      RECT 32.52 6.655 32.845 6.98 ;
      RECT 27.08 6.61 27.43 6.96 ;
      RECT 32.495 6.655 32.845 6.885 ;
      RECT 26.88 6.655 27.43 6.885 ;
      RECT 26.71 6.685 32.845 6.855 ;
      RECT 31.72 2.365 32.04 2.685 ;
      RECT 31.69 2.365 32.04 2.595 ;
      RECT 31.52 2.395 32.04 2.565 ;
      RECT 31.72 6.255 32.04 6.545 ;
      RECT 31.69 6.285 32.04 6.515 ;
      RECT 31.52 6.315 32.04 6.485 ;
      RECT 28.175 2.465 28.465 2.695 ;
      RECT 28.175 2.465 28.63 2.65 ;
      RECT 28.49 2.37 29.11 2.51 ;
      RECT 28.88 2.17 29.2 2.43 ;
      RECT 27.56 2.45 27.88 2.71 ;
      RECT 27.56 2.45 28.025 2.695 ;
      RECT 27.885 2.07 28.025 2.695 ;
      RECT 27.885 2.07 28.15 2.21 ;
      RECT 28.415 1.905 28.705 2.135 ;
      RECT 28.01 1.95 28.705 2.09 ;
      RECT 27.455 3.29 27.745 3.815 ;
      RECT 27.44 3.29 27.76 3.55 ;
      RECT 27.18 1.89 27.5 2.15 ;
      RECT 27.18 1.905 27.745 2.135 ;
      RECT 26.455 3.585 26.745 3.815 ;
      RECT 26.65 2.23 26.79 3.77 ;
      RECT 26.695 2.185 26.985 2.415 ;
      RECT 26.29 2.23 26.985 2.37 ;
      RECT 26.29 2.07 26.43 2.37 ;
      RECT 24.83 2.07 26.43 2.21 ;
      RECT 24.74 1.89 25.06 2.15 ;
      RECT 24.74 1.905 25.305 2.15 ;
      RECT 26.45 7.765 26.74 7.995 ;
      RECT 26.51 7.025 26.68 7.995 ;
      RECT 26.43 7.075 26.8 7.425 ;
      RECT 26.43 7.055 26.74 7.425 ;
      RECT 26.45 7.025 26.74 7.425 ;
      RECT 23.85 2.93 26.43 3.07 ;
      RECT 26.215 2.745 26.505 2.975 ;
      RECT 23.775 2.745 24.44 2.975 ;
      RECT 24.12 2.73 24.44 3.07 ;
      RECT 25.12 2.45 25.44 2.71 ;
      RECT 25.12 2.465 25.545 2.695 ;
      RECT 23.76 2.17 24.08 2.43 ;
      RECT 24.255 2.185 24.545 2.415 ;
      RECT 23.76 2.23 24.545 2.37 ;
      RECT 23.88 3.29 24.2 3.55 ;
      RECT 23.04 3.29 23.36 3.55 ;
      RECT 23.88 3.305 24.305 3.535 ;
      RECT 23.04 3.35 24.305 3.49 ;
      RECT 22.575 3.025 22.865 3.255 ;
      RECT 22.65 1.95 22.79 3.255 ;
      RECT 22.3 2.45 22.79 2.71 ;
      RECT 22.055 2.465 22.79 2.695 ;
      RECT 23.055 1.905 23.345 2.135 ;
      RECT 22.65 1.95 23.345 2.09 ;
      RECT 21.815 3.305 22.105 3.535 ;
      RECT 21.815 3.305 22.27 3.49 ;
      RECT 22.13 2.93 22.27 3.49 ;
      RECT 21.77 2.93 22.27 3.07 ;
      RECT 21.77 1.95 21.91 3.07 ;
      RECT 21.56 1.89 21.88 2.15 ;
      RECT 21.32 3.57 21.64 3.83 ;
      RECT 20.615 3.585 20.905 3.815 ;
      RECT 20.615 3.63 21.64 3.77 ;
      RECT 20.69 3.58 20.95 3.77 ;
      RECT 21.08 2.45 21.4 2.71 ;
      RECT 21.08 2.465 21.625 2.695 ;
      RECT 21.08 3.01 21.4 3.27 ;
      RECT 21.08 3.025 21.625 3.255 ;
      RECT 20.12 3.01 20.44 3.27 ;
      RECT 20.21 1.95 20.35 3.27 ;
      RECT 20.615 1.905 20.905 2.135 ;
      RECT 20.21 1.95 20.905 2.09 ;
      RECT 18.52 7.77 18.81 8 ;
      RECT 18.58 6.29 18.75 8 ;
      RECT 18.575 6.655 18.925 7.005 ;
      RECT 18.52 6.29 18.81 6.52 ;
      RECT 18.115 2.395 18.22 2.965 ;
      RECT 18.115 2.73 18.44 2.96 ;
      RECT 18.115 2.76 18.61 2.93 ;
      RECT 18.115 2.395 18.305 2.96 ;
      RECT 17.53 2.36 17.82 2.59 ;
      RECT 17.53 2.395 18.305 2.565 ;
      RECT 17.59 0.88 17.76 2.59 ;
      RECT 17.53 0.88 17.82 1.11 ;
      RECT 17.53 7.77 17.82 8 ;
      RECT 17.59 6.29 17.76 8 ;
      RECT 17.53 6.29 17.82 6.52 ;
      RECT 17.53 6.325 18.385 6.485 ;
      RECT 18.215 5.92 18.385 6.485 ;
      RECT 17.53 6.32 17.925 6.485 ;
      RECT 18.15 5.92 18.44 6.15 ;
      RECT 18.15 5.95 18.61 6.12 ;
      RECT 17.16 2.73 17.45 2.96 ;
      RECT 17.16 2.76 17.62 2.93 ;
      RECT 17.225 1.655 17.39 2.96 ;
      RECT 15.74 1.625 16.03 1.855 ;
      RECT 15.74 1.655 17.39 1.825 ;
      RECT 15.8 0.885 15.97 1.855 ;
      RECT 15.74 0.885 16.03 1.115 ;
      RECT 15.74 7.765 16.03 7.995 ;
      RECT 15.8 7.025 15.97 7.995 ;
      RECT 15.8 7.12 17.39 7.29 ;
      RECT 17.22 5.92 17.39 7.29 ;
      RECT 15.74 7.025 16.03 7.255 ;
      RECT 17.16 5.92 17.45 6.15 ;
      RECT 17.16 5.95 17.62 6.12 ;
      RECT 16.17 1.965 16.52 2.315 ;
      RECT 13.865 2.025 16.52 2.195 ;
      RECT 13.865 1.46 14.035 2.195 ;
      RECT 13.775 1.46 14.115 1.81 ;
      RECT 16.195 6.655 16.52 6.98 ;
      RECT 11.59 6.605 11.94 6.955 ;
      RECT 16.17 6.655 16.52 6.885 ;
      RECT 10.555 6.655 10.845 6.885 ;
      RECT 10.385 6.685 16.52 6.855 ;
      RECT 15.395 2.365 15.715 2.685 ;
      RECT 15.365 2.365 15.715 2.595 ;
      RECT 15.195 2.395 15.715 2.565 ;
      RECT 15.395 6.255 15.715 6.545 ;
      RECT 15.365 6.285 15.715 6.515 ;
      RECT 15.195 6.315 15.715 6.485 ;
      RECT 11.85 2.465 12.14 2.695 ;
      RECT 11.85 2.465 12.305 2.65 ;
      RECT 12.165 2.37 12.785 2.51 ;
      RECT 12.555 2.17 12.875 2.43 ;
      RECT 11.235 2.45 11.555 2.71 ;
      RECT 11.235 2.45 11.7 2.695 ;
      RECT 11.56 2.07 11.7 2.695 ;
      RECT 11.56 2.07 11.825 2.21 ;
      RECT 12.09 1.905 12.38 2.135 ;
      RECT 11.685 1.95 12.38 2.09 ;
      RECT 11.13 3.29 11.42 3.815 ;
      RECT 11.115 3.29 11.435 3.55 ;
      RECT 10.855 1.89 11.175 2.15 ;
      RECT 10.855 1.905 11.42 2.135 ;
      RECT 10.13 3.585 10.42 3.815 ;
      RECT 10.325 2.23 10.465 3.77 ;
      RECT 10.37 2.185 10.66 2.415 ;
      RECT 9.965 2.23 10.66 2.37 ;
      RECT 9.965 2.07 10.105 2.37 ;
      RECT 8.505 2.07 10.105 2.21 ;
      RECT 8.415 1.89 8.735 2.15 ;
      RECT 8.415 1.905 8.98 2.15 ;
      RECT 10.125 7.765 10.415 7.995 ;
      RECT 10.185 7.025 10.355 7.995 ;
      RECT 10.105 7.075 10.475 7.425 ;
      RECT 10.105 7.055 10.415 7.425 ;
      RECT 10.125 7.025 10.415 7.425 ;
      RECT 7.525 2.93 10.105 3.07 ;
      RECT 9.89 2.745 10.18 2.975 ;
      RECT 7.45 2.745 8.115 2.975 ;
      RECT 7.795 2.73 8.115 3.07 ;
      RECT 8.795 2.45 9.115 2.71 ;
      RECT 8.795 2.465 9.22 2.695 ;
      RECT 7.435 2.17 7.755 2.43 ;
      RECT 7.93 2.185 8.22 2.415 ;
      RECT 7.435 2.23 8.22 2.37 ;
      RECT 7.555 3.29 7.875 3.55 ;
      RECT 6.715 3.29 7.035 3.55 ;
      RECT 7.555 3.305 7.98 3.535 ;
      RECT 6.715 3.35 7.98 3.49 ;
      RECT 6.25 3.025 6.54 3.255 ;
      RECT 6.325 1.95 6.465 3.255 ;
      RECT 5.975 2.45 6.465 2.71 ;
      RECT 5.73 2.465 6.465 2.695 ;
      RECT 6.73 1.905 7.02 2.135 ;
      RECT 6.325 1.95 7.02 2.09 ;
      RECT 5.49 3.305 5.78 3.535 ;
      RECT 5.49 3.305 5.945 3.49 ;
      RECT 5.805 2.93 5.945 3.49 ;
      RECT 5.445 2.93 5.945 3.07 ;
      RECT 5.445 1.95 5.585 3.07 ;
      RECT 5.235 1.89 5.555 2.15 ;
      RECT 4.995 3.57 5.315 3.83 ;
      RECT 4.29 3.585 4.58 3.815 ;
      RECT 4.29 3.63 5.315 3.77 ;
      RECT 4.365 3.58 4.625 3.77 ;
      RECT 4.755 2.45 5.075 2.71 ;
      RECT 4.755 2.465 5.3 2.695 ;
      RECT 4.755 3.01 5.075 3.27 ;
      RECT 4.755 3.025 5.3 3.255 ;
      RECT 3.795 3.01 4.115 3.27 ;
      RECT 3.885 1.95 4.025 3.27 ;
      RECT 4.29 1.905 4.58 2.135 ;
      RECT 3.885 1.95 4.58 2.09 ;
      RECT 1.545 7.765 1.835 7.995 ;
      RECT 1.605 7.025 1.775 7.995 ;
      RECT 1.515 7.025 1.865 7.315 ;
      RECT 1.14 6.285 1.49 6.575 ;
      RECT 1 6.315 1.49 6.485 ;
      RECT 74.695 2.45 75.015 2.71 ;
      RECT 72.255 2.45 72.575 2.71 ;
      RECT 58.37 2.45 58.69 2.71 ;
      RECT 55.93 2.45 56.25 2.71 ;
      RECT 42.045 2.45 42.365 2.71 ;
      RECT 39.605 2.45 39.925 2.71 ;
      RECT 25.72 2.45 26.04 2.71 ;
      RECT 23.28 2.45 23.6 2.71 ;
      RECT 9.395 2.45 9.715 2.71 ;
      RECT 6.955 2.45 7.275 2.71 ;
    LAYER mcon ;
      RECT 83.88 6.32 84.05 6.49 ;
      RECT 83.885 6.315 84.055 6.485 ;
      RECT 67.555 6.32 67.725 6.49 ;
      RECT 67.56 6.315 67.73 6.485 ;
      RECT 51.23 6.32 51.4 6.49 ;
      RECT 51.235 6.315 51.405 6.485 ;
      RECT 34.905 6.32 35.075 6.49 ;
      RECT 34.91 6.315 35.08 6.485 ;
      RECT 18.58 6.32 18.75 6.49 ;
      RECT 18.585 6.315 18.755 6.485 ;
      RECT 83.88 7.8 84.05 7.97 ;
      RECT 83.51 2.76 83.68 2.93 ;
      RECT 83.51 5.95 83.68 6.12 ;
      RECT 82.89 0.91 83.06 1.08 ;
      RECT 82.89 2.39 83.06 2.56 ;
      RECT 82.89 6.32 83.06 6.49 ;
      RECT 82.89 7.8 83.06 7.97 ;
      RECT 82.52 2.76 82.69 2.93 ;
      RECT 82.52 5.95 82.69 6.12 ;
      RECT 81.53 2.025 81.7 2.195 ;
      RECT 81.53 6.685 81.7 6.855 ;
      RECT 81.1 0.915 81.27 1.085 ;
      RECT 81.1 1.655 81.27 1.825 ;
      RECT 81.1 7.055 81.27 7.225 ;
      RECT 81.1 7.795 81.27 7.965 ;
      RECT 80.725 2.395 80.895 2.565 ;
      RECT 80.725 6.315 80.895 6.485 ;
      RECT 77.45 1.935 77.62 2.105 ;
      RECT 77.21 2.495 77.38 2.665 ;
      RECT 76.73 2.495 76.9 2.665 ;
      RECT 76.49 1.935 76.66 2.105 ;
      RECT 76.49 3.615 76.66 3.785 ;
      RECT 75.915 6.685 76.085 6.855 ;
      RECT 75.73 2.215 75.9 2.385 ;
      RECT 75.49 3.615 75.66 3.785 ;
      RECT 75.485 7.055 75.655 7.225 ;
      RECT 75.485 7.795 75.655 7.965 ;
      RECT 75.25 2.775 75.42 2.945 ;
      RECT 74.77 2.495 74.94 2.665 ;
      RECT 74.29 2.495 74.46 2.665 ;
      RECT 74.05 1.935 74.22 2.105 ;
      RECT 73.29 2.215 73.46 2.385 ;
      RECT 73.05 3.335 73.22 3.505 ;
      RECT 72.81 2.775 72.98 2.945 ;
      RECT 72.33 2.495 72.5 2.665 ;
      RECT 72.09 1.935 72.26 2.105 ;
      RECT 72.09 3.335 72.26 3.505 ;
      RECT 71.61 3.055 71.78 3.225 ;
      RECT 71.09 2.495 71.26 2.665 ;
      RECT 70.85 3.335 71.02 3.505 ;
      RECT 70.61 1.935 70.78 2.105 ;
      RECT 70.37 2.495 70.54 2.665 ;
      RECT 70.37 3.055 70.54 3.225 ;
      RECT 69.65 1.935 69.82 2.105 ;
      RECT 69.65 3.615 69.82 3.785 ;
      RECT 69.17 3.055 69.34 3.225 ;
      RECT 67.555 7.8 67.725 7.97 ;
      RECT 67.185 2.76 67.355 2.93 ;
      RECT 67.185 5.95 67.355 6.12 ;
      RECT 66.565 0.91 66.735 1.08 ;
      RECT 66.565 2.39 66.735 2.56 ;
      RECT 66.565 6.32 66.735 6.49 ;
      RECT 66.565 7.8 66.735 7.97 ;
      RECT 66.195 2.76 66.365 2.93 ;
      RECT 66.195 5.95 66.365 6.12 ;
      RECT 65.205 2.025 65.375 2.195 ;
      RECT 65.205 6.685 65.375 6.855 ;
      RECT 64.775 0.915 64.945 1.085 ;
      RECT 64.775 1.655 64.945 1.825 ;
      RECT 64.775 7.055 64.945 7.225 ;
      RECT 64.775 7.795 64.945 7.965 ;
      RECT 64.4 2.395 64.57 2.565 ;
      RECT 64.4 6.315 64.57 6.485 ;
      RECT 61.125 1.935 61.295 2.105 ;
      RECT 60.885 2.495 61.055 2.665 ;
      RECT 60.405 2.495 60.575 2.665 ;
      RECT 60.165 1.935 60.335 2.105 ;
      RECT 60.165 3.615 60.335 3.785 ;
      RECT 59.59 6.685 59.76 6.855 ;
      RECT 59.405 2.215 59.575 2.385 ;
      RECT 59.165 3.615 59.335 3.785 ;
      RECT 59.16 7.055 59.33 7.225 ;
      RECT 59.16 7.795 59.33 7.965 ;
      RECT 58.925 2.775 59.095 2.945 ;
      RECT 58.445 2.495 58.615 2.665 ;
      RECT 57.965 2.495 58.135 2.665 ;
      RECT 57.725 1.935 57.895 2.105 ;
      RECT 56.965 2.215 57.135 2.385 ;
      RECT 56.725 3.335 56.895 3.505 ;
      RECT 56.485 2.775 56.655 2.945 ;
      RECT 56.005 2.495 56.175 2.665 ;
      RECT 55.765 1.935 55.935 2.105 ;
      RECT 55.765 3.335 55.935 3.505 ;
      RECT 55.285 3.055 55.455 3.225 ;
      RECT 54.765 2.495 54.935 2.665 ;
      RECT 54.525 3.335 54.695 3.505 ;
      RECT 54.285 1.935 54.455 2.105 ;
      RECT 54.045 2.495 54.215 2.665 ;
      RECT 54.045 3.055 54.215 3.225 ;
      RECT 53.325 1.935 53.495 2.105 ;
      RECT 53.325 3.615 53.495 3.785 ;
      RECT 52.845 3.055 53.015 3.225 ;
      RECT 51.23 7.8 51.4 7.97 ;
      RECT 50.86 2.76 51.03 2.93 ;
      RECT 50.86 5.95 51.03 6.12 ;
      RECT 50.24 0.91 50.41 1.08 ;
      RECT 50.24 2.39 50.41 2.56 ;
      RECT 50.24 6.32 50.41 6.49 ;
      RECT 50.24 7.8 50.41 7.97 ;
      RECT 49.87 2.76 50.04 2.93 ;
      RECT 49.87 5.95 50.04 6.12 ;
      RECT 48.88 2.025 49.05 2.195 ;
      RECT 48.88 6.685 49.05 6.855 ;
      RECT 48.45 0.915 48.62 1.085 ;
      RECT 48.45 1.655 48.62 1.825 ;
      RECT 48.45 7.055 48.62 7.225 ;
      RECT 48.45 7.795 48.62 7.965 ;
      RECT 48.075 2.395 48.245 2.565 ;
      RECT 48.075 6.315 48.245 6.485 ;
      RECT 44.8 1.935 44.97 2.105 ;
      RECT 44.56 2.495 44.73 2.665 ;
      RECT 44.08 2.495 44.25 2.665 ;
      RECT 43.84 1.935 44.01 2.105 ;
      RECT 43.84 3.615 44.01 3.785 ;
      RECT 43.265 6.685 43.435 6.855 ;
      RECT 43.08 2.215 43.25 2.385 ;
      RECT 42.84 3.615 43.01 3.785 ;
      RECT 42.835 7.055 43.005 7.225 ;
      RECT 42.835 7.795 43.005 7.965 ;
      RECT 42.6 2.775 42.77 2.945 ;
      RECT 42.12 2.495 42.29 2.665 ;
      RECT 41.64 2.495 41.81 2.665 ;
      RECT 41.4 1.935 41.57 2.105 ;
      RECT 40.64 2.215 40.81 2.385 ;
      RECT 40.4 3.335 40.57 3.505 ;
      RECT 40.16 2.775 40.33 2.945 ;
      RECT 39.68 2.495 39.85 2.665 ;
      RECT 39.44 1.935 39.61 2.105 ;
      RECT 39.44 3.335 39.61 3.505 ;
      RECT 38.96 3.055 39.13 3.225 ;
      RECT 38.44 2.495 38.61 2.665 ;
      RECT 38.2 3.335 38.37 3.505 ;
      RECT 37.96 1.935 38.13 2.105 ;
      RECT 37.72 2.495 37.89 2.665 ;
      RECT 37.72 3.055 37.89 3.225 ;
      RECT 37 1.935 37.17 2.105 ;
      RECT 37 3.615 37.17 3.785 ;
      RECT 36.52 3.055 36.69 3.225 ;
      RECT 34.905 7.8 35.075 7.97 ;
      RECT 34.535 2.76 34.705 2.93 ;
      RECT 34.535 5.95 34.705 6.12 ;
      RECT 33.915 0.91 34.085 1.08 ;
      RECT 33.915 2.39 34.085 2.56 ;
      RECT 33.915 6.32 34.085 6.49 ;
      RECT 33.915 7.8 34.085 7.97 ;
      RECT 33.545 2.76 33.715 2.93 ;
      RECT 33.545 5.95 33.715 6.12 ;
      RECT 32.555 2.025 32.725 2.195 ;
      RECT 32.555 6.685 32.725 6.855 ;
      RECT 32.125 0.915 32.295 1.085 ;
      RECT 32.125 1.655 32.295 1.825 ;
      RECT 32.125 7.055 32.295 7.225 ;
      RECT 32.125 7.795 32.295 7.965 ;
      RECT 31.75 2.395 31.92 2.565 ;
      RECT 31.75 6.315 31.92 6.485 ;
      RECT 28.475 1.935 28.645 2.105 ;
      RECT 28.235 2.495 28.405 2.665 ;
      RECT 27.755 2.495 27.925 2.665 ;
      RECT 27.515 1.935 27.685 2.105 ;
      RECT 27.515 3.615 27.685 3.785 ;
      RECT 26.94 6.685 27.11 6.855 ;
      RECT 26.755 2.215 26.925 2.385 ;
      RECT 26.515 3.615 26.685 3.785 ;
      RECT 26.51 7.055 26.68 7.225 ;
      RECT 26.51 7.795 26.68 7.965 ;
      RECT 26.275 2.775 26.445 2.945 ;
      RECT 25.795 2.495 25.965 2.665 ;
      RECT 25.315 2.495 25.485 2.665 ;
      RECT 25.075 1.935 25.245 2.105 ;
      RECT 24.315 2.215 24.485 2.385 ;
      RECT 24.075 3.335 24.245 3.505 ;
      RECT 23.835 2.775 24.005 2.945 ;
      RECT 23.355 2.495 23.525 2.665 ;
      RECT 23.115 1.935 23.285 2.105 ;
      RECT 23.115 3.335 23.285 3.505 ;
      RECT 22.635 3.055 22.805 3.225 ;
      RECT 22.115 2.495 22.285 2.665 ;
      RECT 21.875 3.335 22.045 3.505 ;
      RECT 21.635 1.935 21.805 2.105 ;
      RECT 21.395 2.495 21.565 2.665 ;
      RECT 21.395 3.055 21.565 3.225 ;
      RECT 20.675 1.935 20.845 2.105 ;
      RECT 20.675 3.615 20.845 3.785 ;
      RECT 20.195 3.055 20.365 3.225 ;
      RECT 18.58 7.8 18.75 7.97 ;
      RECT 18.21 2.76 18.38 2.93 ;
      RECT 18.21 5.95 18.38 6.12 ;
      RECT 17.59 0.91 17.76 1.08 ;
      RECT 17.59 2.39 17.76 2.56 ;
      RECT 17.59 6.32 17.76 6.49 ;
      RECT 17.59 7.8 17.76 7.97 ;
      RECT 17.22 2.76 17.39 2.93 ;
      RECT 17.22 5.95 17.39 6.12 ;
      RECT 16.23 2.025 16.4 2.195 ;
      RECT 16.23 6.685 16.4 6.855 ;
      RECT 15.8 0.915 15.97 1.085 ;
      RECT 15.8 1.655 15.97 1.825 ;
      RECT 15.8 7.055 15.97 7.225 ;
      RECT 15.8 7.795 15.97 7.965 ;
      RECT 15.425 2.395 15.595 2.565 ;
      RECT 15.425 6.315 15.595 6.485 ;
      RECT 12.15 1.935 12.32 2.105 ;
      RECT 11.91 2.495 12.08 2.665 ;
      RECT 11.43 2.495 11.6 2.665 ;
      RECT 11.19 1.935 11.36 2.105 ;
      RECT 11.19 3.615 11.36 3.785 ;
      RECT 10.615 6.685 10.785 6.855 ;
      RECT 10.43 2.215 10.6 2.385 ;
      RECT 10.19 3.615 10.36 3.785 ;
      RECT 10.185 7.055 10.355 7.225 ;
      RECT 10.185 7.795 10.355 7.965 ;
      RECT 9.95 2.775 10.12 2.945 ;
      RECT 9.47 2.495 9.64 2.665 ;
      RECT 8.99 2.495 9.16 2.665 ;
      RECT 8.75 1.935 8.92 2.105 ;
      RECT 7.99 2.215 8.16 2.385 ;
      RECT 7.75 3.335 7.92 3.505 ;
      RECT 7.51 2.775 7.68 2.945 ;
      RECT 7.03 2.495 7.2 2.665 ;
      RECT 6.79 1.935 6.96 2.105 ;
      RECT 6.79 3.335 6.96 3.505 ;
      RECT 6.31 3.055 6.48 3.225 ;
      RECT 5.79 2.495 5.96 2.665 ;
      RECT 5.55 3.335 5.72 3.505 ;
      RECT 5.31 1.935 5.48 2.105 ;
      RECT 5.07 2.495 5.24 2.665 ;
      RECT 5.07 3.055 5.24 3.225 ;
      RECT 4.35 1.935 4.52 2.105 ;
      RECT 4.35 3.615 4.52 3.785 ;
      RECT 3.87 3.055 4.04 3.225 ;
      RECT 1.605 7.055 1.775 7.225 ;
      RECT 1.605 7.795 1.775 7.965 ;
      RECT 1.23 6.315 1.4 6.485 ;
    LAYER li1 ;
      RECT 83.88 5.02 84.05 6.49 ;
      RECT 83.88 6.315 84.055 6.485 ;
      RECT 83.51 1.74 83.68 2.93 ;
      RECT 83.51 1.74 83.98 1.91 ;
      RECT 83.51 6.97 83.98 7.14 ;
      RECT 83.51 5.95 83.68 7.14 ;
      RECT 82.52 1.74 82.69 2.93 ;
      RECT 82.52 1.74 82.99 1.91 ;
      RECT 82.52 6.97 82.99 7.14 ;
      RECT 82.52 5.95 82.69 7.14 ;
      RECT 80.67 2.635 80.84 3.865 ;
      RECT 80.725 0.855 80.895 2.805 ;
      RECT 80.67 0.575 80.84 1.025 ;
      RECT 80.67 7.855 80.84 8.305 ;
      RECT 80.725 6.075 80.895 8.025 ;
      RECT 80.67 5.015 80.84 6.245 ;
      RECT 80.15 0.575 80.32 3.865 ;
      RECT 80.15 2.075 80.555 2.405 ;
      RECT 80.15 1.235 80.555 1.565 ;
      RECT 80.15 5.015 80.32 8.305 ;
      RECT 80.15 7.315 80.555 7.645 ;
      RECT 80.15 6.475 80.555 6.805 ;
      RECT 77.45 1.835 77.62 2.105 ;
      RECT 77.45 1.835 78.18 2.005 ;
      RECT 77.37 3.225 77.7 3.395 ;
      RECT 76.61 3.055 77.62 3.225 ;
      RECT 76.61 2.575 76.78 3.225 ;
      RECT 76.73 2.495 76.9 2.825 ;
      RECT 75.89 3.225 76.22 3.395 ;
      RECT 73.97 3.225 75.26 3.395 ;
      RECT 75.01 3.14 76.14 3.31 ;
      RECT 75.73 2.215 76.14 2.385 ;
      RECT 75.97 1.755 76.14 2.385 ;
      RECT 74.535 5.015 74.705 8.305 ;
      RECT 74.535 7.315 74.94 7.645 ;
      RECT 74.535 6.475 74.94 6.805 ;
      RECT 73.21 2.575 74.54 2.745 ;
      RECT 74.29 2.495 74.46 2.745 ;
      RECT 73.29 2.175 73.46 2.385 ;
      RECT 73.29 2.175 73.78 2.345 ;
      RECT 71.97 3.335 72.26 3.505 ;
      RECT 71.97 2.575 72.14 3.505 ;
      RECT 71.77 2.575 72.14 2.745 ;
      RECT 70.77 2.575 71.26 2.745 ;
      RECT 71.09 2.495 71.26 2.745 ;
      RECT 70.85 3.335 71.26 3.505 ;
      RECT 71.09 3.145 71.26 3.505 ;
      RECT 69.89 3.055 70.54 3.225 ;
      RECT 69.89 2.495 70.06 3.225 ;
      RECT 69.53 3.615 69.82 3.785 ;
      RECT 69.53 2.575 69.7 3.785 ;
      RECT 69.33 2.575 69.7 2.745 ;
      RECT 67.555 5.02 67.725 6.49 ;
      RECT 67.555 6.315 67.73 6.485 ;
      RECT 67.185 1.74 67.355 2.93 ;
      RECT 67.185 1.74 67.655 1.91 ;
      RECT 67.185 6.97 67.655 7.14 ;
      RECT 67.185 5.95 67.355 7.14 ;
      RECT 66.195 1.74 66.365 2.93 ;
      RECT 66.195 1.74 66.665 1.91 ;
      RECT 66.195 6.97 66.665 7.14 ;
      RECT 66.195 5.95 66.365 7.14 ;
      RECT 64.345 2.635 64.515 3.865 ;
      RECT 64.4 0.855 64.57 2.805 ;
      RECT 64.345 0.575 64.515 1.025 ;
      RECT 64.345 7.855 64.515 8.305 ;
      RECT 64.4 6.075 64.57 8.025 ;
      RECT 64.345 5.015 64.515 6.245 ;
      RECT 63.825 0.575 63.995 3.865 ;
      RECT 63.825 2.075 64.23 2.405 ;
      RECT 63.825 1.235 64.23 1.565 ;
      RECT 63.825 5.015 63.995 8.305 ;
      RECT 63.825 7.315 64.23 7.645 ;
      RECT 63.825 6.475 64.23 6.805 ;
      RECT 61.125 1.835 61.295 2.105 ;
      RECT 61.125 1.835 61.855 2.005 ;
      RECT 61.045 3.225 61.375 3.395 ;
      RECT 60.285 3.055 61.295 3.225 ;
      RECT 60.285 2.575 60.455 3.225 ;
      RECT 60.405 2.495 60.575 2.825 ;
      RECT 59.565 3.225 59.895 3.395 ;
      RECT 57.645 3.225 58.935 3.395 ;
      RECT 58.685 3.14 59.815 3.31 ;
      RECT 59.405 2.215 59.815 2.385 ;
      RECT 59.645 1.755 59.815 2.385 ;
      RECT 58.21 5.015 58.38 8.305 ;
      RECT 58.21 7.315 58.615 7.645 ;
      RECT 58.21 6.475 58.615 6.805 ;
      RECT 56.885 2.575 58.215 2.745 ;
      RECT 57.965 2.495 58.135 2.745 ;
      RECT 56.965 2.175 57.135 2.385 ;
      RECT 56.965 2.175 57.455 2.345 ;
      RECT 55.645 3.335 55.935 3.505 ;
      RECT 55.645 2.575 55.815 3.505 ;
      RECT 55.445 2.575 55.815 2.745 ;
      RECT 54.445 2.575 54.935 2.745 ;
      RECT 54.765 2.495 54.935 2.745 ;
      RECT 54.525 3.335 54.935 3.505 ;
      RECT 54.765 3.145 54.935 3.505 ;
      RECT 53.565 3.055 54.215 3.225 ;
      RECT 53.565 2.495 53.735 3.225 ;
      RECT 53.205 3.615 53.495 3.785 ;
      RECT 53.205 2.575 53.375 3.785 ;
      RECT 53.005 2.575 53.375 2.745 ;
      RECT 51.23 5.02 51.4 6.49 ;
      RECT 51.23 6.315 51.405 6.485 ;
      RECT 50.86 1.74 51.03 2.93 ;
      RECT 50.86 1.74 51.33 1.91 ;
      RECT 50.86 6.97 51.33 7.14 ;
      RECT 50.86 5.95 51.03 7.14 ;
      RECT 49.87 1.74 50.04 2.93 ;
      RECT 49.87 1.74 50.34 1.91 ;
      RECT 49.87 6.97 50.34 7.14 ;
      RECT 49.87 5.95 50.04 7.14 ;
      RECT 48.02 2.635 48.19 3.865 ;
      RECT 48.075 0.855 48.245 2.805 ;
      RECT 48.02 0.575 48.19 1.025 ;
      RECT 48.02 7.855 48.19 8.305 ;
      RECT 48.075 6.075 48.245 8.025 ;
      RECT 48.02 5.015 48.19 6.245 ;
      RECT 47.5 0.575 47.67 3.865 ;
      RECT 47.5 2.075 47.905 2.405 ;
      RECT 47.5 1.235 47.905 1.565 ;
      RECT 47.5 5.015 47.67 8.305 ;
      RECT 47.5 7.315 47.905 7.645 ;
      RECT 47.5 6.475 47.905 6.805 ;
      RECT 44.8 1.835 44.97 2.105 ;
      RECT 44.8 1.835 45.53 2.005 ;
      RECT 44.72 3.225 45.05 3.395 ;
      RECT 43.96 3.055 44.97 3.225 ;
      RECT 43.96 2.575 44.13 3.225 ;
      RECT 44.08 2.495 44.25 2.825 ;
      RECT 43.24 3.225 43.57 3.395 ;
      RECT 41.32 3.225 42.61 3.395 ;
      RECT 42.36 3.14 43.49 3.31 ;
      RECT 43.08 2.215 43.49 2.385 ;
      RECT 43.32 1.755 43.49 2.385 ;
      RECT 41.885 5.015 42.055 8.305 ;
      RECT 41.885 7.315 42.29 7.645 ;
      RECT 41.885 6.475 42.29 6.805 ;
      RECT 40.56 2.575 41.89 2.745 ;
      RECT 41.64 2.495 41.81 2.745 ;
      RECT 40.64 2.175 40.81 2.385 ;
      RECT 40.64 2.175 41.13 2.345 ;
      RECT 39.32 3.335 39.61 3.505 ;
      RECT 39.32 2.575 39.49 3.505 ;
      RECT 39.12 2.575 39.49 2.745 ;
      RECT 38.12 2.575 38.61 2.745 ;
      RECT 38.44 2.495 38.61 2.745 ;
      RECT 38.2 3.335 38.61 3.505 ;
      RECT 38.44 3.145 38.61 3.505 ;
      RECT 37.24 3.055 37.89 3.225 ;
      RECT 37.24 2.495 37.41 3.225 ;
      RECT 36.88 3.615 37.17 3.785 ;
      RECT 36.88 2.575 37.05 3.785 ;
      RECT 36.68 2.575 37.05 2.745 ;
      RECT 34.905 5.02 35.075 6.49 ;
      RECT 34.905 6.315 35.08 6.485 ;
      RECT 34.535 1.74 34.705 2.93 ;
      RECT 34.535 1.74 35.005 1.91 ;
      RECT 34.535 6.97 35.005 7.14 ;
      RECT 34.535 5.95 34.705 7.14 ;
      RECT 33.545 1.74 33.715 2.93 ;
      RECT 33.545 1.74 34.015 1.91 ;
      RECT 33.545 6.97 34.015 7.14 ;
      RECT 33.545 5.95 33.715 7.14 ;
      RECT 31.695 2.635 31.865 3.865 ;
      RECT 31.75 0.855 31.92 2.805 ;
      RECT 31.695 0.575 31.865 1.025 ;
      RECT 31.695 7.855 31.865 8.305 ;
      RECT 31.75 6.075 31.92 8.025 ;
      RECT 31.695 5.015 31.865 6.245 ;
      RECT 31.175 0.575 31.345 3.865 ;
      RECT 31.175 2.075 31.58 2.405 ;
      RECT 31.175 1.235 31.58 1.565 ;
      RECT 31.175 5.015 31.345 8.305 ;
      RECT 31.175 7.315 31.58 7.645 ;
      RECT 31.175 6.475 31.58 6.805 ;
      RECT 28.475 1.835 28.645 2.105 ;
      RECT 28.475 1.835 29.205 2.005 ;
      RECT 28.395 3.225 28.725 3.395 ;
      RECT 27.635 3.055 28.645 3.225 ;
      RECT 27.635 2.575 27.805 3.225 ;
      RECT 27.755 2.495 27.925 2.825 ;
      RECT 26.915 3.225 27.245 3.395 ;
      RECT 24.995 3.225 26.285 3.395 ;
      RECT 26.035 3.14 27.165 3.31 ;
      RECT 26.755 2.215 27.165 2.385 ;
      RECT 26.995 1.755 27.165 2.385 ;
      RECT 25.56 5.015 25.73 8.305 ;
      RECT 25.56 7.315 25.965 7.645 ;
      RECT 25.56 6.475 25.965 6.805 ;
      RECT 24.235 2.575 25.565 2.745 ;
      RECT 25.315 2.495 25.485 2.745 ;
      RECT 24.315 2.175 24.485 2.385 ;
      RECT 24.315 2.175 24.805 2.345 ;
      RECT 22.995 3.335 23.285 3.505 ;
      RECT 22.995 2.575 23.165 3.505 ;
      RECT 22.795 2.575 23.165 2.745 ;
      RECT 21.795 2.575 22.285 2.745 ;
      RECT 22.115 2.495 22.285 2.745 ;
      RECT 21.875 3.335 22.285 3.505 ;
      RECT 22.115 3.145 22.285 3.505 ;
      RECT 20.915 3.055 21.565 3.225 ;
      RECT 20.915 2.495 21.085 3.225 ;
      RECT 20.555 3.615 20.845 3.785 ;
      RECT 20.555 2.575 20.725 3.785 ;
      RECT 20.355 2.575 20.725 2.745 ;
      RECT 18.58 5.02 18.75 6.49 ;
      RECT 18.58 6.315 18.755 6.485 ;
      RECT 18.21 1.74 18.38 2.93 ;
      RECT 18.21 1.74 18.68 1.91 ;
      RECT 18.21 6.97 18.68 7.14 ;
      RECT 18.21 5.95 18.38 7.14 ;
      RECT 17.22 1.74 17.39 2.93 ;
      RECT 17.22 1.74 17.69 1.91 ;
      RECT 17.22 6.97 17.69 7.14 ;
      RECT 17.22 5.95 17.39 7.14 ;
      RECT 15.37 2.635 15.54 3.865 ;
      RECT 15.425 0.855 15.595 2.805 ;
      RECT 15.37 0.575 15.54 1.025 ;
      RECT 15.37 7.855 15.54 8.305 ;
      RECT 15.425 6.075 15.595 8.025 ;
      RECT 15.37 5.015 15.54 6.245 ;
      RECT 14.85 0.575 15.02 3.865 ;
      RECT 14.85 2.075 15.255 2.405 ;
      RECT 14.85 1.235 15.255 1.565 ;
      RECT 14.85 5.015 15.02 8.305 ;
      RECT 14.85 7.315 15.255 7.645 ;
      RECT 14.85 6.475 15.255 6.805 ;
      RECT 12.15 1.835 12.32 2.105 ;
      RECT 12.15 1.835 12.88 2.005 ;
      RECT 12.07 3.225 12.4 3.395 ;
      RECT 11.31 3.055 12.32 3.225 ;
      RECT 11.31 2.575 11.48 3.225 ;
      RECT 11.43 2.495 11.6 2.825 ;
      RECT 10.59 3.225 10.92 3.395 ;
      RECT 8.67 3.225 9.96 3.395 ;
      RECT 9.71 3.14 10.84 3.31 ;
      RECT 10.43 2.215 10.84 2.385 ;
      RECT 10.67 1.755 10.84 2.385 ;
      RECT 9.235 5.015 9.405 8.305 ;
      RECT 9.235 7.315 9.64 7.645 ;
      RECT 9.235 6.475 9.64 6.805 ;
      RECT 7.91 2.575 9.24 2.745 ;
      RECT 8.99 2.495 9.16 2.745 ;
      RECT 7.99 2.175 8.16 2.385 ;
      RECT 7.99 2.175 8.48 2.345 ;
      RECT 6.67 3.335 6.96 3.505 ;
      RECT 6.67 2.575 6.84 3.505 ;
      RECT 6.47 2.575 6.84 2.745 ;
      RECT 5.47 2.575 5.96 2.745 ;
      RECT 5.79 2.495 5.96 2.745 ;
      RECT 5.55 3.335 5.96 3.505 ;
      RECT 5.79 3.145 5.96 3.505 ;
      RECT 4.59 3.055 5.24 3.225 ;
      RECT 4.59 2.495 4.76 3.225 ;
      RECT 4.23 3.615 4.52 3.785 ;
      RECT 4.23 2.575 4.4 3.785 ;
      RECT 4.03 2.575 4.4 2.745 ;
      RECT 1.175 7.855 1.345 8.305 ;
      RECT 1.23 6.075 1.4 8.025 ;
      RECT 1.175 5.015 1.345 6.245 ;
      RECT 0.655 5.015 0.825 8.305 ;
      RECT 0.655 7.315 1.06 7.645 ;
      RECT 0.655 6.475 1.06 6.805 ;
      RECT 83.88 7.8 84.05 8.31 ;
      RECT 82.89 0.57 83.06 1.08 ;
      RECT 82.89 2.39 83.06 3.86 ;
      RECT 82.89 5.02 83.06 6.49 ;
      RECT 82.89 7.8 83.06 8.31 ;
      RECT 81.53 0.575 81.7 3.865 ;
      RECT 81.53 5.015 81.7 8.305 ;
      RECT 81.1 0.575 81.27 1.085 ;
      RECT 81.1 1.655 81.27 3.865 ;
      RECT 81.1 5.015 81.27 7.225 ;
      RECT 81.1 7.795 81.27 8.305 ;
      RECT 77.21 2.495 77.38 2.825 ;
      RECT 76.49 1.755 76.66 2.105 ;
      RECT 76.49 3.485 76.66 3.815 ;
      RECT 75.915 5.015 76.085 8.305 ;
      RECT 75.49 3.485 75.66 3.815 ;
      RECT 75.485 5.015 75.655 7.225 ;
      RECT 75.485 7.795 75.655 8.305 ;
      RECT 75.25 2.495 75.42 2.945 ;
      RECT 74.77 2.495 74.94 2.825 ;
      RECT 74.05 1.755 74.22 2.105 ;
      RECT 73.05 3.145 73.22 3.505 ;
      RECT 72.81 2.495 72.98 2.945 ;
      RECT 72.33 2.495 72.5 2.825 ;
      RECT 72.09 1.755 72.26 2.105 ;
      RECT 71.61 3.055 71.78 3.475 ;
      RECT 70.61 1.755 70.78 2.105 ;
      RECT 70.37 2.495 70.54 2.825 ;
      RECT 69.65 1.755 69.82 2.105 ;
      RECT 69.17 3.055 69.34 3.475 ;
      RECT 67.555 7.8 67.725 8.31 ;
      RECT 66.565 0.57 66.735 1.08 ;
      RECT 66.565 2.39 66.735 3.86 ;
      RECT 66.565 5.02 66.735 6.49 ;
      RECT 66.565 7.8 66.735 8.31 ;
      RECT 65.205 0.575 65.375 3.865 ;
      RECT 65.205 5.015 65.375 8.305 ;
      RECT 64.775 0.575 64.945 1.085 ;
      RECT 64.775 1.655 64.945 3.865 ;
      RECT 64.775 5.015 64.945 7.225 ;
      RECT 64.775 7.795 64.945 8.305 ;
      RECT 60.885 2.495 61.055 2.825 ;
      RECT 60.165 1.755 60.335 2.105 ;
      RECT 60.165 3.485 60.335 3.815 ;
      RECT 59.59 5.015 59.76 8.305 ;
      RECT 59.165 3.485 59.335 3.815 ;
      RECT 59.16 5.015 59.33 7.225 ;
      RECT 59.16 7.795 59.33 8.305 ;
      RECT 58.925 2.495 59.095 2.945 ;
      RECT 58.445 2.495 58.615 2.825 ;
      RECT 57.725 1.755 57.895 2.105 ;
      RECT 56.725 3.145 56.895 3.505 ;
      RECT 56.485 2.495 56.655 2.945 ;
      RECT 56.005 2.495 56.175 2.825 ;
      RECT 55.765 1.755 55.935 2.105 ;
      RECT 55.285 3.055 55.455 3.475 ;
      RECT 54.285 1.755 54.455 2.105 ;
      RECT 54.045 2.495 54.215 2.825 ;
      RECT 53.325 1.755 53.495 2.105 ;
      RECT 52.845 3.055 53.015 3.475 ;
      RECT 51.23 7.8 51.4 8.31 ;
      RECT 50.24 0.57 50.41 1.08 ;
      RECT 50.24 2.39 50.41 3.86 ;
      RECT 50.24 5.02 50.41 6.49 ;
      RECT 50.24 7.8 50.41 8.31 ;
      RECT 48.88 0.575 49.05 3.865 ;
      RECT 48.88 5.015 49.05 8.305 ;
      RECT 48.45 0.575 48.62 1.085 ;
      RECT 48.45 1.655 48.62 3.865 ;
      RECT 48.45 5.015 48.62 7.225 ;
      RECT 48.45 7.795 48.62 8.305 ;
      RECT 44.56 2.495 44.73 2.825 ;
      RECT 43.84 1.755 44.01 2.105 ;
      RECT 43.84 3.485 44.01 3.815 ;
      RECT 43.265 5.015 43.435 8.305 ;
      RECT 42.84 3.485 43.01 3.815 ;
      RECT 42.835 5.015 43.005 7.225 ;
      RECT 42.835 7.795 43.005 8.305 ;
      RECT 42.6 2.495 42.77 2.945 ;
      RECT 42.12 2.495 42.29 2.825 ;
      RECT 41.4 1.755 41.57 2.105 ;
      RECT 40.4 3.145 40.57 3.505 ;
      RECT 40.16 2.495 40.33 2.945 ;
      RECT 39.68 2.495 39.85 2.825 ;
      RECT 39.44 1.755 39.61 2.105 ;
      RECT 38.96 3.055 39.13 3.475 ;
      RECT 37.96 1.755 38.13 2.105 ;
      RECT 37.72 2.495 37.89 2.825 ;
      RECT 37 1.755 37.17 2.105 ;
      RECT 36.52 3.055 36.69 3.475 ;
      RECT 34.905 7.8 35.075 8.31 ;
      RECT 33.915 0.57 34.085 1.08 ;
      RECT 33.915 2.39 34.085 3.86 ;
      RECT 33.915 5.02 34.085 6.49 ;
      RECT 33.915 7.8 34.085 8.31 ;
      RECT 32.555 0.575 32.725 3.865 ;
      RECT 32.555 5.015 32.725 8.305 ;
      RECT 32.125 0.575 32.295 1.085 ;
      RECT 32.125 1.655 32.295 3.865 ;
      RECT 32.125 5.015 32.295 7.225 ;
      RECT 32.125 7.795 32.295 8.305 ;
      RECT 28.235 2.495 28.405 2.825 ;
      RECT 27.515 1.755 27.685 2.105 ;
      RECT 27.515 3.485 27.685 3.815 ;
      RECT 26.94 5.015 27.11 8.305 ;
      RECT 26.515 3.485 26.685 3.815 ;
      RECT 26.51 5.015 26.68 7.225 ;
      RECT 26.51 7.795 26.68 8.305 ;
      RECT 26.275 2.495 26.445 2.945 ;
      RECT 25.795 2.495 25.965 2.825 ;
      RECT 25.075 1.755 25.245 2.105 ;
      RECT 24.075 3.145 24.245 3.505 ;
      RECT 23.835 2.495 24.005 2.945 ;
      RECT 23.355 2.495 23.525 2.825 ;
      RECT 23.115 1.755 23.285 2.105 ;
      RECT 22.635 3.055 22.805 3.475 ;
      RECT 21.635 1.755 21.805 2.105 ;
      RECT 21.395 2.495 21.565 2.825 ;
      RECT 20.675 1.755 20.845 2.105 ;
      RECT 20.195 3.055 20.365 3.475 ;
      RECT 18.58 7.8 18.75 8.31 ;
      RECT 17.59 0.57 17.76 1.08 ;
      RECT 17.59 2.39 17.76 3.86 ;
      RECT 17.59 5.02 17.76 6.49 ;
      RECT 17.59 7.8 17.76 8.31 ;
      RECT 16.23 0.575 16.4 3.865 ;
      RECT 16.23 5.015 16.4 8.305 ;
      RECT 15.8 0.575 15.97 1.085 ;
      RECT 15.8 1.655 15.97 3.865 ;
      RECT 15.8 5.015 15.97 7.225 ;
      RECT 15.8 7.795 15.97 8.305 ;
      RECT 11.91 2.495 12.08 2.825 ;
      RECT 11.19 1.755 11.36 2.105 ;
      RECT 11.19 3.485 11.36 3.815 ;
      RECT 10.615 5.015 10.785 8.305 ;
      RECT 10.19 3.485 10.36 3.815 ;
      RECT 10.185 5.015 10.355 7.225 ;
      RECT 10.185 7.795 10.355 8.305 ;
      RECT 9.95 2.495 10.12 2.945 ;
      RECT 9.47 2.495 9.64 2.825 ;
      RECT 8.75 1.755 8.92 2.105 ;
      RECT 7.75 3.145 7.92 3.505 ;
      RECT 7.51 2.495 7.68 2.945 ;
      RECT 7.03 2.495 7.2 2.825 ;
      RECT 6.79 1.755 6.96 2.105 ;
      RECT 6.31 3.055 6.48 3.475 ;
      RECT 5.31 1.755 5.48 2.105 ;
      RECT 5.07 2.495 5.24 2.825 ;
      RECT 4.35 1.755 4.52 2.105 ;
      RECT 3.87 3.055 4.04 3.475 ;
      RECT 1.605 5.015 1.775 7.225 ;
      RECT 1.605 7.795 1.775 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r2 ;
  SIZE 84.42 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 18.58 0.915 18.75 1.085 ;
        RECT 18.575 0.91 18.745 1.08 ;
        RECT 18.575 2.39 18.745 2.56 ;
      LAYER li1 ;
        RECT 18.58 0.915 18.75 1.085 ;
        RECT 18.575 0.57 18.745 1.08 ;
        RECT 18.575 2.39 18.745 3.86 ;
      LAYER met1 ;
        RECT 18.515 2.36 18.805 2.59 ;
        RECT 18.515 0.88 18.805 1.11 ;
        RECT 18.575 0.88 18.745 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 34.905 0.915 35.075 1.085 ;
        RECT 34.9 0.91 35.07 1.08 ;
        RECT 34.9 2.39 35.07 2.56 ;
      LAYER li1 ;
        RECT 34.905 0.915 35.075 1.085 ;
        RECT 34.9 0.57 35.07 1.08 ;
        RECT 34.9 2.39 35.07 3.86 ;
      LAYER met1 ;
        RECT 34.84 2.36 35.13 2.59 ;
        RECT 34.84 0.88 35.13 1.11 ;
        RECT 34.9 0.88 35.07 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 51.23 0.915 51.4 1.085 ;
        RECT 51.225 0.91 51.395 1.08 ;
        RECT 51.225 2.39 51.395 2.56 ;
      LAYER li1 ;
        RECT 51.23 0.915 51.4 1.085 ;
        RECT 51.225 0.57 51.395 1.08 ;
        RECT 51.225 2.39 51.395 3.86 ;
      LAYER met1 ;
        RECT 51.165 2.36 51.455 2.59 ;
        RECT 51.165 0.88 51.455 1.11 ;
        RECT 51.225 0.88 51.395 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 67.555 0.915 67.725 1.085 ;
        RECT 67.55 0.91 67.72 1.08 ;
        RECT 67.55 2.39 67.72 2.56 ;
      LAYER li1 ;
        RECT 67.555 0.915 67.725 1.085 ;
        RECT 67.55 0.57 67.72 1.08 ;
        RECT 67.55 2.39 67.72 3.86 ;
      LAYER met1 ;
        RECT 67.49 2.36 67.78 2.59 ;
        RECT 67.49 0.88 67.78 1.11 ;
        RECT 67.55 0.88 67.72 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 83.88 0.915 84.05 1.085 ;
        RECT 83.875 0.91 84.045 1.08 ;
        RECT 83.875 2.39 84.045 2.56 ;
      LAYER li1 ;
        RECT 83.88 0.915 84.05 1.085 ;
        RECT 83.875 0.57 84.045 1.08 ;
        RECT 83.875 2.39 84.045 3.86 ;
      LAYER met1 ;
        RECT 83.815 2.36 84.105 2.59 ;
        RECT 83.815 0.88 84.105 1.11 ;
        RECT 83.875 0.88 84.045 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 14.425 1.66 14.595 2.935 ;
        RECT 14.425 5.945 14.595 7.22 ;
        RECT 8.81 5.945 8.98 7.22 ;
      LAYER met2 ;
        RECT 14.35 2.705 14.69 3.055 ;
        RECT 14.34 5.84 14.68 6.19 ;
        RECT 14.425 2.705 14.595 6.19 ;
      LAYER met1 ;
        RECT 14.35 2.765 14.825 2.935 ;
        RECT 14.35 2.705 14.69 3.055 ;
        RECT 8.75 5.945 14.825 6.115 ;
        RECT 14.34 5.84 14.68 6.19 ;
        RECT 8.75 5.915 9.04 6.145 ;
      LAYER mcon ;
        RECT 8.81 5.945 8.98 6.115 ;
        RECT 14.425 5.945 14.595 6.115 ;
        RECT 14.425 2.765 14.595 2.935 ;
      LAYER via1 ;
        RECT 14.44 5.94 14.59 6.09 ;
        RECT 14.45 2.805 14.6 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 30.75 1.66 30.92 2.935 ;
        RECT 30.75 5.945 30.92 7.22 ;
        RECT 25.135 5.945 25.305 7.22 ;
      LAYER met2 ;
        RECT 30.675 2.705 31.015 3.055 ;
        RECT 30.665 5.84 31.005 6.19 ;
        RECT 30.75 2.705 30.92 6.19 ;
      LAYER met1 ;
        RECT 30.675 2.765 31.15 2.935 ;
        RECT 30.675 2.705 31.015 3.055 ;
        RECT 25.075 5.945 31.15 6.115 ;
        RECT 30.665 5.84 31.005 6.19 ;
        RECT 25.075 5.915 25.365 6.145 ;
      LAYER mcon ;
        RECT 25.135 5.945 25.305 6.115 ;
        RECT 30.75 5.945 30.92 6.115 ;
        RECT 30.75 2.765 30.92 2.935 ;
      LAYER via1 ;
        RECT 30.765 5.94 30.915 6.09 ;
        RECT 30.775 2.805 30.925 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 47.075 1.66 47.245 2.935 ;
        RECT 47.075 5.945 47.245 7.22 ;
        RECT 41.46 5.945 41.63 7.22 ;
      LAYER met2 ;
        RECT 47 2.705 47.34 3.055 ;
        RECT 46.99 5.84 47.33 6.19 ;
        RECT 47.075 2.705 47.245 6.19 ;
      LAYER met1 ;
        RECT 47 2.765 47.475 2.935 ;
        RECT 47 2.705 47.34 3.055 ;
        RECT 41.4 5.945 47.475 6.115 ;
        RECT 46.99 5.84 47.33 6.19 ;
        RECT 41.4 5.915 41.69 6.145 ;
      LAYER mcon ;
        RECT 41.46 5.945 41.63 6.115 ;
        RECT 47.075 5.945 47.245 6.115 ;
        RECT 47.075 2.765 47.245 2.935 ;
      LAYER via1 ;
        RECT 47.09 5.94 47.24 6.09 ;
        RECT 47.1 2.805 47.25 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 63.4 1.66 63.57 2.935 ;
        RECT 63.4 5.945 63.57 7.22 ;
        RECT 57.785 5.945 57.955 7.22 ;
      LAYER met2 ;
        RECT 63.325 2.705 63.665 3.055 ;
        RECT 63.315 5.84 63.655 6.19 ;
        RECT 63.4 2.705 63.57 6.19 ;
      LAYER met1 ;
        RECT 63.325 2.765 63.8 2.935 ;
        RECT 63.325 2.705 63.665 3.055 ;
        RECT 57.725 5.945 63.8 6.115 ;
        RECT 63.315 5.84 63.655 6.19 ;
        RECT 57.725 5.915 58.015 6.145 ;
      LAYER mcon ;
        RECT 57.785 5.945 57.955 6.115 ;
        RECT 63.4 5.945 63.57 6.115 ;
        RECT 63.4 2.765 63.57 2.935 ;
      LAYER via1 ;
        RECT 63.415 5.94 63.565 6.09 ;
        RECT 63.425 2.805 63.575 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 79.725 1.66 79.895 2.935 ;
        RECT 79.725 5.945 79.895 7.22 ;
        RECT 74.11 5.945 74.28 7.22 ;
      LAYER met2 ;
        RECT 79.65 2.705 79.99 3.055 ;
        RECT 79.64 5.84 79.98 6.19 ;
        RECT 79.725 2.705 79.895 6.19 ;
      LAYER met1 ;
        RECT 79.65 2.765 80.125 2.935 ;
        RECT 79.65 2.705 79.99 3.055 ;
        RECT 74.05 5.945 80.125 6.115 ;
        RECT 79.64 5.84 79.98 6.19 ;
        RECT 74.05 5.915 74.34 6.145 ;
      LAYER mcon ;
        RECT 74.11 5.945 74.28 6.115 ;
        RECT 79.725 5.945 79.895 6.115 ;
        RECT 79.725 2.765 79.895 2.935 ;
      LAYER via1 ;
        RECT 79.74 5.94 79.89 6.09 ;
        RECT 79.75 2.805 79.9 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 5.945 0.4 7.22 ;
      LAYER met1 ;
        RECT 0.17 5.945 0.63 6.115 ;
        RECT 0.17 5.915 0.46 6.145 ;
      LAYER mcon ;
        RECT 0.23 5.945 0.4 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.41 4.255 2.215 4.635 ;
      LAYER li1 ;
        RECT 0 4.44 84.42 4.745 ;
        RECT 1.875 4.135 84.42 4.745 ;
        RECT 82.285 4.13 84.265 4.75 ;
        RECT 83.445 3.4 83.615 5.48 ;
        RECT 82.455 3.4 82.625 5.48 ;
        RECT 79.715 3.405 79.885 5.475 ;
        RECT 77.925 3.635 78.095 4.745 ;
        RECT 76.965 3.635 77.135 4.745 ;
        RECT 74.525 3.635 74.695 4.745 ;
        RECT 74.1 4.135 74.27 5.475 ;
        RECT 73.525 3.635 73.695 4.745 ;
        RECT 72.565 3.635 72.735 4.745 ;
        RECT 70.125 3.635 70.295 4.745 ;
        RECT 65.96 4.13 67.94 4.75 ;
        RECT 67.12 3.4 67.29 5.48 ;
        RECT 66.13 3.4 66.3 5.48 ;
        RECT 63.39 3.405 63.56 5.475 ;
        RECT 61.6 3.635 61.77 4.745 ;
        RECT 60.64 3.635 60.81 4.745 ;
        RECT 58.2 3.635 58.37 4.745 ;
        RECT 57.775 4.135 57.945 5.475 ;
        RECT 57.2 3.635 57.37 4.745 ;
        RECT 56.24 3.635 56.41 4.745 ;
        RECT 53.8 3.635 53.97 4.745 ;
        RECT 49.635 4.13 51.615 4.75 ;
        RECT 50.795 3.4 50.965 5.48 ;
        RECT 49.805 3.4 49.975 5.48 ;
        RECT 47.065 3.405 47.235 5.475 ;
        RECT 45.275 3.635 45.445 4.745 ;
        RECT 44.315 3.635 44.485 4.745 ;
        RECT 41.875 3.635 42.045 4.745 ;
        RECT 41.45 4.135 41.62 5.475 ;
        RECT 40.875 3.635 41.045 4.745 ;
        RECT 39.915 3.635 40.085 4.745 ;
        RECT 37.475 3.635 37.645 4.745 ;
        RECT 33.31 4.13 35.29 4.75 ;
        RECT 34.47 3.4 34.64 5.48 ;
        RECT 33.48 3.4 33.65 5.48 ;
        RECT 30.74 3.405 30.91 5.475 ;
        RECT 28.95 3.635 29.12 4.745 ;
        RECT 27.99 3.635 28.16 4.745 ;
        RECT 25.55 3.635 25.72 4.745 ;
        RECT 25.125 4.135 25.295 5.475 ;
        RECT 24.55 3.635 24.72 4.745 ;
        RECT 23.59 3.635 23.76 4.745 ;
        RECT 21.15 3.635 21.32 4.745 ;
        RECT 16.985 4.13 18.965 4.75 ;
        RECT 18.145 3.4 18.315 5.48 ;
        RECT 17.155 3.4 17.325 5.48 ;
        RECT 14.415 3.405 14.585 5.475 ;
        RECT 12.625 3.635 12.795 4.745 ;
        RECT 11.665 3.635 11.835 4.745 ;
        RECT 9.225 3.635 9.395 4.745 ;
        RECT 8.8 4.135 8.97 5.475 ;
        RECT 8.225 3.635 8.395 4.745 ;
        RECT 7.265 3.635 7.435 4.745 ;
        RECT 4.825 3.635 4.995 4.745 ;
        RECT 2.03 4.135 2.2 8.305 ;
        RECT 0 4.135 84.42 4.33 ;
        RECT 0 4.135 1.705 4.745 ;
        RECT 0.22 4.135 0.39 5.475 ;
      LAYER met2 ;
        RECT 1.6 4.255 1.98 4.635 ;
      LAYER met1 ;
        RECT 0 4.135 84.42 4.745 ;
        RECT 82.285 4.13 84.265 4.75 ;
        RECT 68.835 3.98 78.495 4.745 ;
        RECT 65.96 4.13 67.94 4.75 ;
        RECT 52.51 3.98 62.17 4.745 ;
        RECT 49.635 4.13 51.615 4.75 ;
        RECT 36.185 3.98 45.845 4.745 ;
        RECT 33.31 4.13 35.29 4.75 ;
        RECT 19.86 3.98 29.52 4.745 ;
        RECT 16.985 4.13 18.965 4.75 ;
        RECT 3.535 3.98 13.195 4.745 ;
        RECT 1.97 6.655 2.26 6.885 ;
        RECT 1.8 6.685 2.26 6.855 ;
      LAYER via2 ;
        RECT 1.69 4.345 1.89 4.545 ;
      LAYER mcon ;
        RECT 2.03 6.685 2.2 6.855 ;
        RECT 2.34 4.545 2.51 4.715 ;
        RECT 3.68 4.135 3.85 4.305 ;
        RECT 4.14 4.135 4.31 4.305 ;
        RECT 4.6 4.135 4.77 4.305 ;
        RECT 5.06 4.135 5.23 4.305 ;
        RECT 5.52 4.135 5.69 4.305 ;
        RECT 5.98 4.135 6.15 4.305 ;
        RECT 6.44 4.135 6.61 4.305 ;
        RECT 6.9 4.135 7.07 4.305 ;
        RECT 7.36 4.135 7.53 4.305 ;
        RECT 7.82 4.135 7.99 4.305 ;
        RECT 8.28 4.135 8.45 4.305 ;
        RECT 8.74 4.135 8.91 4.305 ;
        RECT 9.2 4.135 9.37 4.305 ;
        RECT 9.66 4.135 9.83 4.305 ;
        RECT 10.12 4.135 10.29 4.305 ;
        RECT 10.58 4.135 10.75 4.305 ;
        RECT 10.92 4.545 11.09 4.715 ;
        RECT 11.04 4.135 11.21 4.305 ;
        RECT 11.5 4.135 11.67 4.305 ;
        RECT 11.96 4.135 12.13 4.305 ;
        RECT 12.42 4.135 12.59 4.305 ;
        RECT 12.88 4.135 13.05 4.305 ;
        RECT 16.535 4.545 16.705 4.715 ;
        RECT 16.535 4.165 16.705 4.335 ;
        RECT 17.235 4.55 17.405 4.72 ;
        RECT 17.235 4.16 17.405 4.33 ;
        RECT 18.225 4.55 18.395 4.72 ;
        RECT 18.225 4.16 18.395 4.33 ;
        RECT 20.005 4.135 20.175 4.305 ;
        RECT 20.465 4.135 20.635 4.305 ;
        RECT 20.925 4.135 21.095 4.305 ;
        RECT 21.385 4.135 21.555 4.305 ;
        RECT 21.845 4.135 22.015 4.305 ;
        RECT 22.305 4.135 22.475 4.305 ;
        RECT 22.765 4.135 22.935 4.305 ;
        RECT 23.225 4.135 23.395 4.305 ;
        RECT 23.685 4.135 23.855 4.305 ;
        RECT 24.145 4.135 24.315 4.305 ;
        RECT 24.605 4.135 24.775 4.305 ;
        RECT 25.065 4.135 25.235 4.305 ;
        RECT 25.525 4.135 25.695 4.305 ;
        RECT 25.985 4.135 26.155 4.305 ;
        RECT 26.445 4.135 26.615 4.305 ;
        RECT 26.905 4.135 27.075 4.305 ;
        RECT 27.245 4.545 27.415 4.715 ;
        RECT 27.365 4.135 27.535 4.305 ;
        RECT 27.825 4.135 27.995 4.305 ;
        RECT 28.285 4.135 28.455 4.305 ;
        RECT 28.745 4.135 28.915 4.305 ;
        RECT 29.205 4.135 29.375 4.305 ;
        RECT 32.86 4.545 33.03 4.715 ;
        RECT 32.86 4.165 33.03 4.335 ;
        RECT 33.56 4.55 33.73 4.72 ;
        RECT 33.56 4.16 33.73 4.33 ;
        RECT 34.55 4.55 34.72 4.72 ;
        RECT 34.55 4.16 34.72 4.33 ;
        RECT 36.33 4.135 36.5 4.305 ;
        RECT 36.79 4.135 36.96 4.305 ;
        RECT 37.25 4.135 37.42 4.305 ;
        RECT 37.71 4.135 37.88 4.305 ;
        RECT 38.17 4.135 38.34 4.305 ;
        RECT 38.63 4.135 38.8 4.305 ;
        RECT 39.09 4.135 39.26 4.305 ;
        RECT 39.55 4.135 39.72 4.305 ;
        RECT 40.01 4.135 40.18 4.305 ;
        RECT 40.47 4.135 40.64 4.305 ;
        RECT 40.93 4.135 41.1 4.305 ;
        RECT 41.39 4.135 41.56 4.305 ;
        RECT 41.85 4.135 42.02 4.305 ;
        RECT 42.31 4.135 42.48 4.305 ;
        RECT 42.77 4.135 42.94 4.305 ;
        RECT 43.23 4.135 43.4 4.305 ;
        RECT 43.57 4.545 43.74 4.715 ;
        RECT 43.69 4.135 43.86 4.305 ;
        RECT 44.15 4.135 44.32 4.305 ;
        RECT 44.61 4.135 44.78 4.305 ;
        RECT 45.07 4.135 45.24 4.305 ;
        RECT 45.53 4.135 45.7 4.305 ;
        RECT 49.185 4.545 49.355 4.715 ;
        RECT 49.185 4.165 49.355 4.335 ;
        RECT 49.885 4.55 50.055 4.72 ;
        RECT 49.885 4.16 50.055 4.33 ;
        RECT 50.875 4.55 51.045 4.72 ;
        RECT 50.875 4.16 51.045 4.33 ;
        RECT 52.655 4.135 52.825 4.305 ;
        RECT 53.115 4.135 53.285 4.305 ;
        RECT 53.575 4.135 53.745 4.305 ;
        RECT 54.035 4.135 54.205 4.305 ;
        RECT 54.495 4.135 54.665 4.305 ;
        RECT 54.955 4.135 55.125 4.305 ;
        RECT 55.415 4.135 55.585 4.305 ;
        RECT 55.875 4.135 56.045 4.305 ;
        RECT 56.335 4.135 56.505 4.305 ;
        RECT 56.795 4.135 56.965 4.305 ;
        RECT 57.255 4.135 57.425 4.305 ;
        RECT 57.715 4.135 57.885 4.305 ;
        RECT 58.175 4.135 58.345 4.305 ;
        RECT 58.635 4.135 58.805 4.305 ;
        RECT 59.095 4.135 59.265 4.305 ;
        RECT 59.555 4.135 59.725 4.305 ;
        RECT 59.895 4.545 60.065 4.715 ;
        RECT 60.015 4.135 60.185 4.305 ;
        RECT 60.475 4.135 60.645 4.305 ;
        RECT 60.935 4.135 61.105 4.305 ;
        RECT 61.395 4.135 61.565 4.305 ;
        RECT 61.855 4.135 62.025 4.305 ;
        RECT 65.51 4.545 65.68 4.715 ;
        RECT 65.51 4.165 65.68 4.335 ;
        RECT 66.21 4.55 66.38 4.72 ;
        RECT 66.21 4.16 66.38 4.33 ;
        RECT 67.2 4.55 67.37 4.72 ;
        RECT 67.2 4.16 67.37 4.33 ;
        RECT 68.98 4.135 69.15 4.305 ;
        RECT 69.44 4.135 69.61 4.305 ;
        RECT 69.9 4.135 70.07 4.305 ;
        RECT 70.36 4.135 70.53 4.305 ;
        RECT 70.82 4.135 70.99 4.305 ;
        RECT 71.28 4.135 71.45 4.305 ;
        RECT 71.74 4.135 71.91 4.305 ;
        RECT 72.2 4.135 72.37 4.305 ;
        RECT 72.66 4.135 72.83 4.305 ;
        RECT 73.12 4.135 73.29 4.305 ;
        RECT 73.58 4.135 73.75 4.305 ;
        RECT 74.04 4.135 74.21 4.305 ;
        RECT 74.5 4.135 74.67 4.305 ;
        RECT 74.96 4.135 75.13 4.305 ;
        RECT 75.42 4.135 75.59 4.305 ;
        RECT 75.88 4.135 76.05 4.305 ;
        RECT 76.22 4.545 76.39 4.715 ;
        RECT 76.34 4.135 76.51 4.305 ;
        RECT 76.8 4.135 76.97 4.305 ;
        RECT 77.26 4.135 77.43 4.305 ;
        RECT 77.72 4.135 77.89 4.305 ;
        RECT 78.18 4.135 78.35 4.305 ;
        RECT 81.835 4.545 82.005 4.715 ;
        RECT 81.835 4.165 82.005 4.335 ;
        RECT 82.535 4.55 82.705 4.72 ;
        RECT 82.535 4.16 82.705 4.33 ;
        RECT 83.525 4.55 83.695 4.72 ;
        RECT 83.525 4.16 83.695 4.33 ;
      LAYER via1 ;
        RECT 1.715 4.37 1.865 4.52 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 77.725 2.975 78.055 3.705 ;
        RECT 61.4 2.975 61.73 3.705 ;
        RECT 45.075 2.975 45.405 3.705 ;
        RECT 28.75 2.975 29.08 3.705 ;
        RECT 12.425 2.975 12.755 3.705 ;
        RECT 0.005 8.5 0.81 8.88 ;
        RECT 0 0 0.805 0.38 ;
      LAYER li1 ;
        RECT 84.24 0 84.42 0.305 ;
        RECT 0.465 0 84.42 0.3 ;
        RECT 83.445 0 83.615 0.93 ;
        RECT 82.455 0 82.625 0.93 ;
        RECT 67.915 0 82.29 0.305 ;
        RECT 79.715 0 79.885 0.935 ;
        RECT 68.835 0 78.65 1.585 ;
        RECT 76.965 0 77.135 2.085 ;
        RECT 75.005 0 75.175 2.085 ;
        RECT 74.935 0 75.175 1.595 ;
        RECT 73.385 0 73.58 1.595 ;
        RECT 72.565 0 72.735 2.085 ;
        RECT 71.605 0 71.775 2.085 ;
        RECT 71.26 0 71.455 1.595 ;
        RECT 71.085 0 71.255 2.085 ;
        RECT 70.125 0 70.295 2.085 ;
        RECT 69.165 0 69.335 2.085 ;
        RECT 68.96 0 69.155 1.595 ;
        RECT 67.12 0 67.29 0.93 ;
        RECT 66.13 0 66.3 0.93 ;
        RECT 51.59 0 65.965 0.305 ;
        RECT 63.39 0 63.56 0.935 ;
        RECT 52.51 0 62.325 1.585 ;
        RECT 60.64 0 60.81 2.085 ;
        RECT 58.68 0 58.85 2.085 ;
        RECT 58.61 0 58.85 1.595 ;
        RECT 57.06 0 57.255 1.595 ;
        RECT 56.24 0 56.41 2.085 ;
        RECT 55.28 0 55.45 2.085 ;
        RECT 54.935 0 55.13 1.595 ;
        RECT 54.76 0 54.93 2.085 ;
        RECT 53.8 0 53.97 2.085 ;
        RECT 52.84 0 53.01 2.085 ;
        RECT 52.635 0 52.83 1.595 ;
        RECT 50.795 0 50.965 0.93 ;
        RECT 49.805 0 49.975 0.93 ;
        RECT 35.265 0 49.64 0.305 ;
        RECT 47.065 0 47.235 0.935 ;
        RECT 36.185 0 46 1.585 ;
        RECT 44.315 0 44.485 2.085 ;
        RECT 42.355 0 42.525 2.085 ;
        RECT 42.285 0 42.525 1.595 ;
        RECT 40.735 0 40.93 1.595 ;
        RECT 39.915 0 40.085 2.085 ;
        RECT 38.955 0 39.125 2.085 ;
        RECT 38.61 0 38.805 1.595 ;
        RECT 38.435 0 38.605 2.085 ;
        RECT 37.475 0 37.645 2.085 ;
        RECT 36.515 0 36.685 2.085 ;
        RECT 36.31 0 36.505 1.595 ;
        RECT 34.47 0 34.64 0.93 ;
        RECT 33.48 0 33.65 0.93 ;
        RECT 18.94 0 33.315 0.305 ;
        RECT 30.74 0 30.91 0.935 ;
        RECT 19.86 0 29.675 1.585 ;
        RECT 27.99 0 28.16 2.085 ;
        RECT 26.03 0 26.2 2.085 ;
        RECT 25.96 0 26.2 1.595 ;
        RECT 24.41 0 24.605 1.595 ;
        RECT 23.59 0 23.76 2.085 ;
        RECT 22.63 0 22.8 2.085 ;
        RECT 22.285 0 22.48 1.595 ;
        RECT 22.11 0 22.28 2.085 ;
        RECT 21.15 0 21.32 2.085 ;
        RECT 20.19 0 20.36 2.085 ;
        RECT 19.985 0 20.18 1.595 ;
        RECT 18.145 0 18.315 0.93 ;
        RECT 17.155 0 17.325 0.93 ;
        RECT 0 0.245 16.99 0.305 ;
        RECT 14.415 0 14.585 0.935 ;
        RECT 3.535 0 13.35 1.585 ;
        RECT 11.665 0 11.835 2.085 ;
        RECT 9.705 0 9.875 2.085 ;
        RECT 9.635 0 9.875 1.595 ;
        RECT 8.085 0 8.28 1.595 ;
        RECT 7.265 0 7.435 2.085 ;
        RECT 6.305 0 6.475 2.085 ;
        RECT 5.96 0 6.155 1.595 ;
        RECT 5.785 0 5.955 2.085 ;
        RECT 4.825 0 4.995 2.085 ;
        RECT 3.865 0 4.035 2.085 ;
        RECT 3.66 0 3.855 1.595 ;
        RECT 0 0.245 0.805 0.315 ;
        RECT 0.295 0.245 0.465 0.335 ;
        RECT 0 0 84.42 0.075 ;
        RECT 0 0 0.295 0.315 ;
        RECT 0 8.58 84.42 8.88 ;
        RECT 84.24 8.575 84.42 8.88 ;
        RECT 83.445 7.95 83.615 8.88 ;
        RECT 82.455 7.95 82.625 8.88 ;
        RECT 67.915 8.575 82.29 8.88 ;
        RECT 79.715 7.945 79.885 8.88 ;
        RECT 74.1 7.945 74.27 8.88 ;
        RECT 67.12 7.95 67.29 8.88 ;
        RECT 66.13 7.95 66.3 8.88 ;
        RECT 51.59 8.575 65.965 8.88 ;
        RECT 63.39 7.945 63.56 8.88 ;
        RECT 57.775 7.945 57.945 8.88 ;
        RECT 50.795 7.95 50.965 8.88 ;
        RECT 49.805 7.95 49.975 8.88 ;
        RECT 35.265 8.575 49.64 8.88 ;
        RECT 47.065 7.945 47.235 8.88 ;
        RECT 41.45 7.945 41.62 8.88 ;
        RECT 34.47 7.95 34.64 8.88 ;
        RECT 33.48 7.95 33.65 8.88 ;
        RECT 18.94 8.575 33.315 8.88 ;
        RECT 30.74 7.945 30.91 8.88 ;
        RECT 25.125 7.945 25.295 8.88 ;
        RECT 18.145 7.95 18.315 8.88 ;
        RECT 17.155 7.95 17.325 8.88 ;
        RECT 0 8.575 16.99 8.88 ;
        RECT 14.415 7.945 14.585 8.88 ;
        RECT 8.8 7.945 8.97 8.88 ;
        RECT 0.005 8.565 0.81 8.88 ;
        RECT 0.22 8.545 0.47 8.88 ;
        RECT 0.22 7.945 0.39 8.88 ;
        RECT 77.925 2.575 78.095 2.945 ;
        RECT 77.605 2.575 78.095 2.745 ;
        RECT 75.965 2.575 76.135 2.945 ;
        RECT 75.645 2.575 76.135 2.745 ;
        RECT 75.105 6.075 75.275 8.025 ;
        RECT 75.05 7.855 75.22 8.305 ;
        RECT 75.05 5.015 75.22 6.245 ;
        RECT 61.6 2.575 61.77 2.945 ;
        RECT 61.28 2.575 61.77 2.745 ;
        RECT 59.64 2.575 59.81 2.945 ;
        RECT 59.32 2.575 59.81 2.745 ;
        RECT 58.78 6.075 58.95 8.025 ;
        RECT 58.725 7.855 58.895 8.305 ;
        RECT 58.725 5.015 58.895 6.245 ;
        RECT 45.275 2.575 45.445 2.945 ;
        RECT 44.955 2.575 45.445 2.745 ;
        RECT 43.315 2.575 43.485 2.945 ;
        RECT 42.995 2.575 43.485 2.745 ;
        RECT 42.455 6.075 42.625 8.025 ;
        RECT 42.4 7.855 42.57 8.305 ;
        RECT 42.4 5.015 42.57 6.245 ;
        RECT 28.95 2.575 29.12 2.945 ;
        RECT 28.63 2.575 29.12 2.745 ;
        RECT 26.99 2.575 27.16 2.945 ;
        RECT 26.67 2.575 27.16 2.745 ;
        RECT 26.13 6.075 26.3 8.025 ;
        RECT 26.075 7.855 26.245 8.305 ;
        RECT 26.075 5.015 26.245 6.245 ;
        RECT 12.625 2.575 12.795 2.945 ;
        RECT 12.305 2.575 12.795 2.745 ;
        RECT 10.665 2.575 10.835 2.945 ;
        RECT 10.345 2.575 10.835 2.745 ;
        RECT 9.805 6.075 9.975 8.025 ;
        RECT 9.75 7.855 9.92 8.305 ;
        RECT 9.75 5.015 9.92 6.245 ;
      LAYER met2 ;
        RECT 77.75 2.955 78.03 3.325 ;
        RECT 77.76 2.7 78.02 3.325 ;
        RECT 61.425 2.955 61.705 3.325 ;
        RECT 61.435 2.7 61.695 3.325 ;
        RECT 45.1 2.955 45.38 3.325 ;
        RECT 45.11 2.7 45.37 3.325 ;
        RECT 28.775 2.955 29.055 3.325 ;
        RECT 28.785 2.7 29.045 3.325 ;
        RECT 12.45 2.955 12.73 3.325 ;
        RECT 12.46 2.7 12.72 3.325 ;
        RECT 0.195 8.5 0.575 8.88 ;
        RECT 0.19 0 0.57 0.38 ;
        RECT 0.235 0 0.375 8.88 ;
      LAYER met1 ;
        RECT 84.24 0 84.42 0.305 ;
        RECT 0 0 84.42 0.3 ;
        RECT 67.915 0 82.29 0.305 ;
        RECT 78.465 0 78.65 2.945 ;
        RECT 77.7 2.79 78.65 2.945 ;
        RECT 77.73 2.76 78.65 2.945 ;
        RECT 68.835 0 78.65 1.74 ;
        RECT 77.73 2.745 78.155 2.975 ;
        RECT 77.73 2.73 78.05 2.99 ;
        RECT 76.24 2.93 78.005 3.055 ;
        RECT 76.24 2.93 77.84 3.07 ;
        RECT 75.905 2.79 76.38 2.975 ;
        RECT 75.905 2.745 76.195 2.975 ;
        RECT 51.59 0 65.965 0.305 ;
        RECT 62.14 0 62.325 2.945 ;
        RECT 61.375 2.79 62.325 2.945 ;
        RECT 61.405 2.76 62.325 2.945 ;
        RECT 52.51 0 62.325 1.74 ;
        RECT 61.405 2.745 61.83 2.975 ;
        RECT 61.405 2.73 61.725 2.99 ;
        RECT 59.915 2.93 61.68 3.055 ;
        RECT 59.915 2.93 61.515 3.07 ;
        RECT 59.58 2.79 60.055 2.975 ;
        RECT 59.58 2.745 59.87 2.975 ;
        RECT 35.265 0 49.64 0.305 ;
        RECT 45.815 0 46 2.945 ;
        RECT 45.05 2.79 46 2.945 ;
        RECT 45.08 2.76 46 2.945 ;
        RECT 36.185 0 46 1.74 ;
        RECT 45.08 2.745 45.505 2.975 ;
        RECT 45.08 2.73 45.4 2.99 ;
        RECT 43.59 2.93 45.355 3.055 ;
        RECT 43.59 2.93 45.19 3.07 ;
        RECT 43.255 2.79 43.73 2.975 ;
        RECT 43.255 2.745 43.545 2.975 ;
        RECT 18.94 0 33.315 0.305 ;
        RECT 29.49 0 29.675 2.945 ;
        RECT 28.725 2.79 29.675 2.945 ;
        RECT 28.755 2.76 29.675 2.945 ;
        RECT 19.86 0 29.675 1.74 ;
        RECT 28.755 2.745 29.18 2.975 ;
        RECT 28.755 2.73 29.075 2.99 ;
        RECT 27.265 2.93 29.03 3.055 ;
        RECT 27.265 2.93 28.865 3.07 ;
        RECT 26.93 2.79 27.405 2.975 ;
        RECT 26.93 2.745 27.22 2.975 ;
        RECT 0 0 16.99 0.305 ;
        RECT 13.165 0 13.35 2.945 ;
        RECT 12.4 2.79 13.35 2.945 ;
        RECT 12.43 2.76 13.35 2.945 ;
        RECT 3.535 0 13.35 1.74 ;
        RECT 12.43 2.745 12.855 2.975 ;
        RECT 12.43 2.73 12.75 2.99 ;
        RECT 10.94 2.93 12.705 3.055 ;
        RECT 10.94 2.93 12.54 3.07 ;
        RECT 10.605 2.79 11.08 2.975 ;
        RECT 10.605 2.745 10.895 2.975 ;
        RECT 0 0 0.805 0.315 ;
        RECT 0.205 0 0.555 0.335 ;
        RECT 0 8.58 84.42 8.88 ;
        RECT 84.24 8.575 84.42 8.88 ;
        RECT 67.915 8.575 82.29 8.88 ;
        RECT 75.045 6.285 75.335 6.515 ;
        RECT 74.67 6.315 75.335 6.485 ;
        RECT 74.67 6.315 74.845 8.88 ;
        RECT 51.59 8.575 65.965 8.88 ;
        RECT 58.72 6.285 59.01 6.515 ;
        RECT 58.345 6.315 59.01 6.485 ;
        RECT 58.345 6.315 58.52 8.88 ;
        RECT 35.265 8.575 49.64 8.88 ;
        RECT 42.395 6.285 42.685 6.515 ;
        RECT 42.02 6.315 42.685 6.485 ;
        RECT 42.02 6.315 42.195 8.88 ;
        RECT 18.94 8.575 33.315 8.88 ;
        RECT 26.07 6.285 26.36 6.515 ;
        RECT 25.695 6.315 26.36 6.485 ;
        RECT 25.695 6.315 25.87 8.88 ;
        RECT 0 8.575 16.99 8.88 ;
        RECT 9.745 6.285 10.035 6.515 ;
        RECT 9.37 6.315 10.035 6.485 ;
        RECT 9.37 6.315 9.545 8.88 ;
        RECT 0.005 8.565 0.81 8.88 ;
        RECT 0.21 8.545 0.56 8.88 ;
      LAYER via2 ;
        RECT 0.28 0.09 0.48 0.29 ;
        RECT 0.285 8.59 0.485 8.79 ;
        RECT 12.49 3.04 12.69 3.24 ;
        RECT 28.815 3.04 29.015 3.24 ;
        RECT 45.14 3.04 45.34 3.24 ;
        RECT 61.465 3.04 61.665 3.24 ;
        RECT 77.79 3.04 77.99 3.24 ;
      LAYER mcon ;
        RECT 0.3 8.605 0.47 8.775 ;
        RECT 0.98 8.605 1.15 8.775 ;
        RECT 1.66 8.605 1.83 8.775 ;
        RECT 2.34 8.605 2.51 8.775 ;
        RECT 3.68 1.415 3.85 1.585 ;
        RECT 4.14 1.415 4.31 1.585 ;
        RECT 4.6 1.415 4.77 1.585 ;
        RECT 5.06 1.415 5.23 1.585 ;
        RECT 5.52 1.415 5.69 1.585 ;
        RECT 5.98 1.415 6.15 1.585 ;
        RECT 6.44 1.415 6.61 1.585 ;
        RECT 6.9 1.415 7.07 1.585 ;
        RECT 7.36 1.415 7.53 1.585 ;
        RECT 7.82 1.415 7.99 1.585 ;
        RECT 8.28 1.415 8.45 1.585 ;
        RECT 8.74 1.415 8.91 1.585 ;
        RECT 8.88 8.605 9.05 8.775 ;
        RECT 9.2 1.415 9.37 1.585 ;
        RECT 9.56 8.605 9.73 8.775 ;
        RECT 9.66 1.415 9.83 1.585 ;
        RECT 9.805 6.315 9.975 6.485 ;
        RECT 10.12 1.415 10.29 1.585 ;
        RECT 10.24 8.605 10.41 8.775 ;
        RECT 10.58 1.415 10.75 1.585 ;
        RECT 10.665 2.775 10.835 2.945 ;
        RECT 10.92 8.605 11.09 8.775 ;
        RECT 11.04 1.415 11.21 1.585 ;
        RECT 11.5 1.415 11.67 1.585 ;
        RECT 11.96 1.415 12.13 1.585 ;
        RECT 12.42 1.415 12.59 1.585 ;
        RECT 12.625 2.775 12.795 2.945 ;
        RECT 12.88 1.415 13.05 1.585 ;
        RECT 14.495 8.605 14.665 8.775 ;
        RECT 14.495 0.105 14.665 0.275 ;
        RECT 15.175 8.605 15.345 8.775 ;
        RECT 15.175 0.105 15.345 0.275 ;
        RECT 15.855 8.605 16.025 8.775 ;
        RECT 15.855 0.105 16.025 0.275 ;
        RECT 16.535 8.605 16.705 8.775 ;
        RECT 16.535 0.105 16.705 0.275 ;
        RECT 17.235 8.61 17.405 8.78 ;
        RECT 17.235 0.1 17.405 0.27 ;
        RECT 18.225 8.61 18.395 8.78 ;
        RECT 18.225 0.1 18.395 0.27 ;
        RECT 20.005 1.415 20.175 1.585 ;
        RECT 20.465 1.415 20.635 1.585 ;
        RECT 20.925 1.415 21.095 1.585 ;
        RECT 21.385 1.415 21.555 1.585 ;
        RECT 21.845 1.415 22.015 1.585 ;
        RECT 22.305 1.415 22.475 1.585 ;
        RECT 22.765 1.415 22.935 1.585 ;
        RECT 23.225 1.415 23.395 1.585 ;
        RECT 23.685 1.415 23.855 1.585 ;
        RECT 24.145 1.415 24.315 1.585 ;
        RECT 24.605 1.415 24.775 1.585 ;
        RECT 25.065 1.415 25.235 1.585 ;
        RECT 25.205 8.605 25.375 8.775 ;
        RECT 25.525 1.415 25.695 1.585 ;
        RECT 25.885 8.605 26.055 8.775 ;
        RECT 25.985 1.415 26.155 1.585 ;
        RECT 26.13 6.315 26.3 6.485 ;
        RECT 26.445 1.415 26.615 1.585 ;
        RECT 26.565 8.605 26.735 8.775 ;
        RECT 26.905 1.415 27.075 1.585 ;
        RECT 26.99 2.775 27.16 2.945 ;
        RECT 27.245 8.605 27.415 8.775 ;
        RECT 27.365 1.415 27.535 1.585 ;
        RECT 27.825 1.415 27.995 1.585 ;
        RECT 28.285 1.415 28.455 1.585 ;
        RECT 28.745 1.415 28.915 1.585 ;
        RECT 28.95 2.775 29.12 2.945 ;
        RECT 29.205 1.415 29.375 1.585 ;
        RECT 30.82 8.605 30.99 8.775 ;
        RECT 30.82 0.105 30.99 0.275 ;
        RECT 31.5 8.605 31.67 8.775 ;
        RECT 31.5 0.105 31.67 0.275 ;
        RECT 32.18 8.605 32.35 8.775 ;
        RECT 32.18 0.105 32.35 0.275 ;
        RECT 32.86 8.605 33.03 8.775 ;
        RECT 32.86 0.105 33.03 0.275 ;
        RECT 33.56 8.61 33.73 8.78 ;
        RECT 33.56 0.1 33.73 0.27 ;
        RECT 34.55 8.61 34.72 8.78 ;
        RECT 34.55 0.1 34.72 0.27 ;
        RECT 36.33 1.415 36.5 1.585 ;
        RECT 36.79 1.415 36.96 1.585 ;
        RECT 37.25 1.415 37.42 1.585 ;
        RECT 37.71 1.415 37.88 1.585 ;
        RECT 38.17 1.415 38.34 1.585 ;
        RECT 38.63 1.415 38.8 1.585 ;
        RECT 39.09 1.415 39.26 1.585 ;
        RECT 39.55 1.415 39.72 1.585 ;
        RECT 40.01 1.415 40.18 1.585 ;
        RECT 40.47 1.415 40.64 1.585 ;
        RECT 40.93 1.415 41.1 1.585 ;
        RECT 41.39 1.415 41.56 1.585 ;
        RECT 41.53 8.605 41.7 8.775 ;
        RECT 41.85 1.415 42.02 1.585 ;
        RECT 42.21 8.605 42.38 8.775 ;
        RECT 42.31 1.415 42.48 1.585 ;
        RECT 42.455 6.315 42.625 6.485 ;
        RECT 42.77 1.415 42.94 1.585 ;
        RECT 42.89 8.605 43.06 8.775 ;
        RECT 43.23 1.415 43.4 1.585 ;
        RECT 43.315 2.775 43.485 2.945 ;
        RECT 43.57 8.605 43.74 8.775 ;
        RECT 43.69 1.415 43.86 1.585 ;
        RECT 44.15 1.415 44.32 1.585 ;
        RECT 44.61 1.415 44.78 1.585 ;
        RECT 45.07 1.415 45.24 1.585 ;
        RECT 45.275 2.775 45.445 2.945 ;
        RECT 45.53 1.415 45.7 1.585 ;
        RECT 47.145 8.605 47.315 8.775 ;
        RECT 47.145 0.105 47.315 0.275 ;
        RECT 47.825 8.605 47.995 8.775 ;
        RECT 47.825 0.105 47.995 0.275 ;
        RECT 48.505 8.605 48.675 8.775 ;
        RECT 48.505 0.105 48.675 0.275 ;
        RECT 49.185 8.605 49.355 8.775 ;
        RECT 49.185 0.105 49.355 0.275 ;
        RECT 49.885 8.61 50.055 8.78 ;
        RECT 49.885 0.1 50.055 0.27 ;
        RECT 50.875 8.61 51.045 8.78 ;
        RECT 50.875 0.1 51.045 0.27 ;
        RECT 52.655 1.415 52.825 1.585 ;
        RECT 53.115 1.415 53.285 1.585 ;
        RECT 53.575 1.415 53.745 1.585 ;
        RECT 54.035 1.415 54.205 1.585 ;
        RECT 54.495 1.415 54.665 1.585 ;
        RECT 54.955 1.415 55.125 1.585 ;
        RECT 55.415 1.415 55.585 1.585 ;
        RECT 55.875 1.415 56.045 1.585 ;
        RECT 56.335 1.415 56.505 1.585 ;
        RECT 56.795 1.415 56.965 1.585 ;
        RECT 57.255 1.415 57.425 1.585 ;
        RECT 57.715 1.415 57.885 1.585 ;
        RECT 57.855 8.605 58.025 8.775 ;
        RECT 58.175 1.415 58.345 1.585 ;
        RECT 58.535 8.605 58.705 8.775 ;
        RECT 58.635 1.415 58.805 1.585 ;
        RECT 58.78 6.315 58.95 6.485 ;
        RECT 59.095 1.415 59.265 1.585 ;
        RECT 59.215 8.605 59.385 8.775 ;
        RECT 59.555 1.415 59.725 1.585 ;
        RECT 59.64 2.775 59.81 2.945 ;
        RECT 59.895 8.605 60.065 8.775 ;
        RECT 60.015 1.415 60.185 1.585 ;
        RECT 60.475 1.415 60.645 1.585 ;
        RECT 60.935 1.415 61.105 1.585 ;
        RECT 61.395 1.415 61.565 1.585 ;
        RECT 61.6 2.775 61.77 2.945 ;
        RECT 61.855 1.415 62.025 1.585 ;
        RECT 63.47 8.605 63.64 8.775 ;
        RECT 63.47 0.105 63.64 0.275 ;
        RECT 64.15 8.605 64.32 8.775 ;
        RECT 64.15 0.105 64.32 0.275 ;
        RECT 64.83 8.605 65 8.775 ;
        RECT 64.83 0.105 65 0.275 ;
        RECT 65.51 8.605 65.68 8.775 ;
        RECT 65.51 0.105 65.68 0.275 ;
        RECT 66.21 8.61 66.38 8.78 ;
        RECT 66.21 0.1 66.38 0.27 ;
        RECT 67.2 8.61 67.37 8.78 ;
        RECT 67.2 0.1 67.37 0.27 ;
        RECT 68.98 1.415 69.15 1.585 ;
        RECT 69.44 1.415 69.61 1.585 ;
        RECT 69.9 1.415 70.07 1.585 ;
        RECT 70.36 1.415 70.53 1.585 ;
        RECT 70.82 1.415 70.99 1.585 ;
        RECT 71.28 1.415 71.45 1.585 ;
        RECT 71.74 1.415 71.91 1.585 ;
        RECT 72.2 1.415 72.37 1.585 ;
        RECT 72.66 1.415 72.83 1.585 ;
        RECT 73.12 1.415 73.29 1.585 ;
        RECT 73.58 1.415 73.75 1.585 ;
        RECT 74.04 1.415 74.21 1.585 ;
        RECT 74.18 8.605 74.35 8.775 ;
        RECT 74.5 1.415 74.67 1.585 ;
        RECT 74.86 8.605 75.03 8.775 ;
        RECT 74.96 1.415 75.13 1.585 ;
        RECT 75.105 6.315 75.275 6.485 ;
        RECT 75.42 1.415 75.59 1.585 ;
        RECT 75.54 8.605 75.71 8.775 ;
        RECT 75.88 1.415 76.05 1.585 ;
        RECT 75.965 2.775 76.135 2.945 ;
        RECT 76.22 8.605 76.39 8.775 ;
        RECT 76.34 1.415 76.51 1.585 ;
        RECT 76.8 1.415 76.97 1.585 ;
        RECT 77.26 1.415 77.43 1.585 ;
        RECT 77.72 1.415 77.89 1.585 ;
        RECT 77.925 2.775 78.095 2.945 ;
        RECT 78.18 1.415 78.35 1.585 ;
        RECT 79.795 8.605 79.965 8.775 ;
        RECT 79.795 0.105 79.965 0.275 ;
        RECT 80.475 8.605 80.645 8.775 ;
        RECT 80.475 0.105 80.645 0.275 ;
        RECT 81.155 8.605 81.325 8.775 ;
        RECT 81.155 0.105 81.325 0.275 ;
        RECT 81.835 8.605 82.005 8.775 ;
        RECT 81.835 0.105 82.005 0.275 ;
        RECT 82.535 8.61 82.705 8.78 ;
        RECT 82.535 0.1 82.705 0.27 ;
        RECT 83.525 8.61 83.695 8.78 ;
        RECT 83.525 0.1 83.695 0.27 ;
      LAYER via1 ;
        RECT 0.305 0.115 0.455 0.265 ;
        RECT 0.31 8.615 0.46 8.765 ;
        RECT 12.515 2.785 12.665 2.935 ;
        RECT 28.84 2.785 28.99 2.935 ;
        RECT 45.165 2.785 45.315 2.935 ;
        RECT 61.49 2.785 61.64 2.935 ;
        RECT 77.815 2.785 77.965 2.935 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 75.4 7.055 75.77 7.425 ;
      RECT 75.4 7.09 77.385 7.39 ;
      RECT 77.085 2.28 77.385 7.39 ;
      RECT 74.085 2.015 74.415 2.745 ;
      RECT 73.205 2.015 73.535 2.745 ;
      RECT 76.285 2.28 77.575 2.58 ;
      RECT 77.245 1.85 77.575 2.58 ;
      RECT 73.205 2.28 75.345 2.58 ;
      RECT 75.045 1.965 75.345 2.58 ;
      RECT 76.285 1.98 76.59 2.58 ;
      RECT 75.045 1.965 76.405 2.275 ;
      RECT 73.705 3.535 74.035 3.865 ;
      RECT 72.5 3.55 74.035 3.85 ;
      RECT 72.5 2.43 72.8 3.85 ;
      RECT 72.245 2.415 72.575 2.745 ;
      RECT 59.075 7.055 59.445 7.425 ;
      RECT 59.075 7.09 61.06 7.39 ;
      RECT 60.76 2.28 61.06 7.39 ;
      RECT 57.76 2.015 58.09 2.745 ;
      RECT 56.88 2.015 57.21 2.745 ;
      RECT 59.96 2.28 61.25 2.58 ;
      RECT 60.92 1.85 61.25 2.58 ;
      RECT 56.88 2.28 59.02 2.58 ;
      RECT 58.72 1.965 59.02 2.58 ;
      RECT 59.96 1.98 60.265 2.58 ;
      RECT 58.72 1.965 60.08 2.275 ;
      RECT 57.38 3.535 57.71 3.865 ;
      RECT 56.175 3.55 57.71 3.85 ;
      RECT 56.175 2.43 56.475 3.85 ;
      RECT 55.92 2.415 56.25 2.745 ;
      RECT 42.75 7.055 43.12 7.425 ;
      RECT 42.75 7.09 44.735 7.39 ;
      RECT 44.435 2.28 44.735 7.39 ;
      RECT 41.435 2.015 41.765 2.745 ;
      RECT 40.555 2.015 40.885 2.745 ;
      RECT 43.635 2.28 44.925 2.58 ;
      RECT 44.595 1.85 44.925 2.58 ;
      RECT 40.555 2.28 42.695 2.58 ;
      RECT 42.395 1.965 42.695 2.58 ;
      RECT 43.635 1.98 43.94 2.58 ;
      RECT 42.395 1.965 43.755 2.275 ;
      RECT 41.055 3.535 41.385 3.865 ;
      RECT 39.85 3.55 41.385 3.85 ;
      RECT 39.85 2.43 40.15 3.85 ;
      RECT 39.595 2.415 39.925 2.745 ;
      RECT 26.425 7.055 26.795 7.425 ;
      RECT 26.425 7.09 28.41 7.39 ;
      RECT 28.11 2.28 28.41 7.39 ;
      RECT 25.11 2.015 25.44 2.745 ;
      RECT 24.23 2.015 24.56 2.745 ;
      RECT 27.31 2.28 28.6 2.58 ;
      RECT 28.27 1.85 28.6 2.58 ;
      RECT 24.23 2.28 26.37 2.58 ;
      RECT 26.07 1.965 26.37 2.58 ;
      RECT 27.31 1.98 27.615 2.58 ;
      RECT 26.07 1.965 27.43 2.275 ;
      RECT 24.73 3.535 25.06 3.865 ;
      RECT 23.525 3.55 25.06 3.85 ;
      RECT 23.525 2.43 23.825 3.85 ;
      RECT 23.27 2.415 23.6 2.745 ;
      RECT 10.1 7.055 10.47 7.425 ;
      RECT 10.1 7.09 12.085 7.39 ;
      RECT 11.785 2.28 12.085 7.39 ;
      RECT 8.785 2.015 9.115 2.745 ;
      RECT 7.905 2.015 8.235 2.745 ;
      RECT 10.985 2.28 12.275 2.58 ;
      RECT 11.945 1.85 12.275 2.58 ;
      RECT 7.905 2.28 10.045 2.58 ;
      RECT 9.745 1.965 10.045 2.58 ;
      RECT 10.985 1.98 11.29 2.58 ;
      RECT 9.745 1.965 11.105 2.275 ;
      RECT 8.405 3.535 8.735 3.865 ;
      RECT 7.2 3.55 8.735 3.85 ;
      RECT 7.2 2.43 7.5 3.85 ;
      RECT 6.945 2.415 7.275 2.745 ;
      RECT 75.645 2.575 75.975 3.305 ;
      RECT 71.525 2.415 71.855 3.145 ;
      RECT 70.525 1.855 70.855 2.585 ;
      RECT 69.085 2.575 69.415 3.305 ;
      RECT 59.32 2.575 59.65 3.305 ;
      RECT 55.2 2.415 55.53 3.145 ;
      RECT 54.2 1.855 54.53 2.585 ;
      RECT 52.76 2.575 53.09 3.305 ;
      RECT 42.995 2.575 43.325 3.305 ;
      RECT 38.875 2.415 39.205 3.145 ;
      RECT 37.875 1.855 38.205 2.585 ;
      RECT 36.435 2.575 36.765 3.305 ;
      RECT 26.67 2.575 27 3.305 ;
      RECT 22.55 2.415 22.88 3.145 ;
      RECT 21.55 1.855 21.88 2.585 ;
      RECT 20.11 2.575 20.44 3.305 ;
      RECT 10.345 2.575 10.675 3.305 ;
      RECT 6.225 2.415 6.555 3.145 ;
      RECT 5.225 1.855 5.555 2.585 ;
      RECT 3.785 2.575 4.115 3.305 ;
    LAYER via2 ;
      RECT 77.31 2.315 77.51 2.515 ;
      RECT 75.71 3.04 75.91 3.24 ;
      RECT 75.485 7.14 75.685 7.34 ;
      RECT 74.15 2.48 74.35 2.68 ;
      RECT 73.77 3.6 73.97 3.8 ;
      RECT 73.27 2.48 73.47 2.68 ;
      RECT 72.31 2.48 72.51 2.68 ;
      RECT 71.59 2.48 71.79 2.68 ;
      RECT 70.59 1.92 70.79 2.12 ;
      RECT 69.15 3.04 69.35 3.24 ;
      RECT 60.985 2.315 61.185 2.515 ;
      RECT 59.385 3.04 59.585 3.24 ;
      RECT 59.16 7.14 59.36 7.34 ;
      RECT 57.825 2.48 58.025 2.68 ;
      RECT 57.445 3.6 57.645 3.8 ;
      RECT 56.945 2.48 57.145 2.68 ;
      RECT 55.985 2.48 56.185 2.68 ;
      RECT 55.265 2.48 55.465 2.68 ;
      RECT 54.265 1.92 54.465 2.12 ;
      RECT 52.825 3.04 53.025 3.24 ;
      RECT 44.66 2.315 44.86 2.515 ;
      RECT 43.06 3.04 43.26 3.24 ;
      RECT 42.835 7.14 43.035 7.34 ;
      RECT 41.5 2.48 41.7 2.68 ;
      RECT 41.12 3.6 41.32 3.8 ;
      RECT 40.62 2.48 40.82 2.68 ;
      RECT 39.66 2.48 39.86 2.68 ;
      RECT 38.94 2.48 39.14 2.68 ;
      RECT 37.94 1.92 38.14 2.12 ;
      RECT 36.5 3.04 36.7 3.24 ;
      RECT 28.335 2.315 28.535 2.515 ;
      RECT 26.735 3.04 26.935 3.24 ;
      RECT 26.51 7.14 26.71 7.34 ;
      RECT 25.175 2.48 25.375 2.68 ;
      RECT 24.795 3.6 24.995 3.8 ;
      RECT 24.295 2.48 24.495 2.68 ;
      RECT 23.335 2.48 23.535 2.68 ;
      RECT 22.615 2.48 22.815 2.68 ;
      RECT 21.615 1.92 21.815 2.12 ;
      RECT 20.175 3.04 20.375 3.24 ;
      RECT 12.01 2.315 12.21 2.515 ;
      RECT 10.41 3.04 10.61 3.24 ;
      RECT 10.185 7.14 10.385 7.34 ;
      RECT 8.85 2.48 9.05 2.68 ;
      RECT 8.47 3.6 8.67 3.8 ;
      RECT 7.97 2.48 8.17 2.68 ;
      RECT 7.01 2.48 7.21 2.68 ;
      RECT 6.29 2.48 6.49 2.68 ;
      RECT 5.29 1.92 5.49 2.12 ;
      RECT 3.85 3.04 4.05 3.24 ;
    LAYER met2 ;
      RECT 1.225 8.4 84.05 8.57 ;
      RECT 83.88 7.275 84.05 8.57 ;
      RECT 1.225 6.255 1.395 8.57 ;
      RECT 83.85 7.275 84.2 7.625 ;
      RECT 1.165 6.255 1.455 6.605 ;
      RECT 80.69 6.22 81.01 6.545 ;
      RECT 80.72 5.695 80.89 6.545 ;
      RECT 80.72 5.695 80.895 6.045 ;
      RECT 80.72 5.695 81.695 5.87 ;
      RECT 81.52 1.965 81.695 5.87 ;
      RECT 81.465 1.965 81.815 2.315 ;
      RECT 81.49 6.655 81.815 6.98 ;
      RECT 80.375 6.745 81.815 6.915 ;
      RECT 80.375 2.395 80.535 6.915 ;
      RECT 80.69 2.365 81.01 2.685 ;
      RECT 80.375 2.395 81.01 2.565 ;
      RECT 69.11 2.955 69.39 3.325 ;
      RECT 69.165 1.29 69.335 3.325 ;
      RECT 79.16 1.29 79.33 1.815 ;
      RECT 79.07 1.46 79.41 1.81 ;
      RECT 69.165 1.29 79.33 1.46 ;
      RECT 75.79 2.395 76.07 2.765 ;
      RECT 74.72 2.42 74.98 2.74 ;
      RECT 77.27 2.23 77.55 2.6 ;
      RECT 77.88 2.14 78.14 2.46 ;
      RECT 74.78 1.58 74.92 2.74 ;
      RECT 75.86 1.58 76 2.765 ;
      RECT 76.98 2.23 78.14 2.37 ;
      RECT 76.98 1.58 77.12 2.37 ;
      RECT 74.78 1.58 77.12 1.72 ;
      RECT 74.81 3.72 76.985 3.885 ;
      RECT 76.84 2.6 76.985 3.885 ;
      RECT 73.73 3.515 74.01 3.885 ;
      RECT 73.73 3.63 74.95 3.77 ;
      RECT 76.56 2.6 76.985 2.74 ;
      RECT 76.56 2.42 76.82 2.74 ;
      RECT 69.9 4 73.56 4.14 ;
      RECT 73.42 3.185 73.56 4.14 ;
      RECT 69.9 3.07 70.04 4.14 ;
      RECT 76.44 3.26 76.7 3.58 ;
      RECT 73.42 3.185 75.95 3.325 ;
      RECT 75.67 2.955 75.95 3.325 ;
      RECT 69.9 3.07 70.35 3.325 ;
      RECT 70.07 2.955 70.35 3.325 ;
      RECT 76.44 3.07 76.64 3.58 ;
      RECT 75.67 3.07 76.64 3.21 ;
      RECT 76.24 1.86 76.38 3.21 ;
      RECT 76.18 1.86 76.44 2.18 ;
      RECT 67.5 6.655 67.85 7.005 ;
      RECT 76.055 6.61 76.405 6.96 ;
      RECT 67.5 6.685 76.405 6.885 ;
      RECT 70.08 2.42 70.34 2.74 ;
      RECT 70.08 2.51 71.12 2.65 ;
      RECT 70.98 1.72 71.12 2.65 ;
      RECT 73.74 1.86 74 2.18 ;
      RECT 70.98 1.72 73.94 1.86 ;
      RECT 73.12 2.7 73.38 3.02 ;
      RECT 73.12 2.7 73.44 2.93 ;
      RECT 73.23 2.395 73.51 2.765 ;
      RECT 72.82 3.26 73.14 3.58 ;
      RECT 72.82 2.14 72.96 3.58 ;
      RECT 72.76 2.14 73.02 2.46 ;
      RECT 70.32 3.54 70.58 3.86 ;
      RECT 70.32 3.63 72 3.77 ;
      RECT 71.86 3.35 72 3.77 ;
      RECT 71.86 3.35 72.3 3.58 ;
      RECT 72.04 3.26 72.3 3.58 ;
      RECT 71.36 2.42 71.76 2.93 ;
      RECT 71.55 2.395 71.83 2.765 ;
      RECT 71.3 2.42 71.83 2.74 ;
      RECT 64.365 6.22 64.685 6.545 ;
      RECT 64.395 5.695 64.565 6.545 ;
      RECT 64.395 5.695 64.57 6.045 ;
      RECT 64.395 5.695 65.37 5.87 ;
      RECT 65.195 1.965 65.37 5.87 ;
      RECT 65.14 1.965 65.49 2.315 ;
      RECT 65.165 6.655 65.49 6.98 ;
      RECT 64.05 6.745 65.49 6.915 ;
      RECT 64.05 2.395 64.21 6.915 ;
      RECT 64.365 2.365 64.685 2.685 ;
      RECT 64.05 2.395 64.685 2.565 ;
      RECT 52.785 2.955 53.065 3.325 ;
      RECT 52.84 1.29 53.01 3.325 ;
      RECT 62.835 1.29 63.005 1.815 ;
      RECT 62.745 1.46 63.085 1.81 ;
      RECT 52.84 1.29 63.005 1.46 ;
      RECT 59.465 2.395 59.745 2.765 ;
      RECT 58.395 2.42 58.655 2.74 ;
      RECT 60.945 2.23 61.225 2.6 ;
      RECT 61.555 2.14 61.815 2.46 ;
      RECT 58.455 1.58 58.595 2.74 ;
      RECT 59.535 1.58 59.675 2.765 ;
      RECT 60.655 2.23 61.815 2.37 ;
      RECT 60.655 1.58 60.795 2.37 ;
      RECT 58.455 1.58 60.795 1.72 ;
      RECT 58.485 3.72 60.66 3.885 ;
      RECT 60.515 2.6 60.66 3.885 ;
      RECT 57.405 3.515 57.685 3.885 ;
      RECT 57.405 3.63 58.625 3.77 ;
      RECT 60.235 2.6 60.66 2.74 ;
      RECT 60.235 2.42 60.495 2.74 ;
      RECT 53.575 4 57.235 4.14 ;
      RECT 57.095 3.185 57.235 4.14 ;
      RECT 53.575 3.07 53.715 4.14 ;
      RECT 60.115 3.26 60.375 3.58 ;
      RECT 57.095 3.185 59.625 3.325 ;
      RECT 59.345 2.955 59.625 3.325 ;
      RECT 53.575 3.07 54.025 3.325 ;
      RECT 53.745 2.955 54.025 3.325 ;
      RECT 60.115 3.07 60.315 3.58 ;
      RECT 59.345 3.07 60.315 3.21 ;
      RECT 59.915 1.86 60.055 3.21 ;
      RECT 59.855 1.86 60.115 2.18 ;
      RECT 51.175 6.655 51.525 7.005 ;
      RECT 59.725 6.61 60.075 6.96 ;
      RECT 51.175 6.685 60.075 6.885 ;
      RECT 53.755 2.42 54.015 2.74 ;
      RECT 53.755 2.51 54.795 2.65 ;
      RECT 54.655 1.72 54.795 2.65 ;
      RECT 57.415 1.86 57.675 2.18 ;
      RECT 54.655 1.72 57.615 1.86 ;
      RECT 56.795 2.7 57.055 3.02 ;
      RECT 56.795 2.7 57.115 2.93 ;
      RECT 56.905 2.395 57.185 2.765 ;
      RECT 56.495 3.26 56.815 3.58 ;
      RECT 56.495 2.14 56.635 3.58 ;
      RECT 56.435 2.14 56.695 2.46 ;
      RECT 53.995 3.54 54.255 3.86 ;
      RECT 53.995 3.63 55.675 3.77 ;
      RECT 55.535 3.35 55.675 3.77 ;
      RECT 55.535 3.35 55.975 3.58 ;
      RECT 55.715 3.26 55.975 3.58 ;
      RECT 55.035 2.42 55.435 2.93 ;
      RECT 55.225 2.395 55.505 2.765 ;
      RECT 54.975 2.42 55.505 2.74 ;
      RECT 48.04 6.22 48.36 6.545 ;
      RECT 48.07 5.695 48.24 6.545 ;
      RECT 48.07 5.695 48.245 6.045 ;
      RECT 48.07 5.695 49.045 5.87 ;
      RECT 48.87 1.965 49.045 5.87 ;
      RECT 48.815 1.965 49.165 2.315 ;
      RECT 48.84 6.655 49.165 6.98 ;
      RECT 47.725 6.745 49.165 6.915 ;
      RECT 47.725 2.395 47.885 6.915 ;
      RECT 48.04 2.365 48.36 2.685 ;
      RECT 47.725 2.395 48.36 2.565 ;
      RECT 36.46 2.955 36.74 3.325 ;
      RECT 36.515 1.29 36.685 3.325 ;
      RECT 46.51 1.29 46.68 1.815 ;
      RECT 46.42 1.46 46.76 1.81 ;
      RECT 36.515 1.29 46.68 1.46 ;
      RECT 43.14 2.395 43.42 2.765 ;
      RECT 42.07 2.42 42.33 2.74 ;
      RECT 44.62 2.23 44.9 2.6 ;
      RECT 45.23 2.14 45.49 2.46 ;
      RECT 42.13 1.58 42.27 2.74 ;
      RECT 43.21 1.58 43.35 2.765 ;
      RECT 44.33 2.23 45.49 2.37 ;
      RECT 44.33 1.58 44.47 2.37 ;
      RECT 42.13 1.58 44.47 1.72 ;
      RECT 42.16 3.72 44.335 3.885 ;
      RECT 44.19 2.6 44.335 3.885 ;
      RECT 41.08 3.515 41.36 3.885 ;
      RECT 41.08 3.63 42.3 3.77 ;
      RECT 43.91 2.6 44.335 2.74 ;
      RECT 43.91 2.42 44.17 2.74 ;
      RECT 37.25 4 40.91 4.14 ;
      RECT 40.77 3.185 40.91 4.14 ;
      RECT 37.25 3.07 37.39 4.14 ;
      RECT 43.79 3.26 44.05 3.58 ;
      RECT 40.77 3.185 43.3 3.325 ;
      RECT 43.02 2.955 43.3 3.325 ;
      RECT 37.25 3.07 37.7 3.325 ;
      RECT 37.42 2.955 37.7 3.325 ;
      RECT 43.79 3.07 43.99 3.58 ;
      RECT 43.02 3.07 43.99 3.21 ;
      RECT 43.59 1.86 43.73 3.21 ;
      RECT 43.53 1.86 43.79 2.18 ;
      RECT 34.895 6.66 35.245 7.01 ;
      RECT 43.4 6.615 43.75 6.965 ;
      RECT 34.895 6.69 43.75 6.89 ;
      RECT 37.43 2.42 37.69 2.74 ;
      RECT 37.43 2.51 38.47 2.65 ;
      RECT 38.33 1.72 38.47 2.65 ;
      RECT 41.09 1.86 41.35 2.18 ;
      RECT 38.33 1.72 41.29 1.86 ;
      RECT 40.47 2.7 40.73 3.02 ;
      RECT 40.47 2.7 40.79 2.93 ;
      RECT 40.58 2.395 40.86 2.765 ;
      RECT 40.17 3.26 40.49 3.58 ;
      RECT 40.17 2.14 40.31 3.58 ;
      RECT 40.11 2.14 40.37 2.46 ;
      RECT 37.67 3.54 37.93 3.86 ;
      RECT 37.67 3.63 39.35 3.77 ;
      RECT 39.21 3.35 39.35 3.77 ;
      RECT 39.21 3.35 39.65 3.58 ;
      RECT 39.39 3.26 39.65 3.58 ;
      RECT 38.71 2.42 39.11 2.93 ;
      RECT 38.9 2.395 39.18 2.765 ;
      RECT 38.65 2.42 39.18 2.74 ;
      RECT 31.715 6.22 32.035 6.545 ;
      RECT 31.745 5.695 31.915 6.545 ;
      RECT 31.745 5.695 31.92 6.045 ;
      RECT 31.745 5.695 32.72 5.87 ;
      RECT 32.545 1.965 32.72 5.87 ;
      RECT 32.49 1.965 32.84 2.315 ;
      RECT 32.515 6.655 32.84 6.98 ;
      RECT 31.4 6.745 32.84 6.915 ;
      RECT 31.4 2.395 31.56 6.915 ;
      RECT 31.715 2.365 32.035 2.685 ;
      RECT 31.4 2.395 32.035 2.565 ;
      RECT 20.135 2.955 20.415 3.325 ;
      RECT 20.19 1.29 20.36 3.325 ;
      RECT 30.185 1.29 30.355 1.815 ;
      RECT 30.095 1.46 30.435 1.81 ;
      RECT 20.19 1.29 30.355 1.46 ;
      RECT 26.815 2.395 27.095 2.765 ;
      RECT 25.745 2.42 26.005 2.74 ;
      RECT 28.295 2.23 28.575 2.6 ;
      RECT 28.905 2.14 29.165 2.46 ;
      RECT 25.805 1.58 25.945 2.74 ;
      RECT 26.885 1.58 27.025 2.765 ;
      RECT 28.005 2.23 29.165 2.37 ;
      RECT 28.005 1.58 28.145 2.37 ;
      RECT 25.805 1.58 28.145 1.72 ;
      RECT 25.835 3.72 28.01 3.885 ;
      RECT 27.865 2.6 28.01 3.885 ;
      RECT 24.755 3.515 25.035 3.885 ;
      RECT 24.755 3.63 25.975 3.77 ;
      RECT 27.585 2.6 28.01 2.74 ;
      RECT 27.585 2.42 27.845 2.74 ;
      RECT 20.925 4 24.585 4.14 ;
      RECT 24.445 3.185 24.585 4.14 ;
      RECT 20.925 3.07 21.065 4.14 ;
      RECT 27.465 3.26 27.725 3.58 ;
      RECT 24.445 3.185 26.975 3.325 ;
      RECT 26.695 2.955 26.975 3.325 ;
      RECT 20.925 3.07 21.375 3.325 ;
      RECT 21.095 2.955 21.375 3.325 ;
      RECT 27.465 3.07 27.665 3.58 ;
      RECT 26.695 3.07 27.665 3.21 ;
      RECT 27.265 1.86 27.405 3.21 ;
      RECT 27.205 1.86 27.465 2.18 ;
      RECT 18.57 6.655 18.92 7.005 ;
      RECT 27.075 6.61 27.425 6.96 ;
      RECT 18.57 6.685 27.425 6.885 ;
      RECT 21.105 2.42 21.365 2.74 ;
      RECT 21.105 2.51 22.145 2.65 ;
      RECT 22.005 1.72 22.145 2.65 ;
      RECT 24.765 1.86 25.025 2.18 ;
      RECT 22.005 1.72 24.965 1.86 ;
      RECT 24.145 2.7 24.405 3.02 ;
      RECT 24.145 2.7 24.465 2.93 ;
      RECT 24.255 2.395 24.535 2.765 ;
      RECT 23.845 3.26 24.165 3.58 ;
      RECT 23.845 2.14 23.985 3.58 ;
      RECT 23.785 2.14 24.045 2.46 ;
      RECT 21.345 3.54 21.605 3.86 ;
      RECT 21.345 3.63 23.025 3.77 ;
      RECT 22.885 3.35 23.025 3.77 ;
      RECT 22.885 3.35 23.325 3.58 ;
      RECT 23.065 3.26 23.325 3.58 ;
      RECT 22.385 2.42 22.785 2.93 ;
      RECT 22.575 2.395 22.855 2.765 ;
      RECT 22.325 2.42 22.855 2.74 ;
      RECT 15.39 6.22 15.71 6.545 ;
      RECT 15.42 5.695 15.59 6.545 ;
      RECT 15.42 5.695 15.595 6.045 ;
      RECT 15.42 5.695 16.395 5.87 ;
      RECT 16.22 1.965 16.395 5.87 ;
      RECT 16.165 1.965 16.515 2.315 ;
      RECT 16.19 6.655 16.515 6.98 ;
      RECT 15.075 6.745 16.515 6.915 ;
      RECT 15.075 2.395 15.235 6.915 ;
      RECT 15.39 2.365 15.71 2.685 ;
      RECT 15.075 2.395 15.71 2.565 ;
      RECT 3.81 2.955 4.09 3.325 ;
      RECT 3.865 1.29 4.035 3.325 ;
      RECT 13.86 1.29 14.03 1.815 ;
      RECT 13.77 1.46 14.11 1.81 ;
      RECT 3.865 1.29 14.03 1.46 ;
      RECT 10.49 2.395 10.77 2.765 ;
      RECT 9.42 2.42 9.68 2.74 ;
      RECT 11.97 2.23 12.25 2.6 ;
      RECT 12.58 2.14 12.84 2.46 ;
      RECT 9.48 1.58 9.62 2.74 ;
      RECT 10.56 1.58 10.7 2.765 ;
      RECT 11.68 2.23 12.84 2.37 ;
      RECT 11.68 1.58 11.82 2.37 ;
      RECT 9.48 1.58 11.82 1.72 ;
      RECT 1.54 6.995 1.83 7.345 ;
      RECT 1.54 7.05 2.88 7.22 ;
      RECT 2.71 6.685 2.88 7.22 ;
      RECT 11.585 6.605 11.935 6.955 ;
      RECT 2.71 6.685 11.935 6.855 ;
      RECT 9.51 3.72 11.685 3.885 ;
      RECT 11.54 2.6 11.685 3.885 ;
      RECT 8.43 3.515 8.71 3.885 ;
      RECT 8.43 3.63 9.65 3.77 ;
      RECT 11.26 2.6 11.685 2.74 ;
      RECT 11.26 2.42 11.52 2.74 ;
      RECT 4.6 4 8.26 4.14 ;
      RECT 8.12 3.185 8.26 4.14 ;
      RECT 4.6 3.07 4.74 4.14 ;
      RECT 11.14 3.26 11.4 3.58 ;
      RECT 8.12 3.185 10.65 3.325 ;
      RECT 10.37 2.955 10.65 3.325 ;
      RECT 4.6 3.07 5.05 3.325 ;
      RECT 4.77 2.955 5.05 3.325 ;
      RECT 11.14 3.07 11.34 3.58 ;
      RECT 10.37 3.07 11.34 3.21 ;
      RECT 10.94 1.86 11.08 3.21 ;
      RECT 10.88 1.86 11.14 2.18 ;
      RECT 4.78 2.42 5.04 2.74 ;
      RECT 4.78 2.51 5.82 2.65 ;
      RECT 5.68 1.72 5.82 2.65 ;
      RECT 8.44 1.86 8.7 2.18 ;
      RECT 5.68 1.72 8.64 1.86 ;
      RECT 7.82 2.7 8.08 3.02 ;
      RECT 7.82 2.7 8.14 2.93 ;
      RECT 7.93 2.395 8.21 2.765 ;
      RECT 7.52 3.26 7.84 3.58 ;
      RECT 7.52 2.14 7.66 3.58 ;
      RECT 7.46 2.14 7.72 2.46 ;
      RECT 5.02 3.54 5.28 3.86 ;
      RECT 5.02 3.63 6.7 3.77 ;
      RECT 6.56 3.35 6.7 3.77 ;
      RECT 6.56 3.35 7 3.58 ;
      RECT 6.74 3.26 7 3.58 ;
      RECT 6.06 2.42 6.46 2.93 ;
      RECT 6.25 2.395 6.53 2.765 ;
      RECT 6 2.42 6.53 2.74 ;
      RECT 75.4 7.055 75.77 7.425 ;
      RECT 74.11 2.395 74.39 2.765 ;
      RECT 72.27 2.395 72.55 2.765 ;
      RECT 70.55 1.835 70.83 2.205 ;
      RECT 59.075 7.055 59.445 7.425 ;
      RECT 57.785 2.395 58.065 2.765 ;
      RECT 55.945 2.395 56.225 2.765 ;
      RECT 54.225 1.835 54.505 2.205 ;
      RECT 42.75 7.055 43.12 7.425 ;
      RECT 41.46 2.395 41.74 2.765 ;
      RECT 39.62 2.395 39.9 2.765 ;
      RECT 37.9 1.835 38.18 2.205 ;
      RECT 26.425 7.055 26.795 7.425 ;
      RECT 25.135 2.395 25.415 2.765 ;
      RECT 23.295 2.395 23.575 2.765 ;
      RECT 21.575 1.835 21.855 2.205 ;
      RECT 10.1 7.055 10.47 7.425 ;
      RECT 8.81 2.395 9.09 2.765 ;
      RECT 6.97 2.395 7.25 2.765 ;
      RECT 5.25 1.835 5.53 2.205 ;
    LAYER via1 ;
      RECT 83.95 7.375 84.1 7.525 ;
      RECT 81.58 6.74 81.73 6.89 ;
      RECT 81.565 2.065 81.715 2.215 ;
      RECT 80.775 2.45 80.925 2.6 ;
      RECT 80.775 6.325 80.925 6.475 ;
      RECT 79.17 1.56 79.32 1.71 ;
      RECT 77.935 2.225 78.085 2.375 ;
      RECT 76.615 2.505 76.765 2.655 ;
      RECT 76.495 3.345 76.645 3.495 ;
      RECT 76.235 1.945 76.385 2.095 ;
      RECT 76.155 6.71 76.305 6.86 ;
      RECT 75.51 7.165 75.66 7.315 ;
      RECT 74.775 2.505 74.925 2.655 ;
      RECT 74.175 2.505 74.325 2.655 ;
      RECT 73.795 1.945 73.945 2.095 ;
      RECT 73.175 2.785 73.325 2.935 ;
      RECT 72.935 3.345 73.085 3.495 ;
      RECT 72.815 2.225 72.965 2.375 ;
      RECT 72.335 2.505 72.485 2.655 ;
      RECT 72.095 3.345 72.245 3.495 ;
      RECT 71.355 2.505 71.505 2.655 ;
      RECT 70.615 1.945 70.765 2.095 ;
      RECT 70.375 3.625 70.525 3.775 ;
      RECT 70.135 2.505 70.285 2.655 ;
      RECT 70.135 3.065 70.285 3.215 ;
      RECT 69.175 3.065 69.325 3.215 ;
      RECT 67.6 6.755 67.75 6.905 ;
      RECT 65.255 6.74 65.405 6.89 ;
      RECT 65.24 2.065 65.39 2.215 ;
      RECT 64.45 2.45 64.6 2.6 ;
      RECT 64.45 6.325 64.6 6.475 ;
      RECT 62.845 1.56 62.995 1.71 ;
      RECT 61.61 2.225 61.76 2.375 ;
      RECT 60.29 2.505 60.44 2.655 ;
      RECT 60.17 3.345 60.32 3.495 ;
      RECT 59.91 1.945 60.06 2.095 ;
      RECT 59.825 6.71 59.975 6.86 ;
      RECT 59.185 7.165 59.335 7.315 ;
      RECT 58.45 2.505 58.6 2.655 ;
      RECT 57.85 2.505 58 2.655 ;
      RECT 57.47 1.945 57.62 2.095 ;
      RECT 56.85 2.785 57 2.935 ;
      RECT 56.61 3.345 56.76 3.495 ;
      RECT 56.49 2.225 56.64 2.375 ;
      RECT 56.01 2.505 56.16 2.655 ;
      RECT 55.77 3.345 55.92 3.495 ;
      RECT 55.03 2.505 55.18 2.655 ;
      RECT 54.29 1.945 54.44 2.095 ;
      RECT 54.05 3.625 54.2 3.775 ;
      RECT 53.81 2.505 53.96 2.655 ;
      RECT 53.81 3.065 53.96 3.215 ;
      RECT 52.85 3.065 53 3.215 ;
      RECT 51.275 6.755 51.425 6.905 ;
      RECT 48.93 6.74 49.08 6.89 ;
      RECT 48.915 2.065 49.065 2.215 ;
      RECT 48.125 2.45 48.275 2.6 ;
      RECT 48.125 6.325 48.275 6.475 ;
      RECT 46.52 1.56 46.67 1.71 ;
      RECT 45.285 2.225 45.435 2.375 ;
      RECT 43.965 2.505 44.115 2.655 ;
      RECT 43.845 3.345 43.995 3.495 ;
      RECT 43.585 1.945 43.735 2.095 ;
      RECT 43.5 6.715 43.65 6.865 ;
      RECT 42.86 7.165 43.01 7.315 ;
      RECT 42.125 2.505 42.275 2.655 ;
      RECT 41.525 2.505 41.675 2.655 ;
      RECT 41.145 1.945 41.295 2.095 ;
      RECT 40.525 2.785 40.675 2.935 ;
      RECT 40.285 3.345 40.435 3.495 ;
      RECT 40.165 2.225 40.315 2.375 ;
      RECT 39.685 2.505 39.835 2.655 ;
      RECT 39.445 3.345 39.595 3.495 ;
      RECT 38.705 2.505 38.855 2.655 ;
      RECT 37.965 1.945 38.115 2.095 ;
      RECT 37.725 3.625 37.875 3.775 ;
      RECT 37.485 2.505 37.635 2.655 ;
      RECT 37.485 3.065 37.635 3.215 ;
      RECT 36.525 3.065 36.675 3.215 ;
      RECT 34.995 6.76 35.145 6.91 ;
      RECT 32.605 6.74 32.755 6.89 ;
      RECT 32.59 2.065 32.74 2.215 ;
      RECT 31.8 2.45 31.95 2.6 ;
      RECT 31.8 6.325 31.95 6.475 ;
      RECT 30.195 1.56 30.345 1.71 ;
      RECT 28.96 2.225 29.11 2.375 ;
      RECT 27.64 2.505 27.79 2.655 ;
      RECT 27.52 3.345 27.67 3.495 ;
      RECT 27.26 1.945 27.41 2.095 ;
      RECT 27.175 6.71 27.325 6.86 ;
      RECT 26.535 7.165 26.685 7.315 ;
      RECT 25.8 2.505 25.95 2.655 ;
      RECT 25.2 2.505 25.35 2.655 ;
      RECT 24.82 1.945 24.97 2.095 ;
      RECT 24.2 2.785 24.35 2.935 ;
      RECT 23.96 3.345 24.11 3.495 ;
      RECT 23.84 2.225 23.99 2.375 ;
      RECT 23.36 2.505 23.51 2.655 ;
      RECT 23.12 3.345 23.27 3.495 ;
      RECT 22.38 2.505 22.53 2.655 ;
      RECT 21.64 1.945 21.79 2.095 ;
      RECT 21.4 3.625 21.55 3.775 ;
      RECT 21.16 2.505 21.31 2.655 ;
      RECT 21.16 3.065 21.31 3.215 ;
      RECT 20.2 3.065 20.35 3.215 ;
      RECT 18.67 6.755 18.82 6.905 ;
      RECT 16.28 6.74 16.43 6.89 ;
      RECT 16.265 2.065 16.415 2.215 ;
      RECT 15.475 2.45 15.625 2.6 ;
      RECT 15.475 6.325 15.625 6.475 ;
      RECT 13.87 1.56 14.02 1.71 ;
      RECT 12.635 2.225 12.785 2.375 ;
      RECT 11.685 6.705 11.835 6.855 ;
      RECT 11.315 2.505 11.465 2.655 ;
      RECT 11.195 3.345 11.345 3.495 ;
      RECT 10.935 1.945 11.085 2.095 ;
      RECT 10.21 7.165 10.36 7.315 ;
      RECT 9.475 2.505 9.625 2.655 ;
      RECT 8.875 2.505 9.025 2.655 ;
      RECT 8.495 1.945 8.645 2.095 ;
      RECT 7.875 2.785 8.025 2.935 ;
      RECT 7.635 3.345 7.785 3.495 ;
      RECT 7.515 2.225 7.665 2.375 ;
      RECT 7.035 2.505 7.185 2.655 ;
      RECT 6.795 3.345 6.945 3.495 ;
      RECT 6.055 2.505 6.205 2.655 ;
      RECT 5.315 1.945 5.465 2.095 ;
      RECT 5.075 3.625 5.225 3.775 ;
      RECT 4.835 2.505 4.985 2.655 ;
      RECT 4.835 3.065 4.985 3.215 ;
      RECT 3.875 3.065 4.025 3.215 ;
      RECT 1.61 7.095 1.76 7.245 ;
      RECT 1.235 6.355 1.385 6.505 ;
    LAYER met1 ;
      RECT 83.815 7.77 84.105 8 ;
      RECT 83.875 6.29 84.045 8 ;
      RECT 83.85 7.275 84.2 7.625 ;
      RECT 83.815 6.29 84.105 6.52 ;
      RECT 83.41 2.395 83.515 2.965 ;
      RECT 83.41 2.73 83.735 2.96 ;
      RECT 83.41 2.76 83.905 2.93 ;
      RECT 83.41 2.395 83.6 2.96 ;
      RECT 82.825 2.36 83.115 2.59 ;
      RECT 82.825 2.395 83.6 2.565 ;
      RECT 82.885 0.88 83.055 2.59 ;
      RECT 82.825 0.88 83.115 1.11 ;
      RECT 82.825 7.77 83.115 8 ;
      RECT 82.885 6.29 83.055 8 ;
      RECT 82.825 6.29 83.115 6.52 ;
      RECT 82.825 6.325 83.68 6.485 ;
      RECT 83.51 5.92 83.68 6.485 ;
      RECT 82.825 6.32 83.22 6.485 ;
      RECT 83.445 5.92 83.735 6.15 ;
      RECT 83.445 5.95 83.905 6.12 ;
      RECT 82.455 2.73 82.745 2.96 ;
      RECT 82.455 2.76 82.915 2.93 ;
      RECT 82.52 1.655 82.685 2.96 ;
      RECT 81.035 1.625 81.325 1.855 ;
      RECT 81.035 1.655 82.685 1.825 ;
      RECT 81.095 0.885 81.265 1.855 ;
      RECT 81.035 0.885 81.325 1.115 ;
      RECT 81.035 7.765 81.325 7.995 ;
      RECT 81.095 7.025 81.265 7.995 ;
      RECT 81.095 7.12 82.685 7.29 ;
      RECT 82.515 5.92 82.685 7.29 ;
      RECT 81.035 7.025 81.325 7.255 ;
      RECT 82.455 5.92 82.745 6.15 ;
      RECT 82.455 5.95 82.915 6.12 ;
      RECT 81.465 1.965 81.815 2.315 ;
      RECT 79.16 2.025 81.815 2.195 ;
      RECT 79.16 1.46 79.33 2.195 ;
      RECT 79.07 1.46 79.41 1.81 ;
      RECT 81.49 6.655 81.815 6.98 ;
      RECT 76.055 6.61 76.405 6.96 ;
      RECT 81.465 6.655 81.815 6.885 ;
      RECT 75.85 6.655 76.405 6.885 ;
      RECT 75.68 6.685 81.815 6.855 ;
      RECT 80.69 2.365 81.01 2.685 ;
      RECT 80.66 2.365 81.01 2.595 ;
      RECT 80.49 2.395 81.01 2.565 ;
      RECT 80.69 6.255 81.01 6.545 ;
      RECT 80.66 6.285 81.01 6.515 ;
      RECT 80.49 6.315 81.01 6.485 ;
      RECT 77.145 2.465 77.435 2.695 ;
      RECT 77.145 2.465 77.6 2.65 ;
      RECT 77.46 2.37 78.08 2.51 ;
      RECT 77.85 2.17 78.17 2.43 ;
      RECT 76.53 2.45 76.85 2.71 ;
      RECT 76.53 2.45 76.995 2.695 ;
      RECT 76.855 2.07 76.995 2.695 ;
      RECT 76.855 2.07 77.12 2.21 ;
      RECT 77.385 1.905 77.675 2.135 ;
      RECT 76.98 1.95 77.675 2.09 ;
      RECT 76.425 3.29 76.715 3.815 ;
      RECT 76.41 3.29 76.73 3.55 ;
      RECT 76.15 1.89 76.47 2.15 ;
      RECT 76.15 1.905 76.715 2.135 ;
      RECT 75.425 3.585 75.715 3.815 ;
      RECT 75.62 2.23 75.76 3.77 ;
      RECT 75.665 2.185 75.955 2.415 ;
      RECT 75.26 2.23 75.955 2.37 ;
      RECT 75.26 2.07 75.4 2.37 ;
      RECT 73.8 2.07 75.4 2.21 ;
      RECT 73.71 1.89 74.03 2.15 ;
      RECT 73.71 1.905 74.275 2.15 ;
      RECT 75.42 7.765 75.71 7.995 ;
      RECT 75.48 7.025 75.65 7.995 ;
      RECT 75.4 7.075 75.77 7.425 ;
      RECT 75.4 7.055 75.71 7.425 ;
      RECT 75.42 7.025 75.71 7.425 ;
      RECT 72.82 2.93 75.4 3.07 ;
      RECT 75.185 2.745 75.475 2.975 ;
      RECT 72.745 2.745 73.41 2.975 ;
      RECT 73.09 2.73 73.41 3.07 ;
      RECT 74.09 2.45 74.41 2.71 ;
      RECT 74.09 2.465 74.515 2.695 ;
      RECT 72.73 2.17 73.05 2.43 ;
      RECT 73.225 2.185 73.515 2.415 ;
      RECT 72.73 2.23 73.515 2.37 ;
      RECT 72.85 3.29 73.17 3.55 ;
      RECT 72.01 3.29 72.33 3.55 ;
      RECT 72.85 3.305 73.275 3.535 ;
      RECT 72.01 3.35 73.275 3.49 ;
      RECT 71.545 3.025 71.835 3.255 ;
      RECT 71.62 1.95 71.76 3.255 ;
      RECT 71.27 2.45 71.76 2.71 ;
      RECT 71.025 2.465 71.76 2.695 ;
      RECT 72.025 1.905 72.315 2.135 ;
      RECT 71.62 1.95 72.315 2.09 ;
      RECT 70.785 3.305 71.075 3.535 ;
      RECT 70.785 3.305 71.24 3.49 ;
      RECT 71.1 2.93 71.24 3.49 ;
      RECT 70.74 2.93 71.24 3.07 ;
      RECT 70.74 1.95 70.88 3.07 ;
      RECT 70.53 1.89 70.85 2.15 ;
      RECT 70.29 3.57 70.61 3.83 ;
      RECT 69.585 3.585 69.875 3.815 ;
      RECT 69.585 3.63 70.61 3.77 ;
      RECT 69.66 3.58 69.92 3.77 ;
      RECT 70.05 2.45 70.37 2.71 ;
      RECT 70.05 2.465 70.595 2.695 ;
      RECT 70.05 3.01 70.37 3.27 ;
      RECT 70.05 3.025 70.595 3.255 ;
      RECT 69.09 3.01 69.41 3.27 ;
      RECT 69.18 1.95 69.32 3.27 ;
      RECT 69.585 1.905 69.875 2.135 ;
      RECT 69.18 1.95 69.875 2.09 ;
      RECT 67.49 7.77 67.78 8 ;
      RECT 67.55 6.29 67.72 8 ;
      RECT 67.5 6.655 67.85 7.005 ;
      RECT 67.49 6.29 67.78 6.52 ;
      RECT 67.085 2.395 67.19 2.965 ;
      RECT 67.085 2.73 67.41 2.96 ;
      RECT 67.085 2.76 67.58 2.93 ;
      RECT 67.085 2.395 67.275 2.96 ;
      RECT 66.5 2.36 66.79 2.59 ;
      RECT 66.5 2.395 67.275 2.565 ;
      RECT 66.56 0.88 66.73 2.59 ;
      RECT 66.5 0.88 66.79 1.11 ;
      RECT 66.5 7.77 66.79 8 ;
      RECT 66.56 6.29 66.73 8 ;
      RECT 66.5 6.29 66.79 6.52 ;
      RECT 66.5 6.325 67.355 6.485 ;
      RECT 67.185 5.92 67.355 6.485 ;
      RECT 66.5 6.32 66.895 6.485 ;
      RECT 67.12 5.92 67.41 6.15 ;
      RECT 67.12 5.95 67.58 6.12 ;
      RECT 66.13 2.73 66.42 2.96 ;
      RECT 66.13 2.76 66.59 2.93 ;
      RECT 66.195 1.655 66.36 2.96 ;
      RECT 64.71 1.625 65 1.855 ;
      RECT 64.71 1.655 66.36 1.825 ;
      RECT 64.77 0.885 64.94 1.855 ;
      RECT 64.71 0.885 65 1.115 ;
      RECT 64.71 7.765 65 7.995 ;
      RECT 64.77 7.025 64.94 7.995 ;
      RECT 64.77 7.12 66.36 7.29 ;
      RECT 66.19 5.92 66.36 7.29 ;
      RECT 64.71 7.025 65 7.255 ;
      RECT 66.13 5.92 66.42 6.15 ;
      RECT 66.13 5.95 66.59 6.12 ;
      RECT 65.14 1.965 65.49 2.315 ;
      RECT 62.835 2.025 65.49 2.195 ;
      RECT 62.835 1.46 63.005 2.195 ;
      RECT 62.745 1.46 63.085 1.81 ;
      RECT 65.165 6.655 65.49 6.98 ;
      RECT 59.725 6.61 60.075 6.96 ;
      RECT 65.14 6.655 65.49 6.885 ;
      RECT 59.525 6.655 60.075 6.885 ;
      RECT 59.355 6.685 65.49 6.855 ;
      RECT 64.365 2.365 64.685 2.685 ;
      RECT 64.335 2.365 64.685 2.595 ;
      RECT 64.165 2.395 64.685 2.565 ;
      RECT 64.365 6.255 64.685 6.545 ;
      RECT 64.335 6.285 64.685 6.515 ;
      RECT 64.165 6.315 64.685 6.485 ;
      RECT 60.82 2.465 61.11 2.695 ;
      RECT 60.82 2.465 61.275 2.65 ;
      RECT 61.135 2.37 61.755 2.51 ;
      RECT 61.525 2.17 61.845 2.43 ;
      RECT 60.205 2.45 60.525 2.71 ;
      RECT 60.205 2.45 60.67 2.695 ;
      RECT 60.53 2.07 60.67 2.695 ;
      RECT 60.53 2.07 60.795 2.21 ;
      RECT 61.06 1.905 61.35 2.135 ;
      RECT 60.655 1.95 61.35 2.09 ;
      RECT 60.1 3.29 60.39 3.815 ;
      RECT 60.085 3.29 60.405 3.55 ;
      RECT 59.825 1.89 60.145 2.15 ;
      RECT 59.825 1.905 60.39 2.135 ;
      RECT 59.1 3.585 59.39 3.815 ;
      RECT 59.295 2.23 59.435 3.77 ;
      RECT 59.34 2.185 59.63 2.415 ;
      RECT 58.935 2.23 59.63 2.37 ;
      RECT 58.935 2.07 59.075 2.37 ;
      RECT 57.475 2.07 59.075 2.21 ;
      RECT 57.385 1.89 57.705 2.15 ;
      RECT 57.385 1.905 57.95 2.15 ;
      RECT 59.095 7.765 59.385 7.995 ;
      RECT 59.155 7.025 59.325 7.995 ;
      RECT 59.075 7.075 59.445 7.425 ;
      RECT 59.075 7.055 59.385 7.425 ;
      RECT 59.095 7.025 59.385 7.425 ;
      RECT 56.495 2.93 59.075 3.07 ;
      RECT 58.86 2.745 59.15 2.975 ;
      RECT 56.42 2.745 57.085 2.975 ;
      RECT 56.765 2.73 57.085 3.07 ;
      RECT 57.765 2.45 58.085 2.71 ;
      RECT 57.765 2.465 58.19 2.695 ;
      RECT 56.405 2.17 56.725 2.43 ;
      RECT 56.9 2.185 57.19 2.415 ;
      RECT 56.405 2.23 57.19 2.37 ;
      RECT 56.525 3.29 56.845 3.55 ;
      RECT 55.685 3.29 56.005 3.55 ;
      RECT 56.525 3.305 56.95 3.535 ;
      RECT 55.685 3.35 56.95 3.49 ;
      RECT 55.22 3.025 55.51 3.255 ;
      RECT 55.295 1.95 55.435 3.255 ;
      RECT 54.945 2.45 55.435 2.71 ;
      RECT 54.7 2.465 55.435 2.695 ;
      RECT 55.7 1.905 55.99 2.135 ;
      RECT 55.295 1.95 55.99 2.09 ;
      RECT 54.46 3.305 54.75 3.535 ;
      RECT 54.46 3.305 54.915 3.49 ;
      RECT 54.775 2.93 54.915 3.49 ;
      RECT 54.415 2.93 54.915 3.07 ;
      RECT 54.415 1.95 54.555 3.07 ;
      RECT 54.205 1.89 54.525 2.15 ;
      RECT 53.965 3.57 54.285 3.83 ;
      RECT 53.26 3.585 53.55 3.815 ;
      RECT 53.26 3.63 54.285 3.77 ;
      RECT 53.335 3.58 53.595 3.77 ;
      RECT 53.725 2.45 54.045 2.71 ;
      RECT 53.725 2.465 54.27 2.695 ;
      RECT 53.725 3.01 54.045 3.27 ;
      RECT 53.725 3.025 54.27 3.255 ;
      RECT 52.765 3.01 53.085 3.27 ;
      RECT 52.855 1.95 52.995 3.27 ;
      RECT 53.26 1.905 53.55 2.135 ;
      RECT 52.855 1.95 53.55 2.09 ;
      RECT 51.165 7.77 51.455 8 ;
      RECT 51.225 6.29 51.395 8 ;
      RECT 51.175 6.655 51.525 7.005 ;
      RECT 51.165 6.29 51.455 6.52 ;
      RECT 50.76 2.395 50.865 2.965 ;
      RECT 50.76 2.73 51.085 2.96 ;
      RECT 50.76 2.76 51.255 2.93 ;
      RECT 50.76 2.395 50.95 2.96 ;
      RECT 50.175 2.36 50.465 2.59 ;
      RECT 50.175 2.395 50.95 2.565 ;
      RECT 50.235 0.88 50.405 2.59 ;
      RECT 50.175 0.88 50.465 1.11 ;
      RECT 50.175 7.77 50.465 8 ;
      RECT 50.235 6.29 50.405 8 ;
      RECT 50.175 6.29 50.465 6.52 ;
      RECT 50.175 6.325 51.03 6.485 ;
      RECT 50.86 5.92 51.03 6.485 ;
      RECT 50.175 6.32 50.57 6.485 ;
      RECT 50.795 5.92 51.085 6.15 ;
      RECT 50.795 5.95 51.255 6.12 ;
      RECT 49.805 2.73 50.095 2.96 ;
      RECT 49.805 2.76 50.265 2.93 ;
      RECT 49.87 1.655 50.035 2.96 ;
      RECT 48.385 1.625 48.675 1.855 ;
      RECT 48.385 1.655 50.035 1.825 ;
      RECT 48.445 0.885 48.615 1.855 ;
      RECT 48.385 0.885 48.675 1.115 ;
      RECT 48.385 7.765 48.675 7.995 ;
      RECT 48.445 7.025 48.615 7.995 ;
      RECT 48.445 7.12 50.035 7.29 ;
      RECT 49.865 5.92 50.035 7.29 ;
      RECT 48.385 7.025 48.675 7.255 ;
      RECT 49.805 5.92 50.095 6.15 ;
      RECT 49.805 5.95 50.265 6.12 ;
      RECT 48.815 1.965 49.165 2.315 ;
      RECT 46.51 2.025 49.165 2.195 ;
      RECT 46.51 1.46 46.68 2.195 ;
      RECT 46.42 1.46 46.76 1.81 ;
      RECT 48.84 6.655 49.165 6.98 ;
      RECT 43.4 6.615 43.75 6.965 ;
      RECT 48.815 6.655 49.165 6.885 ;
      RECT 43.2 6.655 43.75 6.885 ;
      RECT 43.03 6.685 49.165 6.855 ;
      RECT 48.04 2.365 48.36 2.685 ;
      RECT 48.01 2.365 48.36 2.595 ;
      RECT 47.84 2.395 48.36 2.565 ;
      RECT 48.04 6.255 48.36 6.545 ;
      RECT 48.01 6.285 48.36 6.515 ;
      RECT 47.84 6.315 48.36 6.485 ;
      RECT 44.495 2.465 44.785 2.695 ;
      RECT 44.495 2.465 44.95 2.65 ;
      RECT 44.81 2.37 45.43 2.51 ;
      RECT 45.2 2.17 45.52 2.43 ;
      RECT 43.88 2.45 44.2 2.71 ;
      RECT 43.88 2.45 44.345 2.695 ;
      RECT 44.205 2.07 44.345 2.695 ;
      RECT 44.205 2.07 44.47 2.21 ;
      RECT 44.735 1.905 45.025 2.135 ;
      RECT 44.33 1.95 45.025 2.09 ;
      RECT 43.775 3.29 44.065 3.815 ;
      RECT 43.76 3.29 44.08 3.55 ;
      RECT 43.5 1.89 43.82 2.15 ;
      RECT 43.5 1.905 44.065 2.135 ;
      RECT 42.775 3.585 43.065 3.815 ;
      RECT 42.97 2.23 43.11 3.77 ;
      RECT 43.015 2.185 43.305 2.415 ;
      RECT 42.61 2.23 43.305 2.37 ;
      RECT 42.61 2.07 42.75 2.37 ;
      RECT 41.15 2.07 42.75 2.21 ;
      RECT 41.06 1.89 41.38 2.15 ;
      RECT 41.06 1.905 41.625 2.15 ;
      RECT 42.77 7.765 43.06 7.995 ;
      RECT 42.83 7.025 43 7.995 ;
      RECT 42.75 7.075 43.12 7.425 ;
      RECT 42.75 7.055 43.06 7.425 ;
      RECT 42.77 7.025 43.06 7.425 ;
      RECT 40.17 2.93 42.75 3.07 ;
      RECT 42.535 2.745 42.825 2.975 ;
      RECT 40.095 2.745 40.76 2.975 ;
      RECT 40.44 2.73 40.76 3.07 ;
      RECT 41.44 2.45 41.76 2.71 ;
      RECT 41.44 2.465 41.865 2.695 ;
      RECT 40.08 2.17 40.4 2.43 ;
      RECT 40.575 2.185 40.865 2.415 ;
      RECT 40.08 2.23 40.865 2.37 ;
      RECT 40.2 3.29 40.52 3.55 ;
      RECT 39.36 3.29 39.68 3.55 ;
      RECT 40.2 3.305 40.625 3.535 ;
      RECT 39.36 3.35 40.625 3.49 ;
      RECT 38.895 3.025 39.185 3.255 ;
      RECT 38.97 1.95 39.11 3.255 ;
      RECT 38.62 2.45 39.11 2.71 ;
      RECT 38.375 2.465 39.11 2.695 ;
      RECT 39.375 1.905 39.665 2.135 ;
      RECT 38.97 1.95 39.665 2.09 ;
      RECT 38.135 3.305 38.425 3.535 ;
      RECT 38.135 3.305 38.59 3.49 ;
      RECT 38.45 2.93 38.59 3.49 ;
      RECT 38.09 2.93 38.59 3.07 ;
      RECT 38.09 1.95 38.23 3.07 ;
      RECT 37.88 1.89 38.2 2.15 ;
      RECT 37.64 3.57 37.96 3.83 ;
      RECT 36.935 3.585 37.225 3.815 ;
      RECT 36.935 3.63 37.96 3.77 ;
      RECT 37.01 3.58 37.27 3.77 ;
      RECT 37.4 2.45 37.72 2.71 ;
      RECT 37.4 2.465 37.945 2.695 ;
      RECT 37.4 3.01 37.72 3.27 ;
      RECT 37.4 3.025 37.945 3.255 ;
      RECT 36.44 3.01 36.76 3.27 ;
      RECT 36.53 1.95 36.67 3.27 ;
      RECT 36.935 1.905 37.225 2.135 ;
      RECT 36.53 1.95 37.225 2.09 ;
      RECT 34.84 7.77 35.13 8 ;
      RECT 34.9 6.29 35.07 8 ;
      RECT 34.89 6.66 35.245 7.015 ;
      RECT 34.84 6.29 35.13 6.52 ;
      RECT 34.435 2.395 34.54 2.965 ;
      RECT 34.435 2.73 34.76 2.96 ;
      RECT 34.435 2.76 34.93 2.93 ;
      RECT 34.435 2.395 34.625 2.96 ;
      RECT 33.85 2.36 34.14 2.59 ;
      RECT 33.85 2.395 34.625 2.565 ;
      RECT 33.91 0.88 34.08 2.59 ;
      RECT 33.85 0.88 34.14 1.11 ;
      RECT 33.85 7.77 34.14 8 ;
      RECT 33.91 6.29 34.08 8 ;
      RECT 33.85 6.29 34.14 6.52 ;
      RECT 33.85 6.325 34.705 6.485 ;
      RECT 34.535 5.92 34.705 6.485 ;
      RECT 33.85 6.32 34.245 6.485 ;
      RECT 34.47 5.92 34.76 6.15 ;
      RECT 34.47 5.95 34.93 6.12 ;
      RECT 33.48 2.73 33.77 2.96 ;
      RECT 33.48 2.76 33.94 2.93 ;
      RECT 33.545 1.655 33.71 2.96 ;
      RECT 32.06 1.625 32.35 1.855 ;
      RECT 32.06 1.655 33.71 1.825 ;
      RECT 32.12 0.885 32.29 1.855 ;
      RECT 32.06 0.885 32.35 1.115 ;
      RECT 32.06 7.765 32.35 7.995 ;
      RECT 32.12 7.025 32.29 7.995 ;
      RECT 32.12 7.12 33.71 7.29 ;
      RECT 33.54 5.92 33.71 7.29 ;
      RECT 32.06 7.025 32.35 7.255 ;
      RECT 33.48 5.92 33.77 6.15 ;
      RECT 33.48 5.95 33.94 6.12 ;
      RECT 32.49 1.965 32.84 2.315 ;
      RECT 30.185 2.025 32.84 2.195 ;
      RECT 30.185 1.46 30.355 2.195 ;
      RECT 30.095 1.46 30.435 1.81 ;
      RECT 32.515 6.655 32.84 6.98 ;
      RECT 27.075 6.61 27.425 6.96 ;
      RECT 32.49 6.655 32.84 6.885 ;
      RECT 26.875 6.655 27.425 6.885 ;
      RECT 26.705 6.685 32.84 6.855 ;
      RECT 31.715 2.365 32.035 2.685 ;
      RECT 31.685 2.365 32.035 2.595 ;
      RECT 31.515 2.395 32.035 2.565 ;
      RECT 31.715 6.255 32.035 6.545 ;
      RECT 31.685 6.285 32.035 6.515 ;
      RECT 31.515 6.315 32.035 6.485 ;
      RECT 28.17 2.465 28.46 2.695 ;
      RECT 28.17 2.465 28.625 2.65 ;
      RECT 28.485 2.37 29.105 2.51 ;
      RECT 28.875 2.17 29.195 2.43 ;
      RECT 27.555 2.45 27.875 2.71 ;
      RECT 27.555 2.45 28.02 2.695 ;
      RECT 27.88 2.07 28.02 2.695 ;
      RECT 27.88 2.07 28.145 2.21 ;
      RECT 28.41 1.905 28.7 2.135 ;
      RECT 28.005 1.95 28.7 2.09 ;
      RECT 27.45 3.29 27.74 3.815 ;
      RECT 27.435 3.29 27.755 3.55 ;
      RECT 27.175 1.89 27.495 2.15 ;
      RECT 27.175 1.905 27.74 2.135 ;
      RECT 26.45 3.585 26.74 3.815 ;
      RECT 26.645 2.23 26.785 3.77 ;
      RECT 26.69 2.185 26.98 2.415 ;
      RECT 26.285 2.23 26.98 2.37 ;
      RECT 26.285 2.07 26.425 2.37 ;
      RECT 24.825 2.07 26.425 2.21 ;
      RECT 24.735 1.89 25.055 2.15 ;
      RECT 24.735 1.905 25.3 2.15 ;
      RECT 26.445 7.765 26.735 7.995 ;
      RECT 26.505 7.025 26.675 7.995 ;
      RECT 26.425 7.075 26.795 7.425 ;
      RECT 26.425 7.055 26.735 7.425 ;
      RECT 26.445 7.025 26.735 7.425 ;
      RECT 23.845 2.93 26.425 3.07 ;
      RECT 26.21 2.745 26.5 2.975 ;
      RECT 23.77 2.745 24.435 2.975 ;
      RECT 24.115 2.73 24.435 3.07 ;
      RECT 25.115 2.45 25.435 2.71 ;
      RECT 25.115 2.465 25.54 2.695 ;
      RECT 23.755 2.17 24.075 2.43 ;
      RECT 24.25 2.185 24.54 2.415 ;
      RECT 23.755 2.23 24.54 2.37 ;
      RECT 23.875 3.29 24.195 3.55 ;
      RECT 23.035 3.29 23.355 3.55 ;
      RECT 23.875 3.305 24.3 3.535 ;
      RECT 23.035 3.35 24.3 3.49 ;
      RECT 22.57 3.025 22.86 3.255 ;
      RECT 22.645 1.95 22.785 3.255 ;
      RECT 22.295 2.45 22.785 2.71 ;
      RECT 22.05 2.465 22.785 2.695 ;
      RECT 23.05 1.905 23.34 2.135 ;
      RECT 22.645 1.95 23.34 2.09 ;
      RECT 21.81 3.305 22.1 3.535 ;
      RECT 21.81 3.305 22.265 3.49 ;
      RECT 22.125 2.93 22.265 3.49 ;
      RECT 21.765 2.93 22.265 3.07 ;
      RECT 21.765 1.95 21.905 3.07 ;
      RECT 21.555 1.89 21.875 2.15 ;
      RECT 21.315 3.57 21.635 3.83 ;
      RECT 20.61 3.585 20.9 3.815 ;
      RECT 20.61 3.63 21.635 3.77 ;
      RECT 20.685 3.58 20.945 3.77 ;
      RECT 21.075 2.45 21.395 2.71 ;
      RECT 21.075 2.465 21.62 2.695 ;
      RECT 21.075 3.01 21.395 3.27 ;
      RECT 21.075 3.025 21.62 3.255 ;
      RECT 20.115 3.01 20.435 3.27 ;
      RECT 20.205 1.95 20.345 3.27 ;
      RECT 20.61 1.905 20.9 2.135 ;
      RECT 20.205 1.95 20.9 2.09 ;
      RECT 18.515 7.77 18.805 8 ;
      RECT 18.575 6.29 18.745 8 ;
      RECT 18.57 6.655 18.92 7.005 ;
      RECT 18.515 6.29 18.805 6.52 ;
      RECT 18.11 2.395 18.215 2.965 ;
      RECT 18.11 2.73 18.435 2.96 ;
      RECT 18.11 2.76 18.605 2.93 ;
      RECT 18.11 2.395 18.3 2.96 ;
      RECT 17.525 2.36 17.815 2.59 ;
      RECT 17.525 2.395 18.3 2.565 ;
      RECT 17.585 0.88 17.755 2.59 ;
      RECT 17.525 0.88 17.815 1.11 ;
      RECT 17.525 7.77 17.815 8 ;
      RECT 17.585 6.29 17.755 8 ;
      RECT 17.525 6.29 17.815 6.52 ;
      RECT 17.525 6.325 18.38 6.485 ;
      RECT 18.21 5.92 18.38 6.485 ;
      RECT 17.525 6.32 17.92 6.485 ;
      RECT 18.145 5.92 18.435 6.15 ;
      RECT 18.145 5.95 18.605 6.12 ;
      RECT 17.155 2.73 17.445 2.96 ;
      RECT 17.155 2.76 17.615 2.93 ;
      RECT 17.22 1.655 17.385 2.96 ;
      RECT 15.735 1.625 16.025 1.855 ;
      RECT 15.735 1.655 17.385 1.825 ;
      RECT 15.795 0.885 15.965 1.855 ;
      RECT 15.735 0.885 16.025 1.115 ;
      RECT 15.735 7.765 16.025 7.995 ;
      RECT 15.795 7.025 15.965 7.995 ;
      RECT 15.795 7.12 17.385 7.29 ;
      RECT 17.215 5.92 17.385 7.29 ;
      RECT 15.735 7.025 16.025 7.255 ;
      RECT 17.155 5.92 17.445 6.15 ;
      RECT 17.155 5.95 17.615 6.12 ;
      RECT 16.165 1.965 16.515 2.315 ;
      RECT 13.86 2.025 16.515 2.195 ;
      RECT 13.86 1.46 14.03 2.195 ;
      RECT 13.77 1.46 14.11 1.81 ;
      RECT 16.19 6.655 16.515 6.98 ;
      RECT 11.585 6.605 11.935 6.955 ;
      RECT 16.165 6.655 16.515 6.885 ;
      RECT 10.55 6.655 10.84 6.885 ;
      RECT 10.38 6.685 16.515 6.855 ;
      RECT 15.39 2.365 15.71 2.685 ;
      RECT 15.36 2.365 15.71 2.595 ;
      RECT 15.19 2.395 15.71 2.565 ;
      RECT 15.39 6.255 15.71 6.545 ;
      RECT 15.36 6.285 15.71 6.515 ;
      RECT 15.19 6.315 15.71 6.485 ;
      RECT 11.845 2.465 12.135 2.695 ;
      RECT 11.845 2.465 12.3 2.65 ;
      RECT 12.16 2.37 12.78 2.51 ;
      RECT 12.55 2.17 12.87 2.43 ;
      RECT 11.23 2.45 11.55 2.71 ;
      RECT 11.23 2.45 11.695 2.695 ;
      RECT 11.555 2.07 11.695 2.695 ;
      RECT 11.555 2.07 11.82 2.21 ;
      RECT 12.085 1.905 12.375 2.135 ;
      RECT 11.68 1.95 12.375 2.09 ;
      RECT 11.125 3.29 11.415 3.815 ;
      RECT 11.11 3.29 11.43 3.55 ;
      RECT 10.85 1.89 11.17 2.15 ;
      RECT 10.85 1.905 11.415 2.135 ;
      RECT 10.125 3.585 10.415 3.815 ;
      RECT 10.32 2.23 10.46 3.77 ;
      RECT 10.365 2.185 10.655 2.415 ;
      RECT 9.96 2.23 10.655 2.37 ;
      RECT 9.96 2.07 10.1 2.37 ;
      RECT 8.5 2.07 10.1 2.21 ;
      RECT 8.41 1.89 8.73 2.15 ;
      RECT 8.41 1.905 8.975 2.15 ;
      RECT 10.12 7.765 10.41 7.995 ;
      RECT 10.18 7.025 10.35 7.995 ;
      RECT 10.1 7.075 10.47 7.425 ;
      RECT 10.1 7.055 10.41 7.425 ;
      RECT 10.12 7.025 10.41 7.425 ;
      RECT 7.52 2.93 10.1 3.07 ;
      RECT 9.885 2.745 10.175 2.975 ;
      RECT 7.445 2.745 8.11 2.975 ;
      RECT 7.79 2.73 8.11 3.07 ;
      RECT 8.79 2.45 9.11 2.71 ;
      RECT 8.79 2.465 9.215 2.695 ;
      RECT 7.43 2.17 7.75 2.43 ;
      RECT 7.925 2.185 8.215 2.415 ;
      RECT 7.43 2.23 8.215 2.37 ;
      RECT 7.55 3.29 7.87 3.55 ;
      RECT 6.71 3.29 7.03 3.55 ;
      RECT 7.55 3.305 7.975 3.535 ;
      RECT 6.71 3.35 7.975 3.49 ;
      RECT 6.245 3.025 6.535 3.255 ;
      RECT 6.32 1.95 6.46 3.255 ;
      RECT 5.97 2.45 6.46 2.71 ;
      RECT 5.725 2.465 6.46 2.695 ;
      RECT 6.725 1.905 7.015 2.135 ;
      RECT 6.32 1.95 7.015 2.09 ;
      RECT 5.485 3.305 5.775 3.535 ;
      RECT 5.485 3.305 5.94 3.49 ;
      RECT 5.8 2.93 5.94 3.49 ;
      RECT 5.44 2.93 5.94 3.07 ;
      RECT 5.44 1.95 5.58 3.07 ;
      RECT 5.23 1.89 5.55 2.15 ;
      RECT 4.99 3.57 5.31 3.83 ;
      RECT 4.285 3.585 4.575 3.815 ;
      RECT 4.285 3.63 5.31 3.77 ;
      RECT 4.36 3.58 4.62 3.77 ;
      RECT 4.75 2.45 5.07 2.71 ;
      RECT 4.75 2.465 5.295 2.695 ;
      RECT 4.75 3.01 5.07 3.27 ;
      RECT 4.75 3.025 5.295 3.255 ;
      RECT 3.79 3.01 4.11 3.27 ;
      RECT 3.88 1.95 4.02 3.27 ;
      RECT 4.285 1.905 4.575 2.135 ;
      RECT 3.88 1.95 4.575 2.09 ;
      RECT 1.54 7.765 1.83 7.995 ;
      RECT 1.6 7.025 1.77 7.995 ;
      RECT 1.51 7.025 1.86 7.315 ;
      RECT 1.135 6.285 1.485 6.575 ;
      RECT 0.995 6.315 1.485 6.485 ;
      RECT 74.69 2.45 75.01 2.71 ;
      RECT 72.25 2.45 72.57 2.71 ;
      RECT 58.365 2.45 58.685 2.71 ;
      RECT 55.925 2.45 56.245 2.71 ;
      RECT 42.04 2.45 42.36 2.71 ;
      RECT 39.6 2.45 39.92 2.71 ;
      RECT 25.715 2.45 26.035 2.71 ;
      RECT 23.275 2.45 23.595 2.71 ;
      RECT 9.39 2.45 9.71 2.71 ;
      RECT 6.95 2.45 7.27 2.71 ;
    LAYER mcon ;
      RECT 83.875 6.32 84.045 6.49 ;
      RECT 83.88 6.315 84.05 6.485 ;
      RECT 67.55 6.32 67.72 6.49 ;
      RECT 67.555 6.315 67.725 6.485 ;
      RECT 51.225 6.32 51.395 6.49 ;
      RECT 51.23 6.315 51.4 6.485 ;
      RECT 34.9 6.32 35.07 6.49 ;
      RECT 34.905 6.315 35.075 6.485 ;
      RECT 18.575 6.32 18.745 6.49 ;
      RECT 18.58 6.315 18.75 6.485 ;
      RECT 83.875 7.8 84.045 7.97 ;
      RECT 83.505 2.76 83.675 2.93 ;
      RECT 83.505 5.95 83.675 6.12 ;
      RECT 82.885 0.91 83.055 1.08 ;
      RECT 82.885 2.39 83.055 2.56 ;
      RECT 82.885 6.32 83.055 6.49 ;
      RECT 82.885 7.8 83.055 7.97 ;
      RECT 82.515 2.76 82.685 2.93 ;
      RECT 82.515 5.95 82.685 6.12 ;
      RECT 81.525 2.025 81.695 2.195 ;
      RECT 81.525 6.685 81.695 6.855 ;
      RECT 81.095 0.915 81.265 1.085 ;
      RECT 81.095 1.655 81.265 1.825 ;
      RECT 81.095 7.055 81.265 7.225 ;
      RECT 81.095 7.795 81.265 7.965 ;
      RECT 80.72 2.395 80.89 2.565 ;
      RECT 80.72 6.315 80.89 6.485 ;
      RECT 77.445 1.935 77.615 2.105 ;
      RECT 77.205 2.495 77.375 2.665 ;
      RECT 76.725 2.495 76.895 2.665 ;
      RECT 76.485 1.935 76.655 2.105 ;
      RECT 76.485 3.615 76.655 3.785 ;
      RECT 75.91 6.685 76.08 6.855 ;
      RECT 75.725 2.215 75.895 2.385 ;
      RECT 75.485 3.615 75.655 3.785 ;
      RECT 75.48 7.055 75.65 7.225 ;
      RECT 75.48 7.795 75.65 7.965 ;
      RECT 75.245 2.775 75.415 2.945 ;
      RECT 74.765 2.495 74.935 2.665 ;
      RECT 74.285 2.495 74.455 2.665 ;
      RECT 74.045 1.935 74.215 2.105 ;
      RECT 73.285 2.215 73.455 2.385 ;
      RECT 73.045 3.335 73.215 3.505 ;
      RECT 72.805 2.775 72.975 2.945 ;
      RECT 72.325 2.495 72.495 2.665 ;
      RECT 72.085 1.935 72.255 2.105 ;
      RECT 72.085 3.335 72.255 3.505 ;
      RECT 71.605 3.055 71.775 3.225 ;
      RECT 71.085 2.495 71.255 2.665 ;
      RECT 70.845 3.335 71.015 3.505 ;
      RECT 70.605 1.935 70.775 2.105 ;
      RECT 70.365 2.495 70.535 2.665 ;
      RECT 70.365 3.055 70.535 3.225 ;
      RECT 69.645 1.935 69.815 2.105 ;
      RECT 69.645 3.615 69.815 3.785 ;
      RECT 69.165 3.055 69.335 3.225 ;
      RECT 67.55 7.8 67.72 7.97 ;
      RECT 67.18 2.76 67.35 2.93 ;
      RECT 67.18 5.95 67.35 6.12 ;
      RECT 66.56 0.91 66.73 1.08 ;
      RECT 66.56 2.39 66.73 2.56 ;
      RECT 66.56 6.32 66.73 6.49 ;
      RECT 66.56 7.8 66.73 7.97 ;
      RECT 66.19 2.76 66.36 2.93 ;
      RECT 66.19 5.95 66.36 6.12 ;
      RECT 65.2 2.025 65.37 2.195 ;
      RECT 65.2 6.685 65.37 6.855 ;
      RECT 64.77 0.915 64.94 1.085 ;
      RECT 64.77 1.655 64.94 1.825 ;
      RECT 64.77 7.055 64.94 7.225 ;
      RECT 64.77 7.795 64.94 7.965 ;
      RECT 64.395 2.395 64.565 2.565 ;
      RECT 64.395 6.315 64.565 6.485 ;
      RECT 61.12 1.935 61.29 2.105 ;
      RECT 60.88 2.495 61.05 2.665 ;
      RECT 60.4 2.495 60.57 2.665 ;
      RECT 60.16 1.935 60.33 2.105 ;
      RECT 60.16 3.615 60.33 3.785 ;
      RECT 59.585 6.685 59.755 6.855 ;
      RECT 59.4 2.215 59.57 2.385 ;
      RECT 59.16 3.615 59.33 3.785 ;
      RECT 59.155 7.055 59.325 7.225 ;
      RECT 59.155 7.795 59.325 7.965 ;
      RECT 58.92 2.775 59.09 2.945 ;
      RECT 58.44 2.495 58.61 2.665 ;
      RECT 57.96 2.495 58.13 2.665 ;
      RECT 57.72 1.935 57.89 2.105 ;
      RECT 56.96 2.215 57.13 2.385 ;
      RECT 56.72 3.335 56.89 3.505 ;
      RECT 56.48 2.775 56.65 2.945 ;
      RECT 56 2.495 56.17 2.665 ;
      RECT 55.76 1.935 55.93 2.105 ;
      RECT 55.76 3.335 55.93 3.505 ;
      RECT 55.28 3.055 55.45 3.225 ;
      RECT 54.76 2.495 54.93 2.665 ;
      RECT 54.52 3.335 54.69 3.505 ;
      RECT 54.28 1.935 54.45 2.105 ;
      RECT 54.04 2.495 54.21 2.665 ;
      RECT 54.04 3.055 54.21 3.225 ;
      RECT 53.32 1.935 53.49 2.105 ;
      RECT 53.32 3.615 53.49 3.785 ;
      RECT 52.84 3.055 53.01 3.225 ;
      RECT 51.225 7.8 51.395 7.97 ;
      RECT 50.855 2.76 51.025 2.93 ;
      RECT 50.855 5.95 51.025 6.12 ;
      RECT 50.235 0.91 50.405 1.08 ;
      RECT 50.235 2.39 50.405 2.56 ;
      RECT 50.235 6.32 50.405 6.49 ;
      RECT 50.235 7.8 50.405 7.97 ;
      RECT 49.865 2.76 50.035 2.93 ;
      RECT 49.865 5.95 50.035 6.12 ;
      RECT 48.875 2.025 49.045 2.195 ;
      RECT 48.875 6.685 49.045 6.855 ;
      RECT 48.445 0.915 48.615 1.085 ;
      RECT 48.445 1.655 48.615 1.825 ;
      RECT 48.445 7.055 48.615 7.225 ;
      RECT 48.445 7.795 48.615 7.965 ;
      RECT 48.07 2.395 48.24 2.565 ;
      RECT 48.07 6.315 48.24 6.485 ;
      RECT 44.795 1.935 44.965 2.105 ;
      RECT 44.555 2.495 44.725 2.665 ;
      RECT 44.075 2.495 44.245 2.665 ;
      RECT 43.835 1.935 44.005 2.105 ;
      RECT 43.835 3.615 44.005 3.785 ;
      RECT 43.26 6.685 43.43 6.855 ;
      RECT 43.075 2.215 43.245 2.385 ;
      RECT 42.835 3.615 43.005 3.785 ;
      RECT 42.83 7.055 43 7.225 ;
      RECT 42.83 7.795 43 7.965 ;
      RECT 42.595 2.775 42.765 2.945 ;
      RECT 42.115 2.495 42.285 2.665 ;
      RECT 41.635 2.495 41.805 2.665 ;
      RECT 41.395 1.935 41.565 2.105 ;
      RECT 40.635 2.215 40.805 2.385 ;
      RECT 40.395 3.335 40.565 3.505 ;
      RECT 40.155 2.775 40.325 2.945 ;
      RECT 39.675 2.495 39.845 2.665 ;
      RECT 39.435 1.935 39.605 2.105 ;
      RECT 39.435 3.335 39.605 3.505 ;
      RECT 38.955 3.055 39.125 3.225 ;
      RECT 38.435 2.495 38.605 2.665 ;
      RECT 38.195 3.335 38.365 3.505 ;
      RECT 37.955 1.935 38.125 2.105 ;
      RECT 37.715 2.495 37.885 2.665 ;
      RECT 37.715 3.055 37.885 3.225 ;
      RECT 36.995 1.935 37.165 2.105 ;
      RECT 36.995 3.615 37.165 3.785 ;
      RECT 36.515 3.055 36.685 3.225 ;
      RECT 34.9 7.8 35.07 7.97 ;
      RECT 34.53 2.76 34.7 2.93 ;
      RECT 34.53 5.95 34.7 6.12 ;
      RECT 33.91 0.91 34.08 1.08 ;
      RECT 33.91 2.39 34.08 2.56 ;
      RECT 33.91 6.32 34.08 6.49 ;
      RECT 33.91 7.8 34.08 7.97 ;
      RECT 33.54 2.76 33.71 2.93 ;
      RECT 33.54 5.95 33.71 6.12 ;
      RECT 32.55 2.025 32.72 2.195 ;
      RECT 32.55 6.685 32.72 6.855 ;
      RECT 32.12 0.915 32.29 1.085 ;
      RECT 32.12 1.655 32.29 1.825 ;
      RECT 32.12 7.055 32.29 7.225 ;
      RECT 32.12 7.795 32.29 7.965 ;
      RECT 31.745 2.395 31.915 2.565 ;
      RECT 31.745 6.315 31.915 6.485 ;
      RECT 28.47 1.935 28.64 2.105 ;
      RECT 28.23 2.495 28.4 2.665 ;
      RECT 27.75 2.495 27.92 2.665 ;
      RECT 27.51 1.935 27.68 2.105 ;
      RECT 27.51 3.615 27.68 3.785 ;
      RECT 26.935 6.685 27.105 6.855 ;
      RECT 26.75 2.215 26.92 2.385 ;
      RECT 26.51 3.615 26.68 3.785 ;
      RECT 26.505 7.055 26.675 7.225 ;
      RECT 26.505 7.795 26.675 7.965 ;
      RECT 26.27 2.775 26.44 2.945 ;
      RECT 25.79 2.495 25.96 2.665 ;
      RECT 25.31 2.495 25.48 2.665 ;
      RECT 25.07 1.935 25.24 2.105 ;
      RECT 24.31 2.215 24.48 2.385 ;
      RECT 24.07 3.335 24.24 3.505 ;
      RECT 23.83 2.775 24 2.945 ;
      RECT 23.35 2.495 23.52 2.665 ;
      RECT 23.11 1.935 23.28 2.105 ;
      RECT 23.11 3.335 23.28 3.505 ;
      RECT 22.63 3.055 22.8 3.225 ;
      RECT 22.11 2.495 22.28 2.665 ;
      RECT 21.87 3.335 22.04 3.505 ;
      RECT 21.63 1.935 21.8 2.105 ;
      RECT 21.39 2.495 21.56 2.665 ;
      RECT 21.39 3.055 21.56 3.225 ;
      RECT 20.67 1.935 20.84 2.105 ;
      RECT 20.67 3.615 20.84 3.785 ;
      RECT 20.19 3.055 20.36 3.225 ;
      RECT 18.575 7.8 18.745 7.97 ;
      RECT 18.205 2.76 18.375 2.93 ;
      RECT 18.205 5.95 18.375 6.12 ;
      RECT 17.585 0.91 17.755 1.08 ;
      RECT 17.585 2.39 17.755 2.56 ;
      RECT 17.585 6.32 17.755 6.49 ;
      RECT 17.585 7.8 17.755 7.97 ;
      RECT 17.215 2.76 17.385 2.93 ;
      RECT 17.215 5.95 17.385 6.12 ;
      RECT 16.225 2.025 16.395 2.195 ;
      RECT 16.225 6.685 16.395 6.855 ;
      RECT 15.795 0.915 15.965 1.085 ;
      RECT 15.795 1.655 15.965 1.825 ;
      RECT 15.795 7.055 15.965 7.225 ;
      RECT 15.795 7.795 15.965 7.965 ;
      RECT 15.42 2.395 15.59 2.565 ;
      RECT 15.42 6.315 15.59 6.485 ;
      RECT 12.145 1.935 12.315 2.105 ;
      RECT 11.905 2.495 12.075 2.665 ;
      RECT 11.425 2.495 11.595 2.665 ;
      RECT 11.185 1.935 11.355 2.105 ;
      RECT 11.185 3.615 11.355 3.785 ;
      RECT 10.61 6.685 10.78 6.855 ;
      RECT 10.425 2.215 10.595 2.385 ;
      RECT 10.185 3.615 10.355 3.785 ;
      RECT 10.18 7.055 10.35 7.225 ;
      RECT 10.18 7.795 10.35 7.965 ;
      RECT 9.945 2.775 10.115 2.945 ;
      RECT 9.465 2.495 9.635 2.665 ;
      RECT 8.985 2.495 9.155 2.665 ;
      RECT 8.745 1.935 8.915 2.105 ;
      RECT 7.985 2.215 8.155 2.385 ;
      RECT 7.745 3.335 7.915 3.505 ;
      RECT 7.505 2.775 7.675 2.945 ;
      RECT 7.025 2.495 7.195 2.665 ;
      RECT 6.785 1.935 6.955 2.105 ;
      RECT 6.785 3.335 6.955 3.505 ;
      RECT 6.305 3.055 6.475 3.225 ;
      RECT 5.785 2.495 5.955 2.665 ;
      RECT 5.545 3.335 5.715 3.505 ;
      RECT 5.305 1.935 5.475 2.105 ;
      RECT 5.065 2.495 5.235 2.665 ;
      RECT 5.065 3.055 5.235 3.225 ;
      RECT 4.345 1.935 4.515 2.105 ;
      RECT 4.345 3.615 4.515 3.785 ;
      RECT 3.865 3.055 4.035 3.225 ;
      RECT 1.6 7.055 1.77 7.225 ;
      RECT 1.6 7.795 1.77 7.965 ;
      RECT 1.225 6.315 1.395 6.485 ;
    LAYER li1 ;
      RECT 83.875 5.02 84.045 6.49 ;
      RECT 83.875 6.315 84.05 6.485 ;
      RECT 83.505 1.74 83.675 2.93 ;
      RECT 83.505 1.74 83.975 1.91 ;
      RECT 83.505 6.97 83.975 7.14 ;
      RECT 83.505 5.95 83.675 7.14 ;
      RECT 82.515 1.74 82.685 2.93 ;
      RECT 82.515 1.74 82.985 1.91 ;
      RECT 82.515 6.97 82.985 7.14 ;
      RECT 82.515 5.95 82.685 7.14 ;
      RECT 80.665 2.635 80.835 3.865 ;
      RECT 80.72 0.855 80.89 2.805 ;
      RECT 80.665 0.575 80.835 1.025 ;
      RECT 80.665 7.855 80.835 8.305 ;
      RECT 80.72 6.075 80.89 8.025 ;
      RECT 80.665 5.015 80.835 6.245 ;
      RECT 80.145 0.575 80.315 3.865 ;
      RECT 80.145 2.075 80.55 2.405 ;
      RECT 80.145 1.235 80.55 1.565 ;
      RECT 80.145 5.015 80.315 8.305 ;
      RECT 80.145 7.315 80.55 7.645 ;
      RECT 80.145 6.475 80.55 6.805 ;
      RECT 77.445 1.835 77.615 2.105 ;
      RECT 77.445 1.835 78.175 2.005 ;
      RECT 77.365 3.225 77.695 3.395 ;
      RECT 76.605 3.055 77.615 3.225 ;
      RECT 76.605 2.575 76.775 3.225 ;
      RECT 76.725 2.495 76.895 2.825 ;
      RECT 75.885 3.225 76.215 3.395 ;
      RECT 73.965 3.225 75.255 3.395 ;
      RECT 75.005 3.14 76.135 3.31 ;
      RECT 75.725 2.215 76.135 2.385 ;
      RECT 75.965 1.755 76.135 2.385 ;
      RECT 74.53 5.015 74.7 8.305 ;
      RECT 74.53 7.315 74.935 7.645 ;
      RECT 74.53 6.475 74.935 6.805 ;
      RECT 73.205 2.575 74.535 2.745 ;
      RECT 74.285 2.495 74.455 2.745 ;
      RECT 73.285 2.175 73.455 2.385 ;
      RECT 73.285 2.175 73.775 2.345 ;
      RECT 71.965 3.335 72.255 3.505 ;
      RECT 71.965 2.575 72.135 3.505 ;
      RECT 71.765 2.575 72.135 2.745 ;
      RECT 70.765 2.575 71.255 2.745 ;
      RECT 71.085 2.495 71.255 2.745 ;
      RECT 70.845 3.335 71.255 3.505 ;
      RECT 71.085 3.145 71.255 3.505 ;
      RECT 69.885 3.055 70.535 3.225 ;
      RECT 69.885 2.495 70.055 3.225 ;
      RECT 69.525 3.615 69.815 3.785 ;
      RECT 69.525 2.575 69.695 3.785 ;
      RECT 69.325 2.575 69.695 2.745 ;
      RECT 67.55 5.02 67.72 6.49 ;
      RECT 67.55 6.315 67.725 6.485 ;
      RECT 67.18 1.74 67.35 2.93 ;
      RECT 67.18 1.74 67.65 1.91 ;
      RECT 67.18 6.97 67.65 7.14 ;
      RECT 67.18 5.95 67.35 7.14 ;
      RECT 66.19 1.74 66.36 2.93 ;
      RECT 66.19 1.74 66.66 1.91 ;
      RECT 66.19 6.97 66.66 7.14 ;
      RECT 66.19 5.95 66.36 7.14 ;
      RECT 64.34 2.635 64.51 3.865 ;
      RECT 64.395 0.855 64.565 2.805 ;
      RECT 64.34 0.575 64.51 1.025 ;
      RECT 64.34 7.855 64.51 8.305 ;
      RECT 64.395 6.075 64.565 8.025 ;
      RECT 64.34 5.015 64.51 6.245 ;
      RECT 63.82 0.575 63.99 3.865 ;
      RECT 63.82 2.075 64.225 2.405 ;
      RECT 63.82 1.235 64.225 1.565 ;
      RECT 63.82 5.015 63.99 8.305 ;
      RECT 63.82 7.315 64.225 7.645 ;
      RECT 63.82 6.475 64.225 6.805 ;
      RECT 61.12 1.835 61.29 2.105 ;
      RECT 61.12 1.835 61.85 2.005 ;
      RECT 61.04 3.225 61.37 3.395 ;
      RECT 60.28 3.055 61.29 3.225 ;
      RECT 60.28 2.575 60.45 3.225 ;
      RECT 60.4 2.495 60.57 2.825 ;
      RECT 59.56 3.225 59.89 3.395 ;
      RECT 57.64 3.225 58.93 3.395 ;
      RECT 58.68 3.14 59.81 3.31 ;
      RECT 59.4 2.215 59.81 2.385 ;
      RECT 59.64 1.755 59.81 2.385 ;
      RECT 58.205 5.015 58.375 8.305 ;
      RECT 58.205 7.315 58.61 7.645 ;
      RECT 58.205 6.475 58.61 6.805 ;
      RECT 56.88 2.575 58.21 2.745 ;
      RECT 57.96 2.495 58.13 2.745 ;
      RECT 56.96 2.175 57.13 2.385 ;
      RECT 56.96 2.175 57.45 2.345 ;
      RECT 55.64 3.335 55.93 3.505 ;
      RECT 55.64 2.575 55.81 3.505 ;
      RECT 55.44 2.575 55.81 2.745 ;
      RECT 54.44 2.575 54.93 2.745 ;
      RECT 54.76 2.495 54.93 2.745 ;
      RECT 54.52 3.335 54.93 3.505 ;
      RECT 54.76 3.145 54.93 3.505 ;
      RECT 53.56 3.055 54.21 3.225 ;
      RECT 53.56 2.495 53.73 3.225 ;
      RECT 53.2 3.615 53.49 3.785 ;
      RECT 53.2 2.575 53.37 3.785 ;
      RECT 53 2.575 53.37 2.745 ;
      RECT 51.225 5.02 51.395 6.49 ;
      RECT 51.225 6.315 51.4 6.485 ;
      RECT 50.855 1.74 51.025 2.93 ;
      RECT 50.855 1.74 51.325 1.91 ;
      RECT 50.855 6.97 51.325 7.14 ;
      RECT 50.855 5.95 51.025 7.14 ;
      RECT 49.865 1.74 50.035 2.93 ;
      RECT 49.865 1.74 50.335 1.91 ;
      RECT 49.865 6.97 50.335 7.14 ;
      RECT 49.865 5.95 50.035 7.14 ;
      RECT 48.015 2.635 48.185 3.865 ;
      RECT 48.07 0.855 48.24 2.805 ;
      RECT 48.015 0.575 48.185 1.025 ;
      RECT 48.015 7.855 48.185 8.305 ;
      RECT 48.07 6.075 48.24 8.025 ;
      RECT 48.015 5.015 48.185 6.245 ;
      RECT 47.495 0.575 47.665 3.865 ;
      RECT 47.495 2.075 47.9 2.405 ;
      RECT 47.495 1.235 47.9 1.565 ;
      RECT 47.495 5.015 47.665 8.305 ;
      RECT 47.495 7.315 47.9 7.645 ;
      RECT 47.495 6.475 47.9 6.805 ;
      RECT 44.795 1.835 44.965 2.105 ;
      RECT 44.795 1.835 45.525 2.005 ;
      RECT 44.715 3.225 45.045 3.395 ;
      RECT 43.955 3.055 44.965 3.225 ;
      RECT 43.955 2.575 44.125 3.225 ;
      RECT 44.075 2.495 44.245 2.825 ;
      RECT 43.235 3.225 43.565 3.395 ;
      RECT 41.315 3.225 42.605 3.395 ;
      RECT 42.355 3.14 43.485 3.31 ;
      RECT 43.075 2.215 43.485 2.385 ;
      RECT 43.315 1.755 43.485 2.385 ;
      RECT 41.88 5.015 42.05 8.305 ;
      RECT 41.88 7.315 42.285 7.645 ;
      RECT 41.88 6.475 42.285 6.805 ;
      RECT 40.555 2.575 41.885 2.745 ;
      RECT 41.635 2.495 41.805 2.745 ;
      RECT 40.635 2.175 40.805 2.385 ;
      RECT 40.635 2.175 41.125 2.345 ;
      RECT 39.315 3.335 39.605 3.505 ;
      RECT 39.315 2.575 39.485 3.505 ;
      RECT 39.115 2.575 39.485 2.745 ;
      RECT 38.115 2.575 38.605 2.745 ;
      RECT 38.435 2.495 38.605 2.745 ;
      RECT 38.195 3.335 38.605 3.505 ;
      RECT 38.435 3.145 38.605 3.505 ;
      RECT 37.235 3.055 37.885 3.225 ;
      RECT 37.235 2.495 37.405 3.225 ;
      RECT 36.875 3.615 37.165 3.785 ;
      RECT 36.875 2.575 37.045 3.785 ;
      RECT 36.675 2.575 37.045 2.745 ;
      RECT 34.9 5.02 35.07 6.49 ;
      RECT 34.9 6.315 35.075 6.485 ;
      RECT 34.53 1.74 34.7 2.93 ;
      RECT 34.53 1.74 35 1.91 ;
      RECT 34.53 6.97 35 7.14 ;
      RECT 34.53 5.95 34.7 7.14 ;
      RECT 33.54 1.74 33.71 2.93 ;
      RECT 33.54 1.74 34.01 1.91 ;
      RECT 33.54 6.97 34.01 7.14 ;
      RECT 33.54 5.95 33.71 7.14 ;
      RECT 31.69 2.635 31.86 3.865 ;
      RECT 31.745 0.855 31.915 2.805 ;
      RECT 31.69 0.575 31.86 1.025 ;
      RECT 31.69 7.855 31.86 8.305 ;
      RECT 31.745 6.075 31.915 8.025 ;
      RECT 31.69 5.015 31.86 6.245 ;
      RECT 31.17 0.575 31.34 3.865 ;
      RECT 31.17 2.075 31.575 2.405 ;
      RECT 31.17 1.235 31.575 1.565 ;
      RECT 31.17 5.015 31.34 8.305 ;
      RECT 31.17 7.315 31.575 7.645 ;
      RECT 31.17 6.475 31.575 6.805 ;
      RECT 28.47 1.835 28.64 2.105 ;
      RECT 28.47 1.835 29.2 2.005 ;
      RECT 28.39 3.225 28.72 3.395 ;
      RECT 27.63 3.055 28.64 3.225 ;
      RECT 27.63 2.575 27.8 3.225 ;
      RECT 27.75 2.495 27.92 2.825 ;
      RECT 26.91 3.225 27.24 3.395 ;
      RECT 24.99 3.225 26.28 3.395 ;
      RECT 26.03 3.14 27.16 3.31 ;
      RECT 26.75 2.215 27.16 2.385 ;
      RECT 26.99 1.755 27.16 2.385 ;
      RECT 25.555 5.015 25.725 8.305 ;
      RECT 25.555 7.315 25.96 7.645 ;
      RECT 25.555 6.475 25.96 6.805 ;
      RECT 24.23 2.575 25.56 2.745 ;
      RECT 25.31 2.495 25.48 2.745 ;
      RECT 24.31 2.175 24.48 2.385 ;
      RECT 24.31 2.175 24.8 2.345 ;
      RECT 22.99 3.335 23.28 3.505 ;
      RECT 22.99 2.575 23.16 3.505 ;
      RECT 22.79 2.575 23.16 2.745 ;
      RECT 21.79 2.575 22.28 2.745 ;
      RECT 22.11 2.495 22.28 2.745 ;
      RECT 21.87 3.335 22.28 3.505 ;
      RECT 22.11 3.145 22.28 3.505 ;
      RECT 20.91 3.055 21.56 3.225 ;
      RECT 20.91 2.495 21.08 3.225 ;
      RECT 20.55 3.615 20.84 3.785 ;
      RECT 20.55 2.575 20.72 3.785 ;
      RECT 20.35 2.575 20.72 2.745 ;
      RECT 18.575 5.02 18.745 6.49 ;
      RECT 18.575 6.315 18.75 6.485 ;
      RECT 18.205 1.74 18.375 2.93 ;
      RECT 18.205 1.74 18.675 1.91 ;
      RECT 18.205 6.97 18.675 7.14 ;
      RECT 18.205 5.95 18.375 7.14 ;
      RECT 17.215 1.74 17.385 2.93 ;
      RECT 17.215 1.74 17.685 1.91 ;
      RECT 17.215 6.97 17.685 7.14 ;
      RECT 17.215 5.95 17.385 7.14 ;
      RECT 15.365 2.635 15.535 3.865 ;
      RECT 15.42 0.855 15.59 2.805 ;
      RECT 15.365 0.575 15.535 1.025 ;
      RECT 15.365 7.855 15.535 8.305 ;
      RECT 15.42 6.075 15.59 8.025 ;
      RECT 15.365 5.015 15.535 6.245 ;
      RECT 14.845 0.575 15.015 3.865 ;
      RECT 14.845 2.075 15.25 2.405 ;
      RECT 14.845 1.235 15.25 1.565 ;
      RECT 14.845 5.015 15.015 8.305 ;
      RECT 14.845 7.315 15.25 7.645 ;
      RECT 14.845 6.475 15.25 6.805 ;
      RECT 12.145 1.835 12.315 2.105 ;
      RECT 12.145 1.835 12.875 2.005 ;
      RECT 12.065 3.225 12.395 3.395 ;
      RECT 11.305 3.055 12.315 3.225 ;
      RECT 11.305 2.575 11.475 3.225 ;
      RECT 11.425 2.495 11.595 2.825 ;
      RECT 10.585 3.225 10.915 3.395 ;
      RECT 8.665 3.225 9.955 3.395 ;
      RECT 9.705 3.14 10.835 3.31 ;
      RECT 10.425 2.215 10.835 2.385 ;
      RECT 10.665 1.755 10.835 2.385 ;
      RECT 9.23 5.015 9.4 8.305 ;
      RECT 9.23 7.315 9.635 7.645 ;
      RECT 9.23 6.475 9.635 6.805 ;
      RECT 7.905 2.575 9.235 2.745 ;
      RECT 8.985 2.495 9.155 2.745 ;
      RECT 7.985 2.175 8.155 2.385 ;
      RECT 7.985 2.175 8.475 2.345 ;
      RECT 6.665 3.335 6.955 3.505 ;
      RECT 6.665 2.575 6.835 3.505 ;
      RECT 6.465 2.575 6.835 2.745 ;
      RECT 5.465 2.575 5.955 2.745 ;
      RECT 5.785 2.495 5.955 2.745 ;
      RECT 5.545 3.335 5.955 3.505 ;
      RECT 5.785 3.145 5.955 3.505 ;
      RECT 4.585 3.055 5.235 3.225 ;
      RECT 4.585 2.495 4.755 3.225 ;
      RECT 4.225 3.615 4.515 3.785 ;
      RECT 4.225 2.575 4.395 3.785 ;
      RECT 4.025 2.575 4.395 2.745 ;
      RECT 1.17 7.855 1.34 8.305 ;
      RECT 1.225 6.075 1.395 8.025 ;
      RECT 1.17 5.015 1.34 6.245 ;
      RECT 0.65 5.015 0.82 8.305 ;
      RECT 0.65 7.315 1.055 7.645 ;
      RECT 0.65 6.475 1.055 6.805 ;
      RECT 83.875 7.8 84.045 8.31 ;
      RECT 82.885 0.57 83.055 1.08 ;
      RECT 82.885 2.39 83.055 3.86 ;
      RECT 82.885 5.02 83.055 6.49 ;
      RECT 82.885 7.8 83.055 8.31 ;
      RECT 81.525 0.575 81.695 3.865 ;
      RECT 81.525 5.015 81.695 8.305 ;
      RECT 81.095 0.575 81.265 1.085 ;
      RECT 81.095 1.655 81.265 3.865 ;
      RECT 81.095 5.015 81.265 7.225 ;
      RECT 81.095 7.795 81.265 8.305 ;
      RECT 77.205 2.495 77.375 2.825 ;
      RECT 76.485 1.755 76.655 2.105 ;
      RECT 76.485 3.485 76.655 3.815 ;
      RECT 75.91 5.015 76.08 8.305 ;
      RECT 75.485 3.485 75.655 3.815 ;
      RECT 75.48 5.015 75.65 7.225 ;
      RECT 75.48 7.795 75.65 8.305 ;
      RECT 75.245 2.495 75.415 2.945 ;
      RECT 74.765 2.495 74.935 2.825 ;
      RECT 74.045 1.755 74.215 2.105 ;
      RECT 73.045 3.145 73.215 3.505 ;
      RECT 72.805 2.495 72.975 2.945 ;
      RECT 72.325 2.495 72.495 2.825 ;
      RECT 72.085 1.755 72.255 2.105 ;
      RECT 71.605 3.055 71.775 3.475 ;
      RECT 70.605 1.755 70.775 2.105 ;
      RECT 70.365 2.495 70.535 2.825 ;
      RECT 69.645 1.755 69.815 2.105 ;
      RECT 69.165 3.055 69.335 3.475 ;
      RECT 67.55 7.8 67.72 8.31 ;
      RECT 66.56 0.57 66.73 1.08 ;
      RECT 66.56 2.39 66.73 3.86 ;
      RECT 66.56 5.02 66.73 6.49 ;
      RECT 66.56 7.8 66.73 8.31 ;
      RECT 65.2 0.575 65.37 3.865 ;
      RECT 65.2 5.015 65.37 8.305 ;
      RECT 64.77 0.575 64.94 1.085 ;
      RECT 64.77 1.655 64.94 3.865 ;
      RECT 64.77 5.015 64.94 7.225 ;
      RECT 64.77 7.795 64.94 8.305 ;
      RECT 60.88 2.495 61.05 2.825 ;
      RECT 60.16 1.755 60.33 2.105 ;
      RECT 60.16 3.485 60.33 3.815 ;
      RECT 59.585 5.015 59.755 8.305 ;
      RECT 59.16 3.485 59.33 3.815 ;
      RECT 59.155 5.015 59.325 7.225 ;
      RECT 59.155 7.795 59.325 8.305 ;
      RECT 58.92 2.495 59.09 2.945 ;
      RECT 58.44 2.495 58.61 2.825 ;
      RECT 57.72 1.755 57.89 2.105 ;
      RECT 56.72 3.145 56.89 3.505 ;
      RECT 56.48 2.495 56.65 2.945 ;
      RECT 56 2.495 56.17 2.825 ;
      RECT 55.76 1.755 55.93 2.105 ;
      RECT 55.28 3.055 55.45 3.475 ;
      RECT 54.28 1.755 54.45 2.105 ;
      RECT 54.04 2.495 54.21 2.825 ;
      RECT 53.32 1.755 53.49 2.105 ;
      RECT 52.84 3.055 53.01 3.475 ;
      RECT 51.225 7.8 51.395 8.31 ;
      RECT 50.235 0.57 50.405 1.08 ;
      RECT 50.235 2.39 50.405 3.86 ;
      RECT 50.235 5.02 50.405 6.49 ;
      RECT 50.235 7.8 50.405 8.31 ;
      RECT 48.875 0.575 49.045 3.865 ;
      RECT 48.875 5.015 49.045 8.305 ;
      RECT 48.445 0.575 48.615 1.085 ;
      RECT 48.445 1.655 48.615 3.865 ;
      RECT 48.445 5.015 48.615 7.225 ;
      RECT 48.445 7.795 48.615 8.305 ;
      RECT 44.555 2.495 44.725 2.825 ;
      RECT 43.835 1.755 44.005 2.105 ;
      RECT 43.835 3.485 44.005 3.815 ;
      RECT 43.26 5.015 43.43 8.305 ;
      RECT 42.835 3.485 43.005 3.815 ;
      RECT 42.83 5.015 43 7.225 ;
      RECT 42.83 7.795 43 8.305 ;
      RECT 42.595 2.495 42.765 2.945 ;
      RECT 42.115 2.495 42.285 2.825 ;
      RECT 41.395 1.755 41.565 2.105 ;
      RECT 40.395 3.145 40.565 3.505 ;
      RECT 40.155 2.495 40.325 2.945 ;
      RECT 39.675 2.495 39.845 2.825 ;
      RECT 39.435 1.755 39.605 2.105 ;
      RECT 38.955 3.055 39.125 3.475 ;
      RECT 37.955 1.755 38.125 2.105 ;
      RECT 37.715 2.495 37.885 2.825 ;
      RECT 36.995 1.755 37.165 2.105 ;
      RECT 36.515 3.055 36.685 3.475 ;
      RECT 34.9 7.8 35.07 8.31 ;
      RECT 33.91 0.57 34.08 1.08 ;
      RECT 33.91 2.39 34.08 3.86 ;
      RECT 33.91 5.02 34.08 6.49 ;
      RECT 33.91 7.8 34.08 8.31 ;
      RECT 32.55 0.575 32.72 3.865 ;
      RECT 32.55 5.015 32.72 8.305 ;
      RECT 32.12 0.575 32.29 1.085 ;
      RECT 32.12 1.655 32.29 3.865 ;
      RECT 32.12 5.015 32.29 7.225 ;
      RECT 32.12 7.795 32.29 8.305 ;
      RECT 28.23 2.495 28.4 2.825 ;
      RECT 27.51 1.755 27.68 2.105 ;
      RECT 27.51 3.485 27.68 3.815 ;
      RECT 26.935 5.015 27.105 8.305 ;
      RECT 26.51 3.485 26.68 3.815 ;
      RECT 26.505 5.015 26.675 7.225 ;
      RECT 26.505 7.795 26.675 8.305 ;
      RECT 26.27 2.495 26.44 2.945 ;
      RECT 25.79 2.495 25.96 2.825 ;
      RECT 25.07 1.755 25.24 2.105 ;
      RECT 24.07 3.145 24.24 3.505 ;
      RECT 23.83 2.495 24 2.945 ;
      RECT 23.35 2.495 23.52 2.825 ;
      RECT 23.11 1.755 23.28 2.105 ;
      RECT 22.63 3.055 22.8 3.475 ;
      RECT 21.63 1.755 21.8 2.105 ;
      RECT 21.39 2.495 21.56 2.825 ;
      RECT 20.67 1.755 20.84 2.105 ;
      RECT 20.19 3.055 20.36 3.475 ;
      RECT 18.575 7.8 18.745 8.31 ;
      RECT 17.585 0.57 17.755 1.08 ;
      RECT 17.585 2.39 17.755 3.86 ;
      RECT 17.585 5.02 17.755 6.49 ;
      RECT 17.585 7.8 17.755 8.31 ;
      RECT 16.225 0.575 16.395 3.865 ;
      RECT 16.225 5.015 16.395 8.305 ;
      RECT 15.795 0.575 15.965 1.085 ;
      RECT 15.795 1.655 15.965 3.865 ;
      RECT 15.795 5.015 15.965 7.225 ;
      RECT 15.795 7.795 15.965 8.305 ;
      RECT 11.905 2.495 12.075 2.825 ;
      RECT 11.185 1.755 11.355 2.105 ;
      RECT 11.185 3.485 11.355 3.815 ;
      RECT 10.61 5.015 10.78 8.305 ;
      RECT 10.185 3.485 10.355 3.815 ;
      RECT 10.18 5.015 10.35 7.225 ;
      RECT 10.18 7.795 10.35 8.305 ;
      RECT 9.945 2.495 10.115 2.945 ;
      RECT 9.465 2.495 9.635 2.825 ;
      RECT 8.745 1.755 8.915 2.105 ;
      RECT 7.745 3.145 7.915 3.505 ;
      RECT 7.505 2.495 7.675 2.945 ;
      RECT 7.025 2.495 7.195 2.825 ;
      RECT 6.785 1.755 6.955 2.105 ;
      RECT 6.305 3.055 6.475 3.475 ;
      RECT 5.305 1.755 5.475 2.105 ;
      RECT 5.065 2.495 5.235 2.825 ;
      RECT 4.345 1.755 4.515 2.105 ;
      RECT 3.865 3.055 4.035 3.475 ;
      RECT 1.6 5.015 1.77 7.225 ;
      RECT 1.6 7.795 1.77 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r1 ;
  SIZE 95.595 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 20.815 0.915 20.985 1.085 ;
        RECT 20.81 0.91 20.98 1.08 ;
        RECT 20.81 2.39 20.98 2.56 ;
      LAYER li1 ;
        RECT 20.815 0.915 20.985 1.085 ;
        RECT 20.81 0.57 20.98 1.08 ;
        RECT 20.81 2.39 20.98 3.86 ;
      LAYER met1 ;
        RECT 20.75 2.36 21.04 2.59 ;
        RECT 20.75 0.88 21.04 1.11 ;
        RECT 20.81 0.88 20.98 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 39.375 0.915 39.545 1.085 ;
        RECT 39.37 0.91 39.54 1.08 ;
        RECT 39.37 2.39 39.54 2.56 ;
      LAYER li1 ;
        RECT 39.375 0.915 39.545 1.085 ;
        RECT 39.37 0.57 39.54 1.08 ;
        RECT 39.37 2.39 39.54 3.86 ;
      LAYER met1 ;
        RECT 39.31 2.36 39.6 2.59 ;
        RECT 39.31 0.88 39.6 1.11 ;
        RECT 39.37 0.88 39.54 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 57.935 0.915 58.105 1.085 ;
        RECT 57.93 0.91 58.1 1.08 ;
        RECT 57.93 2.39 58.1 2.56 ;
      LAYER li1 ;
        RECT 57.935 0.915 58.105 1.085 ;
        RECT 57.93 0.57 58.1 1.08 ;
        RECT 57.93 2.39 58.1 3.86 ;
      LAYER met1 ;
        RECT 57.87 2.36 58.16 2.59 ;
        RECT 57.87 0.88 58.16 1.11 ;
        RECT 57.93 0.88 58.1 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 76.495 0.915 76.665 1.085 ;
        RECT 76.49 0.91 76.66 1.08 ;
        RECT 76.49 2.39 76.66 2.56 ;
      LAYER li1 ;
        RECT 76.495 0.915 76.665 1.085 ;
        RECT 76.49 0.57 76.66 1.08 ;
        RECT 76.49 2.39 76.66 3.86 ;
      LAYER met1 ;
        RECT 76.43 2.36 76.72 2.59 ;
        RECT 76.43 0.88 76.72 1.11 ;
        RECT 76.49 0.88 76.66 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 95.055 0.915 95.225 1.085 ;
        RECT 95.05 0.91 95.22 1.08 ;
        RECT 95.05 2.39 95.22 2.56 ;
      LAYER li1 ;
        RECT 95.055 0.915 95.225 1.085 ;
        RECT 95.05 0.57 95.22 1.08 ;
        RECT 95.05 2.39 95.22 3.86 ;
      LAYER met1 ;
        RECT 94.99 2.36 95.28 2.59 ;
        RECT 94.99 0.88 95.28 1.11 ;
        RECT 95.05 0.88 95.22 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 16.66 1.66 16.83 2.935 ;
        RECT 16.66 5.945 16.83 7.22 ;
        RECT 11.045 5.945 11.215 7.22 ;
      LAYER met2 ;
        RECT 16.585 2.705 16.925 3.055 ;
        RECT 16.575 5.845 16.915 6.195 ;
        RECT 16.66 2.705 16.83 6.195 ;
      LAYER met1 ;
        RECT 16.585 2.765 17.06 2.935 ;
        RECT 16.585 2.705 16.925 3.055 ;
        RECT 10.985 5.945 17.06 6.115 ;
        RECT 16.575 5.845 16.915 6.195 ;
        RECT 10.985 5.915 11.275 6.145 ;
      LAYER mcon ;
        RECT 11.045 5.945 11.215 6.115 ;
        RECT 16.66 5.945 16.83 6.115 ;
        RECT 16.66 2.765 16.83 2.935 ;
      LAYER via1 ;
        RECT 16.675 5.945 16.825 6.095 ;
        RECT 16.685 2.805 16.835 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 35.22 1.66 35.39 2.935 ;
        RECT 35.22 5.945 35.39 7.22 ;
        RECT 29.605 5.945 29.775 7.22 ;
      LAYER met2 ;
        RECT 35.145 2.705 35.485 3.055 ;
        RECT 35.135 5.845 35.475 6.195 ;
        RECT 35.22 2.705 35.39 6.195 ;
      LAYER met1 ;
        RECT 35.145 2.765 35.62 2.935 ;
        RECT 35.145 2.705 35.485 3.055 ;
        RECT 29.545 5.945 35.62 6.115 ;
        RECT 35.135 5.845 35.475 6.195 ;
        RECT 29.545 5.915 29.835 6.145 ;
      LAYER mcon ;
        RECT 29.605 5.945 29.775 6.115 ;
        RECT 35.22 5.945 35.39 6.115 ;
        RECT 35.22 2.765 35.39 2.935 ;
      LAYER via1 ;
        RECT 35.235 5.945 35.385 6.095 ;
        RECT 35.245 2.805 35.395 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 53.78 1.66 53.95 2.935 ;
        RECT 53.78 5.945 53.95 7.22 ;
        RECT 48.165 5.945 48.335 7.22 ;
      LAYER met2 ;
        RECT 53.705 2.705 54.045 3.055 ;
        RECT 53.695 5.845 54.035 6.195 ;
        RECT 53.78 2.705 53.95 6.195 ;
      LAYER met1 ;
        RECT 53.705 2.765 54.18 2.935 ;
        RECT 53.705 2.705 54.045 3.055 ;
        RECT 48.105 5.945 54.18 6.115 ;
        RECT 53.695 5.845 54.035 6.195 ;
        RECT 48.105 5.915 48.395 6.145 ;
      LAYER mcon ;
        RECT 48.165 5.945 48.335 6.115 ;
        RECT 53.78 5.945 53.95 6.115 ;
        RECT 53.78 2.765 53.95 2.935 ;
      LAYER via1 ;
        RECT 53.795 5.945 53.945 6.095 ;
        RECT 53.805 2.805 53.955 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 72.34 1.66 72.51 2.935 ;
        RECT 72.34 5.945 72.51 7.22 ;
        RECT 66.725 5.945 66.895 7.22 ;
      LAYER met2 ;
        RECT 72.265 2.705 72.605 3.055 ;
        RECT 72.255 5.845 72.595 6.195 ;
        RECT 72.34 2.705 72.51 6.195 ;
      LAYER met1 ;
        RECT 72.265 2.765 72.74 2.935 ;
        RECT 72.265 2.705 72.605 3.055 ;
        RECT 66.665 5.945 72.74 6.115 ;
        RECT 72.255 5.845 72.595 6.195 ;
        RECT 66.665 5.915 66.955 6.145 ;
      LAYER mcon ;
        RECT 66.725 5.945 66.895 6.115 ;
        RECT 72.34 5.945 72.51 6.115 ;
        RECT 72.34 2.765 72.51 2.935 ;
      LAYER via1 ;
        RECT 72.355 5.945 72.505 6.095 ;
        RECT 72.365 2.805 72.515 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 90.9 1.66 91.07 2.935 ;
        RECT 90.9 5.945 91.07 7.22 ;
        RECT 85.285 5.945 85.455 7.22 ;
      LAYER met2 ;
        RECT 90.825 2.705 91.165 3.055 ;
        RECT 90.815 5.845 91.155 6.195 ;
        RECT 90.9 2.705 91.07 6.195 ;
      LAYER met1 ;
        RECT 90.825 2.765 91.3 2.935 ;
        RECT 90.825 2.705 91.165 3.055 ;
        RECT 85.225 5.945 91.3 6.115 ;
        RECT 90.815 5.845 91.155 6.195 ;
        RECT 85.225 5.915 85.515 6.145 ;
      LAYER mcon ;
        RECT 85.285 5.945 85.455 6.115 ;
        RECT 90.9 5.945 91.07 6.115 ;
        RECT 90.9 2.765 91.07 2.935 ;
      LAYER via1 ;
        RECT 90.915 5.945 91.065 6.095 ;
        RECT 90.925 2.805 91.075 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 5.945 0.4 7.22 ;
      LAYER met1 ;
        RECT 0.17 5.945 0.63 6.115 ;
        RECT 0.17 5.915 0.46 6.145 ;
      LAYER mcon ;
        RECT 0.23 5.945 0.4 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 12.315 7.095 13.32 7.395 ;
        RECT 13.02 4.405 13.32 7.395 ;
        RECT 0 4.405 13.32 4.705 ;
        RECT 12.315 7.055 12.69 7.425 ;
        RECT 7.67 2.415 8.4 2.745 ;
        RECT 7.695 2.415 7.995 4.705 ;
        RECT 6.23 2.975 6.96 3.305 ;
        RECT 6.26 2.975 6.56 4.705 ;
        RECT 0 4.145 5.26 4.75 ;
        RECT 4.12 2.415 4.85 2.745 ;
        RECT 3.19 2.42 4.85 2.72 ;
        RECT 3.19 2.42 3.49 4.75 ;
      LAYER li1 ;
        RECT 77.78 4.135 95.595 4.745 ;
        RECT 93.46 4.13 95.44 4.75 ;
        RECT 94.62 3.4 94.79 5.48 ;
        RECT 93.63 3.4 93.8 5.48 ;
        RECT 90.89 3.405 91.06 5.475 ;
        RECT 87.87 3.635 88.04 4.745 ;
        RECT 85.43 3.635 85.6 4.745 ;
        RECT 85.275 4.135 85.445 5.475 ;
        RECT 83.47 3.635 83.64 4.745 ;
        RECT 82.51 3.635 82.68 4.745 ;
        RECT 80.55 3.635 80.72 4.745 ;
        RECT 79.55 3.635 79.72 4.745 ;
        RECT 77.035 4.145 79.5 4.75 ;
        RECT 78.59 3.635 78.76 4.75 ;
        RECT 59.22 4.135 77.035 4.745 ;
        RECT 74.9 4.13 76.88 4.75 ;
        RECT 76.06 3.4 76.23 5.48 ;
        RECT 75.07 3.4 75.24 5.48 ;
        RECT 72.33 3.405 72.5 5.475 ;
        RECT 69.31 3.635 69.48 4.745 ;
        RECT 66.87 3.635 67.04 4.745 ;
        RECT 66.715 4.135 66.885 5.475 ;
        RECT 64.91 3.635 65.08 4.745 ;
        RECT 63.95 3.635 64.12 4.745 ;
        RECT 61.99 3.635 62.16 4.745 ;
        RECT 60.99 3.635 61.16 4.745 ;
        RECT 58.475 4.145 60.94 4.75 ;
        RECT 60.03 3.635 60.2 4.75 ;
        RECT 40.66 4.135 58.475 4.745 ;
        RECT 56.34 4.13 58.32 4.75 ;
        RECT 57.5 3.4 57.67 5.48 ;
        RECT 56.51 3.4 56.68 5.48 ;
        RECT 53.77 3.405 53.94 5.475 ;
        RECT 50.75 3.635 50.92 4.745 ;
        RECT 48.31 3.635 48.48 4.745 ;
        RECT 48.155 4.135 48.325 5.475 ;
        RECT 46.35 3.635 46.52 4.745 ;
        RECT 45.39 3.635 45.56 4.745 ;
        RECT 43.43 3.635 43.6 4.745 ;
        RECT 42.43 3.635 42.6 4.745 ;
        RECT 39.915 4.145 42.38 4.75 ;
        RECT 41.47 3.635 41.64 4.75 ;
        RECT 22.1 4.135 39.915 4.745 ;
        RECT 37.78 4.13 39.76 4.75 ;
        RECT 38.94 3.4 39.11 5.48 ;
        RECT 37.95 3.4 38.12 5.48 ;
        RECT 35.21 3.405 35.38 5.475 ;
        RECT 32.19 3.635 32.36 4.745 ;
        RECT 29.75 3.635 29.92 4.745 ;
        RECT 29.595 4.135 29.765 5.475 ;
        RECT 27.79 3.635 27.96 4.745 ;
        RECT 26.83 3.635 27 4.745 ;
        RECT 24.87 3.635 25.04 4.745 ;
        RECT 23.87 3.635 24.04 4.745 ;
        RECT 21.355 4.145 23.82 4.75 ;
        RECT 22.91 3.635 23.08 4.75 ;
        RECT 3.54 4.135 21.355 4.745 ;
        RECT 19.22 4.13 21.2 4.75 ;
        RECT 20.38 3.4 20.55 5.48 ;
        RECT 19.39 3.4 19.56 5.48 ;
        RECT 16.65 3.405 16.82 5.475 ;
        RECT 13.63 3.635 13.8 4.745 ;
        RECT 11.19 3.635 11.36 4.745 ;
        RECT 11.035 4.135 11.205 5.475 ;
        RECT 9.23 3.635 9.4 4.745 ;
        RECT 8.27 3.635 8.44 4.745 ;
        RECT 6.31 3.635 6.48 4.745 ;
        RECT 5.31 3.635 5.48 4.745 ;
        RECT 0 4.44 5.26 4.75 ;
        RECT 4.35 3.635 4.52 4.75 ;
        RECT 1.955 4.145 95.595 4.745 ;
        RECT 2.03 4.145 2.2 8.305 ;
        RECT 0 4.145 95.595 4.34 ;
        RECT 0 4.145 1.785 4.75 ;
        RECT 0.22 4.145 0.39 5.475 ;
        RECT 12.415 5.015 12.585 7.225 ;
        RECT 12.415 7.795 12.585 8.305 ;
        RECT 8.99 2.495 9.16 2.825 ;
        RECT 8.27 2.575 8.76 2.745 ;
        RECT 8.27 2.575 8.44 3.225 ;
        RECT 7.43 2.575 7.92 2.745 ;
        RECT 7.75 2.495 7.92 2.745 ;
        RECT 6.55 2.495 6.72 2.945 ;
        RECT 5.745 2.575 6.32 2.745 ;
        RECT 5.745 2.495 5.915 2.745 ;
        RECT 4.59 2.495 4.76 2.825 ;
      LAYER met2 ;
        RECT 12.315 7.055 12.69 7.425 ;
        RECT 8.225 2.98 8.485 3.3 ;
        RECT 5.905 3.07 8.485 3.21 ;
        RECT 6.255 2.955 6.535 3.325 ;
        RECT 5.905 2.98 6.535 3.3 ;
        RECT 7.695 2.42 8.225 2.74 ;
        RECT 7.695 2.395 7.975 2.765 ;
        RECT 4.295 2.395 4.575 2.765 ;
        RECT 1.68 4.265 2.06 4.645 ;
      LAYER met1 ;
        RECT 77.78 4.135 95.595 4.745 ;
        RECT 93.46 4.13 95.44 4.75 ;
        RECT 77.78 3.98 89.74 4.745 ;
        RECT 77.035 4.145 79.5 4.75 ;
        RECT 59.22 4.135 77.035 4.745 ;
        RECT 74.9 4.13 76.88 4.75 ;
        RECT 59.22 3.98 71.18 4.745 ;
        RECT 58.475 4.145 60.94 4.75 ;
        RECT 40.66 4.135 58.475 4.745 ;
        RECT 56.34 4.13 58.32 4.75 ;
        RECT 40.66 3.98 52.62 4.745 ;
        RECT 39.915 4.145 42.38 4.75 ;
        RECT 22.1 4.135 39.915 4.745 ;
        RECT 37.78 4.13 39.76 4.75 ;
        RECT 22.1 3.98 34.06 4.745 ;
        RECT 21.355 4.145 23.82 4.75 ;
        RECT 3.54 4.135 21.355 4.745 ;
        RECT 19.22 4.13 21.2 4.75 ;
        RECT 3.54 3.98 15.5 4.745 ;
        RECT 0 4.145 5.26 4.75 ;
        RECT 12.315 7.055 12.695 7.425 ;
        RECT 12.355 7.765 12.645 7.995 ;
        RECT 12.355 7.025 12.645 7.425 ;
        RECT 12.415 7.025 12.585 7.995 ;
        RECT 8.93 2.465 9.22 2.695 ;
        RECT 7.69 2.51 9.22 2.65 ;
        RECT 7.935 2.45 8.255 2.71 ;
        RECT 7.69 2.465 8.255 2.695 ;
        RECT 8.195 3.01 8.515 3.27 ;
        RECT 6.49 2.745 6.78 2.975 ;
        RECT 5.875 3.01 6.705 3.15 ;
        RECT 6.49 2.745 6.705 3.15 ;
        RECT 5.875 3.01 6.195 3.27 ;
        RECT 5.685 2.465 5.975 2.695 ;
        RECT 5.085 2.37 5.725 2.51 ;
        RECT 5.585 2.465 5.975 2.65 ;
        RECT 4.275 2.55 5.225 2.69 ;
        RECT 5.085 2.37 5.225 2.69 ;
        RECT 4.275 2.465 4.82 2.695 ;
        RECT 4.275 2.45 4.595 2.71 ;
        RECT 1.97 6.655 2.26 6.885 ;
        RECT 1.8 6.685 2.26 6.855 ;
      LAYER via2 ;
        RECT 1.77 4.355 1.97 4.555 ;
        RECT 4.335 2.48 4.535 2.68 ;
        RECT 6.295 3.04 6.495 3.24 ;
        RECT 7.735 2.48 7.935 2.68 ;
        RECT 12.4 7.14 12.6 7.34 ;
      LAYER mcon ;
        RECT 2.03 6.685 2.2 6.855 ;
        RECT 2.34 4.545 2.51 4.715 ;
        RECT 3.685 4.135 3.855 4.305 ;
        RECT 4.145 4.135 4.315 4.305 ;
        RECT 4.59 2.495 4.76 2.665 ;
        RECT 4.605 4.135 4.775 4.305 ;
        RECT 5.065 4.135 5.235 4.305 ;
        RECT 5.525 4.135 5.695 4.305 ;
        RECT 5.745 2.495 5.915 2.665 ;
        RECT 5.985 4.135 6.155 4.305 ;
        RECT 6.445 4.135 6.615 4.305 ;
        RECT 6.55 2.775 6.72 2.945 ;
        RECT 6.905 4.135 7.075 4.305 ;
        RECT 7.365 4.135 7.535 4.305 ;
        RECT 7.75 2.495 7.92 2.665 ;
        RECT 7.825 4.135 7.995 4.305 ;
        RECT 8.27 3.055 8.44 3.225 ;
        RECT 8.285 4.135 8.455 4.305 ;
        RECT 8.745 4.135 8.915 4.305 ;
        RECT 8.99 2.495 9.16 2.665 ;
        RECT 9.205 4.135 9.375 4.305 ;
        RECT 9.665 4.135 9.835 4.305 ;
        RECT 10.125 4.135 10.295 4.305 ;
        RECT 10.585 4.135 10.755 4.305 ;
        RECT 11.045 4.135 11.215 4.305 ;
        RECT 11.505 4.135 11.675 4.305 ;
        RECT 11.965 4.135 12.135 4.305 ;
        RECT 12.415 7.795 12.585 7.965 ;
        RECT 12.415 7.055 12.585 7.225 ;
        RECT 12.425 4.135 12.595 4.305 ;
        RECT 12.885 4.135 13.055 4.305 ;
        RECT 13.155 4.545 13.325 4.715 ;
        RECT 13.345 4.135 13.515 4.305 ;
        RECT 13.805 4.135 13.975 4.305 ;
        RECT 14.265 4.135 14.435 4.305 ;
        RECT 14.725 4.135 14.895 4.305 ;
        RECT 15.185 4.135 15.355 4.305 ;
        RECT 18.77 4.545 18.94 4.715 ;
        RECT 18.77 4.165 18.94 4.335 ;
        RECT 19.47 4.55 19.64 4.72 ;
        RECT 19.47 4.16 19.64 4.33 ;
        RECT 20.46 4.55 20.63 4.72 ;
        RECT 20.46 4.16 20.63 4.33 ;
        RECT 22.245 4.135 22.415 4.305 ;
        RECT 22.705 4.135 22.875 4.305 ;
        RECT 23.165 4.135 23.335 4.305 ;
        RECT 23.625 4.135 23.795 4.305 ;
        RECT 24.085 4.135 24.255 4.305 ;
        RECT 24.545 4.135 24.715 4.305 ;
        RECT 25.005 4.135 25.175 4.305 ;
        RECT 25.465 4.135 25.635 4.305 ;
        RECT 25.925 4.135 26.095 4.305 ;
        RECT 26.385 4.135 26.555 4.305 ;
        RECT 26.845 4.135 27.015 4.305 ;
        RECT 27.305 4.135 27.475 4.305 ;
        RECT 27.765 4.135 27.935 4.305 ;
        RECT 28.225 4.135 28.395 4.305 ;
        RECT 28.685 4.135 28.855 4.305 ;
        RECT 29.145 4.135 29.315 4.305 ;
        RECT 29.605 4.135 29.775 4.305 ;
        RECT 30.065 4.135 30.235 4.305 ;
        RECT 30.525 4.135 30.695 4.305 ;
        RECT 30.985 4.135 31.155 4.305 ;
        RECT 31.445 4.135 31.615 4.305 ;
        RECT 31.715 4.545 31.885 4.715 ;
        RECT 31.905 4.135 32.075 4.305 ;
        RECT 32.365 4.135 32.535 4.305 ;
        RECT 32.825 4.135 32.995 4.305 ;
        RECT 33.285 4.135 33.455 4.305 ;
        RECT 33.745 4.135 33.915 4.305 ;
        RECT 37.33 4.545 37.5 4.715 ;
        RECT 37.33 4.165 37.5 4.335 ;
        RECT 38.03 4.55 38.2 4.72 ;
        RECT 38.03 4.16 38.2 4.33 ;
        RECT 39.02 4.55 39.19 4.72 ;
        RECT 39.02 4.16 39.19 4.33 ;
        RECT 40.805 4.135 40.975 4.305 ;
        RECT 41.265 4.135 41.435 4.305 ;
        RECT 41.725 4.135 41.895 4.305 ;
        RECT 42.185 4.135 42.355 4.305 ;
        RECT 42.645 4.135 42.815 4.305 ;
        RECT 43.105 4.135 43.275 4.305 ;
        RECT 43.565 4.135 43.735 4.305 ;
        RECT 44.025 4.135 44.195 4.305 ;
        RECT 44.485 4.135 44.655 4.305 ;
        RECT 44.945 4.135 45.115 4.305 ;
        RECT 45.405 4.135 45.575 4.305 ;
        RECT 45.865 4.135 46.035 4.305 ;
        RECT 46.325 4.135 46.495 4.305 ;
        RECT 46.785 4.135 46.955 4.305 ;
        RECT 47.245 4.135 47.415 4.305 ;
        RECT 47.705 4.135 47.875 4.305 ;
        RECT 48.165 4.135 48.335 4.305 ;
        RECT 48.625 4.135 48.795 4.305 ;
        RECT 49.085 4.135 49.255 4.305 ;
        RECT 49.545 4.135 49.715 4.305 ;
        RECT 50.005 4.135 50.175 4.305 ;
        RECT 50.275 4.545 50.445 4.715 ;
        RECT 50.465 4.135 50.635 4.305 ;
        RECT 50.925 4.135 51.095 4.305 ;
        RECT 51.385 4.135 51.555 4.305 ;
        RECT 51.845 4.135 52.015 4.305 ;
        RECT 52.305 4.135 52.475 4.305 ;
        RECT 55.89 4.545 56.06 4.715 ;
        RECT 55.89 4.165 56.06 4.335 ;
        RECT 56.59 4.55 56.76 4.72 ;
        RECT 56.59 4.16 56.76 4.33 ;
        RECT 57.58 4.55 57.75 4.72 ;
        RECT 57.58 4.16 57.75 4.33 ;
        RECT 59.365 4.135 59.535 4.305 ;
        RECT 59.825 4.135 59.995 4.305 ;
        RECT 60.285 4.135 60.455 4.305 ;
        RECT 60.745 4.135 60.915 4.305 ;
        RECT 61.205 4.135 61.375 4.305 ;
        RECT 61.665 4.135 61.835 4.305 ;
        RECT 62.125 4.135 62.295 4.305 ;
        RECT 62.585 4.135 62.755 4.305 ;
        RECT 63.045 4.135 63.215 4.305 ;
        RECT 63.505 4.135 63.675 4.305 ;
        RECT 63.965 4.135 64.135 4.305 ;
        RECT 64.425 4.135 64.595 4.305 ;
        RECT 64.885 4.135 65.055 4.305 ;
        RECT 65.345 4.135 65.515 4.305 ;
        RECT 65.805 4.135 65.975 4.305 ;
        RECT 66.265 4.135 66.435 4.305 ;
        RECT 66.725 4.135 66.895 4.305 ;
        RECT 67.185 4.135 67.355 4.305 ;
        RECT 67.645 4.135 67.815 4.305 ;
        RECT 68.105 4.135 68.275 4.305 ;
        RECT 68.565 4.135 68.735 4.305 ;
        RECT 68.835 4.545 69.005 4.715 ;
        RECT 69.025 4.135 69.195 4.305 ;
        RECT 69.485 4.135 69.655 4.305 ;
        RECT 69.945 4.135 70.115 4.305 ;
        RECT 70.405 4.135 70.575 4.305 ;
        RECT 70.865 4.135 71.035 4.305 ;
        RECT 74.45 4.545 74.62 4.715 ;
        RECT 74.45 4.165 74.62 4.335 ;
        RECT 75.15 4.55 75.32 4.72 ;
        RECT 75.15 4.16 75.32 4.33 ;
        RECT 76.14 4.55 76.31 4.72 ;
        RECT 76.14 4.16 76.31 4.33 ;
        RECT 77.925 4.135 78.095 4.305 ;
        RECT 78.385 4.135 78.555 4.305 ;
        RECT 78.845 4.135 79.015 4.305 ;
        RECT 79.305 4.135 79.475 4.305 ;
        RECT 79.765 4.135 79.935 4.305 ;
        RECT 80.225 4.135 80.395 4.305 ;
        RECT 80.685 4.135 80.855 4.305 ;
        RECT 81.145 4.135 81.315 4.305 ;
        RECT 81.605 4.135 81.775 4.305 ;
        RECT 82.065 4.135 82.235 4.305 ;
        RECT 82.525 4.135 82.695 4.305 ;
        RECT 82.985 4.135 83.155 4.305 ;
        RECT 83.445 4.135 83.615 4.305 ;
        RECT 83.905 4.135 84.075 4.305 ;
        RECT 84.365 4.135 84.535 4.305 ;
        RECT 84.825 4.135 84.995 4.305 ;
        RECT 85.285 4.135 85.455 4.305 ;
        RECT 85.745 4.135 85.915 4.305 ;
        RECT 86.205 4.135 86.375 4.305 ;
        RECT 86.665 4.135 86.835 4.305 ;
        RECT 87.125 4.135 87.295 4.305 ;
        RECT 87.395 4.545 87.565 4.715 ;
        RECT 87.585 4.135 87.755 4.305 ;
        RECT 88.045 4.135 88.215 4.305 ;
        RECT 88.505 4.135 88.675 4.305 ;
        RECT 88.965 4.135 89.135 4.305 ;
        RECT 89.425 4.135 89.595 4.305 ;
        RECT 93.01 4.545 93.18 4.715 ;
        RECT 93.01 4.165 93.18 4.335 ;
        RECT 93.71 4.55 93.88 4.72 ;
        RECT 93.71 4.16 93.88 4.33 ;
        RECT 94.7 4.55 94.87 4.72 ;
        RECT 94.7 4.16 94.87 4.33 ;
      LAYER via1 ;
        RECT 1.795 4.38 1.945 4.53 ;
        RECT 4.36 2.505 4.51 2.655 ;
        RECT 5.96 3.065 6.11 3.215 ;
        RECT 8.02 2.505 8.17 2.655 ;
        RECT 8.28 3.065 8.43 3.215 ;
        RECT 12.425 7.165 12.575 7.315 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 79.395 2.415 80.125 2.745 ;
        RECT 60.835 2.415 61.565 2.745 ;
        RECT 42.275 2.415 43.005 2.745 ;
        RECT 23.715 2.415 24.445 2.745 ;
        RECT 5.155 2.415 5.885 2.745 ;
        RECT 0.005 8.5 0.81 8.88 ;
        RECT 0 0 0.805 0.38 ;
      LAYER li1 ;
        RECT 95.415 0 95.595 0.305 ;
        RECT 0.465 0 95.595 0.3 ;
        RECT 94.62 0 94.79 0.93 ;
        RECT 93.63 0 93.8 0.93 ;
        RECT 76.855 0 93.465 0.305 ;
        RECT 90.89 0 91.06 0.935 ;
        RECT 77.78 0 89.825 1.585 ;
        RECT 88.83 0 89 2.085 ;
        RECT 87.87 0 88.04 2.085 ;
        RECT 86.91 0 87.08 2.085 ;
        RECT 86.39 0 86.56 2.085 ;
        RECT 86.11 0 86.305 1.595 ;
        RECT 85.43 0 85.6 2.085 ;
        RECT 84.43 0 84.6 2.085 ;
        RECT 83.47 0 83.64 2.085 ;
        RECT 82.435 0 82.63 1.595 ;
        RECT 81.99 0 82.16 2.085 ;
        RECT 80.07 0 80.33 1.595 ;
        RECT 80.07 0 80.24 2.085 ;
        RECT 78.59 0 78.76 2.085 ;
        RECT 76.06 0 76.23 0.93 ;
        RECT 75.07 0 75.24 0.93 ;
        RECT 58.295 0 74.905 0.305 ;
        RECT 72.33 0 72.5 0.935 ;
        RECT 59.22 0 71.265 1.585 ;
        RECT 70.27 0 70.44 2.085 ;
        RECT 69.31 0 69.48 2.085 ;
        RECT 68.35 0 68.52 2.085 ;
        RECT 67.83 0 68 2.085 ;
        RECT 67.55 0 67.745 1.595 ;
        RECT 66.87 0 67.04 2.085 ;
        RECT 65.87 0 66.04 2.085 ;
        RECT 64.91 0 65.08 2.085 ;
        RECT 63.875 0 64.07 1.595 ;
        RECT 63.43 0 63.6 2.085 ;
        RECT 61.51 0 61.77 1.595 ;
        RECT 61.51 0 61.68 2.085 ;
        RECT 60.03 0 60.2 2.085 ;
        RECT 57.5 0 57.67 0.93 ;
        RECT 56.51 0 56.68 0.93 ;
        RECT 39.735 0 56.345 0.305 ;
        RECT 53.77 0 53.94 0.935 ;
        RECT 40.66 0 52.705 1.585 ;
        RECT 51.71 0 51.88 2.085 ;
        RECT 50.75 0 50.92 2.085 ;
        RECT 49.79 0 49.96 2.085 ;
        RECT 49.27 0 49.44 2.085 ;
        RECT 48.99 0 49.185 1.595 ;
        RECT 48.31 0 48.48 2.085 ;
        RECT 47.31 0 47.48 2.085 ;
        RECT 46.35 0 46.52 2.085 ;
        RECT 45.315 0 45.51 1.595 ;
        RECT 44.87 0 45.04 2.085 ;
        RECT 42.95 0 43.21 1.595 ;
        RECT 42.95 0 43.12 2.085 ;
        RECT 41.47 0 41.64 2.085 ;
        RECT 38.94 0 39.11 0.93 ;
        RECT 37.95 0 38.12 0.93 ;
        RECT 21.175 0 37.785 0.305 ;
        RECT 35.21 0 35.38 0.935 ;
        RECT 22.1 0 34.145 1.585 ;
        RECT 33.15 0 33.32 2.085 ;
        RECT 32.19 0 32.36 2.085 ;
        RECT 31.23 0 31.4 2.085 ;
        RECT 30.71 0 30.88 2.085 ;
        RECT 30.43 0 30.625 1.595 ;
        RECT 29.75 0 29.92 2.085 ;
        RECT 28.75 0 28.92 2.085 ;
        RECT 27.79 0 27.96 2.085 ;
        RECT 26.755 0 26.95 1.595 ;
        RECT 26.31 0 26.48 2.085 ;
        RECT 24.39 0 24.65 1.595 ;
        RECT 24.39 0 24.56 2.085 ;
        RECT 22.91 0 23.08 2.085 ;
        RECT 20.38 0 20.55 0.93 ;
        RECT 19.39 0 19.56 0.93 ;
        RECT 0 0.245 19.225 0.305 ;
        RECT 16.65 0 16.82 0.935 ;
        RECT 3.54 0 15.585 1.585 ;
        RECT 14.59 0 14.76 2.085 ;
        RECT 13.63 0 13.8 2.085 ;
        RECT 12.67 0 12.84 2.085 ;
        RECT 12.15 0 12.32 2.085 ;
        RECT 11.87 0 12.065 1.595 ;
        RECT 11.19 0 11.36 2.085 ;
        RECT 10.19 0 10.36 2.085 ;
        RECT 9.23 0 9.4 2.085 ;
        RECT 8.195 0 8.39 1.595 ;
        RECT 7.75 0 7.92 2.085 ;
        RECT 5.83 0 6.09 1.595 ;
        RECT 5.83 0 6 2.085 ;
        RECT 4.35 0 4.52 2.085 ;
        RECT 0 0.245 0.805 0.315 ;
        RECT 0.295 0.245 0.465 0.335 ;
        RECT 0 0 95.595 0.075 ;
        RECT 0 0 0.295 0.315 ;
        RECT 0 8.58 95.595 8.88 ;
        RECT 95.415 8.575 95.595 8.88 ;
        RECT 94.62 7.95 94.79 8.88 ;
        RECT 93.63 7.95 93.8 8.88 ;
        RECT 76.855 8.575 93.465 8.88 ;
        RECT 90.89 7.945 91.06 8.88 ;
        RECT 85.275 7.945 85.445 8.88 ;
        RECT 76.06 7.95 76.23 8.88 ;
        RECT 75.07 7.95 75.24 8.88 ;
        RECT 58.295 8.575 74.905 8.88 ;
        RECT 72.33 7.945 72.5 8.88 ;
        RECT 66.715 7.945 66.885 8.88 ;
        RECT 57.5 7.95 57.67 8.88 ;
        RECT 56.51 7.95 56.68 8.88 ;
        RECT 39.735 8.575 56.345 8.88 ;
        RECT 53.77 7.945 53.94 8.88 ;
        RECT 48.155 7.945 48.325 8.88 ;
        RECT 38.94 7.95 39.11 8.88 ;
        RECT 37.95 7.95 38.12 8.88 ;
        RECT 21.175 8.575 37.785 8.88 ;
        RECT 35.21 7.945 35.38 8.88 ;
        RECT 29.595 7.945 29.765 8.88 ;
        RECT 20.38 7.95 20.55 8.88 ;
        RECT 19.39 7.95 19.56 8.88 ;
        RECT 0 8.575 19.225 8.88 ;
        RECT 16.65 7.945 16.82 8.88 ;
        RECT 11.035 7.945 11.205 8.88 ;
        RECT 0.005 8.565 0.81 8.88 ;
        RECT 0.22 8.545 0.47 8.88 ;
        RECT 0.22 7.945 0.39 8.88 ;
        RECT 86.28 6.075 86.45 8.025 ;
        RECT 86.225 7.855 86.395 8.305 ;
        RECT 86.225 5.015 86.395 6.245 ;
        RECT 81.27 2.495 81.44 2.825 ;
        RECT 79.43 3.055 79.72 3.225 ;
        RECT 79.43 2.575 79.6 3.225 ;
        RECT 79.23 2.575 79.6 2.745 ;
        RECT 67.72 6.075 67.89 8.025 ;
        RECT 67.665 7.855 67.835 8.305 ;
        RECT 67.665 5.015 67.835 6.245 ;
        RECT 62.71 2.495 62.88 2.825 ;
        RECT 60.87 3.055 61.16 3.225 ;
        RECT 60.87 2.575 61.04 3.225 ;
        RECT 60.67 2.575 61.04 2.745 ;
        RECT 49.16 6.075 49.33 8.025 ;
        RECT 49.105 7.855 49.275 8.305 ;
        RECT 49.105 5.015 49.275 6.245 ;
        RECT 44.15 2.495 44.32 2.825 ;
        RECT 42.31 3.055 42.6 3.225 ;
        RECT 42.31 2.575 42.48 3.225 ;
        RECT 42.11 2.575 42.48 2.745 ;
        RECT 30.6 6.075 30.77 8.025 ;
        RECT 30.545 7.855 30.715 8.305 ;
        RECT 30.545 5.015 30.715 6.245 ;
        RECT 25.59 2.495 25.76 2.825 ;
        RECT 23.75 3.055 24.04 3.225 ;
        RECT 23.75 2.575 23.92 3.225 ;
        RECT 23.55 2.575 23.92 2.745 ;
        RECT 12.04 6.075 12.21 8.025 ;
        RECT 11.985 7.855 12.155 8.305 ;
        RECT 11.985 5.015 12.155 6.245 ;
        RECT 7.03 2.495 7.2 2.825 ;
        RECT 5.19 3.055 5.48 3.225 ;
        RECT 5.19 2.575 5.36 3.225 ;
        RECT 4.99 2.575 5.36 2.745 ;
      LAYER met2 ;
        RECT 81.225 2.42 81.485 2.74 ;
        RECT 79.445 2.51 81.485 2.65 ;
        RECT 79.825 1 80.165 1.34 ;
        RECT 79.755 2.395 80.035 2.765 ;
        RECT 79.85 1 80.02 2.765 ;
        RECT 79.505 2.98 79.765 3.3 ;
        RECT 79.445 2.51 79.585 3.21 ;
        RECT 62.665 2.42 62.925 2.74 ;
        RECT 60.885 2.51 62.925 2.65 ;
        RECT 61.265 1 61.605 1.34 ;
        RECT 61.195 2.395 61.475 2.765 ;
        RECT 61.29 1 61.46 2.765 ;
        RECT 60.945 2.98 61.205 3.3 ;
        RECT 60.885 2.51 61.025 3.21 ;
        RECT 44.105 2.42 44.365 2.74 ;
        RECT 42.325 2.51 44.365 2.65 ;
        RECT 42.705 1 43.045 1.34 ;
        RECT 42.635 2.395 42.915 2.765 ;
        RECT 42.73 1 42.9 2.765 ;
        RECT 42.385 2.98 42.645 3.3 ;
        RECT 42.325 2.51 42.465 3.21 ;
        RECT 25.545 2.42 25.805 2.74 ;
        RECT 23.765 2.51 25.805 2.65 ;
        RECT 24.145 1 24.485 1.34 ;
        RECT 24.075 2.395 24.355 2.765 ;
        RECT 24.17 1 24.34 2.765 ;
        RECT 23.825 2.98 24.085 3.3 ;
        RECT 23.765 2.51 23.905 3.21 ;
        RECT 6.985 2.42 7.245 2.74 ;
        RECT 5.205 2.51 7.245 2.65 ;
        RECT 5.585 1 5.925 1.34 ;
        RECT 5.515 2.395 5.795 2.765 ;
        RECT 5.61 1 5.78 2.765 ;
        RECT 5.265 2.98 5.525 3.3 ;
        RECT 5.205 2.51 5.345 3.21 ;
        RECT 0.195 8.5 0.575 8.88 ;
        RECT 0.19 0 0.57 0.38 ;
        RECT 0.235 0 0.405 8.88 ;
      LAYER met1 ;
        RECT 95.415 0 95.595 0.305 ;
        RECT 0 0 95.595 0.3 ;
        RECT 76.855 0 93.465 0.305 ;
        RECT 77.78 0 89.825 1.585 ;
        RECT 77.78 0 89.74 1.74 ;
        RECT 58.295 0 74.905 0.305 ;
        RECT 59.22 0 71.265 1.585 ;
        RECT 59.22 0 71.18 1.74 ;
        RECT 39.735 0 56.345 0.305 ;
        RECT 40.66 0 52.705 1.585 ;
        RECT 40.66 0 52.62 1.74 ;
        RECT 21.175 0 37.785 0.305 ;
        RECT 22.1 0 34.145 1.585 ;
        RECT 22.1 0 34.06 1.74 ;
        RECT 0 0 19.225 0.305 ;
        RECT 3.54 0 15.585 1.585 ;
        RECT 3.54 0 15.5 1.74 ;
        RECT 0 0 0.805 0.315 ;
        RECT 0.205 0 0.555 0.335 ;
        RECT 0 8.58 95.595 8.88 ;
        RECT 95.415 8.575 95.595 8.88 ;
        RECT 76.855 8.575 93.465 8.88 ;
        RECT 86.22 6.285 86.51 6.515 ;
        RECT 85.785 6.315 86.51 6.485 ;
        RECT 85.785 6.315 85.955 8.88 ;
        RECT 58.295 8.575 74.905 8.88 ;
        RECT 67.66 6.285 67.95 6.515 ;
        RECT 67.225 6.315 67.95 6.485 ;
        RECT 67.225 6.315 67.395 8.88 ;
        RECT 39.735 8.575 56.345 8.88 ;
        RECT 49.1 6.285 49.39 6.515 ;
        RECT 48.665 6.315 49.39 6.485 ;
        RECT 48.665 6.315 48.835 8.88 ;
        RECT 21.175 8.575 37.785 8.88 ;
        RECT 30.54 6.285 30.83 6.515 ;
        RECT 30.105 6.315 30.83 6.485 ;
        RECT 30.105 6.315 30.275 8.88 ;
        RECT 0 8.575 19.225 8.88 ;
        RECT 11.98 6.285 12.27 6.515 ;
        RECT 11.545 6.315 12.27 6.485 ;
        RECT 11.545 6.315 11.715 8.88 ;
        RECT 0.005 8.565 0.81 8.88 ;
        RECT 0.21 8.545 0.56 8.88 ;
        RECT 81.21 2.37 81.5 2.74 ;
        RECT 80.445 2.37 81.5 2.51 ;
        RECT 79.475 3.01 79.795 3.27 ;
        RECT 62.65 2.37 62.94 2.74 ;
        RECT 61.885 2.37 62.94 2.51 ;
        RECT 60.915 3.01 61.235 3.27 ;
        RECT 44.09 2.37 44.38 2.74 ;
        RECT 43.325 2.37 44.38 2.51 ;
        RECT 42.355 3.01 42.675 3.27 ;
        RECT 25.53 2.37 25.82 2.74 ;
        RECT 24.765 2.37 25.82 2.51 ;
        RECT 23.795 3.01 24.115 3.27 ;
        RECT 6.97 2.37 7.26 2.74 ;
        RECT 6.205 2.37 7.26 2.51 ;
        RECT 5.235 3.01 5.555 3.27 ;
      LAYER via2 ;
        RECT 0.28 0.09 0.48 0.29 ;
        RECT 0.285 8.59 0.485 8.79 ;
        RECT 5.555 2.48 5.755 2.68 ;
        RECT 24.115 2.48 24.315 2.68 ;
        RECT 42.675 2.48 42.875 2.68 ;
        RECT 61.235 2.48 61.435 2.68 ;
        RECT 79.795 2.48 79.995 2.68 ;
      LAYER mcon ;
        RECT 0.3 8.605 0.47 8.775 ;
        RECT 0.98 8.605 1.15 8.775 ;
        RECT 1.66 8.605 1.83 8.775 ;
        RECT 2.34 8.605 2.51 8.775 ;
        RECT 3.685 1.415 3.855 1.585 ;
        RECT 4.145 1.415 4.315 1.585 ;
        RECT 4.605 1.415 4.775 1.585 ;
        RECT 5.065 1.415 5.235 1.585 ;
        RECT 5.31 3.055 5.48 3.225 ;
        RECT 5.525 1.415 5.695 1.585 ;
        RECT 5.985 1.415 6.155 1.585 ;
        RECT 6.445 1.415 6.615 1.585 ;
        RECT 6.905 1.415 7.075 1.585 ;
        RECT 7.03 2.495 7.2 2.665 ;
        RECT 7.365 1.415 7.535 1.585 ;
        RECT 7.825 1.415 7.995 1.585 ;
        RECT 8.285 1.415 8.455 1.585 ;
        RECT 8.745 1.415 8.915 1.585 ;
        RECT 9.205 1.415 9.375 1.585 ;
        RECT 9.665 1.415 9.835 1.585 ;
        RECT 10.125 1.415 10.295 1.585 ;
        RECT 10.585 1.415 10.755 1.585 ;
        RECT 11.045 1.415 11.215 1.585 ;
        RECT 11.115 8.605 11.285 8.775 ;
        RECT 11.505 1.415 11.675 1.585 ;
        RECT 11.795 8.605 11.965 8.775 ;
        RECT 11.965 1.415 12.135 1.585 ;
        RECT 12.04 6.315 12.21 6.485 ;
        RECT 12.425 1.415 12.595 1.585 ;
        RECT 12.475 8.605 12.645 8.775 ;
        RECT 12.885 1.415 13.055 1.585 ;
        RECT 13.155 8.605 13.325 8.775 ;
        RECT 13.345 1.415 13.515 1.585 ;
        RECT 13.805 1.415 13.975 1.585 ;
        RECT 14.265 1.415 14.435 1.585 ;
        RECT 14.725 1.415 14.895 1.585 ;
        RECT 15.185 1.415 15.355 1.585 ;
        RECT 16.73 8.605 16.9 8.775 ;
        RECT 16.73 0.105 16.9 0.275 ;
        RECT 17.41 8.605 17.58 8.775 ;
        RECT 17.41 0.105 17.58 0.275 ;
        RECT 18.09 8.605 18.26 8.775 ;
        RECT 18.09 0.105 18.26 0.275 ;
        RECT 18.77 8.605 18.94 8.775 ;
        RECT 18.77 0.105 18.94 0.275 ;
        RECT 19.47 8.61 19.64 8.78 ;
        RECT 19.47 0.1 19.64 0.27 ;
        RECT 20.46 8.61 20.63 8.78 ;
        RECT 20.46 0.1 20.63 0.27 ;
        RECT 22.245 1.415 22.415 1.585 ;
        RECT 22.705 1.415 22.875 1.585 ;
        RECT 23.165 1.415 23.335 1.585 ;
        RECT 23.625 1.415 23.795 1.585 ;
        RECT 23.87 3.055 24.04 3.225 ;
        RECT 24.085 1.415 24.255 1.585 ;
        RECT 24.545 1.415 24.715 1.585 ;
        RECT 25.005 1.415 25.175 1.585 ;
        RECT 25.465 1.415 25.635 1.585 ;
        RECT 25.59 2.495 25.76 2.665 ;
        RECT 25.925 1.415 26.095 1.585 ;
        RECT 26.385 1.415 26.555 1.585 ;
        RECT 26.845 1.415 27.015 1.585 ;
        RECT 27.305 1.415 27.475 1.585 ;
        RECT 27.765 1.415 27.935 1.585 ;
        RECT 28.225 1.415 28.395 1.585 ;
        RECT 28.685 1.415 28.855 1.585 ;
        RECT 29.145 1.415 29.315 1.585 ;
        RECT 29.605 1.415 29.775 1.585 ;
        RECT 29.675 8.605 29.845 8.775 ;
        RECT 30.065 1.415 30.235 1.585 ;
        RECT 30.355 8.605 30.525 8.775 ;
        RECT 30.525 1.415 30.695 1.585 ;
        RECT 30.6 6.315 30.77 6.485 ;
        RECT 30.985 1.415 31.155 1.585 ;
        RECT 31.035 8.605 31.205 8.775 ;
        RECT 31.445 1.415 31.615 1.585 ;
        RECT 31.715 8.605 31.885 8.775 ;
        RECT 31.905 1.415 32.075 1.585 ;
        RECT 32.365 1.415 32.535 1.585 ;
        RECT 32.825 1.415 32.995 1.585 ;
        RECT 33.285 1.415 33.455 1.585 ;
        RECT 33.745 1.415 33.915 1.585 ;
        RECT 35.29 8.605 35.46 8.775 ;
        RECT 35.29 0.105 35.46 0.275 ;
        RECT 35.97 8.605 36.14 8.775 ;
        RECT 35.97 0.105 36.14 0.275 ;
        RECT 36.65 8.605 36.82 8.775 ;
        RECT 36.65 0.105 36.82 0.275 ;
        RECT 37.33 8.605 37.5 8.775 ;
        RECT 37.33 0.105 37.5 0.275 ;
        RECT 38.03 8.61 38.2 8.78 ;
        RECT 38.03 0.1 38.2 0.27 ;
        RECT 39.02 8.61 39.19 8.78 ;
        RECT 39.02 0.1 39.19 0.27 ;
        RECT 40.805 1.415 40.975 1.585 ;
        RECT 41.265 1.415 41.435 1.585 ;
        RECT 41.725 1.415 41.895 1.585 ;
        RECT 42.185 1.415 42.355 1.585 ;
        RECT 42.43 3.055 42.6 3.225 ;
        RECT 42.645 1.415 42.815 1.585 ;
        RECT 43.105 1.415 43.275 1.585 ;
        RECT 43.565 1.415 43.735 1.585 ;
        RECT 44.025 1.415 44.195 1.585 ;
        RECT 44.15 2.495 44.32 2.665 ;
        RECT 44.485 1.415 44.655 1.585 ;
        RECT 44.945 1.415 45.115 1.585 ;
        RECT 45.405 1.415 45.575 1.585 ;
        RECT 45.865 1.415 46.035 1.585 ;
        RECT 46.325 1.415 46.495 1.585 ;
        RECT 46.785 1.415 46.955 1.585 ;
        RECT 47.245 1.415 47.415 1.585 ;
        RECT 47.705 1.415 47.875 1.585 ;
        RECT 48.165 1.415 48.335 1.585 ;
        RECT 48.235 8.605 48.405 8.775 ;
        RECT 48.625 1.415 48.795 1.585 ;
        RECT 48.915 8.605 49.085 8.775 ;
        RECT 49.085 1.415 49.255 1.585 ;
        RECT 49.16 6.315 49.33 6.485 ;
        RECT 49.545 1.415 49.715 1.585 ;
        RECT 49.595 8.605 49.765 8.775 ;
        RECT 50.005 1.415 50.175 1.585 ;
        RECT 50.275 8.605 50.445 8.775 ;
        RECT 50.465 1.415 50.635 1.585 ;
        RECT 50.925 1.415 51.095 1.585 ;
        RECT 51.385 1.415 51.555 1.585 ;
        RECT 51.845 1.415 52.015 1.585 ;
        RECT 52.305 1.415 52.475 1.585 ;
        RECT 53.85 8.605 54.02 8.775 ;
        RECT 53.85 0.105 54.02 0.275 ;
        RECT 54.53 8.605 54.7 8.775 ;
        RECT 54.53 0.105 54.7 0.275 ;
        RECT 55.21 8.605 55.38 8.775 ;
        RECT 55.21 0.105 55.38 0.275 ;
        RECT 55.89 8.605 56.06 8.775 ;
        RECT 55.89 0.105 56.06 0.275 ;
        RECT 56.59 8.61 56.76 8.78 ;
        RECT 56.59 0.1 56.76 0.27 ;
        RECT 57.58 8.61 57.75 8.78 ;
        RECT 57.58 0.1 57.75 0.27 ;
        RECT 59.365 1.415 59.535 1.585 ;
        RECT 59.825 1.415 59.995 1.585 ;
        RECT 60.285 1.415 60.455 1.585 ;
        RECT 60.745 1.415 60.915 1.585 ;
        RECT 60.99 3.055 61.16 3.225 ;
        RECT 61.205 1.415 61.375 1.585 ;
        RECT 61.665 1.415 61.835 1.585 ;
        RECT 62.125 1.415 62.295 1.585 ;
        RECT 62.585 1.415 62.755 1.585 ;
        RECT 62.71 2.495 62.88 2.665 ;
        RECT 63.045 1.415 63.215 1.585 ;
        RECT 63.505 1.415 63.675 1.585 ;
        RECT 63.965 1.415 64.135 1.585 ;
        RECT 64.425 1.415 64.595 1.585 ;
        RECT 64.885 1.415 65.055 1.585 ;
        RECT 65.345 1.415 65.515 1.585 ;
        RECT 65.805 1.415 65.975 1.585 ;
        RECT 66.265 1.415 66.435 1.585 ;
        RECT 66.725 1.415 66.895 1.585 ;
        RECT 66.795 8.605 66.965 8.775 ;
        RECT 67.185 1.415 67.355 1.585 ;
        RECT 67.475 8.605 67.645 8.775 ;
        RECT 67.645 1.415 67.815 1.585 ;
        RECT 67.72 6.315 67.89 6.485 ;
        RECT 68.105 1.415 68.275 1.585 ;
        RECT 68.155 8.605 68.325 8.775 ;
        RECT 68.565 1.415 68.735 1.585 ;
        RECT 68.835 8.605 69.005 8.775 ;
        RECT 69.025 1.415 69.195 1.585 ;
        RECT 69.485 1.415 69.655 1.585 ;
        RECT 69.945 1.415 70.115 1.585 ;
        RECT 70.405 1.415 70.575 1.585 ;
        RECT 70.865 1.415 71.035 1.585 ;
        RECT 72.41 8.605 72.58 8.775 ;
        RECT 72.41 0.105 72.58 0.275 ;
        RECT 73.09 8.605 73.26 8.775 ;
        RECT 73.09 0.105 73.26 0.275 ;
        RECT 73.77 8.605 73.94 8.775 ;
        RECT 73.77 0.105 73.94 0.275 ;
        RECT 74.45 8.605 74.62 8.775 ;
        RECT 74.45 0.105 74.62 0.275 ;
        RECT 75.15 8.61 75.32 8.78 ;
        RECT 75.15 0.1 75.32 0.27 ;
        RECT 76.14 8.61 76.31 8.78 ;
        RECT 76.14 0.1 76.31 0.27 ;
        RECT 77.925 1.415 78.095 1.585 ;
        RECT 78.385 1.415 78.555 1.585 ;
        RECT 78.845 1.415 79.015 1.585 ;
        RECT 79.305 1.415 79.475 1.585 ;
        RECT 79.55 3.055 79.72 3.225 ;
        RECT 79.765 1.415 79.935 1.585 ;
        RECT 80.225 1.415 80.395 1.585 ;
        RECT 80.685 1.415 80.855 1.585 ;
        RECT 81.145 1.415 81.315 1.585 ;
        RECT 81.27 2.495 81.44 2.665 ;
        RECT 81.605 1.415 81.775 1.585 ;
        RECT 82.065 1.415 82.235 1.585 ;
        RECT 82.525 1.415 82.695 1.585 ;
        RECT 82.985 1.415 83.155 1.585 ;
        RECT 83.445 1.415 83.615 1.585 ;
        RECT 83.905 1.415 84.075 1.585 ;
        RECT 84.365 1.415 84.535 1.585 ;
        RECT 84.825 1.415 84.995 1.585 ;
        RECT 85.285 1.415 85.455 1.585 ;
        RECT 85.355 8.605 85.525 8.775 ;
        RECT 85.745 1.415 85.915 1.585 ;
        RECT 86.035 8.605 86.205 8.775 ;
        RECT 86.205 1.415 86.375 1.585 ;
        RECT 86.28 6.315 86.45 6.485 ;
        RECT 86.665 1.415 86.835 1.585 ;
        RECT 86.715 8.605 86.885 8.775 ;
        RECT 87.125 1.415 87.295 1.585 ;
        RECT 87.395 8.605 87.565 8.775 ;
        RECT 87.585 1.415 87.755 1.585 ;
        RECT 88.045 1.415 88.215 1.585 ;
        RECT 88.505 1.415 88.675 1.585 ;
        RECT 88.965 1.415 89.135 1.585 ;
        RECT 89.425 1.415 89.595 1.585 ;
        RECT 90.97 8.605 91.14 8.775 ;
        RECT 90.97 0.105 91.14 0.275 ;
        RECT 91.65 8.605 91.82 8.775 ;
        RECT 91.65 0.105 91.82 0.275 ;
        RECT 92.33 8.605 92.5 8.775 ;
        RECT 92.33 0.105 92.5 0.275 ;
        RECT 93.01 8.605 93.18 8.775 ;
        RECT 93.01 0.105 93.18 0.275 ;
        RECT 93.71 8.61 93.88 8.78 ;
        RECT 93.71 0.1 93.88 0.27 ;
        RECT 94.7 8.61 94.87 8.78 ;
        RECT 94.7 0.1 94.87 0.27 ;
      LAYER via1 ;
        RECT 0.305 0.115 0.455 0.265 ;
        RECT 0.31 8.615 0.46 8.765 ;
        RECT 5.32 3.065 5.47 3.215 ;
        RECT 5.68 1.095 5.83 1.245 ;
        RECT 7.04 2.505 7.19 2.655 ;
        RECT 23.88 3.065 24.03 3.215 ;
        RECT 24.24 1.095 24.39 1.245 ;
        RECT 25.6 2.505 25.75 2.655 ;
        RECT 42.44 3.065 42.59 3.215 ;
        RECT 42.8 1.095 42.95 1.245 ;
        RECT 44.16 2.505 44.31 2.655 ;
        RECT 61 3.065 61.15 3.215 ;
        RECT 61.36 1.095 61.51 1.245 ;
        RECT 62.72 2.505 62.87 2.655 ;
        RECT 79.56 3.065 79.71 3.215 ;
        RECT 79.92 1.095 80.07 1.245 ;
        RECT 81.28 2.505 81.43 2.655 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 87.085 3.535 87.64 3.865 ;
      RECT 87.085 1.87 87.385 3.865 ;
      RECT 83.15 2.975 83.705 3.305 ;
      RECT 83.405 1.87 83.705 3.305 ;
      RECT 83.405 1.87 87.385 2.17 ;
      RECT 86.555 7.055 86.93 7.425 ;
      RECT 86.555 7.095 87.56 7.395 ;
      RECT 87.26 4.405 87.56 7.395 ;
      RECT 77.43 4.405 87.56 4.705 ;
      RECT 81.935 2.415 82.235 4.705 ;
      RECT 80.5 2.975 80.8 4.705 ;
      RECT 77.43 2.42 77.73 4.705 ;
      RECT 80.47 2.975 81.2 3.305 ;
      RECT 81.91 2.415 82.64 2.745 ;
      RECT 78.36 2.415 79.09 2.745 ;
      RECT 77.43 2.42 79.09 2.72 ;
      RECT 68.525 3.535 69.08 3.865 ;
      RECT 68.525 1.87 68.825 3.865 ;
      RECT 64.59 2.975 65.145 3.305 ;
      RECT 64.845 1.87 65.145 3.305 ;
      RECT 64.845 1.87 68.825 2.17 ;
      RECT 67.995 7.055 68.37 7.425 ;
      RECT 67.995 7.095 69 7.395 ;
      RECT 68.7 4.405 69 7.395 ;
      RECT 58.87 4.405 69 4.705 ;
      RECT 63.375 2.415 63.675 4.705 ;
      RECT 61.94 2.975 62.24 4.705 ;
      RECT 58.87 2.42 59.17 4.705 ;
      RECT 61.91 2.975 62.64 3.305 ;
      RECT 63.35 2.415 64.08 2.745 ;
      RECT 59.8 2.415 60.53 2.745 ;
      RECT 58.87 2.42 60.53 2.72 ;
      RECT 49.965 3.535 50.52 3.865 ;
      RECT 49.965 1.87 50.265 3.865 ;
      RECT 46.03 2.975 46.585 3.305 ;
      RECT 46.285 1.87 46.585 3.305 ;
      RECT 46.285 1.87 50.265 2.17 ;
      RECT 49.435 7.055 49.81 7.425 ;
      RECT 49.435 7.095 50.44 7.395 ;
      RECT 50.14 4.405 50.44 7.395 ;
      RECT 40.31 4.405 50.44 4.705 ;
      RECT 44.815 2.415 45.115 4.705 ;
      RECT 43.38 2.975 43.68 4.705 ;
      RECT 40.31 2.42 40.61 4.705 ;
      RECT 43.35 2.975 44.08 3.305 ;
      RECT 44.79 2.415 45.52 2.745 ;
      RECT 41.24 2.415 41.97 2.745 ;
      RECT 40.31 2.42 41.97 2.72 ;
      RECT 31.405 3.535 31.96 3.865 ;
      RECT 31.405 1.87 31.705 3.865 ;
      RECT 27.47 2.975 28.025 3.305 ;
      RECT 27.725 1.87 28.025 3.305 ;
      RECT 27.725 1.87 31.705 2.17 ;
      RECT 30.875 7.055 31.25 7.425 ;
      RECT 30.875 7.095 31.88 7.395 ;
      RECT 31.58 4.405 31.88 7.395 ;
      RECT 21.75 4.405 31.88 4.705 ;
      RECT 26.255 2.415 26.555 4.705 ;
      RECT 24.82 2.975 25.12 4.705 ;
      RECT 21.75 2.42 22.05 4.705 ;
      RECT 24.79 2.975 25.52 3.305 ;
      RECT 26.23 2.415 26.96 2.745 ;
      RECT 22.68 2.415 23.41 2.745 ;
      RECT 21.75 2.42 23.41 2.72 ;
      RECT 12.845 3.535 13.4 3.865 ;
      RECT 12.845 1.87 13.145 3.865 ;
      RECT 8.91 2.975 9.465 3.305 ;
      RECT 9.165 1.87 9.465 3.305 ;
      RECT 9.165 1.87 13.145 2.17 ;
      RECT 88.27 1.855 89 2.185 ;
      RECT 86.05 3.535 86.78 3.865 ;
      RECT 84.35 3.535 85.08 3.865 ;
      RECT 78.03 3.535 78.76 3.865 ;
      RECT 69.71 1.855 70.44 2.185 ;
      RECT 67.49 3.535 68.22 3.865 ;
      RECT 65.79 3.535 66.52 3.865 ;
      RECT 59.47 3.535 60.2 3.865 ;
      RECT 51.15 1.855 51.88 2.185 ;
      RECT 48.93 3.535 49.66 3.865 ;
      RECT 47.23 3.535 47.96 3.865 ;
      RECT 40.91 3.535 41.64 3.865 ;
      RECT 32.59 1.855 33.32 2.185 ;
      RECT 30.37 3.535 31.1 3.865 ;
      RECT 28.67 3.535 29.4 3.865 ;
      RECT 22.35 3.535 23.08 3.865 ;
      RECT 14.03 1.855 14.76 2.185 ;
      RECT 11.81 3.535 12.54 3.865 ;
      RECT 10.11 3.535 10.84 3.865 ;
      RECT 3.79 3.535 4.52 3.865 ;
    LAYER via2 ;
      RECT 88.335 1.92 88.535 2.12 ;
      RECT 87.375 3.6 87.575 3.8 ;
      RECT 86.64 7.14 86.84 7.34 ;
      RECT 86.375 3.6 86.575 3.8 ;
      RECT 84.415 3.6 84.615 3.8 ;
      RECT 83.215 3.04 83.415 3.24 ;
      RECT 81.975 2.48 82.175 2.68 ;
      RECT 80.535 3.04 80.735 3.24 ;
      RECT 78.575 2.48 78.775 2.68 ;
      RECT 78.095 3.6 78.295 3.8 ;
      RECT 69.775 1.92 69.975 2.12 ;
      RECT 68.815 3.6 69.015 3.8 ;
      RECT 68.08 7.14 68.28 7.34 ;
      RECT 67.815 3.6 68.015 3.8 ;
      RECT 65.855 3.6 66.055 3.8 ;
      RECT 64.655 3.04 64.855 3.24 ;
      RECT 63.415 2.48 63.615 2.68 ;
      RECT 61.975 3.04 62.175 3.24 ;
      RECT 60.015 2.48 60.215 2.68 ;
      RECT 59.535 3.6 59.735 3.8 ;
      RECT 51.215 1.92 51.415 2.12 ;
      RECT 50.255 3.6 50.455 3.8 ;
      RECT 49.52 7.14 49.72 7.34 ;
      RECT 49.255 3.6 49.455 3.8 ;
      RECT 47.295 3.6 47.495 3.8 ;
      RECT 46.095 3.04 46.295 3.24 ;
      RECT 44.855 2.48 45.055 2.68 ;
      RECT 43.415 3.04 43.615 3.24 ;
      RECT 41.455 2.48 41.655 2.68 ;
      RECT 40.975 3.6 41.175 3.8 ;
      RECT 32.655 1.92 32.855 2.12 ;
      RECT 31.695 3.6 31.895 3.8 ;
      RECT 30.96 7.14 31.16 7.34 ;
      RECT 30.695 3.6 30.895 3.8 ;
      RECT 28.735 3.6 28.935 3.8 ;
      RECT 27.535 3.04 27.735 3.24 ;
      RECT 26.295 2.48 26.495 2.68 ;
      RECT 24.855 3.04 25.055 3.24 ;
      RECT 22.895 2.48 23.095 2.68 ;
      RECT 22.415 3.6 22.615 3.8 ;
      RECT 14.095 1.92 14.295 2.12 ;
      RECT 13.135 3.6 13.335 3.8 ;
      RECT 12.135 3.6 12.335 3.8 ;
      RECT 10.175 3.6 10.375 3.8 ;
      RECT 8.975 3.04 9.175 3.24 ;
      RECT 3.855 3.6 4.055 3.8 ;
    LAYER met2 ;
      RECT 1.23 8.4 95.225 8.57 ;
      RECT 95.055 7.275 95.225 8.57 ;
      RECT 1.23 6.255 1.4 8.57 ;
      RECT 95.025 7.275 95.375 7.625 ;
      RECT 1.165 6.255 1.455 6.605 ;
      RECT 91.865 6.22 92.185 6.545 ;
      RECT 91.895 5.695 92.065 6.545 ;
      RECT 91.895 5.695 92.07 6.045 ;
      RECT 91.895 5.695 92.87 5.87 ;
      RECT 92.695 1.965 92.87 5.87 ;
      RECT 92.64 1.965 92.99 2.315 ;
      RECT 92.665 6.655 92.99 6.98 ;
      RECT 91.55 6.745 92.99 6.915 ;
      RECT 91.55 2.395 91.71 6.915 ;
      RECT 91.865 2.365 92.185 2.685 ;
      RECT 91.55 2.395 92.185 2.565 ;
      RECT 86.385 4.135 90.52 4.325 ;
      RECT 90.35 3.145 90.52 4.325 ;
      RECT 90.33 3.15 90.52 4.325 ;
      RECT 86.385 3.515 86.575 4.325 ;
      RECT 86.335 3.515 86.615 3.885 ;
      RECT 90.26 3.15 90.6 3.5 ;
      RECT 76.44 6.655 76.79 7.005 ;
      RECT 87.225 6.61 87.575 6.96 ;
      RECT 76.44 6.685 87.575 6.885 ;
      RECT 86.865 2.98 87.125 3.3 ;
      RECT 86.925 1.86 87.065 3.3 ;
      RECT 86.865 1.86 87.125 2.18 ;
      RECT 85.865 3.54 86.125 3.86 ;
      RECT 85.865 2.955 86.065 3.86 ;
      RECT 85.805 1.86 85.945 3.49 ;
      RECT 85.805 2.955 86.305 3.325 ;
      RECT 85.745 1.86 86.005 2.18 ;
      RECT 85.385 3.54 85.645 3.86 ;
      RECT 85.445 1.95 85.585 3.86 ;
      RECT 85.145 1.95 85.585 2.18 ;
      RECT 85.145 1.86 85.405 2.18 ;
      RECT 84.905 2.42 85.165 2.74 ;
      RECT 84.325 2.51 85.165 2.65 ;
      RECT 84.325 1.57 84.465 2.65 ;
      RECT 80.985 1.86 81.245 2.18 ;
      RECT 80.985 1.95 82.025 2.09 ;
      RECT 81.885 1.57 82.025 2.09 ;
      RECT 81.885 1.57 84.465 1.71 ;
      RECT 84.375 3.515 84.655 3.885 ;
      RECT 84.445 3.07 84.585 3.885 ;
      RECT 84.255 2.955 84.535 3.325 ;
      RECT 83.965 3.07 84.585 3.21 ;
      RECT 83.965 1.86 84.105 3.21 ;
      RECT 83.905 1.86 84.165 2.18 ;
      RECT 83.175 2.955 83.455 3.325 ;
      RECT 83.245 1.86 83.385 3.325 ;
      RECT 83.185 1.86 83.445 2.18 ;
      RECT 82.825 3.54 83.085 3.86 ;
      RECT 82.885 1.95 83.025 3.86 ;
      RECT 82.465 1.86 82.725 2.18 ;
      RECT 82.465 1.95 83.025 2.09 ;
      RECT 80.495 2.955 80.775 3.325 ;
      RECT 82.465 2.98 82.725 3.3 ;
      RECT 80.145 2.98 80.775 3.3 ;
      RECT 80.145 3.07 82.725 3.21 ;
      RECT 81.935 2.395 82.215 2.765 ;
      RECT 81.935 2.42 82.465 2.74 ;
      RECT 79.025 2.98 79.285 3.3 ;
      RECT 79.085 1.86 79.225 3.3 ;
      RECT 79.025 1.86 79.285 2.18 ;
      RECT 78.055 3.515 78.335 3.885 ;
      RECT 78.065 3.26 78.325 3.885 ;
      RECT 73.305 6.22 73.625 6.545 ;
      RECT 73.335 5.695 73.505 6.545 ;
      RECT 73.335 5.695 73.51 6.045 ;
      RECT 73.335 5.695 74.31 5.87 ;
      RECT 74.135 1.965 74.31 5.87 ;
      RECT 74.08 1.965 74.43 2.315 ;
      RECT 74.105 6.655 74.43 6.98 ;
      RECT 72.99 6.745 74.43 6.915 ;
      RECT 72.99 2.395 73.15 6.915 ;
      RECT 73.305 2.365 73.625 2.685 ;
      RECT 72.99 2.395 73.625 2.565 ;
      RECT 67.825 4.135 71.96 4.325 ;
      RECT 71.79 3.145 71.96 4.325 ;
      RECT 71.77 3.15 71.96 4.325 ;
      RECT 67.825 3.515 68.015 4.325 ;
      RECT 67.775 3.515 68.055 3.885 ;
      RECT 71.7 3.15 72.04 3.5 ;
      RECT 57.88 6.655 58.23 7.005 ;
      RECT 68.665 6.61 69.015 6.96 ;
      RECT 57.88 6.685 69.015 6.885 ;
      RECT 68.305 2.98 68.565 3.3 ;
      RECT 68.365 1.86 68.505 3.3 ;
      RECT 68.305 1.86 68.565 2.18 ;
      RECT 67.305 3.54 67.565 3.86 ;
      RECT 67.305 2.955 67.505 3.86 ;
      RECT 67.245 1.86 67.385 3.49 ;
      RECT 67.245 2.955 67.745 3.325 ;
      RECT 67.185 1.86 67.445 2.18 ;
      RECT 66.825 3.54 67.085 3.86 ;
      RECT 66.885 1.95 67.025 3.86 ;
      RECT 66.585 1.95 67.025 2.18 ;
      RECT 66.585 1.86 66.845 2.18 ;
      RECT 66.345 2.42 66.605 2.74 ;
      RECT 65.765 2.51 66.605 2.65 ;
      RECT 65.765 1.57 65.905 2.65 ;
      RECT 62.425 1.86 62.685 2.18 ;
      RECT 62.425 1.95 63.465 2.09 ;
      RECT 63.325 1.57 63.465 2.09 ;
      RECT 63.325 1.57 65.905 1.71 ;
      RECT 65.815 3.515 66.095 3.885 ;
      RECT 65.885 3.07 66.025 3.885 ;
      RECT 65.695 2.955 65.975 3.325 ;
      RECT 65.405 3.07 66.025 3.21 ;
      RECT 65.405 1.86 65.545 3.21 ;
      RECT 65.345 1.86 65.605 2.18 ;
      RECT 64.615 2.955 64.895 3.325 ;
      RECT 64.685 1.86 64.825 3.325 ;
      RECT 64.625 1.86 64.885 2.18 ;
      RECT 64.265 3.54 64.525 3.86 ;
      RECT 64.325 1.95 64.465 3.86 ;
      RECT 63.905 1.86 64.165 2.18 ;
      RECT 63.905 1.95 64.465 2.09 ;
      RECT 61.935 2.955 62.215 3.325 ;
      RECT 63.905 2.98 64.165 3.3 ;
      RECT 61.585 2.98 62.215 3.3 ;
      RECT 61.585 3.07 64.165 3.21 ;
      RECT 63.375 2.395 63.655 2.765 ;
      RECT 63.375 2.42 63.905 2.74 ;
      RECT 60.465 2.98 60.725 3.3 ;
      RECT 60.525 1.86 60.665 3.3 ;
      RECT 60.465 1.86 60.725 2.18 ;
      RECT 59.495 3.515 59.775 3.885 ;
      RECT 59.505 3.26 59.765 3.885 ;
      RECT 54.745 6.22 55.065 6.545 ;
      RECT 54.775 5.695 54.945 6.545 ;
      RECT 54.775 5.695 54.95 6.045 ;
      RECT 54.775 5.695 55.75 5.87 ;
      RECT 55.575 1.965 55.75 5.87 ;
      RECT 55.52 1.965 55.87 2.315 ;
      RECT 55.545 6.655 55.87 6.98 ;
      RECT 54.43 6.745 55.87 6.915 ;
      RECT 54.43 2.395 54.59 6.915 ;
      RECT 54.745 2.365 55.065 2.685 ;
      RECT 54.43 2.395 55.065 2.565 ;
      RECT 49.265 4.135 53.4 4.325 ;
      RECT 53.23 3.145 53.4 4.325 ;
      RECT 53.21 3.15 53.4 4.325 ;
      RECT 49.265 3.515 49.455 4.325 ;
      RECT 49.215 3.515 49.495 3.885 ;
      RECT 53.14 3.15 53.48 3.5 ;
      RECT 39.365 6.66 39.715 7.01 ;
      RECT 50.105 6.615 50.455 6.965 ;
      RECT 39.365 6.69 50.455 6.89 ;
      RECT 49.745 2.98 50.005 3.3 ;
      RECT 49.805 1.86 49.945 3.3 ;
      RECT 49.745 1.86 50.005 2.18 ;
      RECT 48.745 3.54 49.005 3.86 ;
      RECT 48.745 2.955 48.945 3.86 ;
      RECT 48.685 1.86 48.825 3.49 ;
      RECT 48.685 2.955 49.185 3.325 ;
      RECT 48.625 1.86 48.885 2.18 ;
      RECT 48.265 3.54 48.525 3.86 ;
      RECT 48.325 1.95 48.465 3.86 ;
      RECT 48.025 1.95 48.465 2.18 ;
      RECT 48.025 1.86 48.285 2.18 ;
      RECT 47.785 2.42 48.045 2.74 ;
      RECT 47.205 2.51 48.045 2.65 ;
      RECT 47.205 1.57 47.345 2.65 ;
      RECT 43.865 1.86 44.125 2.18 ;
      RECT 43.865 1.95 44.905 2.09 ;
      RECT 44.765 1.57 44.905 2.09 ;
      RECT 44.765 1.57 47.345 1.71 ;
      RECT 47.255 3.515 47.535 3.885 ;
      RECT 47.325 3.07 47.465 3.885 ;
      RECT 47.135 2.955 47.415 3.325 ;
      RECT 46.845 3.07 47.465 3.21 ;
      RECT 46.845 1.86 46.985 3.21 ;
      RECT 46.785 1.86 47.045 2.18 ;
      RECT 46.055 2.955 46.335 3.325 ;
      RECT 46.125 1.86 46.265 3.325 ;
      RECT 46.065 1.86 46.325 2.18 ;
      RECT 45.705 3.54 45.965 3.86 ;
      RECT 45.765 1.95 45.905 3.86 ;
      RECT 45.345 1.86 45.605 2.18 ;
      RECT 45.345 1.95 45.905 2.09 ;
      RECT 43.375 2.955 43.655 3.325 ;
      RECT 45.345 2.98 45.605 3.3 ;
      RECT 43.025 2.98 43.655 3.3 ;
      RECT 43.025 3.07 45.605 3.21 ;
      RECT 44.815 2.395 45.095 2.765 ;
      RECT 44.815 2.42 45.345 2.74 ;
      RECT 41.905 2.98 42.165 3.3 ;
      RECT 41.965 1.86 42.105 3.3 ;
      RECT 41.905 1.86 42.165 2.18 ;
      RECT 40.935 3.515 41.215 3.885 ;
      RECT 40.945 3.26 41.205 3.885 ;
      RECT 36.185 6.22 36.505 6.545 ;
      RECT 36.215 5.695 36.385 6.545 ;
      RECT 36.215 5.695 36.39 6.045 ;
      RECT 36.215 5.695 37.19 5.87 ;
      RECT 37.015 1.965 37.19 5.87 ;
      RECT 36.96 1.965 37.31 2.315 ;
      RECT 36.985 6.655 37.31 6.98 ;
      RECT 35.87 6.745 37.31 6.915 ;
      RECT 35.87 2.395 36.03 6.915 ;
      RECT 36.185 2.365 36.505 2.685 ;
      RECT 35.87 2.395 36.505 2.565 ;
      RECT 30.705 4.135 34.84 4.325 ;
      RECT 34.67 3.145 34.84 4.325 ;
      RECT 34.65 3.15 34.84 4.325 ;
      RECT 30.705 3.515 30.895 4.325 ;
      RECT 30.655 3.515 30.935 3.885 ;
      RECT 34.58 3.15 34.92 3.5 ;
      RECT 20.805 6.655 21.155 7.005 ;
      RECT 31.55 6.61 31.9 6.96 ;
      RECT 20.805 6.685 31.9 6.885 ;
      RECT 31.185 2.98 31.445 3.3 ;
      RECT 31.245 1.86 31.385 3.3 ;
      RECT 31.185 1.86 31.445 2.18 ;
      RECT 30.185 3.54 30.445 3.86 ;
      RECT 30.185 2.955 30.385 3.86 ;
      RECT 30.125 1.86 30.265 3.49 ;
      RECT 30.125 2.955 30.625 3.325 ;
      RECT 30.065 1.86 30.325 2.18 ;
      RECT 29.705 3.54 29.965 3.86 ;
      RECT 29.765 1.95 29.905 3.86 ;
      RECT 29.465 1.95 29.905 2.18 ;
      RECT 29.465 1.86 29.725 2.18 ;
      RECT 29.225 2.42 29.485 2.74 ;
      RECT 28.645 2.51 29.485 2.65 ;
      RECT 28.645 1.57 28.785 2.65 ;
      RECT 25.305 1.86 25.565 2.18 ;
      RECT 25.305 1.95 26.345 2.09 ;
      RECT 26.205 1.57 26.345 2.09 ;
      RECT 26.205 1.57 28.785 1.71 ;
      RECT 28.695 3.515 28.975 3.885 ;
      RECT 28.765 3.07 28.905 3.885 ;
      RECT 28.575 2.955 28.855 3.325 ;
      RECT 28.285 3.07 28.905 3.21 ;
      RECT 28.285 1.86 28.425 3.21 ;
      RECT 28.225 1.86 28.485 2.18 ;
      RECT 27.495 2.955 27.775 3.325 ;
      RECT 27.565 1.86 27.705 3.325 ;
      RECT 27.505 1.86 27.765 2.18 ;
      RECT 27.145 3.54 27.405 3.86 ;
      RECT 27.205 1.95 27.345 3.86 ;
      RECT 26.785 1.86 27.045 2.18 ;
      RECT 26.785 1.95 27.345 2.09 ;
      RECT 24.815 2.955 25.095 3.325 ;
      RECT 26.785 2.98 27.045 3.3 ;
      RECT 24.465 2.98 25.095 3.3 ;
      RECT 24.465 3.07 27.045 3.21 ;
      RECT 26.255 2.395 26.535 2.765 ;
      RECT 26.255 2.42 26.785 2.74 ;
      RECT 23.345 2.98 23.605 3.3 ;
      RECT 23.405 1.86 23.545 3.3 ;
      RECT 23.345 1.86 23.605 2.18 ;
      RECT 22.375 3.515 22.655 3.885 ;
      RECT 22.385 3.26 22.645 3.885 ;
      RECT 17.625 6.22 17.945 6.545 ;
      RECT 17.655 5.695 17.825 6.545 ;
      RECT 17.655 5.695 17.83 6.045 ;
      RECT 17.655 5.695 18.63 5.87 ;
      RECT 18.455 1.965 18.63 5.87 ;
      RECT 18.4 1.965 18.75 2.315 ;
      RECT 18.425 6.655 18.75 6.98 ;
      RECT 17.31 6.745 18.75 6.915 ;
      RECT 17.31 2.395 17.47 6.915 ;
      RECT 17.625 2.365 17.945 2.685 ;
      RECT 17.31 2.395 17.945 2.565 ;
      RECT 12.145 4.135 16.28 4.325 ;
      RECT 16.11 3.145 16.28 4.325 ;
      RECT 16.09 3.15 16.28 4.325 ;
      RECT 12.145 3.515 12.335 4.325 ;
      RECT 12.095 3.515 12.375 3.885 ;
      RECT 16.02 3.15 16.36 3.5 ;
      RECT 1.54 6.995 1.83 7.345 ;
      RECT 1.54 7.05 2.855 7.22 ;
      RECT 2.685 6.685 2.855 7.22 ;
      RECT 12.99 6.605 13.34 6.955 ;
      RECT 2.685 6.685 13.34 6.855 ;
      RECT 12.625 2.98 12.885 3.3 ;
      RECT 12.685 1.86 12.825 3.3 ;
      RECT 12.625 1.86 12.885 2.18 ;
      RECT 11.625 3.54 11.885 3.86 ;
      RECT 11.625 2.955 11.825 3.86 ;
      RECT 11.565 1.86 11.705 3.49 ;
      RECT 11.565 2.955 12.065 3.325 ;
      RECT 11.505 1.86 11.765 2.18 ;
      RECT 11.145 3.54 11.405 3.86 ;
      RECT 11.205 1.95 11.345 3.86 ;
      RECT 10.905 1.95 11.345 2.18 ;
      RECT 10.905 1.86 11.165 2.18 ;
      RECT 10.665 2.42 10.925 2.74 ;
      RECT 10.085 2.51 10.925 2.65 ;
      RECT 10.085 1.57 10.225 2.65 ;
      RECT 6.745 1.86 7.005 2.18 ;
      RECT 6.745 1.95 7.785 2.09 ;
      RECT 7.645 1.57 7.785 2.09 ;
      RECT 7.645 1.57 10.225 1.71 ;
      RECT 10.135 3.515 10.415 3.885 ;
      RECT 10.205 3.07 10.345 3.885 ;
      RECT 10.015 2.955 10.295 3.325 ;
      RECT 9.725 3.07 10.345 3.21 ;
      RECT 9.725 1.86 9.865 3.21 ;
      RECT 9.665 1.86 9.925 2.18 ;
      RECT 8.935 2.955 9.215 3.325 ;
      RECT 9.005 1.86 9.145 3.325 ;
      RECT 8.945 1.86 9.205 2.18 ;
      RECT 8.585 3.54 8.845 3.86 ;
      RECT 8.645 1.95 8.785 3.86 ;
      RECT 8.225 1.86 8.485 2.18 ;
      RECT 8.225 1.95 8.785 2.09 ;
      RECT 4.785 2.98 5.045 3.3 ;
      RECT 4.845 1.86 4.985 3.3 ;
      RECT 4.785 1.86 5.045 2.18 ;
      RECT 3.815 3.515 4.095 3.885 ;
      RECT 3.825 3.26 4.085 3.885 ;
      RECT 88.295 1.835 88.575 2.205 ;
      RECT 87.335 3.515 87.615 3.885 ;
      RECT 86.555 7.055 86.93 7.425 ;
      RECT 78.535 2.395 78.815 2.765 ;
      RECT 69.735 1.835 70.015 2.205 ;
      RECT 68.775 3.515 69.055 3.885 ;
      RECT 67.995 7.055 68.37 7.425 ;
      RECT 59.975 2.395 60.255 2.765 ;
      RECT 51.175 1.835 51.455 2.205 ;
      RECT 50.215 3.515 50.495 3.885 ;
      RECT 49.435 7.055 49.81 7.425 ;
      RECT 41.415 2.395 41.695 2.765 ;
      RECT 32.615 1.835 32.895 2.205 ;
      RECT 31.655 3.515 31.935 3.885 ;
      RECT 30.875 7.055 31.25 7.425 ;
      RECT 22.855 2.395 23.135 2.765 ;
      RECT 14.055 1.835 14.335 2.205 ;
      RECT 13.095 3.515 13.375 3.885 ;
    LAYER via1 ;
      RECT 95.125 7.375 95.275 7.525 ;
      RECT 92.755 6.74 92.905 6.89 ;
      RECT 92.74 2.065 92.89 2.215 ;
      RECT 91.95 2.45 92.1 2.6 ;
      RECT 91.95 6.325 92.1 6.475 ;
      RECT 90.36 3.25 90.51 3.4 ;
      RECT 88.36 1.945 88.51 2.095 ;
      RECT 87.4 3.625 87.55 3.775 ;
      RECT 87.325 6.71 87.475 6.86 ;
      RECT 86.92 1.945 87.07 2.095 ;
      RECT 86.92 3.065 87.07 3.215 ;
      RECT 86.665 7.165 86.815 7.315 ;
      RECT 86.4 3.625 86.55 3.775 ;
      RECT 85.92 3.625 86.07 3.775 ;
      RECT 85.8 1.945 85.95 2.095 ;
      RECT 85.44 3.625 85.59 3.775 ;
      RECT 85.2 1.945 85.35 2.095 ;
      RECT 84.96 2.505 85.11 2.655 ;
      RECT 84.44 3.625 84.59 3.775 ;
      RECT 83.96 1.945 84.11 2.095 ;
      RECT 83.24 1.945 83.39 2.095 ;
      RECT 83.24 3.065 83.39 3.215 ;
      RECT 82.88 3.625 83.03 3.775 ;
      RECT 82.52 1.945 82.67 2.095 ;
      RECT 82.52 3.065 82.67 3.215 ;
      RECT 82.26 2.505 82.41 2.655 ;
      RECT 81.04 1.945 81.19 2.095 ;
      RECT 80.2 3.065 80.35 3.215 ;
      RECT 79.08 1.945 79.23 2.095 ;
      RECT 79.08 3.065 79.23 3.215 ;
      RECT 78.6 2.505 78.75 2.655 ;
      RECT 78.12 3.345 78.27 3.495 ;
      RECT 76.54 6.755 76.69 6.905 ;
      RECT 74.195 6.74 74.345 6.89 ;
      RECT 74.18 2.065 74.33 2.215 ;
      RECT 73.39 2.45 73.54 2.6 ;
      RECT 73.39 6.325 73.54 6.475 ;
      RECT 71.8 3.25 71.95 3.4 ;
      RECT 69.8 1.945 69.95 2.095 ;
      RECT 68.84 3.625 68.99 3.775 ;
      RECT 68.765 6.71 68.915 6.86 ;
      RECT 68.36 1.945 68.51 2.095 ;
      RECT 68.36 3.065 68.51 3.215 ;
      RECT 68.105 7.165 68.255 7.315 ;
      RECT 67.84 3.625 67.99 3.775 ;
      RECT 67.36 3.625 67.51 3.775 ;
      RECT 67.24 1.945 67.39 2.095 ;
      RECT 66.88 3.625 67.03 3.775 ;
      RECT 66.64 1.945 66.79 2.095 ;
      RECT 66.4 2.505 66.55 2.655 ;
      RECT 65.88 3.625 66.03 3.775 ;
      RECT 65.4 1.945 65.55 2.095 ;
      RECT 64.68 1.945 64.83 2.095 ;
      RECT 64.68 3.065 64.83 3.215 ;
      RECT 64.32 3.625 64.47 3.775 ;
      RECT 63.96 1.945 64.11 2.095 ;
      RECT 63.96 3.065 64.11 3.215 ;
      RECT 63.7 2.505 63.85 2.655 ;
      RECT 62.48 1.945 62.63 2.095 ;
      RECT 61.64 3.065 61.79 3.215 ;
      RECT 60.52 1.945 60.67 2.095 ;
      RECT 60.52 3.065 60.67 3.215 ;
      RECT 60.04 2.505 60.19 2.655 ;
      RECT 59.56 3.345 59.71 3.495 ;
      RECT 57.98 6.755 58.13 6.905 ;
      RECT 55.635 6.74 55.785 6.89 ;
      RECT 55.62 2.065 55.77 2.215 ;
      RECT 54.83 2.45 54.98 2.6 ;
      RECT 54.83 6.325 54.98 6.475 ;
      RECT 53.24 3.25 53.39 3.4 ;
      RECT 51.24 1.945 51.39 2.095 ;
      RECT 50.28 3.625 50.43 3.775 ;
      RECT 50.205 6.715 50.355 6.865 ;
      RECT 49.8 1.945 49.95 2.095 ;
      RECT 49.8 3.065 49.95 3.215 ;
      RECT 49.545 7.165 49.695 7.315 ;
      RECT 49.28 3.625 49.43 3.775 ;
      RECT 48.8 3.625 48.95 3.775 ;
      RECT 48.68 1.945 48.83 2.095 ;
      RECT 48.32 3.625 48.47 3.775 ;
      RECT 48.08 1.945 48.23 2.095 ;
      RECT 47.84 2.505 47.99 2.655 ;
      RECT 47.32 3.625 47.47 3.775 ;
      RECT 46.84 1.945 46.99 2.095 ;
      RECT 46.12 1.945 46.27 2.095 ;
      RECT 46.12 3.065 46.27 3.215 ;
      RECT 45.76 3.625 45.91 3.775 ;
      RECT 45.4 1.945 45.55 2.095 ;
      RECT 45.4 3.065 45.55 3.215 ;
      RECT 45.14 2.505 45.29 2.655 ;
      RECT 43.92 1.945 44.07 2.095 ;
      RECT 43.08 3.065 43.23 3.215 ;
      RECT 41.96 1.945 42.11 2.095 ;
      RECT 41.96 3.065 42.11 3.215 ;
      RECT 41.48 2.505 41.63 2.655 ;
      RECT 41 3.345 41.15 3.495 ;
      RECT 39.465 6.76 39.615 6.91 ;
      RECT 37.075 6.74 37.225 6.89 ;
      RECT 37.06 2.065 37.21 2.215 ;
      RECT 36.27 2.45 36.42 2.6 ;
      RECT 36.27 6.325 36.42 6.475 ;
      RECT 34.68 3.25 34.83 3.4 ;
      RECT 32.68 1.945 32.83 2.095 ;
      RECT 31.72 3.625 31.87 3.775 ;
      RECT 31.65 6.71 31.8 6.86 ;
      RECT 31.24 1.945 31.39 2.095 ;
      RECT 31.24 3.065 31.39 3.215 ;
      RECT 30.985 7.165 31.135 7.315 ;
      RECT 30.72 3.625 30.87 3.775 ;
      RECT 30.24 3.625 30.39 3.775 ;
      RECT 30.12 1.945 30.27 2.095 ;
      RECT 29.76 3.625 29.91 3.775 ;
      RECT 29.52 1.945 29.67 2.095 ;
      RECT 29.28 2.505 29.43 2.655 ;
      RECT 28.76 3.625 28.91 3.775 ;
      RECT 28.28 1.945 28.43 2.095 ;
      RECT 27.56 1.945 27.71 2.095 ;
      RECT 27.56 3.065 27.71 3.215 ;
      RECT 27.2 3.625 27.35 3.775 ;
      RECT 26.84 1.945 26.99 2.095 ;
      RECT 26.84 3.065 26.99 3.215 ;
      RECT 26.58 2.505 26.73 2.655 ;
      RECT 25.36 1.945 25.51 2.095 ;
      RECT 24.52 3.065 24.67 3.215 ;
      RECT 23.4 1.945 23.55 2.095 ;
      RECT 23.4 3.065 23.55 3.215 ;
      RECT 22.92 2.505 23.07 2.655 ;
      RECT 22.44 3.345 22.59 3.495 ;
      RECT 20.905 6.755 21.055 6.905 ;
      RECT 18.515 6.74 18.665 6.89 ;
      RECT 18.5 2.065 18.65 2.215 ;
      RECT 17.71 2.45 17.86 2.6 ;
      RECT 17.71 6.325 17.86 6.475 ;
      RECT 16.12 3.25 16.27 3.4 ;
      RECT 14.12 1.945 14.27 2.095 ;
      RECT 13.16 3.625 13.31 3.775 ;
      RECT 13.09 6.705 13.24 6.855 ;
      RECT 12.68 1.945 12.83 2.095 ;
      RECT 12.68 3.065 12.83 3.215 ;
      RECT 12.16 3.625 12.31 3.775 ;
      RECT 11.68 3.625 11.83 3.775 ;
      RECT 11.56 1.945 11.71 2.095 ;
      RECT 11.2 3.625 11.35 3.775 ;
      RECT 10.96 1.945 11.11 2.095 ;
      RECT 10.72 2.505 10.87 2.655 ;
      RECT 10.2 3.625 10.35 3.775 ;
      RECT 9.72 1.945 9.87 2.095 ;
      RECT 9 1.945 9.15 2.095 ;
      RECT 9 3.065 9.15 3.215 ;
      RECT 8.64 3.625 8.79 3.775 ;
      RECT 8.28 1.945 8.43 2.095 ;
      RECT 6.8 1.945 6.95 2.095 ;
      RECT 4.84 1.945 4.99 2.095 ;
      RECT 4.84 3.065 4.99 3.215 ;
      RECT 3.88 3.345 4.03 3.495 ;
      RECT 1.61 7.095 1.76 7.245 ;
      RECT 1.235 6.355 1.385 6.505 ;
    LAYER met1 ;
      RECT 94.99 7.77 95.28 8 ;
      RECT 95.05 6.29 95.22 8 ;
      RECT 95.025 7.275 95.375 7.625 ;
      RECT 94.99 6.29 95.28 6.52 ;
      RECT 94.585 2.395 94.69 2.965 ;
      RECT 94.585 2.73 94.91 2.96 ;
      RECT 94.585 2.76 95.08 2.93 ;
      RECT 94.585 2.395 94.775 2.96 ;
      RECT 94 2.36 94.29 2.59 ;
      RECT 94 2.395 94.775 2.565 ;
      RECT 94.06 0.88 94.23 2.59 ;
      RECT 94 0.88 94.29 1.11 ;
      RECT 94 7.77 94.29 8 ;
      RECT 94.06 6.29 94.23 8 ;
      RECT 94 6.29 94.29 6.52 ;
      RECT 94 6.325 94.855 6.485 ;
      RECT 94.685 5.92 94.855 6.485 ;
      RECT 94 6.32 94.395 6.485 ;
      RECT 94.62 5.92 94.91 6.15 ;
      RECT 94.62 5.95 95.08 6.12 ;
      RECT 93.63 2.73 93.92 2.96 ;
      RECT 93.63 2.76 94.09 2.93 ;
      RECT 93.695 1.655 93.86 2.96 ;
      RECT 92.21 1.625 92.5 1.855 ;
      RECT 92.21 1.655 93.86 1.825 ;
      RECT 92.27 0.885 92.44 1.855 ;
      RECT 92.21 0.885 92.5 1.115 ;
      RECT 92.21 7.765 92.5 7.995 ;
      RECT 92.27 7.025 92.44 7.995 ;
      RECT 92.27 7.12 93.86 7.29 ;
      RECT 93.69 5.92 93.86 7.29 ;
      RECT 92.21 7.025 92.5 7.255 ;
      RECT 93.63 5.92 93.92 6.15 ;
      RECT 93.63 5.95 94.09 6.12 ;
      RECT 90.26 3.15 90.6 3.5 ;
      RECT 90.35 2.025 90.52 3.5 ;
      RECT 92.64 1.965 92.99 2.315 ;
      RECT 90.35 2.025 92.99 2.195 ;
      RECT 92.665 6.655 92.99 6.98 ;
      RECT 87.225 6.61 87.575 6.96 ;
      RECT 92.64 6.655 92.99 6.885 ;
      RECT 87.025 6.655 87.575 6.885 ;
      RECT 86.855 6.685 92.99 6.855 ;
      RECT 91.865 2.365 92.185 2.685 ;
      RECT 91.835 2.365 92.185 2.595 ;
      RECT 91.665 2.395 92.185 2.565 ;
      RECT 91.865 6.255 92.185 6.545 ;
      RECT 91.835 6.285 92.185 6.515 ;
      RECT 91.665 6.315 92.185 6.485 ;
      RECT 87.315 3.57 87.635 3.83 ;
      RECT 88.605 2.745 88.745 3.605 ;
      RECT 87.405 3.465 88.745 3.605 ;
      RECT 87.405 3.025 87.545 3.83 ;
      RECT 87.33 3.025 87.62 3.255 ;
      RECT 88.53 2.745 88.82 2.975 ;
      RECT 88.05 3.025 88.34 3.255 ;
      RECT 88.245 1.95 88.385 3.21 ;
      RECT 88.275 1.89 88.595 2.15 ;
      RECT 84.875 2.45 85.195 2.71 ;
      RECT 87.57 2.465 87.86 2.695 ;
      RECT 84.965 2.37 87.785 2.51 ;
      RECT 86.835 1.89 87.155 2.15 ;
      RECT 87.33 1.905 87.62 2.135 ;
      RECT 86.835 1.95 87.62 2.09 ;
      RECT 86.835 3.01 87.155 3.27 ;
      RECT 86.835 2.79 87.065 3.27 ;
      RECT 86.33 2.745 86.62 2.975 ;
      RECT 86.33 2.79 87.065 2.93 ;
      RECT 86.595 7.765 86.885 7.995 ;
      RECT 86.655 7.025 86.825 7.995 ;
      RECT 86.555 7.055 86.935 7.425 ;
      RECT 86.595 7.025 86.885 7.425 ;
      RECT 85.355 3.57 85.675 3.83 ;
      RECT 84.89 3.585 85.18 3.815 ;
      RECT 84.89 3.63 85.675 3.77 ;
      RECT 83.65 2.465 83.94 2.695 ;
      RECT 83.65 2.51 84.585 2.65 ;
      RECT 84.445 1.95 84.585 2.65 ;
      RECT 85.115 1.89 85.435 2.15 ;
      RECT 84.89 1.905 85.435 2.135 ;
      RECT 84.445 1.95 85.435 2.09 ;
      RECT 82.795 3.57 83.115 3.83 ;
      RECT 82.795 3.63 83.865 3.77 ;
      RECT 83.725 3.07 83.865 3.77 ;
      RECT 84.89 3.025 85.18 3.255 ;
      RECT 83.725 3.07 85.18 3.21 ;
      RECT 83.155 1.89 83.475 2.15 ;
      RECT 82.93 1.905 83.475 2.135 ;
      RECT 82.175 2.45 82.495 2.71 ;
      RECT 83.17 2.465 83.46 2.695 ;
      RECT 81.93 2.465 82.495 2.695 ;
      RECT 81.93 2.51 83.46 2.65 ;
      RECT 81.45 3.025 81.74 3.255 ;
      RECT 81.645 1.95 81.785 3.21 ;
      RECT 82.435 1.89 82.755 2.15 ;
      RECT 81.45 1.905 81.74 2.135 ;
      RECT 81.45 1.95 82.755 2.09 ;
      RECT 81.045 3.465 82.145 3.605 ;
      RECT 81.93 3.305 82.22 3.535 ;
      RECT 80.97 3.305 81.26 3.535 ;
      RECT 80.955 1.89 81.275 2.15 ;
      RECT 78.995 1.89 79.315 2.15 ;
      RECT 78.995 1.95 81.275 2.09 ;
      RECT 80.115 3.01 80.435 3.27 ;
      RECT 80.115 3.01 80.945 3.15 ;
      RECT 80.73 2.745 80.945 3.15 ;
      RECT 80.73 2.745 81.02 2.975 ;
      RECT 78.515 2.45 78.835 2.71 ;
      RECT 79.925 2.465 80.215 2.695 ;
      RECT 78.515 2.465 79.06 2.695 ;
      RECT 78.515 2.55 79.465 2.69 ;
      RECT 79.325 2.37 79.465 2.69 ;
      RECT 79.825 2.465 80.215 2.65 ;
      RECT 79.325 2.37 79.965 2.51 ;
      RECT 78.035 3.26 78.355 3.675 ;
      RECT 78.115 1.905 78.27 3.675 ;
      RECT 78.05 1.905 78.34 2.135 ;
      RECT 76.43 7.77 76.72 8 ;
      RECT 76.49 6.29 76.66 8 ;
      RECT 76.44 6.655 76.79 7.005 ;
      RECT 76.43 6.29 76.72 6.52 ;
      RECT 76.025 2.395 76.13 2.965 ;
      RECT 76.025 2.73 76.35 2.96 ;
      RECT 76.025 2.76 76.52 2.93 ;
      RECT 76.025 2.395 76.215 2.96 ;
      RECT 75.44 2.36 75.73 2.59 ;
      RECT 75.44 2.395 76.215 2.565 ;
      RECT 75.5 0.88 75.67 2.59 ;
      RECT 75.44 0.88 75.73 1.11 ;
      RECT 75.44 7.77 75.73 8 ;
      RECT 75.5 6.29 75.67 8 ;
      RECT 75.44 6.29 75.73 6.52 ;
      RECT 75.44 6.325 76.295 6.485 ;
      RECT 76.125 5.92 76.295 6.485 ;
      RECT 75.44 6.32 75.835 6.485 ;
      RECT 76.06 5.92 76.35 6.15 ;
      RECT 76.06 5.95 76.52 6.12 ;
      RECT 75.07 2.73 75.36 2.96 ;
      RECT 75.07 2.76 75.53 2.93 ;
      RECT 75.135 1.655 75.3 2.96 ;
      RECT 73.65 1.625 73.94 1.855 ;
      RECT 73.65 1.655 75.3 1.825 ;
      RECT 73.71 0.885 73.88 1.855 ;
      RECT 73.65 0.885 73.94 1.115 ;
      RECT 73.65 7.765 73.94 7.995 ;
      RECT 73.71 7.025 73.88 7.995 ;
      RECT 73.71 7.12 75.3 7.29 ;
      RECT 75.13 5.92 75.3 7.29 ;
      RECT 73.65 7.025 73.94 7.255 ;
      RECT 75.07 5.92 75.36 6.15 ;
      RECT 75.07 5.95 75.53 6.12 ;
      RECT 71.7 3.15 72.04 3.5 ;
      RECT 71.79 2.025 71.96 3.5 ;
      RECT 74.08 1.965 74.43 2.315 ;
      RECT 71.79 2.025 74.43 2.195 ;
      RECT 74.105 6.655 74.43 6.98 ;
      RECT 68.665 6.61 69.015 6.96 ;
      RECT 74.08 6.655 74.43 6.885 ;
      RECT 68.465 6.655 69.015 6.885 ;
      RECT 68.295 6.685 74.43 6.855 ;
      RECT 73.305 2.365 73.625 2.685 ;
      RECT 73.275 2.365 73.625 2.595 ;
      RECT 73.105 2.395 73.625 2.565 ;
      RECT 73.305 6.255 73.625 6.545 ;
      RECT 73.275 6.285 73.625 6.515 ;
      RECT 73.105 6.315 73.625 6.485 ;
      RECT 68.755 3.57 69.075 3.83 ;
      RECT 70.045 2.745 70.185 3.605 ;
      RECT 68.845 3.465 70.185 3.605 ;
      RECT 68.845 3.025 68.985 3.83 ;
      RECT 68.77 3.025 69.06 3.255 ;
      RECT 69.97 2.745 70.26 2.975 ;
      RECT 69.49 3.025 69.78 3.255 ;
      RECT 69.685 1.95 69.825 3.21 ;
      RECT 69.715 1.89 70.035 2.15 ;
      RECT 66.315 2.45 66.635 2.71 ;
      RECT 69.01 2.465 69.3 2.695 ;
      RECT 66.405 2.37 69.225 2.51 ;
      RECT 68.275 1.89 68.595 2.15 ;
      RECT 68.77 1.905 69.06 2.135 ;
      RECT 68.275 1.95 69.06 2.09 ;
      RECT 68.275 3.01 68.595 3.27 ;
      RECT 68.275 2.79 68.505 3.27 ;
      RECT 67.77 2.745 68.06 2.975 ;
      RECT 67.77 2.79 68.505 2.93 ;
      RECT 68.035 7.765 68.325 7.995 ;
      RECT 68.095 7.025 68.265 7.995 ;
      RECT 67.995 7.055 68.375 7.425 ;
      RECT 68.035 7.025 68.325 7.425 ;
      RECT 66.795 3.57 67.115 3.83 ;
      RECT 66.33 3.585 66.62 3.815 ;
      RECT 66.33 3.63 67.115 3.77 ;
      RECT 65.09 2.465 65.38 2.695 ;
      RECT 65.09 2.51 66.025 2.65 ;
      RECT 65.885 1.95 66.025 2.65 ;
      RECT 66.555 1.89 66.875 2.15 ;
      RECT 66.33 1.905 66.875 2.135 ;
      RECT 65.885 1.95 66.875 2.09 ;
      RECT 64.235 3.57 64.555 3.83 ;
      RECT 64.235 3.63 65.305 3.77 ;
      RECT 65.165 3.07 65.305 3.77 ;
      RECT 66.33 3.025 66.62 3.255 ;
      RECT 65.165 3.07 66.62 3.21 ;
      RECT 64.595 1.89 64.915 2.15 ;
      RECT 64.37 1.905 64.915 2.135 ;
      RECT 63.615 2.45 63.935 2.71 ;
      RECT 64.61 2.465 64.9 2.695 ;
      RECT 63.37 2.465 63.935 2.695 ;
      RECT 63.37 2.51 64.9 2.65 ;
      RECT 62.89 3.025 63.18 3.255 ;
      RECT 63.085 1.95 63.225 3.21 ;
      RECT 63.875 1.89 64.195 2.15 ;
      RECT 62.89 1.905 63.18 2.135 ;
      RECT 62.89 1.95 64.195 2.09 ;
      RECT 62.485 3.465 63.585 3.605 ;
      RECT 63.37 3.305 63.66 3.535 ;
      RECT 62.41 3.305 62.7 3.535 ;
      RECT 62.395 1.89 62.715 2.15 ;
      RECT 60.435 1.89 60.755 2.15 ;
      RECT 60.435 1.95 62.715 2.09 ;
      RECT 61.555 3.01 61.875 3.27 ;
      RECT 61.555 3.01 62.385 3.15 ;
      RECT 62.17 2.745 62.385 3.15 ;
      RECT 62.17 2.745 62.46 2.975 ;
      RECT 59.955 2.45 60.275 2.71 ;
      RECT 61.365 2.465 61.655 2.695 ;
      RECT 59.955 2.465 60.5 2.695 ;
      RECT 59.955 2.55 60.905 2.69 ;
      RECT 60.765 2.37 60.905 2.69 ;
      RECT 61.265 2.465 61.655 2.65 ;
      RECT 60.765 2.37 61.405 2.51 ;
      RECT 59.475 3.26 59.795 3.675 ;
      RECT 59.555 1.905 59.71 3.675 ;
      RECT 59.49 1.905 59.78 2.135 ;
      RECT 57.87 7.77 58.16 8 ;
      RECT 57.93 6.29 58.1 8 ;
      RECT 57.88 6.655 58.23 7.005 ;
      RECT 57.87 6.29 58.16 6.52 ;
      RECT 57.465 2.395 57.57 2.965 ;
      RECT 57.465 2.73 57.79 2.96 ;
      RECT 57.465 2.76 57.96 2.93 ;
      RECT 57.465 2.395 57.655 2.96 ;
      RECT 56.88 2.36 57.17 2.59 ;
      RECT 56.88 2.395 57.655 2.565 ;
      RECT 56.94 0.88 57.11 2.59 ;
      RECT 56.88 0.88 57.17 1.11 ;
      RECT 56.88 7.77 57.17 8 ;
      RECT 56.94 6.29 57.11 8 ;
      RECT 56.88 6.29 57.17 6.52 ;
      RECT 56.88 6.325 57.735 6.485 ;
      RECT 57.565 5.92 57.735 6.485 ;
      RECT 56.88 6.32 57.275 6.485 ;
      RECT 57.5 5.92 57.79 6.15 ;
      RECT 57.5 5.95 57.96 6.12 ;
      RECT 56.51 2.73 56.8 2.96 ;
      RECT 56.51 2.76 56.97 2.93 ;
      RECT 56.575 1.655 56.74 2.96 ;
      RECT 55.09 1.625 55.38 1.855 ;
      RECT 55.09 1.655 56.74 1.825 ;
      RECT 55.15 0.885 55.32 1.855 ;
      RECT 55.09 0.885 55.38 1.115 ;
      RECT 55.09 7.765 55.38 7.995 ;
      RECT 55.15 7.025 55.32 7.995 ;
      RECT 55.15 7.12 56.74 7.29 ;
      RECT 56.57 5.92 56.74 7.29 ;
      RECT 55.09 7.025 55.38 7.255 ;
      RECT 56.51 5.92 56.8 6.15 ;
      RECT 56.51 5.95 56.97 6.12 ;
      RECT 53.14 3.15 53.48 3.5 ;
      RECT 53.23 2.025 53.4 3.5 ;
      RECT 55.52 1.965 55.87 2.315 ;
      RECT 53.23 2.025 55.87 2.195 ;
      RECT 55.545 6.655 55.87 6.98 ;
      RECT 50.105 6.615 50.455 6.965 ;
      RECT 55.52 6.655 55.87 6.885 ;
      RECT 49.905 6.655 50.455 6.885 ;
      RECT 49.735 6.685 55.87 6.855 ;
      RECT 54.745 2.365 55.065 2.685 ;
      RECT 54.715 2.365 55.065 2.595 ;
      RECT 54.545 2.395 55.065 2.565 ;
      RECT 54.745 6.255 55.065 6.545 ;
      RECT 54.715 6.285 55.065 6.515 ;
      RECT 54.545 6.315 55.065 6.485 ;
      RECT 50.195 3.57 50.515 3.83 ;
      RECT 51.485 2.745 51.625 3.605 ;
      RECT 50.285 3.465 51.625 3.605 ;
      RECT 50.285 3.025 50.425 3.83 ;
      RECT 50.21 3.025 50.5 3.255 ;
      RECT 51.41 2.745 51.7 2.975 ;
      RECT 50.93 3.025 51.22 3.255 ;
      RECT 51.125 1.95 51.265 3.21 ;
      RECT 51.155 1.89 51.475 2.15 ;
      RECT 47.755 2.45 48.075 2.71 ;
      RECT 50.45 2.465 50.74 2.695 ;
      RECT 47.845 2.37 50.665 2.51 ;
      RECT 49.715 1.89 50.035 2.15 ;
      RECT 50.21 1.905 50.5 2.135 ;
      RECT 49.715 1.95 50.5 2.09 ;
      RECT 49.715 3.01 50.035 3.27 ;
      RECT 49.715 2.79 49.945 3.27 ;
      RECT 49.21 2.745 49.5 2.975 ;
      RECT 49.21 2.79 49.945 2.93 ;
      RECT 49.475 7.765 49.765 7.995 ;
      RECT 49.535 7.025 49.705 7.995 ;
      RECT 49.435 7.055 49.815 7.425 ;
      RECT 49.475 7.025 49.765 7.425 ;
      RECT 48.235 3.57 48.555 3.83 ;
      RECT 47.77 3.585 48.06 3.815 ;
      RECT 47.77 3.63 48.555 3.77 ;
      RECT 46.53 2.465 46.82 2.695 ;
      RECT 46.53 2.51 47.465 2.65 ;
      RECT 47.325 1.95 47.465 2.65 ;
      RECT 47.995 1.89 48.315 2.15 ;
      RECT 47.77 1.905 48.315 2.135 ;
      RECT 47.325 1.95 48.315 2.09 ;
      RECT 45.675 3.57 45.995 3.83 ;
      RECT 45.675 3.63 46.745 3.77 ;
      RECT 46.605 3.07 46.745 3.77 ;
      RECT 47.77 3.025 48.06 3.255 ;
      RECT 46.605 3.07 48.06 3.21 ;
      RECT 46.035 1.89 46.355 2.15 ;
      RECT 45.81 1.905 46.355 2.135 ;
      RECT 45.055 2.45 45.375 2.71 ;
      RECT 46.05 2.465 46.34 2.695 ;
      RECT 44.81 2.465 45.375 2.695 ;
      RECT 44.81 2.51 46.34 2.65 ;
      RECT 44.33 3.025 44.62 3.255 ;
      RECT 44.525 1.95 44.665 3.21 ;
      RECT 45.315 1.89 45.635 2.15 ;
      RECT 44.33 1.905 44.62 2.135 ;
      RECT 44.33 1.95 45.635 2.09 ;
      RECT 43.925 3.465 45.025 3.605 ;
      RECT 44.81 3.305 45.1 3.535 ;
      RECT 43.85 3.305 44.14 3.535 ;
      RECT 43.835 1.89 44.155 2.15 ;
      RECT 41.875 1.89 42.195 2.15 ;
      RECT 41.875 1.95 44.155 2.09 ;
      RECT 42.995 3.01 43.315 3.27 ;
      RECT 42.995 3.01 43.825 3.15 ;
      RECT 43.61 2.745 43.825 3.15 ;
      RECT 43.61 2.745 43.9 2.975 ;
      RECT 41.395 2.45 41.715 2.71 ;
      RECT 42.805 2.465 43.095 2.695 ;
      RECT 41.395 2.465 41.94 2.695 ;
      RECT 41.395 2.55 42.345 2.69 ;
      RECT 42.205 2.37 42.345 2.69 ;
      RECT 42.705 2.465 43.095 2.65 ;
      RECT 42.205 2.37 42.845 2.51 ;
      RECT 40.915 3.26 41.235 3.675 ;
      RECT 40.995 1.905 41.15 3.675 ;
      RECT 40.93 1.905 41.22 2.135 ;
      RECT 39.31 7.77 39.6 8 ;
      RECT 39.37 6.29 39.54 8 ;
      RECT 39.36 6.66 39.715 7.015 ;
      RECT 39.31 6.29 39.6 6.52 ;
      RECT 38.905 2.395 39.01 2.965 ;
      RECT 38.905 2.73 39.23 2.96 ;
      RECT 38.905 2.76 39.4 2.93 ;
      RECT 38.905 2.395 39.095 2.96 ;
      RECT 38.32 2.36 38.61 2.59 ;
      RECT 38.32 2.395 39.095 2.565 ;
      RECT 38.38 0.88 38.55 2.59 ;
      RECT 38.32 0.88 38.61 1.11 ;
      RECT 38.32 7.77 38.61 8 ;
      RECT 38.38 6.29 38.55 8 ;
      RECT 38.32 6.29 38.61 6.52 ;
      RECT 38.32 6.325 39.175 6.485 ;
      RECT 39.005 5.92 39.175 6.485 ;
      RECT 38.32 6.32 38.715 6.485 ;
      RECT 38.94 5.92 39.23 6.15 ;
      RECT 38.94 5.95 39.4 6.12 ;
      RECT 37.95 2.73 38.24 2.96 ;
      RECT 37.95 2.76 38.41 2.93 ;
      RECT 38.015 1.655 38.18 2.96 ;
      RECT 36.53 1.625 36.82 1.855 ;
      RECT 36.53 1.655 38.18 1.825 ;
      RECT 36.59 0.885 36.76 1.855 ;
      RECT 36.53 0.885 36.82 1.115 ;
      RECT 36.53 7.765 36.82 7.995 ;
      RECT 36.59 7.025 36.76 7.995 ;
      RECT 36.59 7.12 38.18 7.29 ;
      RECT 38.01 5.92 38.18 7.29 ;
      RECT 36.53 7.025 36.82 7.255 ;
      RECT 37.95 5.92 38.24 6.15 ;
      RECT 37.95 5.95 38.41 6.12 ;
      RECT 34.58 3.15 34.92 3.5 ;
      RECT 34.67 2.025 34.84 3.5 ;
      RECT 36.96 1.965 37.31 2.315 ;
      RECT 34.67 2.025 37.31 2.195 ;
      RECT 36.985 6.655 37.31 6.98 ;
      RECT 31.55 6.61 31.9 6.96 ;
      RECT 36.96 6.655 37.31 6.885 ;
      RECT 31.345 6.655 31.9 6.885 ;
      RECT 31.175 6.685 37.31 6.855 ;
      RECT 36.185 2.365 36.505 2.685 ;
      RECT 36.155 2.365 36.505 2.595 ;
      RECT 35.985 2.395 36.505 2.565 ;
      RECT 36.185 6.255 36.505 6.545 ;
      RECT 36.155 6.285 36.505 6.515 ;
      RECT 35.985 6.315 36.505 6.485 ;
      RECT 31.635 3.57 31.955 3.83 ;
      RECT 32.925 2.745 33.065 3.605 ;
      RECT 31.725 3.465 33.065 3.605 ;
      RECT 31.725 3.025 31.865 3.83 ;
      RECT 31.65 3.025 31.94 3.255 ;
      RECT 32.85 2.745 33.14 2.975 ;
      RECT 32.37 3.025 32.66 3.255 ;
      RECT 32.565 1.95 32.705 3.21 ;
      RECT 32.595 1.89 32.915 2.15 ;
      RECT 29.195 2.45 29.515 2.71 ;
      RECT 31.89 2.465 32.18 2.695 ;
      RECT 29.285 2.37 32.105 2.51 ;
      RECT 31.155 1.89 31.475 2.15 ;
      RECT 31.65 1.905 31.94 2.135 ;
      RECT 31.155 1.95 31.94 2.09 ;
      RECT 31.155 3.01 31.475 3.27 ;
      RECT 31.155 2.79 31.385 3.27 ;
      RECT 30.65 2.745 30.94 2.975 ;
      RECT 30.65 2.79 31.385 2.93 ;
      RECT 30.915 7.765 31.205 7.995 ;
      RECT 30.975 7.025 31.145 7.995 ;
      RECT 30.875 7.055 31.255 7.425 ;
      RECT 30.915 7.025 31.205 7.425 ;
      RECT 29.675 3.57 29.995 3.83 ;
      RECT 29.21 3.585 29.5 3.815 ;
      RECT 29.21 3.63 29.995 3.77 ;
      RECT 27.97 2.465 28.26 2.695 ;
      RECT 27.97 2.51 28.905 2.65 ;
      RECT 28.765 1.95 28.905 2.65 ;
      RECT 29.435 1.89 29.755 2.15 ;
      RECT 29.21 1.905 29.755 2.135 ;
      RECT 28.765 1.95 29.755 2.09 ;
      RECT 27.115 3.57 27.435 3.83 ;
      RECT 27.115 3.63 28.185 3.77 ;
      RECT 28.045 3.07 28.185 3.77 ;
      RECT 29.21 3.025 29.5 3.255 ;
      RECT 28.045 3.07 29.5 3.21 ;
      RECT 27.475 1.89 27.795 2.15 ;
      RECT 27.25 1.905 27.795 2.135 ;
      RECT 26.495 2.45 26.815 2.71 ;
      RECT 27.49 2.465 27.78 2.695 ;
      RECT 26.25 2.465 26.815 2.695 ;
      RECT 26.25 2.51 27.78 2.65 ;
      RECT 25.77 3.025 26.06 3.255 ;
      RECT 25.965 1.95 26.105 3.21 ;
      RECT 26.755 1.89 27.075 2.15 ;
      RECT 25.77 1.905 26.06 2.135 ;
      RECT 25.77 1.95 27.075 2.09 ;
      RECT 25.365 3.465 26.465 3.605 ;
      RECT 26.25 3.305 26.54 3.535 ;
      RECT 25.29 3.305 25.58 3.535 ;
      RECT 25.275 1.89 25.595 2.15 ;
      RECT 23.315 1.89 23.635 2.15 ;
      RECT 23.315 1.95 25.595 2.09 ;
      RECT 24.435 3.01 24.755 3.27 ;
      RECT 24.435 3.01 25.265 3.15 ;
      RECT 25.05 2.745 25.265 3.15 ;
      RECT 25.05 2.745 25.34 2.975 ;
      RECT 22.835 2.45 23.155 2.71 ;
      RECT 24.245 2.465 24.535 2.695 ;
      RECT 22.835 2.465 23.38 2.695 ;
      RECT 22.835 2.55 23.785 2.69 ;
      RECT 23.645 2.37 23.785 2.69 ;
      RECT 24.145 2.465 24.535 2.65 ;
      RECT 23.645 2.37 24.285 2.51 ;
      RECT 22.355 3.26 22.675 3.675 ;
      RECT 22.435 1.905 22.59 3.675 ;
      RECT 22.37 1.905 22.66 2.135 ;
      RECT 20.75 7.77 21.04 8 ;
      RECT 20.81 6.29 20.98 8 ;
      RECT 20.805 6.655 21.155 7.005 ;
      RECT 20.75 6.29 21.04 6.52 ;
      RECT 20.345 2.395 20.45 2.965 ;
      RECT 20.345 2.73 20.67 2.96 ;
      RECT 20.345 2.76 20.84 2.93 ;
      RECT 20.345 2.395 20.535 2.96 ;
      RECT 19.76 2.36 20.05 2.59 ;
      RECT 19.76 2.395 20.535 2.565 ;
      RECT 19.82 0.88 19.99 2.59 ;
      RECT 19.76 0.88 20.05 1.11 ;
      RECT 19.76 7.77 20.05 8 ;
      RECT 19.82 6.29 19.99 8 ;
      RECT 19.76 6.29 20.05 6.52 ;
      RECT 19.76 6.325 20.615 6.485 ;
      RECT 20.445 5.92 20.615 6.485 ;
      RECT 19.76 6.32 20.155 6.485 ;
      RECT 20.38 5.92 20.67 6.15 ;
      RECT 20.38 5.95 20.84 6.12 ;
      RECT 19.39 2.73 19.68 2.96 ;
      RECT 19.39 2.76 19.85 2.93 ;
      RECT 19.455 1.655 19.62 2.96 ;
      RECT 17.97 1.625 18.26 1.855 ;
      RECT 17.97 1.655 19.62 1.825 ;
      RECT 18.03 0.885 18.2 1.855 ;
      RECT 17.97 0.885 18.26 1.115 ;
      RECT 17.97 7.765 18.26 7.995 ;
      RECT 18.03 7.025 18.2 7.995 ;
      RECT 18.03 7.12 19.62 7.29 ;
      RECT 19.45 5.92 19.62 7.29 ;
      RECT 17.97 7.025 18.26 7.255 ;
      RECT 19.39 5.92 19.68 6.15 ;
      RECT 19.39 5.95 19.85 6.12 ;
      RECT 16.02 3.15 16.36 3.5 ;
      RECT 16.11 2.025 16.28 3.5 ;
      RECT 18.4 1.965 18.75 2.315 ;
      RECT 16.11 2.025 18.75 2.195 ;
      RECT 18.425 6.655 18.75 6.98 ;
      RECT 12.99 6.605 13.34 6.955 ;
      RECT 18.4 6.655 18.75 6.885 ;
      RECT 12.785 6.655 13.34 6.885 ;
      RECT 12.615 6.685 18.75 6.855 ;
      RECT 17.625 2.365 17.945 2.685 ;
      RECT 17.595 2.365 17.945 2.595 ;
      RECT 17.425 2.395 17.945 2.565 ;
      RECT 17.625 6.255 17.945 6.545 ;
      RECT 17.595 6.285 17.945 6.515 ;
      RECT 17.425 6.315 17.945 6.485 ;
      RECT 13.075 3.57 13.395 3.83 ;
      RECT 14.365 2.745 14.505 3.605 ;
      RECT 13.165 3.465 14.505 3.605 ;
      RECT 13.165 3.025 13.305 3.83 ;
      RECT 13.09 3.025 13.38 3.255 ;
      RECT 14.29 2.745 14.58 2.975 ;
      RECT 13.81 3.025 14.1 3.255 ;
      RECT 14.005 1.95 14.145 3.21 ;
      RECT 14.035 1.89 14.355 2.15 ;
      RECT 10.635 2.45 10.955 2.71 ;
      RECT 13.33 2.465 13.62 2.695 ;
      RECT 10.725 2.37 13.545 2.51 ;
      RECT 12.595 1.89 12.915 2.15 ;
      RECT 13.09 1.905 13.38 2.135 ;
      RECT 12.595 1.95 13.38 2.09 ;
      RECT 12.595 3.01 12.915 3.27 ;
      RECT 12.595 2.79 12.825 3.27 ;
      RECT 12.09 2.745 12.38 2.975 ;
      RECT 12.09 2.79 12.825 2.93 ;
      RECT 11.115 3.57 11.435 3.83 ;
      RECT 10.65 3.585 10.94 3.815 ;
      RECT 10.65 3.63 11.435 3.77 ;
      RECT 9.41 2.465 9.7 2.695 ;
      RECT 9.41 2.51 10.345 2.65 ;
      RECT 10.205 1.95 10.345 2.65 ;
      RECT 10.875 1.89 11.195 2.15 ;
      RECT 10.65 1.905 11.195 2.135 ;
      RECT 10.205 1.95 11.195 2.09 ;
      RECT 8.555 3.57 8.875 3.83 ;
      RECT 8.555 3.63 9.625 3.77 ;
      RECT 9.485 3.07 9.625 3.77 ;
      RECT 10.65 3.025 10.94 3.255 ;
      RECT 9.485 3.07 10.94 3.21 ;
      RECT 8.915 1.89 9.235 2.15 ;
      RECT 8.69 1.905 9.235 2.135 ;
      RECT 7.21 3.025 7.5 3.255 ;
      RECT 7.405 1.95 7.545 3.21 ;
      RECT 8.195 1.89 8.515 2.15 ;
      RECT 7.21 1.905 7.5 2.135 ;
      RECT 7.21 1.95 8.515 2.09 ;
      RECT 6.805 3.465 7.905 3.605 ;
      RECT 7.69 3.305 7.98 3.535 ;
      RECT 6.73 3.305 7.02 3.535 ;
      RECT 6.715 1.89 7.035 2.15 ;
      RECT 4.755 1.89 5.075 2.15 ;
      RECT 4.755 1.95 7.035 2.09 ;
      RECT 3.795 3.26 4.115 3.675 ;
      RECT 3.875 1.905 4.03 3.675 ;
      RECT 3.81 1.905 4.1 2.135 ;
      RECT 1.54 7.765 1.83 7.995 ;
      RECT 1.6 7.025 1.77 7.995 ;
      RECT 1.51 7.025 1.86 7.315 ;
      RECT 1.135 6.285 1.485 6.575 ;
      RECT 0.995 6.315 1.485 6.485 ;
      RECT 86.315 3.57 86.635 3.83 ;
      RECT 85.715 1.89 86.395 2.15 ;
      RECT 85.835 3.57 86.155 3.83 ;
      RECT 84.355 3.57 84.675 3.83 ;
      RECT 83.875 1.89 84.195 2.15 ;
      RECT 83.155 3.01 83.475 3.27 ;
      RECT 82.435 3.01 82.755 3.27 ;
      RECT 78.995 3.01 79.315 3.27 ;
      RECT 67.755 3.57 68.075 3.83 ;
      RECT 67.155 1.89 67.835 2.15 ;
      RECT 67.275 3.57 67.595 3.83 ;
      RECT 65.795 3.57 66.115 3.83 ;
      RECT 65.315 1.89 65.635 2.15 ;
      RECT 64.595 3.01 64.915 3.27 ;
      RECT 63.875 3.01 64.195 3.27 ;
      RECT 60.435 3.01 60.755 3.27 ;
      RECT 49.195 3.57 49.515 3.83 ;
      RECT 48.595 1.89 49.275 2.15 ;
      RECT 48.715 3.57 49.035 3.83 ;
      RECT 47.235 3.57 47.555 3.83 ;
      RECT 46.755 1.89 47.075 2.15 ;
      RECT 46.035 3.01 46.355 3.27 ;
      RECT 45.315 3.01 45.635 3.27 ;
      RECT 41.875 3.01 42.195 3.27 ;
      RECT 30.635 3.57 30.955 3.83 ;
      RECT 30.035 1.89 30.715 2.15 ;
      RECT 30.155 3.57 30.475 3.83 ;
      RECT 28.675 3.57 28.995 3.83 ;
      RECT 28.195 1.89 28.515 2.15 ;
      RECT 27.475 3.01 27.795 3.27 ;
      RECT 26.755 3.01 27.075 3.27 ;
      RECT 23.315 3.01 23.635 3.27 ;
      RECT 12.075 3.57 12.395 3.83 ;
      RECT 11.475 1.89 12.155 2.15 ;
      RECT 11.595 3.57 11.915 3.83 ;
      RECT 10.115 3.57 10.435 3.83 ;
      RECT 9.635 1.89 9.955 2.15 ;
      RECT 8.915 3.01 9.235 3.27 ;
      RECT 4.755 3.01 5.075 3.27 ;
    LAYER mcon ;
      RECT 95.05 6.32 95.22 6.49 ;
      RECT 95.055 6.315 95.225 6.485 ;
      RECT 76.49 6.32 76.66 6.49 ;
      RECT 76.495 6.315 76.665 6.485 ;
      RECT 57.93 6.32 58.1 6.49 ;
      RECT 57.935 6.315 58.105 6.485 ;
      RECT 39.37 6.32 39.54 6.49 ;
      RECT 39.375 6.315 39.545 6.485 ;
      RECT 20.81 6.32 20.98 6.49 ;
      RECT 20.815 6.315 20.985 6.485 ;
      RECT 95.05 7.8 95.22 7.97 ;
      RECT 94.68 2.76 94.85 2.93 ;
      RECT 94.68 5.95 94.85 6.12 ;
      RECT 94.06 0.91 94.23 1.08 ;
      RECT 94.06 2.39 94.23 2.56 ;
      RECT 94.06 6.32 94.23 6.49 ;
      RECT 94.06 7.8 94.23 7.97 ;
      RECT 93.69 2.76 93.86 2.93 ;
      RECT 93.69 5.95 93.86 6.12 ;
      RECT 92.7 2.025 92.87 2.195 ;
      RECT 92.7 6.685 92.87 6.855 ;
      RECT 92.27 0.915 92.44 1.085 ;
      RECT 92.27 1.655 92.44 1.825 ;
      RECT 92.27 7.055 92.44 7.225 ;
      RECT 92.27 7.795 92.44 7.965 ;
      RECT 91.895 2.395 92.065 2.565 ;
      RECT 91.895 6.315 92.065 6.485 ;
      RECT 88.59 2.775 88.76 2.945 ;
      RECT 88.35 1.935 88.52 2.105 ;
      RECT 88.11 3.055 88.28 3.225 ;
      RECT 87.63 2.495 87.8 2.665 ;
      RECT 87.39 1.935 87.56 2.105 ;
      RECT 87.39 3.055 87.56 3.225 ;
      RECT 87.39 3.615 87.56 3.785 ;
      RECT 87.085 6.685 87.255 6.855 ;
      RECT 86.91 3.055 87.08 3.225 ;
      RECT 86.655 7.055 86.825 7.225 ;
      RECT 86.655 7.795 86.825 7.965 ;
      RECT 86.39 2.775 86.56 2.945 ;
      RECT 86.39 3.615 86.56 3.785 ;
      RECT 85.91 1.935 86.08 2.105 ;
      RECT 85.91 3.615 86.08 3.785 ;
      RECT 84.95 1.935 85.12 2.105 ;
      RECT 84.95 2.495 85.12 2.665 ;
      RECT 84.95 3.055 85.12 3.225 ;
      RECT 84.95 3.615 85.12 3.785 ;
      RECT 84.43 3.615 84.6 3.785 ;
      RECT 83.95 1.935 84.12 2.105 ;
      RECT 83.71 2.495 83.88 2.665 ;
      RECT 83.23 2.495 83.4 2.665 ;
      RECT 83.23 3.055 83.4 3.225 ;
      RECT 82.99 1.935 83.16 2.105 ;
      RECT 82.51 3.055 82.68 3.225 ;
      RECT 81.99 2.495 82.16 2.665 ;
      RECT 81.99 3.335 82.16 3.505 ;
      RECT 81.51 1.935 81.68 2.105 ;
      RECT 81.51 3.055 81.68 3.225 ;
      RECT 81.03 3.335 81.2 3.505 ;
      RECT 80.79 2.775 80.96 2.945 ;
      RECT 79.985 2.495 80.155 2.665 ;
      RECT 79.07 1.935 79.24 2.105 ;
      RECT 79.07 3.055 79.24 3.225 ;
      RECT 78.83 2.495 79 2.665 ;
      RECT 78.11 1.935 78.28 2.105 ;
      RECT 78.11 3.475 78.28 3.645 ;
      RECT 76.49 7.8 76.66 7.97 ;
      RECT 76.12 2.76 76.29 2.93 ;
      RECT 76.12 5.95 76.29 6.12 ;
      RECT 75.5 0.91 75.67 1.08 ;
      RECT 75.5 2.39 75.67 2.56 ;
      RECT 75.5 6.32 75.67 6.49 ;
      RECT 75.5 7.8 75.67 7.97 ;
      RECT 75.13 2.76 75.3 2.93 ;
      RECT 75.13 5.95 75.3 6.12 ;
      RECT 74.14 2.025 74.31 2.195 ;
      RECT 74.14 6.685 74.31 6.855 ;
      RECT 73.71 0.915 73.88 1.085 ;
      RECT 73.71 1.655 73.88 1.825 ;
      RECT 73.71 7.055 73.88 7.225 ;
      RECT 73.71 7.795 73.88 7.965 ;
      RECT 73.335 2.395 73.505 2.565 ;
      RECT 73.335 6.315 73.505 6.485 ;
      RECT 70.03 2.775 70.2 2.945 ;
      RECT 69.79 1.935 69.96 2.105 ;
      RECT 69.55 3.055 69.72 3.225 ;
      RECT 69.07 2.495 69.24 2.665 ;
      RECT 68.83 1.935 69 2.105 ;
      RECT 68.83 3.055 69 3.225 ;
      RECT 68.83 3.615 69 3.785 ;
      RECT 68.525 6.685 68.695 6.855 ;
      RECT 68.35 3.055 68.52 3.225 ;
      RECT 68.095 7.055 68.265 7.225 ;
      RECT 68.095 7.795 68.265 7.965 ;
      RECT 67.83 2.775 68 2.945 ;
      RECT 67.83 3.615 68 3.785 ;
      RECT 67.35 1.935 67.52 2.105 ;
      RECT 67.35 3.615 67.52 3.785 ;
      RECT 66.39 1.935 66.56 2.105 ;
      RECT 66.39 2.495 66.56 2.665 ;
      RECT 66.39 3.055 66.56 3.225 ;
      RECT 66.39 3.615 66.56 3.785 ;
      RECT 65.87 3.615 66.04 3.785 ;
      RECT 65.39 1.935 65.56 2.105 ;
      RECT 65.15 2.495 65.32 2.665 ;
      RECT 64.67 2.495 64.84 2.665 ;
      RECT 64.67 3.055 64.84 3.225 ;
      RECT 64.43 1.935 64.6 2.105 ;
      RECT 63.95 3.055 64.12 3.225 ;
      RECT 63.43 2.495 63.6 2.665 ;
      RECT 63.43 3.335 63.6 3.505 ;
      RECT 62.95 1.935 63.12 2.105 ;
      RECT 62.95 3.055 63.12 3.225 ;
      RECT 62.47 3.335 62.64 3.505 ;
      RECT 62.23 2.775 62.4 2.945 ;
      RECT 61.425 2.495 61.595 2.665 ;
      RECT 60.51 1.935 60.68 2.105 ;
      RECT 60.51 3.055 60.68 3.225 ;
      RECT 60.27 2.495 60.44 2.665 ;
      RECT 59.55 1.935 59.72 2.105 ;
      RECT 59.55 3.475 59.72 3.645 ;
      RECT 57.93 7.8 58.1 7.97 ;
      RECT 57.56 2.76 57.73 2.93 ;
      RECT 57.56 5.95 57.73 6.12 ;
      RECT 56.94 0.91 57.11 1.08 ;
      RECT 56.94 2.39 57.11 2.56 ;
      RECT 56.94 6.32 57.11 6.49 ;
      RECT 56.94 7.8 57.11 7.97 ;
      RECT 56.57 2.76 56.74 2.93 ;
      RECT 56.57 5.95 56.74 6.12 ;
      RECT 55.58 2.025 55.75 2.195 ;
      RECT 55.58 6.685 55.75 6.855 ;
      RECT 55.15 0.915 55.32 1.085 ;
      RECT 55.15 1.655 55.32 1.825 ;
      RECT 55.15 7.055 55.32 7.225 ;
      RECT 55.15 7.795 55.32 7.965 ;
      RECT 54.775 2.395 54.945 2.565 ;
      RECT 54.775 6.315 54.945 6.485 ;
      RECT 51.47 2.775 51.64 2.945 ;
      RECT 51.23 1.935 51.4 2.105 ;
      RECT 50.99 3.055 51.16 3.225 ;
      RECT 50.51 2.495 50.68 2.665 ;
      RECT 50.27 1.935 50.44 2.105 ;
      RECT 50.27 3.055 50.44 3.225 ;
      RECT 50.27 3.615 50.44 3.785 ;
      RECT 49.965 6.685 50.135 6.855 ;
      RECT 49.79 3.055 49.96 3.225 ;
      RECT 49.535 7.055 49.705 7.225 ;
      RECT 49.535 7.795 49.705 7.965 ;
      RECT 49.27 2.775 49.44 2.945 ;
      RECT 49.27 3.615 49.44 3.785 ;
      RECT 48.79 1.935 48.96 2.105 ;
      RECT 48.79 3.615 48.96 3.785 ;
      RECT 47.83 1.935 48 2.105 ;
      RECT 47.83 2.495 48 2.665 ;
      RECT 47.83 3.055 48 3.225 ;
      RECT 47.83 3.615 48 3.785 ;
      RECT 47.31 3.615 47.48 3.785 ;
      RECT 46.83 1.935 47 2.105 ;
      RECT 46.59 2.495 46.76 2.665 ;
      RECT 46.11 2.495 46.28 2.665 ;
      RECT 46.11 3.055 46.28 3.225 ;
      RECT 45.87 1.935 46.04 2.105 ;
      RECT 45.39 3.055 45.56 3.225 ;
      RECT 44.87 2.495 45.04 2.665 ;
      RECT 44.87 3.335 45.04 3.505 ;
      RECT 44.39 1.935 44.56 2.105 ;
      RECT 44.39 3.055 44.56 3.225 ;
      RECT 43.91 3.335 44.08 3.505 ;
      RECT 43.67 2.775 43.84 2.945 ;
      RECT 42.865 2.495 43.035 2.665 ;
      RECT 41.95 1.935 42.12 2.105 ;
      RECT 41.95 3.055 42.12 3.225 ;
      RECT 41.71 2.495 41.88 2.665 ;
      RECT 40.99 1.935 41.16 2.105 ;
      RECT 40.99 3.475 41.16 3.645 ;
      RECT 39.37 7.8 39.54 7.97 ;
      RECT 39 2.76 39.17 2.93 ;
      RECT 39 5.95 39.17 6.12 ;
      RECT 38.38 0.91 38.55 1.08 ;
      RECT 38.38 2.39 38.55 2.56 ;
      RECT 38.38 6.32 38.55 6.49 ;
      RECT 38.38 7.8 38.55 7.97 ;
      RECT 38.01 2.76 38.18 2.93 ;
      RECT 38.01 5.95 38.18 6.12 ;
      RECT 37.02 2.025 37.19 2.195 ;
      RECT 37.02 6.685 37.19 6.855 ;
      RECT 36.59 0.915 36.76 1.085 ;
      RECT 36.59 1.655 36.76 1.825 ;
      RECT 36.59 7.055 36.76 7.225 ;
      RECT 36.59 7.795 36.76 7.965 ;
      RECT 36.215 2.395 36.385 2.565 ;
      RECT 36.215 6.315 36.385 6.485 ;
      RECT 32.91 2.775 33.08 2.945 ;
      RECT 32.67 1.935 32.84 2.105 ;
      RECT 32.43 3.055 32.6 3.225 ;
      RECT 31.95 2.495 32.12 2.665 ;
      RECT 31.71 1.935 31.88 2.105 ;
      RECT 31.71 3.055 31.88 3.225 ;
      RECT 31.71 3.615 31.88 3.785 ;
      RECT 31.405 6.685 31.575 6.855 ;
      RECT 31.23 3.055 31.4 3.225 ;
      RECT 30.975 7.055 31.145 7.225 ;
      RECT 30.975 7.795 31.145 7.965 ;
      RECT 30.71 2.775 30.88 2.945 ;
      RECT 30.71 3.615 30.88 3.785 ;
      RECT 30.23 1.935 30.4 2.105 ;
      RECT 30.23 3.615 30.4 3.785 ;
      RECT 29.27 1.935 29.44 2.105 ;
      RECT 29.27 2.495 29.44 2.665 ;
      RECT 29.27 3.055 29.44 3.225 ;
      RECT 29.27 3.615 29.44 3.785 ;
      RECT 28.75 3.615 28.92 3.785 ;
      RECT 28.27 1.935 28.44 2.105 ;
      RECT 28.03 2.495 28.2 2.665 ;
      RECT 27.55 2.495 27.72 2.665 ;
      RECT 27.55 3.055 27.72 3.225 ;
      RECT 27.31 1.935 27.48 2.105 ;
      RECT 26.83 3.055 27 3.225 ;
      RECT 26.31 2.495 26.48 2.665 ;
      RECT 26.31 3.335 26.48 3.505 ;
      RECT 25.83 1.935 26 2.105 ;
      RECT 25.83 3.055 26 3.225 ;
      RECT 25.35 3.335 25.52 3.505 ;
      RECT 25.11 2.775 25.28 2.945 ;
      RECT 24.305 2.495 24.475 2.665 ;
      RECT 23.39 1.935 23.56 2.105 ;
      RECT 23.39 3.055 23.56 3.225 ;
      RECT 23.15 2.495 23.32 2.665 ;
      RECT 22.43 1.935 22.6 2.105 ;
      RECT 22.43 3.475 22.6 3.645 ;
      RECT 20.81 7.8 20.98 7.97 ;
      RECT 20.44 2.76 20.61 2.93 ;
      RECT 20.44 5.95 20.61 6.12 ;
      RECT 19.82 0.91 19.99 1.08 ;
      RECT 19.82 2.39 19.99 2.56 ;
      RECT 19.82 6.32 19.99 6.49 ;
      RECT 19.82 7.8 19.99 7.97 ;
      RECT 19.45 2.76 19.62 2.93 ;
      RECT 19.45 5.95 19.62 6.12 ;
      RECT 18.46 2.025 18.63 2.195 ;
      RECT 18.46 6.685 18.63 6.855 ;
      RECT 18.03 0.915 18.2 1.085 ;
      RECT 18.03 1.655 18.2 1.825 ;
      RECT 18.03 7.055 18.2 7.225 ;
      RECT 18.03 7.795 18.2 7.965 ;
      RECT 17.655 2.395 17.825 2.565 ;
      RECT 17.655 6.315 17.825 6.485 ;
      RECT 14.35 2.775 14.52 2.945 ;
      RECT 14.11 1.935 14.28 2.105 ;
      RECT 13.87 3.055 14.04 3.225 ;
      RECT 13.39 2.495 13.56 2.665 ;
      RECT 13.15 1.935 13.32 2.105 ;
      RECT 13.15 3.055 13.32 3.225 ;
      RECT 13.15 3.615 13.32 3.785 ;
      RECT 12.845 6.685 13.015 6.855 ;
      RECT 12.67 3.055 12.84 3.225 ;
      RECT 12.15 2.775 12.32 2.945 ;
      RECT 12.15 3.615 12.32 3.785 ;
      RECT 11.67 1.935 11.84 2.105 ;
      RECT 11.67 3.615 11.84 3.785 ;
      RECT 10.71 1.935 10.88 2.105 ;
      RECT 10.71 2.495 10.88 2.665 ;
      RECT 10.71 3.055 10.88 3.225 ;
      RECT 10.71 3.615 10.88 3.785 ;
      RECT 10.19 3.615 10.36 3.785 ;
      RECT 9.71 1.935 9.88 2.105 ;
      RECT 9.47 2.495 9.64 2.665 ;
      RECT 8.99 3.055 9.16 3.225 ;
      RECT 8.75 1.935 8.92 2.105 ;
      RECT 7.75 3.335 7.92 3.505 ;
      RECT 7.27 1.935 7.44 2.105 ;
      RECT 7.27 3.055 7.44 3.225 ;
      RECT 6.79 3.335 6.96 3.505 ;
      RECT 4.83 1.935 5 2.105 ;
      RECT 4.83 3.055 5 3.225 ;
      RECT 3.87 1.935 4.04 2.105 ;
      RECT 3.87 3.475 4.04 3.645 ;
      RECT 1.6 7.055 1.77 7.225 ;
      RECT 1.6 7.795 1.77 7.965 ;
      RECT 1.225 6.315 1.395 6.485 ;
    LAYER li1 ;
      RECT 95.05 5.02 95.22 6.49 ;
      RECT 95.05 6.315 95.225 6.485 ;
      RECT 94.68 1.74 94.85 2.93 ;
      RECT 94.68 1.74 95.15 1.91 ;
      RECT 94.68 6.97 95.15 7.14 ;
      RECT 94.68 5.95 94.85 7.14 ;
      RECT 93.69 1.74 93.86 2.93 ;
      RECT 93.69 1.74 94.16 1.91 ;
      RECT 93.69 6.97 94.16 7.14 ;
      RECT 93.69 5.95 93.86 7.14 ;
      RECT 91.84 2.635 92.01 3.865 ;
      RECT 91.895 0.855 92.065 2.805 ;
      RECT 91.84 0.575 92.01 1.025 ;
      RECT 91.84 7.855 92.01 8.305 ;
      RECT 91.895 6.075 92.065 8.025 ;
      RECT 91.84 5.015 92.01 6.245 ;
      RECT 91.32 0.575 91.49 3.865 ;
      RECT 91.32 2.075 91.725 2.405 ;
      RECT 91.32 1.235 91.725 1.565 ;
      RECT 91.32 5.015 91.49 8.305 ;
      RECT 91.32 7.315 91.725 7.645 ;
      RECT 91.32 6.475 91.725 6.805 ;
      RECT 88.11 3.225 89.08 3.395 ;
      RECT 88.11 3.055 88.28 3.395 ;
      RECT 87.63 2.495 87.8 2.825 ;
      RECT 87.63 2.575 88.36 2.745 ;
      RECT 87.27 3.615 87.56 3.785 ;
      RECT 87.27 2.575 87.44 3.785 ;
      RECT 87.27 3.055 87.56 3.225 ;
      RECT 87.07 2.575 87.44 2.745 ;
      RECT 86.39 2.675 86.56 2.945 ;
      RECT 86.15 2.675 86.56 2.845 ;
      RECT 86.07 2.575 86.4 2.745 ;
      RECT 85.91 3.615 86.56 3.785 ;
      RECT 86.39 3.145 86.56 3.785 ;
      RECT 86.27 3.225 86.56 3.785 ;
      RECT 85.705 5.015 85.875 8.305 ;
      RECT 85.705 7.315 86.11 7.645 ;
      RECT 85.705 6.475 86.11 6.805 ;
      RECT 84.95 2.915 85.12 3.225 ;
      RECT 84.95 2.915 85.84 3.085 ;
      RECT 85.67 2.495 85.84 3.085 ;
      RECT 84.95 2.575 85.44 2.745 ;
      RECT 84.95 2.495 85.12 2.745 ;
      RECT 82.91 3.225 83.4 3.395 ;
      RECT 84.07 2.575 84.24 3.225 ;
      RECT 83.23 3.055 84.24 3.225 ;
      RECT 84.19 2.495 84.36 2.825 ;
      RECT 82.99 1.835 83.16 2.105 ;
      RECT 82.43 1.835 83.16 2.005 ;
      RECT 82.51 2.575 82.68 3.225 ;
      RECT 82.51 2.575 83 2.745 ;
      RECT 81.67 2.575 82.16 2.745 ;
      RECT 81.99 2.495 82.16 2.745 ;
      RECT 81.51 1.835 81.68 2.105 ;
      RECT 80.95 1.835 81.68 2.005 ;
      RECT 81.03 3.225 81.2 3.505 ;
      RECT 79.99 3.225 81.28 3.395 ;
      RECT 79.985 2.575 80.56 2.745 ;
      RECT 79.985 2.495 80.155 2.745 ;
      RECT 79.07 1.835 79.24 2.105 ;
      RECT 79.07 1.835 79.8 2.005 ;
      RECT 79.07 3.055 79.24 3.475 ;
      RECT 78.45 3.14 79.24 3.31 ;
      RECT 78.45 2.915 78.62 3.31 ;
      RECT 78.35 2.495 78.52 3.085 ;
      RECT 78.11 2.575 78.52 2.845 ;
      RECT 76.49 5.02 76.66 6.49 ;
      RECT 76.49 6.315 76.665 6.485 ;
      RECT 76.12 1.74 76.29 2.93 ;
      RECT 76.12 1.74 76.59 1.91 ;
      RECT 76.12 6.97 76.59 7.14 ;
      RECT 76.12 5.95 76.29 7.14 ;
      RECT 75.13 1.74 75.3 2.93 ;
      RECT 75.13 1.74 75.6 1.91 ;
      RECT 75.13 6.97 75.6 7.14 ;
      RECT 75.13 5.95 75.3 7.14 ;
      RECT 73.28 2.635 73.45 3.865 ;
      RECT 73.335 0.855 73.505 2.805 ;
      RECT 73.28 0.575 73.45 1.025 ;
      RECT 73.28 7.855 73.45 8.305 ;
      RECT 73.335 6.075 73.505 8.025 ;
      RECT 73.28 5.015 73.45 6.245 ;
      RECT 72.76 0.575 72.93 3.865 ;
      RECT 72.76 2.075 73.165 2.405 ;
      RECT 72.76 1.235 73.165 1.565 ;
      RECT 72.76 5.015 72.93 8.305 ;
      RECT 72.76 7.315 73.165 7.645 ;
      RECT 72.76 6.475 73.165 6.805 ;
      RECT 69.55 3.225 70.52 3.395 ;
      RECT 69.55 3.055 69.72 3.395 ;
      RECT 69.07 2.495 69.24 2.825 ;
      RECT 69.07 2.575 69.8 2.745 ;
      RECT 68.71 3.615 69 3.785 ;
      RECT 68.71 2.575 68.88 3.785 ;
      RECT 68.71 3.055 69 3.225 ;
      RECT 68.51 2.575 68.88 2.745 ;
      RECT 67.83 2.675 68 2.945 ;
      RECT 67.59 2.675 68 2.845 ;
      RECT 67.51 2.575 67.84 2.745 ;
      RECT 67.35 3.615 68 3.785 ;
      RECT 67.83 3.145 68 3.785 ;
      RECT 67.71 3.225 68 3.785 ;
      RECT 67.145 5.015 67.315 8.305 ;
      RECT 67.145 7.315 67.55 7.645 ;
      RECT 67.145 6.475 67.55 6.805 ;
      RECT 66.39 2.915 66.56 3.225 ;
      RECT 66.39 2.915 67.28 3.085 ;
      RECT 67.11 2.495 67.28 3.085 ;
      RECT 66.39 2.575 66.88 2.745 ;
      RECT 66.39 2.495 66.56 2.745 ;
      RECT 64.35 3.225 64.84 3.395 ;
      RECT 65.51 2.575 65.68 3.225 ;
      RECT 64.67 3.055 65.68 3.225 ;
      RECT 65.63 2.495 65.8 2.825 ;
      RECT 64.43 1.835 64.6 2.105 ;
      RECT 63.87 1.835 64.6 2.005 ;
      RECT 63.95 2.575 64.12 3.225 ;
      RECT 63.95 2.575 64.44 2.745 ;
      RECT 63.11 2.575 63.6 2.745 ;
      RECT 63.43 2.495 63.6 2.745 ;
      RECT 62.95 1.835 63.12 2.105 ;
      RECT 62.39 1.835 63.12 2.005 ;
      RECT 62.47 3.225 62.64 3.505 ;
      RECT 61.43 3.225 62.72 3.395 ;
      RECT 61.425 2.575 62 2.745 ;
      RECT 61.425 2.495 61.595 2.745 ;
      RECT 60.51 1.835 60.68 2.105 ;
      RECT 60.51 1.835 61.24 2.005 ;
      RECT 60.51 3.055 60.68 3.475 ;
      RECT 59.89 3.14 60.68 3.31 ;
      RECT 59.89 2.915 60.06 3.31 ;
      RECT 59.79 2.495 59.96 3.085 ;
      RECT 59.55 2.575 59.96 2.845 ;
      RECT 57.93 5.02 58.1 6.49 ;
      RECT 57.93 6.315 58.105 6.485 ;
      RECT 57.56 1.74 57.73 2.93 ;
      RECT 57.56 1.74 58.03 1.91 ;
      RECT 57.56 6.97 58.03 7.14 ;
      RECT 57.56 5.95 57.73 7.14 ;
      RECT 56.57 1.74 56.74 2.93 ;
      RECT 56.57 1.74 57.04 1.91 ;
      RECT 56.57 6.97 57.04 7.14 ;
      RECT 56.57 5.95 56.74 7.14 ;
      RECT 54.72 2.635 54.89 3.865 ;
      RECT 54.775 0.855 54.945 2.805 ;
      RECT 54.72 0.575 54.89 1.025 ;
      RECT 54.72 7.855 54.89 8.305 ;
      RECT 54.775 6.075 54.945 8.025 ;
      RECT 54.72 5.015 54.89 6.245 ;
      RECT 54.2 0.575 54.37 3.865 ;
      RECT 54.2 2.075 54.605 2.405 ;
      RECT 54.2 1.235 54.605 1.565 ;
      RECT 54.2 5.015 54.37 8.305 ;
      RECT 54.2 7.315 54.605 7.645 ;
      RECT 54.2 6.475 54.605 6.805 ;
      RECT 50.99 3.225 51.96 3.395 ;
      RECT 50.99 3.055 51.16 3.395 ;
      RECT 50.51 2.495 50.68 2.825 ;
      RECT 50.51 2.575 51.24 2.745 ;
      RECT 50.15 3.615 50.44 3.785 ;
      RECT 50.15 2.575 50.32 3.785 ;
      RECT 50.15 3.055 50.44 3.225 ;
      RECT 49.95 2.575 50.32 2.745 ;
      RECT 49.27 2.675 49.44 2.945 ;
      RECT 49.03 2.675 49.44 2.845 ;
      RECT 48.95 2.575 49.28 2.745 ;
      RECT 48.79 3.615 49.44 3.785 ;
      RECT 49.27 3.145 49.44 3.785 ;
      RECT 49.15 3.225 49.44 3.785 ;
      RECT 48.585 5.015 48.755 8.305 ;
      RECT 48.585 7.315 48.99 7.645 ;
      RECT 48.585 6.475 48.99 6.805 ;
      RECT 47.83 2.915 48 3.225 ;
      RECT 47.83 2.915 48.72 3.085 ;
      RECT 48.55 2.495 48.72 3.085 ;
      RECT 47.83 2.575 48.32 2.745 ;
      RECT 47.83 2.495 48 2.745 ;
      RECT 45.79 3.225 46.28 3.395 ;
      RECT 46.95 2.575 47.12 3.225 ;
      RECT 46.11 3.055 47.12 3.225 ;
      RECT 47.07 2.495 47.24 2.825 ;
      RECT 45.87 1.835 46.04 2.105 ;
      RECT 45.31 1.835 46.04 2.005 ;
      RECT 45.39 2.575 45.56 3.225 ;
      RECT 45.39 2.575 45.88 2.745 ;
      RECT 44.55 2.575 45.04 2.745 ;
      RECT 44.87 2.495 45.04 2.745 ;
      RECT 44.39 1.835 44.56 2.105 ;
      RECT 43.83 1.835 44.56 2.005 ;
      RECT 43.91 3.225 44.08 3.505 ;
      RECT 42.87 3.225 44.16 3.395 ;
      RECT 42.865 2.575 43.44 2.745 ;
      RECT 42.865 2.495 43.035 2.745 ;
      RECT 41.95 1.835 42.12 2.105 ;
      RECT 41.95 1.835 42.68 2.005 ;
      RECT 41.95 3.055 42.12 3.475 ;
      RECT 41.33 3.14 42.12 3.31 ;
      RECT 41.33 2.915 41.5 3.31 ;
      RECT 41.23 2.495 41.4 3.085 ;
      RECT 40.99 2.575 41.4 2.845 ;
      RECT 39.37 5.02 39.54 6.49 ;
      RECT 39.37 6.315 39.545 6.485 ;
      RECT 39 1.74 39.17 2.93 ;
      RECT 39 1.74 39.47 1.91 ;
      RECT 39 6.97 39.47 7.14 ;
      RECT 39 5.95 39.17 7.14 ;
      RECT 38.01 1.74 38.18 2.93 ;
      RECT 38.01 1.74 38.48 1.91 ;
      RECT 38.01 6.97 38.48 7.14 ;
      RECT 38.01 5.95 38.18 7.14 ;
      RECT 36.16 2.635 36.33 3.865 ;
      RECT 36.215 0.855 36.385 2.805 ;
      RECT 36.16 0.575 36.33 1.025 ;
      RECT 36.16 7.855 36.33 8.305 ;
      RECT 36.215 6.075 36.385 8.025 ;
      RECT 36.16 5.015 36.33 6.245 ;
      RECT 35.64 0.575 35.81 3.865 ;
      RECT 35.64 2.075 36.045 2.405 ;
      RECT 35.64 1.235 36.045 1.565 ;
      RECT 35.64 5.015 35.81 8.305 ;
      RECT 35.64 7.315 36.045 7.645 ;
      RECT 35.64 6.475 36.045 6.805 ;
      RECT 32.43 3.225 33.4 3.395 ;
      RECT 32.43 3.055 32.6 3.395 ;
      RECT 31.95 2.495 32.12 2.825 ;
      RECT 31.95 2.575 32.68 2.745 ;
      RECT 31.59 3.615 31.88 3.785 ;
      RECT 31.59 2.575 31.76 3.785 ;
      RECT 31.59 3.055 31.88 3.225 ;
      RECT 31.39 2.575 31.76 2.745 ;
      RECT 30.71 2.675 30.88 2.945 ;
      RECT 30.47 2.675 30.88 2.845 ;
      RECT 30.39 2.575 30.72 2.745 ;
      RECT 30.23 3.615 30.88 3.785 ;
      RECT 30.71 3.145 30.88 3.785 ;
      RECT 30.59 3.225 30.88 3.785 ;
      RECT 30.025 5.015 30.195 8.305 ;
      RECT 30.025 7.315 30.43 7.645 ;
      RECT 30.025 6.475 30.43 6.805 ;
      RECT 29.27 2.915 29.44 3.225 ;
      RECT 29.27 2.915 30.16 3.085 ;
      RECT 29.99 2.495 30.16 3.085 ;
      RECT 29.27 2.575 29.76 2.745 ;
      RECT 29.27 2.495 29.44 2.745 ;
      RECT 27.23 3.225 27.72 3.395 ;
      RECT 28.39 2.575 28.56 3.225 ;
      RECT 27.55 3.055 28.56 3.225 ;
      RECT 28.51 2.495 28.68 2.825 ;
      RECT 27.31 1.835 27.48 2.105 ;
      RECT 26.75 1.835 27.48 2.005 ;
      RECT 26.83 2.575 27 3.225 ;
      RECT 26.83 2.575 27.32 2.745 ;
      RECT 25.99 2.575 26.48 2.745 ;
      RECT 26.31 2.495 26.48 2.745 ;
      RECT 25.83 1.835 26 2.105 ;
      RECT 25.27 1.835 26 2.005 ;
      RECT 25.35 3.225 25.52 3.505 ;
      RECT 24.31 3.225 25.6 3.395 ;
      RECT 24.305 2.575 24.88 2.745 ;
      RECT 24.305 2.495 24.475 2.745 ;
      RECT 23.39 1.835 23.56 2.105 ;
      RECT 23.39 1.835 24.12 2.005 ;
      RECT 23.39 3.055 23.56 3.475 ;
      RECT 22.77 3.14 23.56 3.31 ;
      RECT 22.77 2.915 22.94 3.31 ;
      RECT 22.67 2.495 22.84 3.085 ;
      RECT 22.43 2.575 22.84 2.845 ;
      RECT 20.81 5.02 20.98 6.49 ;
      RECT 20.81 6.315 20.985 6.485 ;
      RECT 20.44 1.74 20.61 2.93 ;
      RECT 20.44 1.74 20.91 1.91 ;
      RECT 20.44 6.97 20.91 7.14 ;
      RECT 20.44 5.95 20.61 7.14 ;
      RECT 19.45 1.74 19.62 2.93 ;
      RECT 19.45 1.74 19.92 1.91 ;
      RECT 19.45 6.97 19.92 7.14 ;
      RECT 19.45 5.95 19.62 7.14 ;
      RECT 17.6 2.635 17.77 3.865 ;
      RECT 17.655 0.855 17.825 2.805 ;
      RECT 17.6 0.575 17.77 1.025 ;
      RECT 17.6 7.855 17.77 8.305 ;
      RECT 17.655 6.075 17.825 8.025 ;
      RECT 17.6 5.015 17.77 6.245 ;
      RECT 17.08 0.575 17.25 3.865 ;
      RECT 17.08 2.075 17.485 2.405 ;
      RECT 17.08 1.235 17.485 1.565 ;
      RECT 17.08 5.015 17.25 8.305 ;
      RECT 17.08 7.315 17.485 7.645 ;
      RECT 17.08 6.475 17.485 6.805 ;
      RECT 13.87 3.225 14.84 3.395 ;
      RECT 13.87 3.055 14.04 3.395 ;
      RECT 13.39 2.495 13.56 2.825 ;
      RECT 13.39 2.575 14.12 2.745 ;
      RECT 13.03 3.615 13.32 3.785 ;
      RECT 13.03 2.575 13.2 3.785 ;
      RECT 13.03 3.055 13.32 3.225 ;
      RECT 12.83 2.575 13.2 2.745 ;
      RECT 12.15 2.675 12.32 2.945 ;
      RECT 11.91 2.675 12.32 2.845 ;
      RECT 11.83 2.575 12.16 2.745 ;
      RECT 11.67 3.615 12.32 3.785 ;
      RECT 12.15 3.145 12.32 3.785 ;
      RECT 12.03 3.225 12.32 3.785 ;
      RECT 11.465 5.015 11.635 8.305 ;
      RECT 11.465 7.315 11.87 7.645 ;
      RECT 11.465 6.475 11.87 6.805 ;
      RECT 10.71 2.915 10.88 3.225 ;
      RECT 10.71 2.915 11.6 3.085 ;
      RECT 11.43 2.495 11.6 3.085 ;
      RECT 10.71 2.575 11.2 2.745 ;
      RECT 10.71 2.495 10.88 2.745 ;
      RECT 8.67 3.225 9.16 3.395 ;
      RECT 9.83 2.575 10 3.225 ;
      RECT 8.99 3.055 10 3.225 ;
      RECT 9.95 2.495 10.12 2.825 ;
      RECT 8.75 1.835 8.92 2.105 ;
      RECT 8.19 1.835 8.92 2.005 ;
      RECT 7.27 1.835 7.44 2.105 ;
      RECT 6.71 1.835 7.44 2.005 ;
      RECT 6.79 3.225 6.96 3.505 ;
      RECT 5.75 3.225 7.04 3.395 ;
      RECT 4.83 1.835 5 2.105 ;
      RECT 4.83 1.835 5.56 2.005 ;
      RECT 4.83 3.055 5 3.475 ;
      RECT 4.21 3.14 5 3.31 ;
      RECT 4.21 2.915 4.38 3.31 ;
      RECT 4.11 2.495 4.28 3.085 ;
      RECT 3.87 2.575 4.28 2.845 ;
      RECT 1.17 7.855 1.34 8.305 ;
      RECT 1.225 6.075 1.395 8.025 ;
      RECT 1.17 5.015 1.34 6.245 ;
      RECT 0.65 5.015 0.82 8.305 ;
      RECT 0.65 7.315 1.055 7.645 ;
      RECT 0.65 6.475 1.055 6.805 ;
      RECT 95.05 7.8 95.22 8.31 ;
      RECT 94.06 0.57 94.23 1.08 ;
      RECT 94.06 2.39 94.23 3.86 ;
      RECT 94.06 5.02 94.23 6.49 ;
      RECT 94.06 7.8 94.23 8.31 ;
      RECT 92.7 0.575 92.87 3.865 ;
      RECT 92.7 5.015 92.87 8.305 ;
      RECT 92.27 0.575 92.44 1.085 ;
      RECT 92.27 1.655 92.44 3.865 ;
      RECT 92.27 5.015 92.44 7.225 ;
      RECT 92.27 7.795 92.44 8.305 ;
      RECT 88.59 2.495 88.76 2.945 ;
      RECT 88.35 1.755 88.52 2.105 ;
      RECT 87.39 1.755 87.56 2.105 ;
      RECT 87.085 5.015 87.255 8.305 ;
      RECT 86.91 3.055 87.08 3.475 ;
      RECT 86.655 5.015 86.825 7.225 ;
      RECT 86.655 7.795 86.825 8.305 ;
      RECT 85.91 1.755 86.08 2.105 ;
      RECT 84.95 1.755 85.12 2.105 ;
      RECT 84.95 3.485 85.12 3.815 ;
      RECT 84.43 3.145 84.6 3.785 ;
      RECT 83.95 1.755 84.12 2.105 ;
      RECT 83.71 2.495 83.88 2.825 ;
      RECT 83.23 2.495 83.4 2.825 ;
      RECT 81.99 3.145 82.16 3.505 ;
      RECT 81.51 3.055 81.68 3.475 ;
      RECT 80.79 2.495 80.96 2.945 ;
      RECT 78.83 2.495 79 2.825 ;
      RECT 78.11 1.755 78.28 2.105 ;
      RECT 78.11 3.285 78.28 3.645 ;
      RECT 76.49 7.8 76.66 8.31 ;
      RECT 75.5 0.57 75.67 1.08 ;
      RECT 75.5 2.39 75.67 3.86 ;
      RECT 75.5 5.02 75.67 6.49 ;
      RECT 75.5 7.8 75.67 8.31 ;
      RECT 74.14 0.575 74.31 3.865 ;
      RECT 74.14 5.015 74.31 8.305 ;
      RECT 73.71 0.575 73.88 1.085 ;
      RECT 73.71 1.655 73.88 3.865 ;
      RECT 73.71 5.015 73.88 7.225 ;
      RECT 73.71 7.795 73.88 8.305 ;
      RECT 70.03 2.495 70.2 2.945 ;
      RECT 69.79 1.755 69.96 2.105 ;
      RECT 68.83 1.755 69 2.105 ;
      RECT 68.525 5.015 68.695 8.305 ;
      RECT 68.35 3.055 68.52 3.475 ;
      RECT 68.095 5.015 68.265 7.225 ;
      RECT 68.095 7.795 68.265 8.305 ;
      RECT 67.35 1.755 67.52 2.105 ;
      RECT 66.39 1.755 66.56 2.105 ;
      RECT 66.39 3.485 66.56 3.815 ;
      RECT 65.87 3.145 66.04 3.785 ;
      RECT 65.39 1.755 65.56 2.105 ;
      RECT 65.15 2.495 65.32 2.825 ;
      RECT 64.67 2.495 64.84 2.825 ;
      RECT 63.43 3.145 63.6 3.505 ;
      RECT 62.95 3.055 63.12 3.475 ;
      RECT 62.23 2.495 62.4 2.945 ;
      RECT 60.27 2.495 60.44 2.825 ;
      RECT 59.55 1.755 59.72 2.105 ;
      RECT 59.55 3.285 59.72 3.645 ;
      RECT 57.93 7.8 58.1 8.31 ;
      RECT 56.94 0.57 57.11 1.08 ;
      RECT 56.94 2.39 57.11 3.86 ;
      RECT 56.94 5.02 57.11 6.49 ;
      RECT 56.94 7.8 57.11 8.31 ;
      RECT 55.58 0.575 55.75 3.865 ;
      RECT 55.58 5.015 55.75 8.305 ;
      RECT 55.15 0.575 55.32 1.085 ;
      RECT 55.15 1.655 55.32 3.865 ;
      RECT 55.15 5.015 55.32 7.225 ;
      RECT 55.15 7.795 55.32 8.305 ;
      RECT 51.47 2.495 51.64 2.945 ;
      RECT 51.23 1.755 51.4 2.105 ;
      RECT 50.27 1.755 50.44 2.105 ;
      RECT 49.965 5.015 50.135 8.305 ;
      RECT 49.79 3.055 49.96 3.475 ;
      RECT 49.535 5.015 49.705 7.225 ;
      RECT 49.535 7.795 49.705 8.305 ;
      RECT 48.79 1.755 48.96 2.105 ;
      RECT 47.83 1.755 48 2.105 ;
      RECT 47.83 3.485 48 3.815 ;
      RECT 47.31 3.145 47.48 3.785 ;
      RECT 46.83 1.755 47 2.105 ;
      RECT 46.59 2.495 46.76 2.825 ;
      RECT 46.11 2.495 46.28 2.825 ;
      RECT 44.87 3.145 45.04 3.505 ;
      RECT 44.39 3.055 44.56 3.475 ;
      RECT 43.67 2.495 43.84 2.945 ;
      RECT 41.71 2.495 41.88 2.825 ;
      RECT 40.99 1.755 41.16 2.105 ;
      RECT 40.99 3.285 41.16 3.645 ;
      RECT 39.37 7.8 39.54 8.31 ;
      RECT 38.38 0.57 38.55 1.08 ;
      RECT 38.38 2.39 38.55 3.86 ;
      RECT 38.38 5.02 38.55 6.49 ;
      RECT 38.38 7.8 38.55 8.31 ;
      RECT 37.02 0.575 37.19 3.865 ;
      RECT 37.02 5.015 37.19 8.305 ;
      RECT 36.59 0.575 36.76 1.085 ;
      RECT 36.59 1.655 36.76 3.865 ;
      RECT 36.59 5.015 36.76 7.225 ;
      RECT 36.59 7.795 36.76 8.305 ;
      RECT 32.91 2.495 33.08 2.945 ;
      RECT 32.67 1.755 32.84 2.105 ;
      RECT 31.71 1.755 31.88 2.105 ;
      RECT 31.405 5.015 31.575 8.305 ;
      RECT 31.23 3.055 31.4 3.475 ;
      RECT 30.975 5.015 31.145 7.225 ;
      RECT 30.975 7.795 31.145 8.305 ;
      RECT 30.23 1.755 30.4 2.105 ;
      RECT 29.27 1.755 29.44 2.105 ;
      RECT 29.27 3.485 29.44 3.815 ;
      RECT 28.75 3.145 28.92 3.785 ;
      RECT 28.27 1.755 28.44 2.105 ;
      RECT 28.03 2.495 28.2 2.825 ;
      RECT 27.55 2.495 27.72 2.825 ;
      RECT 26.31 3.145 26.48 3.505 ;
      RECT 25.83 3.055 26 3.475 ;
      RECT 25.11 2.495 25.28 2.945 ;
      RECT 23.15 2.495 23.32 2.825 ;
      RECT 22.43 1.755 22.6 2.105 ;
      RECT 22.43 3.285 22.6 3.645 ;
      RECT 20.81 7.8 20.98 8.31 ;
      RECT 19.82 0.57 19.99 1.08 ;
      RECT 19.82 2.39 19.99 3.86 ;
      RECT 19.82 5.02 19.99 6.49 ;
      RECT 19.82 7.8 19.99 8.31 ;
      RECT 18.46 0.575 18.63 3.865 ;
      RECT 18.46 5.015 18.63 8.305 ;
      RECT 18.03 0.575 18.2 1.085 ;
      RECT 18.03 1.655 18.2 3.865 ;
      RECT 18.03 5.015 18.2 7.225 ;
      RECT 18.03 7.795 18.2 8.305 ;
      RECT 14.35 2.495 14.52 2.945 ;
      RECT 14.11 1.755 14.28 2.105 ;
      RECT 13.15 1.755 13.32 2.105 ;
      RECT 12.845 5.015 13.015 8.305 ;
      RECT 12.67 3.055 12.84 3.475 ;
      RECT 11.67 1.755 11.84 2.105 ;
      RECT 10.71 1.755 10.88 2.105 ;
      RECT 10.71 3.485 10.88 3.815 ;
      RECT 10.19 3.145 10.36 3.785 ;
      RECT 9.71 1.755 9.88 2.105 ;
      RECT 9.47 2.495 9.64 2.825 ;
      RECT 7.75 3.145 7.92 3.505 ;
      RECT 7.27 3.055 7.44 3.475 ;
      RECT 3.87 1.755 4.04 2.105 ;
      RECT 3.87 3.285 4.04 3.645 ;
      RECT 1.6 5.015 1.77 7.225 ;
      RECT 1.6 7.795 1.77 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r2 ;
  SIZE 95.595 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 20.815 0.915 20.985 1.085 ;
        RECT 20.81 0.91 20.98 1.08 ;
        RECT 20.81 2.39 20.98 2.56 ;
      LAYER li1 ;
        RECT 20.815 0.915 20.985 1.085 ;
        RECT 20.81 0.57 20.98 1.08 ;
        RECT 20.81 2.39 20.98 3.86 ;
      LAYER met1 ;
        RECT 20.75 2.36 21.04 2.59 ;
        RECT 20.75 0.88 21.04 1.11 ;
        RECT 20.81 0.88 20.98 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 39.375 0.915 39.545 1.085 ;
        RECT 39.37 0.91 39.54 1.08 ;
        RECT 39.37 2.39 39.54 2.56 ;
      LAYER li1 ;
        RECT 39.375 0.915 39.545 1.085 ;
        RECT 39.37 0.57 39.54 1.08 ;
        RECT 39.37 2.39 39.54 3.86 ;
      LAYER met1 ;
        RECT 39.31 2.36 39.6 2.59 ;
        RECT 39.31 0.88 39.6 1.11 ;
        RECT 39.37 0.88 39.54 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 57.935 0.915 58.105 1.085 ;
        RECT 57.93 0.91 58.1 1.08 ;
        RECT 57.93 2.39 58.1 2.56 ;
      LAYER li1 ;
        RECT 57.935 0.915 58.105 1.085 ;
        RECT 57.93 0.57 58.1 1.08 ;
        RECT 57.93 2.39 58.1 3.86 ;
      LAYER met1 ;
        RECT 57.87 2.36 58.16 2.59 ;
        RECT 57.87 0.88 58.16 1.11 ;
        RECT 57.93 0.88 58.1 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 76.495 0.915 76.665 1.085 ;
        RECT 76.49 0.91 76.66 1.08 ;
        RECT 76.49 2.39 76.66 2.56 ;
      LAYER li1 ;
        RECT 76.495 0.915 76.665 1.085 ;
        RECT 76.49 0.57 76.66 1.08 ;
        RECT 76.49 2.39 76.66 3.86 ;
      LAYER met1 ;
        RECT 76.43 2.36 76.72 2.59 ;
        RECT 76.43 0.88 76.72 1.11 ;
        RECT 76.49 0.88 76.66 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 95.055 0.915 95.225 1.085 ;
        RECT 95.05 0.91 95.22 1.08 ;
        RECT 95.05 2.39 95.22 2.56 ;
      LAYER li1 ;
        RECT 95.055 0.915 95.225 1.085 ;
        RECT 95.05 0.57 95.22 1.08 ;
        RECT 95.05 2.39 95.22 3.86 ;
      LAYER met1 ;
        RECT 94.99 2.36 95.28 2.59 ;
        RECT 94.99 0.88 95.28 1.11 ;
        RECT 95.05 0.88 95.22 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 16.66 1.66 16.83 2.935 ;
        RECT 16.66 5.945 16.83 7.22 ;
        RECT 11.045 5.945 11.215 7.22 ;
      LAYER met2 ;
        RECT 16.585 2.705 16.925 3.055 ;
        RECT 16.575 5.845 16.915 6.195 ;
        RECT 16.66 2.705 16.83 6.195 ;
      LAYER met1 ;
        RECT 16.585 2.765 17.06 2.935 ;
        RECT 16.585 2.705 16.925 3.055 ;
        RECT 10.985 5.945 17.06 6.115 ;
        RECT 16.575 5.845 16.915 6.195 ;
        RECT 10.985 5.915 11.275 6.145 ;
      LAYER mcon ;
        RECT 11.045 5.945 11.215 6.115 ;
        RECT 16.66 5.945 16.83 6.115 ;
        RECT 16.66 2.765 16.83 2.935 ;
      LAYER via1 ;
        RECT 16.675 5.945 16.825 6.095 ;
        RECT 16.685 2.805 16.835 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 35.22 1.66 35.39 2.935 ;
        RECT 35.22 5.945 35.39 7.22 ;
        RECT 29.605 5.945 29.775 7.22 ;
      LAYER met2 ;
        RECT 35.145 2.705 35.485 3.055 ;
        RECT 35.135 5.845 35.475 6.195 ;
        RECT 35.22 2.705 35.39 6.195 ;
      LAYER met1 ;
        RECT 35.145 2.765 35.62 2.935 ;
        RECT 35.145 2.705 35.485 3.055 ;
        RECT 29.545 5.945 35.62 6.115 ;
        RECT 35.135 5.845 35.475 6.195 ;
        RECT 29.545 5.915 29.835 6.145 ;
      LAYER mcon ;
        RECT 29.605 5.945 29.775 6.115 ;
        RECT 35.22 5.945 35.39 6.115 ;
        RECT 35.22 2.765 35.39 2.935 ;
      LAYER via1 ;
        RECT 35.235 5.945 35.385 6.095 ;
        RECT 35.245 2.805 35.395 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 53.78 1.66 53.95 2.935 ;
        RECT 53.78 5.945 53.95 7.22 ;
        RECT 48.165 5.945 48.335 7.22 ;
      LAYER met2 ;
        RECT 53.705 2.705 54.045 3.055 ;
        RECT 53.695 5.845 54.035 6.195 ;
        RECT 53.78 2.705 53.95 6.195 ;
      LAYER met1 ;
        RECT 53.705 2.765 54.18 2.935 ;
        RECT 53.705 2.705 54.045 3.055 ;
        RECT 48.105 5.945 54.18 6.115 ;
        RECT 53.695 5.845 54.035 6.195 ;
        RECT 48.105 5.915 48.395 6.145 ;
      LAYER mcon ;
        RECT 48.165 5.945 48.335 6.115 ;
        RECT 53.78 5.945 53.95 6.115 ;
        RECT 53.78 2.765 53.95 2.935 ;
      LAYER via1 ;
        RECT 53.795 5.945 53.945 6.095 ;
        RECT 53.805 2.805 53.955 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 72.34 1.66 72.51 2.935 ;
        RECT 72.34 5.945 72.51 7.22 ;
        RECT 66.725 5.945 66.895 7.22 ;
      LAYER met2 ;
        RECT 72.265 2.705 72.605 3.055 ;
        RECT 72.255 5.845 72.595 6.195 ;
        RECT 72.34 2.705 72.51 6.195 ;
      LAYER met1 ;
        RECT 72.265 2.765 72.74 2.935 ;
        RECT 72.265 2.705 72.605 3.055 ;
        RECT 66.665 5.945 72.74 6.115 ;
        RECT 72.255 5.845 72.595 6.195 ;
        RECT 66.665 5.915 66.955 6.145 ;
      LAYER mcon ;
        RECT 66.725 5.945 66.895 6.115 ;
        RECT 72.34 5.945 72.51 6.115 ;
        RECT 72.34 2.765 72.51 2.935 ;
      LAYER via1 ;
        RECT 72.355 5.945 72.505 6.095 ;
        RECT 72.365 2.805 72.515 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 90.9 1.66 91.07 2.935 ;
        RECT 90.9 5.945 91.07 7.22 ;
        RECT 85.285 5.945 85.455 7.22 ;
      LAYER met2 ;
        RECT 90.825 2.705 91.165 3.055 ;
        RECT 90.815 5.845 91.155 6.195 ;
        RECT 90.9 2.705 91.07 6.195 ;
      LAYER met1 ;
        RECT 90.825 2.765 91.3 2.935 ;
        RECT 90.825 2.705 91.165 3.055 ;
        RECT 85.225 5.945 91.3 6.115 ;
        RECT 90.815 5.845 91.155 6.195 ;
        RECT 85.225 5.915 85.515 6.145 ;
      LAYER mcon ;
        RECT 85.285 5.945 85.455 6.115 ;
        RECT 90.9 5.945 91.07 6.115 ;
        RECT 90.9 2.765 91.07 2.935 ;
      LAYER via1 ;
        RECT 90.915 5.945 91.065 6.095 ;
        RECT 90.925 2.805 91.075 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 5.945 0.4 7.22 ;
      LAYER met1 ;
        RECT 0.14 5.945 0.63 6.115 ;
        RECT 0.14 5.905 0.48 6.165 ;
      LAYER mcon ;
        RECT 0.23 5.945 0.4 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.435 4.25 2.24 4.63 ;
      LAYER li1 ;
        RECT 77.78 4.135 95.595 4.745 ;
        RECT 93.46 4.13 95.44 4.75 ;
        RECT 94.62 3.4 94.79 5.48 ;
        RECT 93.63 3.4 93.8 5.48 ;
        RECT 90.89 3.405 91.06 5.475 ;
        RECT 87.87 3.635 88.04 4.745 ;
        RECT 85.43 3.635 85.6 4.745 ;
        RECT 85.275 4.135 85.445 5.475 ;
        RECT 83.47 3.635 83.64 4.745 ;
        RECT 82.51 3.635 82.68 4.745 ;
        RECT 80.55 3.635 80.72 4.745 ;
        RECT 79.55 3.635 79.72 4.745 ;
        RECT 77.035 4.145 79.5 4.75 ;
        RECT 78.59 3.635 78.76 4.75 ;
        RECT 59.22 4.135 77.035 4.745 ;
        RECT 74.9 4.13 76.88 4.75 ;
        RECT 76.06 3.4 76.23 5.48 ;
        RECT 75.07 3.4 75.24 5.48 ;
        RECT 72.33 3.405 72.5 5.475 ;
        RECT 69.31 3.635 69.48 4.745 ;
        RECT 66.87 3.635 67.04 4.745 ;
        RECT 66.715 4.135 66.885 5.475 ;
        RECT 64.91 3.635 65.08 4.745 ;
        RECT 63.95 3.635 64.12 4.745 ;
        RECT 61.99 3.635 62.16 4.745 ;
        RECT 60.99 3.635 61.16 4.745 ;
        RECT 58.475 4.145 60.94 4.75 ;
        RECT 60.03 3.635 60.2 4.75 ;
        RECT 40.66 4.135 58.475 4.745 ;
        RECT 56.34 4.13 58.32 4.75 ;
        RECT 57.5 3.4 57.67 5.48 ;
        RECT 56.51 3.4 56.68 5.48 ;
        RECT 53.77 3.405 53.94 5.475 ;
        RECT 50.75 3.635 50.92 4.745 ;
        RECT 48.31 3.635 48.48 4.745 ;
        RECT 48.155 4.135 48.325 5.475 ;
        RECT 46.35 3.635 46.52 4.745 ;
        RECT 45.39 3.635 45.56 4.745 ;
        RECT 43.43 3.635 43.6 4.745 ;
        RECT 42.43 3.635 42.6 4.745 ;
        RECT 39.915 4.145 42.38 4.75 ;
        RECT 41.47 3.635 41.64 4.75 ;
        RECT 22.1 4.135 39.915 4.745 ;
        RECT 37.78 4.13 39.76 4.75 ;
        RECT 38.94 3.4 39.11 5.48 ;
        RECT 37.95 3.4 38.12 5.48 ;
        RECT 35.21 3.405 35.38 5.475 ;
        RECT 32.19 3.635 32.36 4.745 ;
        RECT 29.75 3.635 29.92 4.745 ;
        RECT 29.595 4.135 29.765 5.475 ;
        RECT 27.79 3.635 27.96 4.745 ;
        RECT 26.83 3.635 27 4.745 ;
        RECT 24.87 3.635 25.04 4.745 ;
        RECT 23.87 3.635 24.04 4.745 ;
        RECT 21.355 4.145 23.82 4.75 ;
        RECT 22.91 3.635 23.08 4.75 ;
        RECT 3.54 4.135 21.355 4.745 ;
        RECT 19.22 4.13 21.2 4.75 ;
        RECT 20.38 3.4 20.55 5.48 ;
        RECT 19.39 3.4 19.56 5.48 ;
        RECT 16.65 3.405 16.82 5.475 ;
        RECT 13.63 3.635 13.8 4.745 ;
        RECT 11.19 3.635 11.36 4.745 ;
        RECT 11.035 4.135 11.205 5.475 ;
        RECT 9.23 3.635 9.4 4.745 ;
        RECT 8.27 3.635 8.44 4.745 ;
        RECT 6.31 3.635 6.48 4.745 ;
        RECT 5.31 3.635 5.48 4.745 ;
        RECT 0 4.44 5.26 4.75 ;
        RECT 4.35 3.635 4.52 4.75 ;
        RECT 1.9 4.145 95.595 4.745 ;
        RECT 2.03 4.145 2.2 8.305 ;
        RECT 0 4.145 95.595 4.325 ;
        RECT 0 4.145 1.73 4.75 ;
        RECT 0.22 4.145 0.39 5.475 ;
      LAYER met2 ;
        RECT 1.625 4.25 2.005 4.63 ;
      LAYER met1 ;
        RECT 77.78 4.135 95.595 4.745 ;
        RECT 93.46 4.13 95.44 4.75 ;
        RECT 77.78 3.98 89.74 4.745 ;
        RECT 77.035 4.145 79.5 4.75 ;
        RECT 59.22 4.135 77.035 4.745 ;
        RECT 74.9 4.13 76.88 4.75 ;
        RECT 59.22 3.98 71.18 4.745 ;
        RECT 58.475 4.145 60.94 4.75 ;
        RECT 40.66 4.135 58.475 4.745 ;
        RECT 56.34 4.13 58.32 4.75 ;
        RECT 40.66 3.98 52.62 4.745 ;
        RECT 39.915 4.145 42.38 4.75 ;
        RECT 22.1 4.135 39.915 4.745 ;
        RECT 37.78 4.13 39.76 4.75 ;
        RECT 22.1 3.98 34.06 4.745 ;
        RECT 21.355 4.145 23.82 4.75 ;
        RECT 3.54 4.135 21.355 4.745 ;
        RECT 19.22 4.13 21.2 4.75 ;
        RECT 3.54 3.98 15.5 4.745 ;
        RECT 0 4.145 5.26 4.75 ;
        RECT 1.97 6.655 2.26 6.885 ;
        RECT 1.8 6.685 2.26 6.855 ;
      LAYER via2 ;
        RECT 1.715 4.34 1.915 4.54 ;
      LAYER mcon ;
        RECT 2.03 6.685 2.2 6.855 ;
        RECT 2.34 4.545 2.51 4.715 ;
        RECT 3.685 4.135 3.855 4.305 ;
        RECT 4.145 4.135 4.315 4.305 ;
        RECT 4.605 4.135 4.775 4.305 ;
        RECT 5.065 4.135 5.235 4.305 ;
        RECT 5.525 4.135 5.695 4.305 ;
        RECT 5.985 4.135 6.155 4.305 ;
        RECT 6.445 4.135 6.615 4.305 ;
        RECT 6.905 4.135 7.075 4.305 ;
        RECT 7.365 4.135 7.535 4.305 ;
        RECT 7.825 4.135 7.995 4.305 ;
        RECT 8.285 4.135 8.455 4.305 ;
        RECT 8.745 4.135 8.915 4.305 ;
        RECT 9.205 4.135 9.375 4.305 ;
        RECT 9.665 4.135 9.835 4.305 ;
        RECT 10.125 4.135 10.295 4.305 ;
        RECT 10.585 4.135 10.755 4.305 ;
        RECT 11.045 4.135 11.215 4.305 ;
        RECT 11.505 4.135 11.675 4.305 ;
        RECT 11.965 4.135 12.135 4.305 ;
        RECT 12.425 4.135 12.595 4.305 ;
        RECT 12.885 4.135 13.055 4.305 ;
        RECT 13.155 4.545 13.325 4.715 ;
        RECT 13.345 4.135 13.515 4.305 ;
        RECT 13.805 4.135 13.975 4.305 ;
        RECT 14.265 4.135 14.435 4.305 ;
        RECT 14.725 4.135 14.895 4.305 ;
        RECT 15.185 4.135 15.355 4.305 ;
        RECT 18.77 4.545 18.94 4.715 ;
        RECT 18.77 4.165 18.94 4.335 ;
        RECT 19.47 4.55 19.64 4.72 ;
        RECT 19.47 4.16 19.64 4.33 ;
        RECT 20.46 4.55 20.63 4.72 ;
        RECT 20.46 4.16 20.63 4.33 ;
        RECT 22.245 4.135 22.415 4.305 ;
        RECT 22.705 4.135 22.875 4.305 ;
        RECT 23.165 4.135 23.335 4.305 ;
        RECT 23.625 4.135 23.795 4.305 ;
        RECT 24.085 4.135 24.255 4.305 ;
        RECT 24.545 4.135 24.715 4.305 ;
        RECT 25.005 4.135 25.175 4.305 ;
        RECT 25.465 4.135 25.635 4.305 ;
        RECT 25.925 4.135 26.095 4.305 ;
        RECT 26.385 4.135 26.555 4.305 ;
        RECT 26.845 4.135 27.015 4.305 ;
        RECT 27.305 4.135 27.475 4.305 ;
        RECT 27.765 4.135 27.935 4.305 ;
        RECT 28.225 4.135 28.395 4.305 ;
        RECT 28.685 4.135 28.855 4.305 ;
        RECT 29.145 4.135 29.315 4.305 ;
        RECT 29.605 4.135 29.775 4.305 ;
        RECT 30.065 4.135 30.235 4.305 ;
        RECT 30.525 4.135 30.695 4.305 ;
        RECT 30.985 4.135 31.155 4.305 ;
        RECT 31.445 4.135 31.615 4.305 ;
        RECT 31.715 4.545 31.885 4.715 ;
        RECT 31.905 4.135 32.075 4.305 ;
        RECT 32.365 4.135 32.535 4.305 ;
        RECT 32.825 4.135 32.995 4.305 ;
        RECT 33.285 4.135 33.455 4.305 ;
        RECT 33.745 4.135 33.915 4.305 ;
        RECT 37.33 4.545 37.5 4.715 ;
        RECT 37.33 4.165 37.5 4.335 ;
        RECT 38.03 4.55 38.2 4.72 ;
        RECT 38.03 4.16 38.2 4.33 ;
        RECT 39.02 4.55 39.19 4.72 ;
        RECT 39.02 4.16 39.19 4.33 ;
        RECT 40.805 4.135 40.975 4.305 ;
        RECT 41.265 4.135 41.435 4.305 ;
        RECT 41.725 4.135 41.895 4.305 ;
        RECT 42.185 4.135 42.355 4.305 ;
        RECT 42.645 4.135 42.815 4.305 ;
        RECT 43.105 4.135 43.275 4.305 ;
        RECT 43.565 4.135 43.735 4.305 ;
        RECT 44.025 4.135 44.195 4.305 ;
        RECT 44.485 4.135 44.655 4.305 ;
        RECT 44.945 4.135 45.115 4.305 ;
        RECT 45.405 4.135 45.575 4.305 ;
        RECT 45.865 4.135 46.035 4.305 ;
        RECT 46.325 4.135 46.495 4.305 ;
        RECT 46.785 4.135 46.955 4.305 ;
        RECT 47.245 4.135 47.415 4.305 ;
        RECT 47.705 4.135 47.875 4.305 ;
        RECT 48.165 4.135 48.335 4.305 ;
        RECT 48.625 4.135 48.795 4.305 ;
        RECT 49.085 4.135 49.255 4.305 ;
        RECT 49.545 4.135 49.715 4.305 ;
        RECT 50.005 4.135 50.175 4.305 ;
        RECT 50.275 4.545 50.445 4.715 ;
        RECT 50.465 4.135 50.635 4.305 ;
        RECT 50.925 4.135 51.095 4.305 ;
        RECT 51.385 4.135 51.555 4.305 ;
        RECT 51.845 4.135 52.015 4.305 ;
        RECT 52.305 4.135 52.475 4.305 ;
        RECT 55.89 4.545 56.06 4.715 ;
        RECT 55.89 4.165 56.06 4.335 ;
        RECT 56.59 4.55 56.76 4.72 ;
        RECT 56.59 4.16 56.76 4.33 ;
        RECT 57.58 4.55 57.75 4.72 ;
        RECT 57.58 4.16 57.75 4.33 ;
        RECT 59.365 4.135 59.535 4.305 ;
        RECT 59.825 4.135 59.995 4.305 ;
        RECT 60.285 4.135 60.455 4.305 ;
        RECT 60.745 4.135 60.915 4.305 ;
        RECT 61.205 4.135 61.375 4.305 ;
        RECT 61.665 4.135 61.835 4.305 ;
        RECT 62.125 4.135 62.295 4.305 ;
        RECT 62.585 4.135 62.755 4.305 ;
        RECT 63.045 4.135 63.215 4.305 ;
        RECT 63.505 4.135 63.675 4.305 ;
        RECT 63.965 4.135 64.135 4.305 ;
        RECT 64.425 4.135 64.595 4.305 ;
        RECT 64.885 4.135 65.055 4.305 ;
        RECT 65.345 4.135 65.515 4.305 ;
        RECT 65.805 4.135 65.975 4.305 ;
        RECT 66.265 4.135 66.435 4.305 ;
        RECT 66.725 4.135 66.895 4.305 ;
        RECT 67.185 4.135 67.355 4.305 ;
        RECT 67.645 4.135 67.815 4.305 ;
        RECT 68.105 4.135 68.275 4.305 ;
        RECT 68.565 4.135 68.735 4.305 ;
        RECT 68.835 4.545 69.005 4.715 ;
        RECT 69.025 4.135 69.195 4.305 ;
        RECT 69.485 4.135 69.655 4.305 ;
        RECT 69.945 4.135 70.115 4.305 ;
        RECT 70.405 4.135 70.575 4.305 ;
        RECT 70.865 4.135 71.035 4.305 ;
        RECT 74.45 4.545 74.62 4.715 ;
        RECT 74.45 4.165 74.62 4.335 ;
        RECT 75.15 4.55 75.32 4.72 ;
        RECT 75.15 4.16 75.32 4.33 ;
        RECT 76.14 4.55 76.31 4.72 ;
        RECT 76.14 4.16 76.31 4.33 ;
        RECT 77.925 4.135 78.095 4.305 ;
        RECT 78.385 4.135 78.555 4.305 ;
        RECT 78.845 4.135 79.015 4.305 ;
        RECT 79.305 4.135 79.475 4.305 ;
        RECT 79.765 4.135 79.935 4.305 ;
        RECT 80.225 4.135 80.395 4.305 ;
        RECT 80.685 4.135 80.855 4.305 ;
        RECT 81.145 4.135 81.315 4.305 ;
        RECT 81.605 4.135 81.775 4.305 ;
        RECT 82.065 4.135 82.235 4.305 ;
        RECT 82.525 4.135 82.695 4.305 ;
        RECT 82.985 4.135 83.155 4.305 ;
        RECT 83.445 4.135 83.615 4.305 ;
        RECT 83.905 4.135 84.075 4.305 ;
        RECT 84.365 4.135 84.535 4.305 ;
        RECT 84.825 4.135 84.995 4.305 ;
        RECT 85.285 4.135 85.455 4.305 ;
        RECT 85.745 4.135 85.915 4.305 ;
        RECT 86.205 4.135 86.375 4.305 ;
        RECT 86.665 4.135 86.835 4.305 ;
        RECT 87.125 4.135 87.295 4.305 ;
        RECT 87.395 4.545 87.565 4.715 ;
        RECT 87.585 4.135 87.755 4.305 ;
        RECT 88.045 4.135 88.215 4.305 ;
        RECT 88.505 4.135 88.675 4.305 ;
        RECT 88.965 4.135 89.135 4.305 ;
        RECT 89.425 4.135 89.595 4.305 ;
        RECT 93.01 4.545 93.18 4.715 ;
        RECT 93.01 4.165 93.18 4.335 ;
        RECT 93.71 4.55 93.88 4.72 ;
        RECT 93.71 4.16 93.88 4.33 ;
        RECT 94.7 4.55 94.87 4.72 ;
        RECT 94.7 4.16 94.87 4.33 ;
      LAYER via1 ;
        RECT 1.74 4.365 1.89 4.515 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 79.395 2.415 80.125 2.745 ;
        RECT 60.835 2.415 61.565 2.745 ;
        RECT 42.275 2.415 43.005 2.745 ;
        RECT 23.715 2.415 24.445 2.745 ;
        RECT 5.155 2.415 5.885 2.745 ;
        RECT 0.005 8.5 0.81 8.88 ;
        RECT 0 0 0.805 0.38 ;
      LAYER li1 ;
        RECT 95.415 0 95.595 0.305 ;
        RECT 0.465 0 95.595 0.3 ;
        RECT 94.62 0 94.79 0.93 ;
        RECT 93.63 0 93.8 0.93 ;
        RECT 76.855 0 93.465 0.305 ;
        RECT 90.89 0 91.06 0.935 ;
        RECT 77.78 0 89.825 1.585 ;
        RECT 88.83 0 89 2.085 ;
        RECT 87.87 0 88.04 2.085 ;
        RECT 86.91 0 87.08 2.085 ;
        RECT 86.39 0 86.56 2.085 ;
        RECT 86.11 0 86.305 1.595 ;
        RECT 85.43 0 85.6 2.085 ;
        RECT 84.43 0 84.6 2.085 ;
        RECT 83.47 0 83.64 2.085 ;
        RECT 82.435 0 82.63 1.595 ;
        RECT 81.99 0 82.16 2.085 ;
        RECT 80.07 0 80.33 1.595 ;
        RECT 80.07 0 80.24 2.085 ;
        RECT 78.59 0 78.76 2.085 ;
        RECT 76.06 0 76.23 0.93 ;
        RECT 75.07 0 75.24 0.93 ;
        RECT 58.295 0 74.905 0.305 ;
        RECT 72.33 0 72.5 0.935 ;
        RECT 59.22 0 71.265 1.585 ;
        RECT 70.27 0 70.44 2.085 ;
        RECT 69.31 0 69.48 2.085 ;
        RECT 68.35 0 68.52 2.085 ;
        RECT 67.83 0 68 2.085 ;
        RECT 67.55 0 67.745 1.595 ;
        RECT 66.87 0 67.04 2.085 ;
        RECT 65.87 0 66.04 2.085 ;
        RECT 64.91 0 65.08 2.085 ;
        RECT 63.875 0 64.07 1.595 ;
        RECT 63.43 0 63.6 2.085 ;
        RECT 61.51 0 61.77 1.595 ;
        RECT 61.51 0 61.68 2.085 ;
        RECT 60.03 0 60.2 2.085 ;
        RECT 57.5 0 57.67 0.93 ;
        RECT 56.51 0 56.68 0.93 ;
        RECT 39.735 0 56.345 0.305 ;
        RECT 53.77 0 53.94 0.935 ;
        RECT 40.66 0 52.705 1.585 ;
        RECT 51.71 0 51.88 2.085 ;
        RECT 50.75 0 50.92 2.085 ;
        RECT 49.79 0 49.96 2.085 ;
        RECT 49.27 0 49.44 2.085 ;
        RECT 48.99 0 49.185 1.595 ;
        RECT 48.31 0 48.48 2.085 ;
        RECT 47.31 0 47.48 2.085 ;
        RECT 46.35 0 46.52 2.085 ;
        RECT 45.315 0 45.51 1.595 ;
        RECT 44.87 0 45.04 2.085 ;
        RECT 42.95 0 43.21 1.595 ;
        RECT 42.95 0 43.12 2.085 ;
        RECT 41.47 0 41.64 2.085 ;
        RECT 38.94 0 39.11 0.93 ;
        RECT 37.95 0 38.12 0.93 ;
        RECT 21.175 0 37.785 0.305 ;
        RECT 35.21 0 35.38 0.935 ;
        RECT 22.1 0 34.145 1.585 ;
        RECT 33.15 0 33.32 2.085 ;
        RECT 32.19 0 32.36 2.085 ;
        RECT 31.23 0 31.4 2.085 ;
        RECT 30.71 0 30.88 2.085 ;
        RECT 30.43 0 30.625 1.595 ;
        RECT 29.75 0 29.92 2.085 ;
        RECT 28.75 0 28.92 2.085 ;
        RECT 27.79 0 27.96 2.085 ;
        RECT 26.755 0 26.95 1.595 ;
        RECT 26.31 0 26.48 2.085 ;
        RECT 24.39 0 24.65 1.595 ;
        RECT 24.39 0 24.56 2.085 ;
        RECT 22.91 0 23.08 2.085 ;
        RECT 20.38 0 20.55 0.93 ;
        RECT 19.39 0 19.56 0.93 ;
        RECT 0 0.245 19.225 0.305 ;
        RECT 16.65 0 16.82 0.935 ;
        RECT 3.54 0 15.585 1.585 ;
        RECT 14.59 0 14.76 2.085 ;
        RECT 13.63 0 13.8 2.085 ;
        RECT 12.67 0 12.84 2.085 ;
        RECT 12.15 0 12.32 2.085 ;
        RECT 11.87 0 12.065 1.595 ;
        RECT 11.19 0 11.36 2.085 ;
        RECT 10.19 0 10.36 2.085 ;
        RECT 9.23 0 9.4 2.085 ;
        RECT 8.195 0 8.39 1.595 ;
        RECT 7.75 0 7.92 2.085 ;
        RECT 5.83 0 6.09 1.595 ;
        RECT 5.83 0 6 2.085 ;
        RECT 4.35 0 4.52 2.085 ;
        RECT 0 0.245 0.805 0.315 ;
        RECT 0.295 0.245 0.465 0.335 ;
        RECT 0 0 95.595 0.075 ;
        RECT 0 0 0.295 0.315 ;
        RECT 0 8.58 95.595 8.88 ;
        RECT 95.415 8.575 95.595 8.88 ;
        RECT 94.62 7.95 94.79 8.88 ;
        RECT 93.63 7.95 93.8 8.88 ;
        RECT 76.855 8.575 93.465 8.88 ;
        RECT 90.89 7.945 91.06 8.88 ;
        RECT 85.275 7.945 85.445 8.88 ;
        RECT 76.06 7.95 76.23 8.88 ;
        RECT 75.07 7.95 75.24 8.88 ;
        RECT 58.295 8.575 74.905 8.88 ;
        RECT 72.33 7.945 72.5 8.88 ;
        RECT 66.715 7.945 66.885 8.88 ;
        RECT 57.5 7.95 57.67 8.88 ;
        RECT 56.51 7.95 56.68 8.88 ;
        RECT 39.735 8.575 56.345 8.88 ;
        RECT 53.77 7.945 53.94 8.88 ;
        RECT 48.155 7.945 48.325 8.88 ;
        RECT 38.94 7.95 39.11 8.88 ;
        RECT 37.95 7.95 38.12 8.88 ;
        RECT 21.175 8.575 37.785 8.88 ;
        RECT 35.21 7.945 35.38 8.88 ;
        RECT 29.595 7.945 29.765 8.88 ;
        RECT 20.38 7.95 20.55 8.88 ;
        RECT 19.39 7.95 19.56 8.88 ;
        RECT 0 8.575 19.225 8.88 ;
        RECT 16.65 7.945 16.82 8.88 ;
        RECT 11.035 7.945 11.205 8.88 ;
        RECT 0.005 8.565 0.81 8.88 ;
        RECT 0.22 8.545 0.47 8.88 ;
        RECT 0.22 7.945 0.39 8.88 ;
        RECT 86.28 6.075 86.45 8.025 ;
        RECT 86.225 7.855 86.395 8.305 ;
        RECT 86.225 5.015 86.395 6.245 ;
        RECT 81.27 2.495 81.44 2.825 ;
        RECT 79.43 3.055 79.72 3.225 ;
        RECT 79.43 2.575 79.6 3.225 ;
        RECT 79.23 2.575 79.6 2.745 ;
        RECT 67.72 6.075 67.89 8.025 ;
        RECT 67.665 7.855 67.835 8.305 ;
        RECT 67.665 5.015 67.835 6.245 ;
        RECT 62.71 2.495 62.88 2.825 ;
        RECT 60.87 3.055 61.16 3.225 ;
        RECT 60.87 2.575 61.04 3.225 ;
        RECT 60.67 2.575 61.04 2.745 ;
        RECT 49.16 6.075 49.33 8.025 ;
        RECT 49.105 7.855 49.275 8.305 ;
        RECT 49.105 5.015 49.275 6.245 ;
        RECT 44.15 2.495 44.32 2.825 ;
        RECT 42.31 3.055 42.6 3.225 ;
        RECT 42.31 2.575 42.48 3.225 ;
        RECT 42.11 2.575 42.48 2.745 ;
        RECT 30.6 6.075 30.77 8.025 ;
        RECT 30.545 7.855 30.715 8.305 ;
        RECT 30.545 5.015 30.715 6.245 ;
        RECT 25.59 2.495 25.76 2.825 ;
        RECT 23.75 3.055 24.04 3.225 ;
        RECT 23.75 2.575 23.92 3.225 ;
        RECT 23.55 2.575 23.92 2.745 ;
        RECT 12.04 6.075 12.21 8.025 ;
        RECT 11.985 7.855 12.155 8.305 ;
        RECT 11.985 5.015 12.155 6.245 ;
        RECT 7.03 2.495 7.2 2.825 ;
        RECT 5.19 3.055 5.48 3.225 ;
        RECT 5.19 2.575 5.36 3.225 ;
        RECT 4.99 2.575 5.36 2.745 ;
      LAYER met2 ;
        RECT 81.225 2.42 81.485 2.74 ;
        RECT 79.445 2.51 81.485 2.65 ;
        RECT 79.825 1 80.165 1.34 ;
        RECT 79.755 2.395 80.035 2.765 ;
        RECT 79.85 1 80.02 2.765 ;
        RECT 79.505 2.98 79.765 3.3 ;
        RECT 79.445 2.51 79.585 3.21 ;
        RECT 62.665 2.42 62.925 2.74 ;
        RECT 60.885 2.51 62.925 2.65 ;
        RECT 61.265 1 61.605 1.34 ;
        RECT 61.195 2.395 61.475 2.765 ;
        RECT 61.29 1 61.46 2.765 ;
        RECT 60.945 2.98 61.205 3.3 ;
        RECT 60.885 2.51 61.025 3.21 ;
        RECT 44.105 2.42 44.365 2.74 ;
        RECT 42.325 2.51 44.365 2.65 ;
        RECT 42.705 1 43.045 1.34 ;
        RECT 42.635 2.395 42.915 2.765 ;
        RECT 42.73 1 42.9 2.765 ;
        RECT 42.385 2.98 42.645 3.3 ;
        RECT 42.325 2.51 42.465 3.21 ;
        RECT 25.545 2.42 25.805 2.74 ;
        RECT 23.765 2.51 25.805 2.65 ;
        RECT 24.145 1 24.485 1.34 ;
        RECT 24.075 2.395 24.355 2.765 ;
        RECT 24.17 1 24.34 2.765 ;
        RECT 23.825 2.98 24.085 3.3 ;
        RECT 23.765 2.51 23.905 3.21 ;
        RECT 6.985 2.42 7.245 2.74 ;
        RECT 5.205 2.51 7.245 2.65 ;
        RECT 5.585 1 5.925 1.34 ;
        RECT 5.515 2.395 5.795 2.765 ;
        RECT 5.61 1 5.78 2.765 ;
        RECT 5.265 2.98 5.525 3.3 ;
        RECT 5.205 2.51 5.345 3.21 ;
        RECT 0.195 8.5 0.575 8.88 ;
        RECT 0.19 0 0.57 0.38 ;
        RECT 0.235 0 0.395 8.88 ;
      LAYER met1 ;
        RECT 95.415 0 95.595 0.305 ;
        RECT 0 0 95.595 0.3 ;
        RECT 76.855 0 93.465 0.305 ;
        RECT 77.78 0 89.825 1.585 ;
        RECT 77.78 0 89.74 1.74 ;
        RECT 58.295 0 74.905 0.305 ;
        RECT 59.22 0 71.265 1.585 ;
        RECT 59.22 0 71.18 1.74 ;
        RECT 39.735 0 56.345 0.305 ;
        RECT 40.66 0 52.705 1.585 ;
        RECT 40.66 0 52.62 1.74 ;
        RECT 21.175 0 37.785 0.305 ;
        RECT 22.1 0 34.145 1.585 ;
        RECT 22.1 0 34.06 1.74 ;
        RECT 0 0 19.225 0.305 ;
        RECT 3.54 0 15.585 1.585 ;
        RECT 3.54 0 15.5 1.74 ;
        RECT 0 0 0.805 0.315 ;
        RECT 0.205 0 0.555 0.335 ;
        RECT 0 8.58 95.595 8.88 ;
        RECT 95.415 8.575 95.595 8.88 ;
        RECT 76.855 8.575 93.465 8.88 ;
        RECT 86.22 6.285 86.51 6.515 ;
        RECT 85.785 6.315 86.51 6.485 ;
        RECT 85.785 6.315 85.955 8.88 ;
        RECT 58.295 8.575 74.905 8.88 ;
        RECT 67.66 6.285 67.95 6.515 ;
        RECT 67.225 6.315 67.95 6.485 ;
        RECT 67.225 6.315 67.395 8.88 ;
        RECT 39.735 8.575 56.345 8.88 ;
        RECT 49.1 6.285 49.39 6.515 ;
        RECT 48.665 6.315 49.39 6.485 ;
        RECT 48.665 6.315 48.835 8.88 ;
        RECT 21.175 8.575 37.785 8.88 ;
        RECT 30.54 6.285 30.83 6.515 ;
        RECT 30.105 6.315 30.83 6.485 ;
        RECT 30.105 6.315 30.275 8.88 ;
        RECT 0 8.575 19.225 8.88 ;
        RECT 11.98 6.285 12.27 6.515 ;
        RECT 11.545 6.315 12.27 6.485 ;
        RECT 11.545 6.315 11.715 8.88 ;
        RECT 0.005 8.565 0.81 8.88 ;
        RECT 0.21 8.545 0.56 8.88 ;
        RECT 81.21 2.37 81.5 2.74 ;
        RECT 80.445 2.37 81.5 2.51 ;
        RECT 79.475 3.01 79.795 3.27 ;
        RECT 62.65 2.37 62.94 2.74 ;
        RECT 61.885 2.37 62.94 2.51 ;
        RECT 60.915 3.01 61.235 3.27 ;
        RECT 44.09 2.37 44.38 2.74 ;
        RECT 43.325 2.37 44.38 2.51 ;
        RECT 42.355 3.01 42.675 3.27 ;
        RECT 25.53 2.37 25.82 2.74 ;
        RECT 24.765 2.37 25.82 2.51 ;
        RECT 23.795 3.01 24.115 3.27 ;
        RECT 6.97 2.37 7.26 2.74 ;
        RECT 6.205 2.37 7.26 2.51 ;
        RECT 5.235 3.01 5.555 3.27 ;
      LAYER via2 ;
        RECT 0.28 0.09 0.48 0.29 ;
        RECT 0.285 8.59 0.485 8.79 ;
        RECT 5.555 2.48 5.755 2.68 ;
        RECT 24.115 2.48 24.315 2.68 ;
        RECT 42.675 2.48 42.875 2.68 ;
        RECT 61.235 2.48 61.435 2.68 ;
        RECT 79.795 2.48 79.995 2.68 ;
      LAYER mcon ;
        RECT 0.3 8.605 0.47 8.775 ;
        RECT 0.98 8.605 1.15 8.775 ;
        RECT 1.66 8.605 1.83 8.775 ;
        RECT 2.34 8.605 2.51 8.775 ;
        RECT 3.685 1.415 3.855 1.585 ;
        RECT 4.145 1.415 4.315 1.585 ;
        RECT 4.605 1.415 4.775 1.585 ;
        RECT 5.065 1.415 5.235 1.585 ;
        RECT 5.31 3.055 5.48 3.225 ;
        RECT 5.525 1.415 5.695 1.585 ;
        RECT 5.985 1.415 6.155 1.585 ;
        RECT 6.445 1.415 6.615 1.585 ;
        RECT 6.905 1.415 7.075 1.585 ;
        RECT 7.03 2.495 7.2 2.665 ;
        RECT 7.365 1.415 7.535 1.585 ;
        RECT 7.825 1.415 7.995 1.585 ;
        RECT 8.285 1.415 8.455 1.585 ;
        RECT 8.745 1.415 8.915 1.585 ;
        RECT 9.205 1.415 9.375 1.585 ;
        RECT 9.665 1.415 9.835 1.585 ;
        RECT 10.125 1.415 10.295 1.585 ;
        RECT 10.585 1.415 10.755 1.585 ;
        RECT 11.045 1.415 11.215 1.585 ;
        RECT 11.115 8.605 11.285 8.775 ;
        RECT 11.505 1.415 11.675 1.585 ;
        RECT 11.795 8.605 11.965 8.775 ;
        RECT 11.965 1.415 12.135 1.585 ;
        RECT 12.04 6.315 12.21 6.485 ;
        RECT 12.425 1.415 12.595 1.585 ;
        RECT 12.475 8.605 12.645 8.775 ;
        RECT 12.885 1.415 13.055 1.585 ;
        RECT 13.155 8.605 13.325 8.775 ;
        RECT 13.345 1.415 13.515 1.585 ;
        RECT 13.805 1.415 13.975 1.585 ;
        RECT 14.265 1.415 14.435 1.585 ;
        RECT 14.725 1.415 14.895 1.585 ;
        RECT 15.185 1.415 15.355 1.585 ;
        RECT 16.73 8.605 16.9 8.775 ;
        RECT 16.73 0.105 16.9 0.275 ;
        RECT 17.41 8.605 17.58 8.775 ;
        RECT 17.41 0.105 17.58 0.275 ;
        RECT 18.09 8.605 18.26 8.775 ;
        RECT 18.09 0.105 18.26 0.275 ;
        RECT 18.77 8.605 18.94 8.775 ;
        RECT 18.77 0.105 18.94 0.275 ;
        RECT 19.47 8.61 19.64 8.78 ;
        RECT 19.47 0.1 19.64 0.27 ;
        RECT 20.46 8.61 20.63 8.78 ;
        RECT 20.46 0.1 20.63 0.27 ;
        RECT 22.245 1.415 22.415 1.585 ;
        RECT 22.705 1.415 22.875 1.585 ;
        RECT 23.165 1.415 23.335 1.585 ;
        RECT 23.625 1.415 23.795 1.585 ;
        RECT 23.87 3.055 24.04 3.225 ;
        RECT 24.085 1.415 24.255 1.585 ;
        RECT 24.545 1.415 24.715 1.585 ;
        RECT 25.005 1.415 25.175 1.585 ;
        RECT 25.465 1.415 25.635 1.585 ;
        RECT 25.59 2.495 25.76 2.665 ;
        RECT 25.925 1.415 26.095 1.585 ;
        RECT 26.385 1.415 26.555 1.585 ;
        RECT 26.845 1.415 27.015 1.585 ;
        RECT 27.305 1.415 27.475 1.585 ;
        RECT 27.765 1.415 27.935 1.585 ;
        RECT 28.225 1.415 28.395 1.585 ;
        RECT 28.685 1.415 28.855 1.585 ;
        RECT 29.145 1.415 29.315 1.585 ;
        RECT 29.605 1.415 29.775 1.585 ;
        RECT 29.675 8.605 29.845 8.775 ;
        RECT 30.065 1.415 30.235 1.585 ;
        RECT 30.355 8.605 30.525 8.775 ;
        RECT 30.525 1.415 30.695 1.585 ;
        RECT 30.6 6.315 30.77 6.485 ;
        RECT 30.985 1.415 31.155 1.585 ;
        RECT 31.035 8.605 31.205 8.775 ;
        RECT 31.445 1.415 31.615 1.585 ;
        RECT 31.715 8.605 31.885 8.775 ;
        RECT 31.905 1.415 32.075 1.585 ;
        RECT 32.365 1.415 32.535 1.585 ;
        RECT 32.825 1.415 32.995 1.585 ;
        RECT 33.285 1.415 33.455 1.585 ;
        RECT 33.745 1.415 33.915 1.585 ;
        RECT 35.29 8.605 35.46 8.775 ;
        RECT 35.29 0.105 35.46 0.275 ;
        RECT 35.97 8.605 36.14 8.775 ;
        RECT 35.97 0.105 36.14 0.275 ;
        RECT 36.65 8.605 36.82 8.775 ;
        RECT 36.65 0.105 36.82 0.275 ;
        RECT 37.33 8.605 37.5 8.775 ;
        RECT 37.33 0.105 37.5 0.275 ;
        RECT 38.03 8.61 38.2 8.78 ;
        RECT 38.03 0.1 38.2 0.27 ;
        RECT 39.02 8.61 39.19 8.78 ;
        RECT 39.02 0.1 39.19 0.27 ;
        RECT 40.805 1.415 40.975 1.585 ;
        RECT 41.265 1.415 41.435 1.585 ;
        RECT 41.725 1.415 41.895 1.585 ;
        RECT 42.185 1.415 42.355 1.585 ;
        RECT 42.43 3.055 42.6 3.225 ;
        RECT 42.645 1.415 42.815 1.585 ;
        RECT 43.105 1.415 43.275 1.585 ;
        RECT 43.565 1.415 43.735 1.585 ;
        RECT 44.025 1.415 44.195 1.585 ;
        RECT 44.15 2.495 44.32 2.665 ;
        RECT 44.485 1.415 44.655 1.585 ;
        RECT 44.945 1.415 45.115 1.585 ;
        RECT 45.405 1.415 45.575 1.585 ;
        RECT 45.865 1.415 46.035 1.585 ;
        RECT 46.325 1.415 46.495 1.585 ;
        RECT 46.785 1.415 46.955 1.585 ;
        RECT 47.245 1.415 47.415 1.585 ;
        RECT 47.705 1.415 47.875 1.585 ;
        RECT 48.165 1.415 48.335 1.585 ;
        RECT 48.235 8.605 48.405 8.775 ;
        RECT 48.625 1.415 48.795 1.585 ;
        RECT 48.915 8.605 49.085 8.775 ;
        RECT 49.085 1.415 49.255 1.585 ;
        RECT 49.16 6.315 49.33 6.485 ;
        RECT 49.545 1.415 49.715 1.585 ;
        RECT 49.595 8.605 49.765 8.775 ;
        RECT 50.005 1.415 50.175 1.585 ;
        RECT 50.275 8.605 50.445 8.775 ;
        RECT 50.465 1.415 50.635 1.585 ;
        RECT 50.925 1.415 51.095 1.585 ;
        RECT 51.385 1.415 51.555 1.585 ;
        RECT 51.845 1.415 52.015 1.585 ;
        RECT 52.305 1.415 52.475 1.585 ;
        RECT 53.85 8.605 54.02 8.775 ;
        RECT 53.85 0.105 54.02 0.275 ;
        RECT 54.53 8.605 54.7 8.775 ;
        RECT 54.53 0.105 54.7 0.275 ;
        RECT 55.21 8.605 55.38 8.775 ;
        RECT 55.21 0.105 55.38 0.275 ;
        RECT 55.89 8.605 56.06 8.775 ;
        RECT 55.89 0.105 56.06 0.275 ;
        RECT 56.59 8.61 56.76 8.78 ;
        RECT 56.59 0.1 56.76 0.27 ;
        RECT 57.58 8.61 57.75 8.78 ;
        RECT 57.58 0.1 57.75 0.27 ;
        RECT 59.365 1.415 59.535 1.585 ;
        RECT 59.825 1.415 59.995 1.585 ;
        RECT 60.285 1.415 60.455 1.585 ;
        RECT 60.745 1.415 60.915 1.585 ;
        RECT 60.99 3.055 61.16 3.225 ;
        RECT 61.205 1.415 61.375 1.585 ;
        RECT 61.665 1.415 61.835 1.585 ;
        RECT 62.125 1.415 62.295 1.585 ;
        RECT 62.585 1.415 62.755 1.585 ;
        RECT 62.71 2.495 62.88 2.665 ;
        RECT 63.045 1.415 63.215 1.585 ;
        RECT 63.505 1.415 63.675 1.585 ;
        RECT 63.965 1.415 64.135 1.585 ;
        RECT 64.425 1.415 64.595 1.585 ;
        RECT 64.885 1.415 65.055 1.585 ;
        RECT 65.345 1.415 65.515 1.585 ;
        RECT 65.805 1.415 65.975 1.585 ;
        RECT 66.265 1.415 66.435 1.585 ;
        RECT 66.725 1.415 66.895 1.585 ;
        RECT 66.795 8.605 66.965 8.775 ;
        RECT 67.185 1.415 67.355 1.585 ;
        RECT 67.475 8.605 67.645 8.775 ;
        RECT 67.645 1.415 67.815 1.585 ;
        RECT 67.72 6.315 67.89 6.485 ;
        RECT 68.105 1.415 68.275 1.585 ;
        RECT 68.155 8.605 68.325 8.775 ;
        RECT 68.565 1.415 68.735 1.585 ;
        RECT 68.835 8.605 69.005 8.775 ;
        RECT 69.025 1.415 69.195 1.585 ;
        RECT 69.485 1.415 69.655 1.585 ;
        RECT 69.945 1.415 70.115 1.585 ;
        RECT 70.405 1.415 70.575 1.585 ;
        RECT 70.865 1.415 71.035 1.585 ;
        RECT 72.41 8.605 72.58 8.775 ;
        RECT 72.41 0.105 72.58 0.275 ;
        RECT 73.09 8.605 73.26 8.775 ;
        RECT 73.09 0.105 73.26 0.275 ;
        RECT 73.77 8.605 73.94 8.775 ;
        RECT 73.77 0.105 73.94 0.275 ;
        RECT 74.45 8.605 74.62 8.775 ;
        RECT 74.45 0.105 74.62 0.275 ;
        RECT 75.15 8.61 75.32 8.78 ;
        RECT 75.15 0.1 75.32 0.27 ;
        RECT 76.14 8.61 76.31 8.78 ;
        RECT 76.14 0.1 76.31 0.27 ;
        RECT 77.925 1.415 78.095 1.585 ;
        RECT 78.385 1.415 78.555 1.585 ;
        RECT 78.845 1.415 79.015 1.585 ;
        RECT 79.305 1.415 79.475 1.585 ;
        RECT 79.55 3.055 79.72 3.225 ;
        RECT 79.765 1.415 79.935 1.585 ;
        RECT 80.225 1.415 80.395 1.585 ;
        RECT 80.685 1.415 80.855 1.585 ;
        RECT 81.145 1.415 81.315 1.585 ;
        RECT 81.27 2.495 81.44 2.665 ;
        RECT 81.605 1.415 81.775 1.585 ;
        RECT 82.065 1.415 82.235 1.585 ;
        RECT 82.525 1.415 82.695 1.585 ;
        RECT 82.985 1.415 83.155 1.585 ;
        RECT 83.445 1.415 83.615 1.585 ;
        RECT 83.905 1.415 84.075 1.585 ;
        RECT 84.365 1.415 84.535 1.585 ;
        RECT 84.825 1.415 84.995 1.585 ;
        RECT 85.285 1.415 85.455 1.585 ;
        RECT 85.355 8.605 85.525 8.775 ;
        RECT 85.745 1.415 85.915 1.585 ;
        RECT 86.035 8.605 86.205 8.775 ;
        RECT 86.205 1.415 86.375 1.585 ;
        RECT 86.28 6.315 86.45 6.485 ;
        RECT 86.665 1.415 86.835 1.585 ;
        RECT 86.715 8.605 86.885 8.775 ;
        RECT 87.125 1.415 87.295 1.585 ;
        RECT 87.395 8.605 87.565 8.775 ;
        RECT 87.585 1.415 87.755 1.585 ;
        RECT 88.045 1.415 88.215 1.585 ;
        RECT 88.505 1.415 88.675 1.585 ;
        RECT 88.965 1.415 89.135 1.585 ;
        RECT 89.425 1.415 89.595 1.585 ;
        RECT 90.97 8.605 91.14 8.775 ;
        RECT 90.97 0.105 91.14 0.275 ;
        RECT 91.65 8.605 91.82 8.775 ;
        RECT 91.65 0.105 91.82 0.275 ;
        RECT 92.33 8.605 92.5 8.775 ;
        RECT 92.33 0.105 92.5 0.275 ;
        RECT 93.01 8.605 93.18 8.775 ;
        RECT 93.01 0.105 93.18 0.275 ;
        RECT 93.71 8.61 93.88 8.78 ;
        RECT 93.71 0.1 93.88 0.27 ;
        RECT 94.7 8.61 94.87 8.78 ;
        RECT 94.7 0.1 94.87 0.27 ;
      LAYER via1 ;
        RECT 0.305 0.115 0.455 0.265 ;
        RECT 0.31 8.615 0.46 8.765 ;
        RECT 5.32 3.065 5.47 3.215 ;
        RECT 5.68 1.095 5.83 1.245 ;
        RECT 7.04 2.505 7.19 2.655 ;
        RECT 23.88 3.065 24.03 3.215 ;
        RECT 24.24 1.095 24.39 1.245 ;
        RECT 25.6 2.505 25.75 2.655 ;
        RECT 42.44 3.065 42.59 3.215 ;
        RECT 42.8 1.095 42.95 1.245 ;
        RECT 44.16 2.505 44.31 2.655 ;
        RECT 61 3.065 61.15 3.215 ;
        RECT 61.36 1.095 61.51 1.245 ;
        RECT 62.72 2.505 62.87 2.655 ;
        RECT 79.56 3.065 79.71 3.215 ;
        RECT 79.92 1.095 80.07 1.245 ;
        RECT 81.28 2.505 81.43 2.655 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 87.085 3.535 87.64 3.865 ;
      RECT 87.085 1.87 87.385 3.865 ;
      RECT 83.15 2.975 83.705 3.305 ;
      RECT 83.405 1.87 83.705 3.305 ;
      RECT 83.405 1.87 87.385 2.17 ;
      RECT 86.555 7.055 86.93 7.425 ;
      RECT 86.555 7.095 87.56 7.395 ;
      RECT 87.26 4.405 87.56 7.395 ;
      RECT 77.43 4.405 87.56 4.705 ;
      RECT 81.935 2.415 82.235 4.705 ;
      RECT 80.5 2.975 80.8 4.705 ;
      RECT 77.43 2.42 77.73 4.705 ;
      RECT 80.47 2.975 81.2 3.305 ;
      RECT 81.91 2.415 82.64 2.745 ;
      RECT 78.36 2.415 79.09 2.745 ;
      RECT 77.43 2.42 79.09 2.72 ;
      RECT 68.525 3.535 69.08 3.865 ;
      RECT 68.525 1.87 68.825 3.865 ;
      RECT 64.59 2.975 65.145 3.305 ;
      RECT 64.845 1.87 65.145 3.305 ;
      RECT 64.845 1.87 68.825 2.17 ;
      RECT 67.995 7.055 68.37 7.425 ;
      RECT 67.995 7.095 69 7.395 ;
      RECT 68.7 4.405 69 7.395 ;
      RECT 58.87 4.405 69 4.705 ;
      RECT 63.375 2.415 63.675 4.705 ;
      RECT 61.94 2.975 62.24 4.705 ;
      RECT 58.87 2.42 59.17 4.705 ;
      RECT 61.91 2.975 62.64 3.305 ;
      RECT 63.35 2.415 64.08 2.745 ;
      RECT 59.8 2.415 60.53 2.745 ;
      RECT 58.87 2.42 60.53 2.72 ;
      RECT 49.965 3.535 50.52 3.865 ;
      RECT 49.965 1.87 50.265 3.865 ;
      RECT 46.03 2.975 46.585 3.305 ;
      RECT 46.285 1.87 46.585 3.305 ;
      RECT 46.285 1.87 50.265 2.17 ;
      RECT 49.435 7.055 49.81 7.425 ;
      RECT 49.435 7.095 50.44 7.395 ;
      RECT 50.14 4.405 50.44 7.395 ;
      RECT 40.31 4.405 50.44 4.705 ;
      RECT 44.815 2.415 45.115 4.705 ;
      RECT 43.38 2.975 43.68 4.705 ;
      RECT 40.31 2.42 40.61 4.705 ;
      RECT 43.35 2.975 44.08 3.305 ;
      RECT 44.79 2.415 45.52 2.745 ;
      RECT 41.24 2.415 41.97 2.745 ;
      RECT 40.31 2.42 41.97 2.72 ;
      RECT 31.405 3.535 31.96 3.865 ;
      RECT 31.405 1.87 31.705 3.865 ;
      RECT 27.47 2.975 28.025 3.305 ;
      RECT 27.725 1.87 28.025 3.305 ;
      RECT 27.725 1.87 31.705 2.17 ;
      RECT 30.875 7.055 31.25 7.425 ;
      RECT 30.875 7.095 31.88 7.395 ;
      RECT 31.58 4.405 31.88 7.395 ;
      RECT 21.75 4.405 31.88 4.705 ;
      RECT 26.255 2.415 26.555 4.705 ;
      RECT 24.82 2.975 25.12 4.705 ;
      RECT 21.75 2.42 22.05 4.705 ;
      RECT 24.79 2.975 25.52 3.305 ;
      RECT 26.23 2.415 26.96 2.745 ;
      RECT 22.68 2.415 23.41 2.745 ;
      RECT 21.75 2.42 23.41 2.72 ;
      RECT 12.845 3.535 13.4 3.865 ;
      RECT 12.845 1.87 13.145 3.865 ;
      RECT 8.91 2.975 9.465 3.305 ;
      RECT 9.165 1.87 9.465 3.305 ;
      RECT 9.165 1.87 13.145 2.17 ;
      RECT 12.315 7.055 12.69 7.425 ;
      RECT 12.315 7.095 13.32 7.395 ;
      RECT 13.02 4.405 13.32 7.395 ;
      RECT 3.19 4.405 13.32 4.705 ;
      RECT 7.695 2.415 7.995 4.705 ;
      RECT 6.26 2.975 6.56 4.705 ;
      RECT 3.19 2.42 3.49 4.705 ;
      RECT 6.23 2.975 6.96 3.305 ;
      RECT 7.67 2.415 8.4 2.745 ;
      RECT 4.12 2.415 4.85 2.745 ;
      RECT 3.19 2.42 4.85 2.72 ;
      RECT 88.27 1.855 89 2.185 ;
      RECT 86.05 3.535 86.78 3.865 ;
      RECT 84.35 3.535 85.08 3.865 ;
      RECT 78.03 3.535 78.76 3.865 ;
      RECT 69.71 1.855 70.44 2.185 ;
      RECT 67.49 3.535 68.22 3.865 ;
      RECT 65.79 3.535 66.52 3.865 ;
      RECT 59.47 3.535 60.2 3.865 ;
      RECT 51.15 1.855 51.88 2.185 ;
      RECT 48.93 3.535 49.66 3.865 ;
      RECT 47.23 3.535 47.96 3.865 ;
      RECT 40.91 3.535 41.64 3.865 ;
      RECT 32.59 1.855 33.32 2.185 ;
      RECT 30.37 3.535 31.1 3.865 ;
      RECT 28.67 3.535 29.4 3.865 ;
      RECT 22.35 3.535 23.08 3.865 ;
      RECT 14.03 1.855 14.76 2.185 ;
      RECT 11.81 3.535 12.54 3.865 ;
      RECT 10.11 3.535 10.84 3.865 ;
      RECT 3.79 3.535 4.52 3.865 ;
    LAYER via2 ;
      RECT 88.335 1.92 88.535 2.12 ;
      RECT 87.375 3.6 87.575 3.8 ;
      RECT 86.64 7.14 86.84 7.34 ;
      RECT 86.375 3.6 86.575 3.8 ;
      RECT 84.415 3.6 84.615 3.8 ;
      RECT 83.215 3.04 83.415 3.24 ;
      RECT 81.975 2.48 82.175 2.68 ;
      RECT 80.535 3.04 80.735 3.24 ;
      RECT 78.575 2.48 78.775 2.68 ;
      RECT 78.095 3.6 78.295 3.8 ;
      RECT 69.775 1.92 69.975 2.12 ;
      RECT 68.815 3.6 69.015 3.8 ;
      RECT 68.08 7.14 68.28 7.34 ;
      RECT 67.815 3.6 68.015 3.8 ;
      RECT 65.855 3.6 66.055 3.8 ;
      RECT 64.655 3.04 64.855 3.24 ;
      RECT 63.415 2.48 63.615 2.68 ;
      RECT 61.975 3.04 62.175 3.24 ;
      RECT 60.015 2.48 60.215 2.68 ;
      RECT 59.535 3.6 59.735 3.8 ;
      RECT 51.215 1.92 51.415 2.12 ;
      RECT 50.255 3.6 50.455 3.8 ;
      RECT 49.52 7.14 49.72 7.34 ;
      RECT 49.255 3.6 49.455 3.8 ;
      RECT 47.295 3.6 47.495 3.8 ;
      RECT 46.095 3.04 46.295 3.24 ;
      RECT 44.855 2.48 45.055 2.68 ;
      RECT 43.415 3.04 43.615 3.24 ;
      RECT 41.455 2.48 41.655 2.68 ;
      RECT 40.975 3.6 41.175 3.8 ;
      RECT 32.655 1.92 32.855 2.12 ;
      RECT 31.695 3.6 31.895 3.8 ;
      RECT 30.96 7.14 31.16 7.34 ;
      RECT 30.695 3.6 30.895 3.8 ;
      RECT 28.735 3.6 28.935 3.8 ;
      RECT 27.535 3.04 27.735 3.24 ;
      RECT 26.295 2.48 26.495 2.68 ;
      RECT 24.855 3.04 25.055 3.24 ;
      RECT 22.895 2.48 23.095 2.68 ;
      RECT 22.415 3.6 22.615 3.8 ;
      RECT 14.095 1.92 14.295 2.12 ;
      RECT 13.135 3.6 13.335 3.8 ;
      RECT 12.4 7.14 12.6 7.34 ;
      RECT 12.135 3.6 12.335 3.8 ;
      RECT 10.175 3.6 10.375 3.8 ;
      RECT 8.975 3.04 9.175 3.24 ;
      RECT 7.735 2.48 7.935 2.68 ;
      RECT 6.295 3.04 6.495 3.24 ;
      RECT 4.335 2.48 4.535 2.68 ;
      RECT 3.855 3.6 4.055 3.8 ;
    LAYER met2 ;
      RECT 1.225 8.4 95.225 8.57 ;
      RECT 95.055 7.275 95.225 8.57 ;
      RECT 1.225 6.255 1.395 8.57 ;
      RECT 95.025 7.275 95.375 7.625 ;
      RECT 1.165 6.255 1.455 6.605 ;
      RECT 91.865 6.22 92.185 6.545 ;
      RECT 91.895 5.695 92.065 6.545 ;
      RECT 91.895 5.695 92.07 6.045 ;
      RECT 91.895 5.695 92.87 5.87 ;
      RECT 92.695 1.965 92.87 5.87 ;
      RECT 92.64 1.965 92.99 2.315 ;
      RECT 92.665 6.655 92.99 6.98 ;
      RECT 91.55 6.745 92.99 6.915 ;
      RECT 91.55 2.395 91.71 6.915 ;
      RECT 91.865 2.365 92.185 2.685 ;
      RECT 91.55 2.395 92.185 2.565 ;
      RECT 84.43 4.135 90.52 4.325 ;
      RECT 90.35 3.145 90.52 4.325 ;
      RECT 90.33 3.15 90.52 4.325 ;
      RECT 84.43 3.515 84.6 4.325 ;
      RECT 84.375 3.515 84.655 3.885 ;
      RECT 84.445 3.07 84.585 4.325 ;
      RECT 90.26 3.15 90.6 3.5 ;
      RECT 84.255 2.955 84.535 3.325 ;
      RECT 83.965 3.07 84.585 3.21 ;
      RECT 83.965 1.86 84.105 3.21 ;
      RECT 83.905 1.86 84.165 2.18 ;
      RECT 76.44 6.655 76.79 7.005 ;
      RECT 87.225 6.61 87.575 6.96 ;
      RECT 76.44 6.685 87.575 6.885 ;
      RECT 86.865 2.98 87.125 3.3 ;
      RECT 86.925 1.86 87.065 3.3 ;
      RECT 86.865 1.86 87.125 2.18 ;
      RECT 85.865 3.54 86.125 3.86 ;
      RECT 85.865 2.955 86.065 3.86 ;
      RECT 85.805 1.86 85.945 3.49 ;
      RECT 85.805 2.955 86.305 3.325 ;
      RECT 85.745 1.86 86.005 2.18 ;
      RECT 85.385 3.54 85.645 3.86 ;
      RECT 85.445 1.95 85.585 3.86 ;
      RECT 85.145 1.95 85.585 2.18 ;
      RECT 85.145 1.86 85.405 2.18 ;
      RECT 84.905 2.42 85.165 2.74 ;
      RECT 84.325 2.51 85.165 2.65 ;
      RECT 84.325 1.57 84.465 2.65 ;
      RECT 80.985 1.86 81.245 2.18 ;
      RECT 80.985 1.95 82.025 2.09 ;
      RECT 81.885 1.57 82.025 2.09 ;
      RECT 81.885 1.57 84.465 1.71 ;
      RECT 83.175 2.955 83.455 3.325 ;
      RECT 83.245 1.86 83.385 3.325 ;
      RECT 83.185 1.86 83.445 2.18 ;
      RECT 82.825 3.54 83.085 3.86 ;
      RECT 82.885 1.95 83.025 3.86 ;
      RECT 82.465 1.86 82.725 2.18 ;
      RECT 82.465 1.95 83.025 2.09 ;
      RECT 80.495 2.955 80.775 3.325 ;
      RECT 82.465 2.98 82.725 3.3 ;
      RECT 80.145 2.98 80.775 3.3 ;
      RECT 80.145 3.07 82.725 3.21 ;
      RECT 81.935 2.395 82.215 2.765 ;
      RECT 81.935 2.42 82.465 2.74 ;
      RECT 79.025 2.98 79.285 3.3 ;
      RECT 79.085 1.86 79.225 3.3 ;
      RECT 79.025 1.86 79.285 2.18 ;
      RECT 78.055 3.515 78.335 3.885 ;
      RECT 78.065 3.26 78.325 3.885 ;
      RECT 73.305 6.22 73.625 6.545 ;
      RECT 73.335 5.695 73.505 6.545 ;
      RECT 73.335 5.695 73.51 6.045 ;
      RECT 73.335 5.695 74.31 5.87 ;
      RECT 74.135 1.965 74.31 5.87 ;
      RECT 74.08 1.965 74.43 2.315 ;
      RECT 74.105 6.655 74.43 6.98 ;
      RECT 72.99 6.745 74.43 6.915 ;
      RECT 72.99 2.395 73.15 6.915 ;
      RECT 73.305 2.365 73.625 2.685 ;
      RECT 72.99 2.395 73.625 2.565 ;
      RECT 65.87 4.135 71.96 4.325 ;
      RECT 71.79 3.145 71.96 4.325 ;
      RECT 71.77 3.15 71.96 4.325 ;
      RECT 65.87 3.515 66.04 4.325 ;
      RECT 65.815 3.515 66.095 3.885 ;
      RECT 65.885 3.07 66.025 4.325 ;
      RECT 71.7 3.15 72.04 3.5 ;
      RECT 65.695 2.955 65.975 3.325 ;
      RECT 65.405 3.07 66.025 3.21 ;
      RECT 65.405 1.86 65.545 3.21 ;
      RECT 65.345 1.86 65.605 2.18 ;
      RECT 57.88 6.655 58.23 7.005 ;
      RECT 68.665 6.61 69.015 6.96 ;
      RECT 57.88 6.685 69.015 6.885 ;
      RECT 68.305 2.98 68.565 3.3 ;
      RECT 68.365 1.86 68.505 3.3 ;
      RECT 68.305 1.86 68.565 2.18 ;
      RECT 67.305 3.54 67.565 3.86 ;
      RECT 67.305 2.955 67.505 3.86 ;
      RECT 67.245 1.86 67.385 3.49 ;
      RECT 67.245 2.955 67.745 3.325 ;
      RECT 67.185 1.86 67.445 2.18 ;
      RECT 66.825 3.54 67.085 3.86 ;
      RECT 66.885 1.95 67.025 3.86 ;
      RECT 66.585 1.95 67.025 2.18 ;
      RECT 66.585 1.86 66.845 2.18 ;
      RECT 66.345 2.42 66.605 2.74 ;
      RECT 65.765 2.51 66.605 2.65 ;
      RECT 65.765 1.57 65.905 2.65 ;
      RECT 62.425 1.86 62.685 2.18 ;
      RECT 62.425 1.95 63.465 2.09 ;
      RECT 63.325 1.57 63.465 2.09 ;
      RECT 63.325 1.57 65.905 1.71 ;
      RECT 64.615 2.955 64.895 3.325 ;
      RECT 64.685 1.86 64.825 3.325 ;
      RECT 64.625 1.86 64.885 2.18 ;
      RECT 64.265 3.54 64.525 3.86 ;
      RECT 64.325 1.95 64.465 3.86 ;
      RECT 63.905 1.86 64.165 2.18 ;
      RECT 63.905 1.95 64.465 2.09 ;
      RECT 61.935 2.955 62.215 3.325 ;
      RECT 63.905 2.98 64.165 3.3 ;
      RECT 61.585 2.98 62.215 3.3 ;
      RECT 61.585 3.07 64.165 3.21 ;
      RECT 63.375 2.395 63.655 2.765 ;
      RECT 63.375 2.42 63.905 2.74 ;
      RECT 60.465 2.98 60.725 3.3 ;
      RECT 60.525 1.86 60.665 3.3 ;
      RECT 60.465 1.86 60.725 2.18 ;
      RECT 59.495 3.515 59.775 3.885 ;
      RECT 59.505 3.26 59.765 3.885 ;
      RECT 54.745 6.22 55.065 6.545 ;
      RECT 54.775 5.695 54.945 6.545 ;
      RECT 54.775 5.695 54.95 6.045 ;
      RECT 54.775 5.695 55.75 5.87 ;
      RECT 55.575 1.965 55.75 5.87 ;
      RECT 55.52 1.965 55.87 2.315 ;
      RECT 55.545 6.655 55.87 6.98 ;
      RECT 54.43 6.745 55.87 6.915 ;
      RECT 54.43 2.395 54.59 6.915 ;
      RECT 54.745 2.365 55.065 2.685 ;
      RECT 54.43 2.395 55.065 2.565 ;
      RECT 47.31 4.135 53.4 4.325 ;
      RECT 53.23 3.145 53.4 4.325 ;
      RECT 53.21 3.15 53.4 4.325 ;
      RECT 47.31 3.515 47.48 4.325 ;
      RECT 47.255 3.515 47.535 3.885 ;
      RECT 47.325 3.07 47.465 4.325 ;
      RECT 53.14 3.15 53.48 3.5 ;
      RECT 47.135 2.955 47.415 3.325 ;
      RECT 46.845 3.07 47.465 3.21 ;
      RECT 46.845 1.86 46.985 3.21 ;
      RECT 46.785 1.86 47.045 2.18 ;
      RECT 39.365 6.66 39.715 7.01 ;
      RECT 50.105 6.615 50.455 6.965 ;
      RECT 39.365 6.69 50.455 6.89 ;
      RECT 49.745 2.98 50.005 3.3 ;
      RECT 49.805 1.86 49.945 3.3 ;
      RECT 49.745 1.86 50.005 2.18 ;
      RECT 48.745 3.54 49.005 3.86 ;
      RECT 48.745 2.955 48.945 3.86 ;
      RECT 48.685 1.86 48.825 3.49 ;
      RECT 48.685 2.955 49.185 3.325 ;
      RECT 48.625 1.86 48.885 2.18 ;
      RECT 48.265 3.54 48.525 3.86 ;
      RECT 48.325 1.95 48.465 3.86 ;
      RECT 48.025 1.95 48.465 2.18 ;
      RECT 48.025 1.86 48.285 2.18 ;
      RECT 47.785 2.42 48.045 2.74 ;
      RECT 47.205 2.51 48.045 2.65 ;
      RECT 47.205 1.57 47.345 2.65 ;
      RECT 43.865 1.86 44.125 2.18 ;
      RECT 43.865 1.95 44.905 2.09 ;
      RECT 44.765 1.57 44.905 2.09 ;
      RECT 44.765 1.57 47.345 1.71 ;
      RECT 46.055 2.955 46.335 3.325 ;
      RECT 46.125 1.86 46.265 3.325 ;
      RECT 46.065 1.86 46.325 2.18 ;
      RECT 45.705 3.54 45.965 3.86 ;
      RECT 45.765 1.95 45.905 3.86 ;
      RECT 45.345 1.86 45.605 2.18 ;
      RECT 45.345 1.95 45.905 2.09 ;
      RECT 43.375 2.955 43.655 3.325 ;
      RECT 45.345 2.98 45.605 3.3 ;
      RECT 43.025 2.98 43.655 3.3 ;
      RECT 43.025 3.07 45.605 3.21 ;
      RECT 44.815 2.395 45.095 2.765 ;
      RECT 44.815 2.42 45.345 2.74 ;
      RECT 41.905 2.98 42.165 3.3 ;
      RECT 41.965 1.86 42.105 3.3 ;
      RECT 41.905 1.86 42.165 2.18 ;
      RECT 40.935 3.515 41.215 3.885 ;
      RECT 40.945 3.26 41.205 3.885 ;
      RECT 36.185 6.22 36.505 6.545 ;
      RECT 36.215 5.695 36.385 6.545 ;
      RECT 36.215 5.695 36.39 6.045 ;
      RECT 36.215 5.695 37.19 5.87 ;
      RECT 37.015 1.965 37.19 5.87 ;
      RECT 36.96 1.965 37.31 2.315 ;
      RECT 36.985 6.655 37.31 6.98 ;
      RECT 35.87 6.745 37.31 6.915 ;
      RECT 35.87 2.395 36.03 6.915 ;
      RECT 36.185 2.365 36.505 2.685 ;
      RECT 35.87 2.395 36.505 2.565 ;
      RECT 28.75 4.135 34.84 4.325 ;
      RECT 34.67 3.145 34.84 4.325 ;
      RECT 34.65 3.15 34.84 4.325 ;
      RECT 28.75 3.515 28.92 4.325 ;
      RECT 28.695 3.515 28.975 3.885 ;
      RECT 28.765 3.07 28.905 4.325 ;
      RECT 34.58 3.15 34.92 3.5 ;
      RECT 28.575 2.955 28.855 3.325 ;
      RECT 28.285 3.07 28.905 3.21 ;
      RECT 28.285 1.86 28.425 3.21 ;
      RECT 28.225 1.86 28.485 2.18 ;
      RECT 20.805 6.655 21.155 7.005 ;
      RECT 31.55 6.61 31.9 6.96 ;
      RECT 20.805 6.685 31.9 6.885 ;
      RECT 31.185 2.98 31.445 3.3 ;
      RECT 31.245 1.86 31.385 3.3 ;
      RECT 31.185 1.86 31.445 2.18 ;
      RECT 30.185 3.54 30.445 3.86 ;
      RECT 30.185 2.955 30.385 3.86 ;
      RECT 30.125 1.86 30.265 3.49 ;
      RECT 30.125 2.955 30.625 3.325 ;
      RECT 30.065 1.86 30.325 2.18 ;
      RECT 29.705 3.54 29.965 3.86 ;
      RECT 29.765 1.95 29.905 3.86 ;
      RECT 29.465 1.95 29.905 2.18 ;
      RECT 29.465 1.86 29.725 2.18 ;
      RECT 29.225 2.42 29.485 2.74 ;
      RECT 28.645 2.51 29.485 2.65 ;
      RECT 28.645 1.57 28.785 2.65 ;
      RECT 25.305 1.86 25.565 2.18 ;
      RECT 25.305 1.95 26.345 2.09 ;
      RECT 26.205 1.57 26.345 2.09 ;
      RECT 26.205 1.57 28.785 1.71 ;
      RECT 27.495 2.955 27.775 3.325 ;
      RECT 27.565 1.86 27.705 3.325 ;
      RECT 27.505 1.86 27.765 2.18 ;
      RECT 27.145 3.54 27.405 3.86 ;
      RECT 27.205 1.95 27.345 3.86 ;
      RECT 26.785 1.86 27.045 2.18 ;
      RECT 26.785 1.95 27.345 2.09 ;
      RECT 24.815 2.955 25.095 3.325 ;
      RECT 26.785 2.98 27.045 3.3 ;
      RECT 24.465 2.98 25.095 3.3 ;
      RECT 24.465 3.07 27.045 3.21 ;
      RECT 26.255 2.395 26.535 2.765 ;
      RECT 26.255 2.42 26.785 2.74 ;
      RECT 23.345 2.98 23.605 3.3 ;
      RECT 23.405 1.86 23.545 3.3 ;
      RECT 23.345 1.86 23.605 2.18 ;
      RECT 22.375 3.515 22.655 3.885 ;
      RECT 22.385 3.26 22.645 3.885 ;
      RECT 17.625 6.22 17.945 6.545 ;
      RECT 17.655 5.695 17.825 6.545 ;
      RECT 17.655 5.695 17.83 6.045 ;
      RECT 17.655 5.695 18.63 5.87 ;
      RECT 18.455 1.965 18.63 5.87 ;
      RECT 18.4 1.965 18.75 2.315 ;
      RECT 18.425 6.655 18.75 6.98 ;
      RECT 17.31 6.745 18.75 6.915 ;
      RECT 17.31 2.395 17.47 6.915 ;
      RECT 17.625 2.365 17.945 2.685 ;
      RECT 17.31 2.395 17.945 2.565 ;
      RECT 10.19 4.135 16.28 4.325 ;
      RECT 16.11 3.145 16.28 4.325 ;
      RECT 16.09 3.15 16.28 4.325 ;
      RECT 10.19 3.515 10.36 4.325 ;
      RECT 10.135 3.515 10.415 3.885 ;
      RECT 10.205 3.07 10.345 4.325 ;
      RECT 16.02 3.15 16.36 3.5 ;
      RECT 10.015 2.955 10.295 3.325 ;
      RECT 9.725 3.07 10.345 3.21 ;
      RECT 9.725 1.86 9.865 3.21 ;
      RECT 9.665 1.86 9.925 2.18 ;
      RECT 1.54 6.995 1.83 7.345 ;
      RECT 1.54 7.055 2.73 7.225 ;
      RECT 2.56 6.685 2.73 7.225 ;
      RECT 12.99 6.605 13.34 6.955 ;
      RECT 2.56 6.685 13.34 6.855 ;
      RECT 12.625 2.98 12.885 3.3 ;
      RECT 12.685 1.86 12.825 3.3 ;
      RECT 12.625 1.86 12.885 2.18 ;
      RECT 11.625 3.54 11.885 3.86 ;
      RECT 11.625 2.955 11.825 3.86 ;
      RECT 11.565 1.86 11.705 3.49 ;
      RECT 11.565 2.955 12.065 3.325 ;
      RECT 11.505 1.86 11.765 2.18 ;
      RECT 11.145 3.54 11.405 3.86 ;
      RECT 11.205 1.95 11.345 3.86 ;
      RECT 10.905 1.95 11.345 2.18 ;
      RECT 10.905 1.86 11.165 2.18 ;
      RECT 10.665 2.42 10.925 2.74 ;
      RECT 10.085 2.51 10.925 2.65 ;
      RECT 10.085 1.57 10.225 2.65 ;
      RECT 6.745 1.86 7.005 2.18 ;
      RECT 6.745 1.95 7.785 2.09 ;
      RECT 7.645 1.57 7.785 2.09 ;
      RECT 7.645 1.57 10.225 1.71 ;
      RECT 8.935 2.955 9.215 3.325 ;
      RECT 9.005 1.86 9.145 3.325 ;
      RECT 8.945 1.86 9.205 2.18 ;
      RECT 8.585 3.54 8.845 3.86 ;
      RECT 8.645 1.95 8.785 3.86 ;
      RECT 8.225 1.86 8.485 2.18 ;
      RECT 8.225 1.95 8.785 2.09 ;
      RECT 6.255 2.955 6.535 3.325 ;
      RECT 8.225 2.98 8.485 3.3 ;
      RECT 5.905 2.98 6.535 3.3 ;
      RECT 5.905 3.07 8.485 3.21 ;
      RECT 7.695 2.395 7.975 2.765 ;
      RECT 7.695 2.42 8.225 2.74 ;
      RECT 4.785 2.98 5.045 3.3 ;
      RECT 4.845 1.86 4.985 3.3 ;
      RECT 4.785 1.86 5.045 2.18 ;
      RECT 3.815 3.515 4.095 3.885 ;
      RECT 3.825 3.26 4.085 3.885 ;
      RECT 88.295 1.835 88.575 2.205 ;
      RECT 87.335 3.515 87.615 3.885 ;
      RECT 86.555 7.055 86.93 7.425 ;
      RECT 86.335 3.515 86.615 3.885 ;
      RECT 78.535 2.395 78.815 2.765 ;
      RECT 69.735 1.835 70.015 2.205 ;
      RECT 68.775 3.515 69.055 3.885 ;
      RECT 67.995 7.055 68.37 7.425 ;
      RECT 67.775 3.515 68.055 3.885 ;
      RECT 59.975 2.395 60.255 2.765 ;
      RECT 51.175 1.835 51.455 2.205 ;
      RECT 50.215 3.515 50.495 3.885 ;
      RECT 49.435 7.055 49.81 7.425 ;
      RECT 49.215 3.515 49.495 3.885 ;
      RECT 41.415 2.395 41.695 2.765 ;
      RECT 32.615 1.835 32.895 2.205 ;
      RECT 31.655 3.515 31.935 3.885 ;
      RECT 30.875 7.055 31.25 7.425 ;
      RECT 30.655 3.515 30.935 3.885 ;
      RECT 22.855 2.395 23.135 2.765 ;
      RECT 14.055 1.835 14.335 2.205 ;
      RECT 13.095 3.515 13.375 3.885 ;
      RECT 12.315 7.055 12.69 7.425 ;
      RECT 12.095 3.515 12.375 3.885 ;
      RECT 4.295 2.395 4.575 2.765 ;
    LAYER via1 ;
      RECT 95.125 7.375 95.275 7.525 ;
      RECT 92.755 6.74 92.905 6.89 ;
      RECT 92.74 2.065 92.89 2.215 ;
      RECT 91.95 2.45 92.1 2.6 ;
      RECT 91.95 6.325 92.1 6.475 ;
      RECT 90.36 3.25 90.51 3.4 ;
      RECT 88.36 1.945 88.51 2.095 ;
      RECT 87.4 3.625 87.55 3.775 ;
      RECT 87.325 6.71 87.475 6.86 ;
      RECT 86.92 1.945 87.07 2.095 ;
      RECT 86.92 3.065 87.07 3.215 ;
      RECT 86.665 7.165 86.815 7.315 ;
      RECT 86.4 3.625 86.55 3.775 ;
      RECT 85.92 3.625 86.07 3.775 ;
      RECT 85.8 1.945 85.95 2.095 ;
      RECT 85.44 3.625 85.59 3.775 ;
      RECT 85.2 1.945 85.35 2.095 ;
      RECT 84.96 2.505 85.11 2.655 ;
      RECT 84.44 3.625 84.59 3.775 ;
      RECT 83.96 1.945 84.11 2.095 ;
      RECT 83.24 1.945 83.39 2.095 ;
      RECT 83.24 3.065 83.39 3.215 ;
      RECT 82.88 3.625 83.03 3.775 ;
      RECT 82.52 1.945 82.67 2.095 ;
      RECT 82.52 3.065 82.67 3.215 ;
      RECT 82.26 2.505 82.41 2.655 ;
      RECT 81.04 1.945 81.19 2.095 ;
      RECT 80.2 3.065 80.35 3.215 ;
      RECT 79.08 1.945 79.23 2.095 ;
      RECT 79.08 3.065 79.23 3.215 ;
      RECT 78.6 2.505 78.75 2.655 ;
      RECT 78.12 3.345 78.27 3.495 ;
      RECT 76.54 6.755 76.69 6.905 ;
      RECT 74.195 6.74 74.345 6.89 ;
      RECT 74.18 2.065 74.33 2.215 ;
      RECT 73.39 2.45 73.54 2.6 ;
      RECT 73.39 6.325 73.54 6.475 ;
      RECT 71.8 3.25 71.95 3.4 ;
      RECT 69.8 1.945 69.95 2.095 ;
      RECT 68.84 3.625 68.99 3.775 ;
      RECT 68.765 6.71 68.915 6.86 ;
      RECT 68.36 1.945 68.51 2.095 ;
      RECT 68.36 3.065 68.51 3.215 ;
      RECT 68.105 7.165 68.255 7.315 ;
      RECT 67.84 3.625 67.99 3.775 ;
      RECT 67.36 3.625 67.51 3.775 ;
      RECT 67.24 1.945 67.39 2.095 ;
      RECT 66.88 3.625 67.03 3.775 ;
      RECT 66.64 1.945 66.79 2.095 ;
      RECT 66.4 2.505 66.55 2.655 ;
      RECT 65.88 3.625 66.03 3.775 ;
      RECT 65.4 1.945 65.55 2.095 ;
      RECT 64.68 1.945 64.83 2.095 ;
      RECT 64.68 3.065 64.83 3.215 ;
      RECT 64.32 3.625 64.47 3.775 ;
      RECT 63.96 1.945 64.11 2.095 ;
      RECT 63.96 3.065 64.11 3.215 ;
      RECT 63.7 2.505 63.85 2.655 ;
      RECT 62.48 1.945 62.63 2.095 ;
      RECT 61.64 3.065 61.79 3.215 ;
      RECT 60.52 1.945 60.67 2.095 ;
      RECT 60.52 3.065 60.67 3.215 ;
      RECT 60.04 2.505 60.19 2.655 ;
      RECT 59.56 3.345 59.71 3.495 ;
      RECT 57.98 6.755 58.13 6.905 ;
      RECT 55.635 6.74 55.785 6.89 ;
      RECT 55.62 2.065 55.77 2.215 ;
      RECT 54.83 2.45 54.98 2.6 ;
      RECT 54.83 6.325 54.98 6.475 ;
      RECT 53.24 3.25 53.39 3.4 ;
      RECT 51.24 1.945 51.39 2.095 ;
      RECT 50.28 3.625 50.43 3.775 ;
      RECT 50.205 6.715 50.355 6.865 ;
      RECT 49.8 1.945 49.95 2.095 ;
      RECT 49.8 3.065 49.95 3.215 ;
      RECT 49.545 7.165 49.695 7.315 ;
      RECT 49.28 3.625 49.43 3.775 ;
      RECT 48.8 3.625 48.95 3.775 ;
      RECT 48.68 1.945 48.83 2.095 ;
      RECT 48.32 3.625 48.47 3.775 ;
      RECT 48.08 1.945 48.23 2.095 ;
      RECT 47.84 2.505 47.99 2.655 ;
      RECT 47.32 3.625 47.47 3.775 ;
      RECT 46.84 1.945 46.99 2.095 ;
      RECT 46.12 1.945 46.27 2.095 ;
      RECT 46.12 3.065 46.27 3.215 ;
      RECT 45.76 3.625 45.91 3.775 ;
      RECT 45.4 1.945 45.55 2.095 ;
      RECT 45.4 3.065 45.55 3.215 ;
      RECT 45.14 2.505 45.29 2.655 ;
      RECT 43.92 1.945 44.07 2.095 ;
      RECT 43.08 3.065 43.23 3.215 ;
      RECT 41.96 1.945 42.11 2.095 ;
      RECT 41.96 3.065 42.11 3.215 ;
      RECT 41.48 2.505 41.63 2.655 ;
      RECT 41 3.345 41.15 3.495 ;
      RECT 39.465 6.76 39.615 6.91 ;
      RECT 37.075 6.74 37.225 6.89 ;
      RECT 37.06 2.065 37.21 2.215 ;
      RECT 36.27 2.45 36.42 2.6 ;
      RECT 36.27 6.325 36.42 6.475 ;
      RECT 34.68 3.25 34.83 3.4 ;
      RECT 32.68 1.945 32.83 2.095 ;
      RECT 31.72 3.625 31.87 3.775 ;
      RECT 31.65 6.71 31.8 6.86 ;
      RECT 31.24 1.945 31.39 2.095 ;
      RECT 31.24 3.065 31.39 3.215 ;
      RECT 30.985 7.165 31.135 7.315 ;
      RECT 30.72 3.625 30.87 3.775 ;
      RECT 30.24 3.625 30.39 3.775 ;
      RECT 30.12 1.945 30.27 2.095 ;
      RECT 29.76 3.625 29.91 3.775 ;
      RECT 29.52 1.945 29.67 2.095 ;
      RECT 29.28 2.505 29.43 2.655 ;
      RECT 28.76 3.625 28.91 3.775 ;
      RECT 28.28 1.945 28.43 2.095 ;
      RECT 27.56 1.945 27.71 2.095 ;
      RECT 27.56 3.065 27.71 3.215 ;
      RECT 27.2 3.625 27.35 3.775 ;
      RECT 26.84 1.945 26.99 2.095 ;
      RECT 26.84 3.065 26.99 3.215 ;
      RECT 26.58 2.505 26.73 2.655 ;
      RECT 25.36 1.945 25.51 2.095 ;
      RECT 24.52 3.065 24.67 3.215 ;
      RECT 23.4 1.945 23.55 2.095 ;
      RECT 23.4 3.065 23.55 3.215 ;
      RECT 22.92 2.505 23.07 2.655 ;
      RECT 22.44 3.345 22.59 3.495 ;
      RECT 20.905 6.755 21.055 6.905 ;
      RECT 18.515 6.74 18.665 6.89 ;
      RECT 18.5 2.065 18.65 2.215 ;
      RECT 17.71 2.45 17.86 2.6 ;
      RECT 17.71 6.325 17.86 6.475 ;
      RECT 16.12 3.25 16.27 3.4 ;
      RECT 14.12 1.945 14.27 2.095 ;
      RECT 13.16 3.625 13.31 3.775 ;
      RECT 13.09 6.705 13.24 6.855 ;
      RECT 12.68 1.945 12.83 2.095 ;
      RECT 12.68 3.065 12.83 3.215 ;
      RECT 12.425 7.165 12.575 7.315 ;
      RECT 12.16 3.625 12.31 3.775 ;
      RECT 11.68 3.625 11.83 3.775 ;
      RECT 11.56 1.945 11.71 2.095 ;
      RECT 11.2 3.625 11.35 3.775 ;
      RECT 10.96 1.945 11.11 2.095 ;
      RECT 10.72 2.505 10.87 2.655 ;
      RECT 10.2 3.625 10.35 3.775 ;
      RECT 9.72 1.945 9.87 2.095 ;
      RECT 9 1.945 9.15 2.095 ;
      RECT 9 3.065 9.15 3.215 ;
      RECT 8.64 3.625 8.79 3.775 ;
      RECT 8.28 1.945 8.43 2.095 ;
      RECT 8.28 3.065 8.43 3.215 ;
      RECT 8.02 2.505 8.17 2.655 ;
      RECT 6.8 1.945 6.95 2.095 ;
      RECT 5.96 3.065 6.11 3.215 ;
      RECT 4.84 1.945 4.99 2.095 ;
      RECT 4.84 3.065 4.99 3.215 ;
      RECT 4.36 2.505 4.51 2.655 ;
      RECT 3.88 3.345 4.03 3.495 ;
      RECT 1.61 7.095 1.76 7.245 ;
      RECT 1.235 6.355 1.385 6.505 ;
    LAYER met1 ;
      RECT 94.99 7.77 95.28 8 ;
      RECT 95.05 6.29 95.22 8 ;
      RECT 95.025 7.275 95.375 7.625 ;
      RECT 94.99 6.29 95.28 6.52 ;
      RECT 94.585 2.395 94.69 2.965 ;
      RECT 94.585 2.73 94.91 2.96 ;
      RECT 94.585 2.76 95.08 2.93 ;
      RECT 94.585 2.395 94.775 2.96 ;
      RECT 94 2.36 94.29 2.59 ;
      RECT 94 2.395 94.775 2.565 ;
      RECT 94.06 0.88 94.23 2.59 ;
      RECT 94 0.88 94.29 1.11 ;
      RECT 94 7.77 94.29 8 ;
      RECT 94.06 6.29 94.23 8 ;
      RECT 94 6.29 94.29 6.52 ;
      RECT 94 6.325 94.855 6.485 ;
      RECT 94.685 5.92 94.855 6.485 ;
      RECT 94 6.32 94.395 6.485 ;
      RECT 94.62 5.92 94.91 6.15 ;
      RECT 94.62 5.95 95.08 6.12 ;
      RECT 93.63 2.73 93.92 2.96 ;
      RECT 93.63 2.76 94.09 2.93 ;
      RECT 93.695 1.655 93.86 2.96 ;
      RECT 92.21 1.625 92.5 1.855 ;
      RECT 92.21 1.655 93.86 1.825 ;
      RECT 92.27 0.885 92.44 1.855 ;
      RECT 92.21 0.885 92.5 1.115 ;
      RECT 92.21 7.765 92.5 7.995 ;
      RECT 92.27 7.025 92.44 7.995 ;
      RECT 92.27 7.12 93.86 7.29 ;
      RECT 93.69 5.92 93.86 7.29 ;
      RECT 92.21 7.025 92.5 7.255 ;
      RECT 93.63 5.92 93.92 6.15 ;
      RECT 93.63 5.95 94.09 6.12 ;
      RECT 90.26 3.15 90.6 3.5 ;
      RECT 90.35 2.025 90.52 3.5 ;
      RECT 92.64 1.965 92.99 2.315 ;
      RECT 90.35 2.025 92.99 2.195 ;
      RECT 92.665 6.655 92.99 6.98 ;
      RECT 87.225 6.61 87.575 6.96 ;
      RECT 92.64 6.655 92.99 6.885 ;
      RECT 87.025 6.655 87.575 6.885 ;
      RECT 86.855 6.685 92.99 6.855 ;
      RECT 91.865 2.365 92.185 2.685 ;
      RECT 91.835 2.365 92.185 2.595 ;
      RECT 91.665 2.395 92.185 2.565 ;
      RECT 91.865 6.255 92.185 6.545 ;
      RECT 91.835 6.285 92.185 6.515 ;
      RECT 91.665 6.315 92.185 6.485 ;
      RECT 87.315 3.57 87.635 3.83 ;
      RECT 88.605 2.745 88.745 3.605 ;
      RECT 87.405 3.465 88.745 3.605 ;
      RECT 87.405 3.025 87.545 3.83 ;
      RECT 87.33 3.025 87.62 3.255 ;
      RECT 88.53 2.745 88.82 2.975 ;
      RECT 88.05 3.025 88.34 3.255 ;
      RECT 88.245 1.95 88.385 3.21 ;
      RECT 88.275 1.89 88.595 2.15 ;
      RECT 84.875 2.45 85.195 2.71 ;
      RECT 87.57 2.465 87.86 2.695 ;
      RECT 84.965 2.37 87.785 2.51 ;
      RECT 86.835 1.89 87.155 2.15 ;
      RECT 87.33 1.905 87.62 2.135 ;
      RECT 86.835 1.95 87.62 2.09 ;
      RECT 86.835 3.01 87.155 3.27 ;
      RECT 86.835 2.79 87.065 3.27 ;
      RECT 86.33 2.745 86.62 2.975 ;
      RECT 86.33 2.79 87.065 2.93 ;
      RECT 86.595 7.765 86.885 7.995 ;
      RECT 86.655 7.025 86.825 7.995 ;
      RECT 86.555 7.055 86.935 7.425 ;
      RECT 86.595 7.025 86.885 7.425 ;
      RECT 85.355 3.57 85.675 3.83 ;
      RECT 84.89 3.585 85.18 3.815 ;
      RECT 84.89 3.63 85.675 3.77 ;
      RECT 83.65 2.465 83.94 2.695 ;
      RECT 83.65 2.51 84.585 2.65 ;
      RECT 84.445 1.95 84.585 2.65 ;
      RECT 85.115 1.89 85.435 2.15 ;
      RECT 84.89 1.905 85.435 2.135 ;
      RECT 84.445 1.95 85.435 2.09 ;
      RECT 82.795 3.57 83.115 3.83 ;
      RECT 82.795 3.63 83.865 3.77 ;
      RECT 83.725 3.07 83.865 3.77 ;
      RECT 84.89 3.025 85.18 3.255 ;
      RECT 83.725 3.07 85.18 3.21 ;
      RECT 83.155 1.89 83.475 2.15 ;
      RECT 82.93 1.905 83.475 2.135 ;
      RECT 82.175 2.45 82.495 2.71 ;
      RECT 83.17 2.465 83.46 2.695 ;
      RECT 81.93 2.465 82.495 2.695 ;
      RECT 81.93 2.51 83.46 2.65 ;
      RECT 81.45 3.025 81.74 3.255 ;
      RECT 81.645 1.95 81.785 3.21 ;
      RECT 82.435 1.89 82.755 2.15 ;
      RECT 81.45 1.905 81.74 2.135 ;
      RECT 81.45 1.95 82.755 2.09 ;
      RECT 81.045 3.465 82.145 3.605 ;
      RECT 81.93 3.305 82.22 3.535 ;
      RECT 80.97 3.305 81.26 3.535 ;
      RECT 80.955 1.89 81.275 2.15 ;
      RECT 78.995 1.89 79.315 2.15 ;
      RECT 78.995 1.95 81.275 2.09 ;
      RECT 80.115 3.01 80.435 3.27 ;
      RECT 80.115 3.01 80.945 3.15 ;
      RECT 80.73 2.745 80.945 3.15 ;
      RECT 80.73 2.745 81.02 2.975 ;
      RECT 78.515 2.45 78.835 2.71 ;
      RECT 79.925 2.465 80.215 2.695 ;
      RECT 78.515 2.465 79.06 2.695 ;
      RECT 78.515 2.55 79.465 2.69 ;
      RECT 79.325 2.37 79.465 2.69 ;
      RECT 79.825 2.465 80.215 2.65 ;
      RECT 79.325 2.37 79.965 2.51 ;
      RECT 78.035 3.26 78.355 3.675 ;
      RECT 78.115 1.905 78.27 3.675 ;
      RECT 78.05 1.905 78.34 2.135 ;
      RECT 76.43 7.77 76.72 8 ;
      RECT 76.49 6.29 76.66 8 ;
      RECT 76.44 6.655 76.79 7.005 ;
      RECT 76.43 6.29 76.72 6.52 ;
      RECT 76.025 2.395 76.13 2.965 ;
      RECT 76.025 2.73 76.35 2.96 ;
      RECT 76.025 2.76 76.52 2.93 ;
      RECT 76.025 2.395 76.215 2.96 ;
      RECT 75.44 2.36 75.73 2.59 ;
      RECT 75.44 2.395 76.215 2.565 ;
      RECT 75.5 0.88 75.67 2.59 ;
      RECT 75.44 0.88 75.73 1.11 ;
      RECT 75.44 7.77 75.73 8 ;
      RECT 75.5 6.29 75.67 8 ;
      RECT 75.44 6.29 75.73 6.52 ;
      RECT 75.44 6.325 76.295 6.485 ;
      RECT 76.125 5.92 76.295 6.485 ;
      RECT 75.44 6.32 75.835 6.485 ;
      RECT 76.06 5.92 76.35 6.15 ;
      RECT 76.06 5.95 76.52 6.12 ;
      RECT 75.07 2.73 75.36 2.96 ;
      RECT 75.07 2.76 75.53 2.93 ;
      RECT 75.135 1.655 75.3 2.96 ;
      RECT 73.65 1.625 73.94 1.855 ;
      RECT 73.65 1.655 75.3 1.825 ;
      RECT 73.71 0.885 73.88 1.855 ;
      RECT 73.65 0.885 73.94 1.115 ;
      RECT 73.65 7.765 73.94 7.995 ;
      RECT 73.71 7.025 73.88 7.995 ;
      RECT 73.71 7.12 75.3 7.29 ;
      RECT 75.13 5.92 75.3 7.29 ;
      RECT 73.65 7.025 73.94 7.255 ;
      RECT 75.07 5.92 75.36 6.15 ;
      RECT 75.07 5.95 75.53 6.12 ;
      RECT 71.7 3.15 72.04 3.5 ;
      RECT 71.79 2.025 71.96 3.5 ;
      RECT 74.08 1.965 74.43 2.315 ;
      RECT 71.79 2.025 74.43 2.195 ;
      RECT 74.105 6.655 74.43 6.98 ;
      RECT 68.665 6.61 69.015 6.96 ;
      RECT 74.08 6.655 74.43 6.885 ;
      RECT 68.465 6.655 69.015 6.885 ;
      RECT 68.295 6.685 74.43 6.855 ;
      RECT 73.305 2.365 73.625 2.685 ;
      RECT 73.275 2.365 73.625 2.595 ;
      RECT 73.105 2.395 73.625 2.565 ;
      RECT 73.305 6.255 73.625 6.545 ;
      RECT 73.275 6.285 73.625 6.515 ;
      RECT 73.105 6.315 73.625 6.485 ;
      RECT 68.755 3.57 69.075 3.83 ;
      RECT 70.045 2.745 70.185 3.605 ;
      RECT 68.845 3.465 70.185 3.605 ;
      RECT 68.845 3.025 68.985 3.83 ;
      RECT 68.77 3.025 69.06 3.255 ;
      RECT 69.97 2.745 70.26 2.975 ;
      RECT 69.49 3.025 69.78 3.255 ;
      RECT 69.685 1.95 69.825 3.21 ;
      RECT 69.715 1.89 70.035 2.15 ;
      RECT 66.315 2.45 66.635 2.71 ;
      RECT 69.01 2.465 69.3 2.695 ;
      RECT 66.405 2.37 69.225 2.51 ;
      RECT 68.275 1.89 68.595 2.15 ;
      RECT 68.77 1.905 69.06 2.135 ;
      RECT 68.275 1.95 69.06 2.09 ;
      RECT 68.275 3.01 68.595 3.27 ;
      RECT 68.275 2.79 68.505 3.27 ;
      RECT 67.77 2.745 68.06 2.975 ;
      RECT 67.77 2.79 68.505 2.93 ;
      RECT 68.035 7.765 68.325 7.995 ;
      RECT 68.095 7.025 68.265 7.995 ;
      RECT 67.995 7.055 68.375 7.425 ;
      RECT 68.035 7.025 68.325 7.425 ;
      RECT 66.795 3.57 67.115 3.83 ;
      RECT 66.33 3.585 66.62 3.815 ;
      RECT 66.33 3.63 67.115 3.77 ;
      RECT 65.09 2.465 65.38 2.695 ;
      RECT 65.09 2.51 66.025 2.65 ;
      RECT 65.885 1.95 66.025 2.65 ;
      RECT 66.555 1.89 66.875 2.15 ;
      RECT 66.33 1.905 66.875 2.135 ;
      RECT 65.885 1.95 66.875 2.09 ;
      RECT 64.235 3.57 64.555 3.83 ;
      RECT 64.235 3.63 65.305 3.77 ;
      RECT 65.165 3.07 65.305 3.77 ;
      RECT 66.33 3.025 66.62 3.255 ;
      RECT 65.165 3.07 66.62 3.21 ;
      RECT 64.595 1.89 64.915 2.15 ;
      RECT 64.37 1.905 64.915 2.135 ;
      RECT 63.615 2.45 63.935 2.71 ;
      RECT 64.61 2.465 64.9 2.695 ;
      RECT 63.37 2.465 63.935 2.695 ;
      RECT 63.37 2.51 64.9 2.65 ;
      RECT 62.89 3.025 63.18 3.255 ;
      RECT 63.085 1.95 63.225 3.21 ;
      RECT 63.875 1.89 64.195 2.15 ;
      RECT 62.89 1.905 63.18 2.135 ;
      RECT 62.89 1.95 64.195 2.09 ;
      RECT 62.485 3.465 63.585 3.605 ;
      RECT 63.37 3.305 63.66 3.535 ;
      RECT 62.41 3.305 62.7 3.535 ;
      RECT 62.395 1.89 62.715 2.15 ;
      RECT 60.435 1.89 60.755 2.15 ;
      RECT 60.435 1.95 62.715 2.09 ;
      RECT 61.555 3.01 61.875 3.27 ;
      RECT 61.555 3.01 62.385 3.15 ;
      RECT 62.17 2.745 62.385 3.15 ;
      RECT 62.17 2.745 62.46 2.975 ;
      RECT 59.955 2.45 60.275 2.71 ;
      RECT 61.365 2.465 61.655 2.695 ;
      RECT 59.955 2.465 60.5 2.695 ;
      RECT 59.955 2.55 60.905 2.69 ;
      RECT 60.765 2.37 60.905 2.69 ;
      RECT 61.265 2.465 61.655 2.65 ;
      RECT 60.765 2.37 61.405 2.51 ;
      RECT 59.475 3.26 59.795 3.675 ;
      RECT 59.555 1.905 59.71 3.675 ;
      RECT 59.49 1.905 59.78 2.135 ;
      RECT 57.87 7.77 58.16 8 ;
      RECT 57.93 6.29 58.1 8 ;
      RECT 57.88 6.655 58.23 7.005 ;
      RECT 57.87 6.29 58.16 6.52 ;
      RECT 57.465 2.395 57.57 2.965 ;
      RECT 57.465 2.73 57.79 2.96 ;
      RECT 57.465 2.76 57.96 2.93 ;
      RECT 57.465 2.395 57.655 2.96 ;
      RECT 56.88 2.36 57.17 2.59 ;
      RECT 56.88 2.395 57.655 2.565 ;
      RECT 56.94 0.88 57.11 2.59 ;
      RECT 56.88 0.88 57.17 1.11 ;
      RECT 56.88 7.77 57.17 8 ;
      RECT 56.94 6.29 57.11 8 ;
      RECT 56.88 6.29 57.17 6.52 ;
      RECT 56.88 6.325 57.735 6.485 ;
      RECT 57.565 5.92 57.735 6.485 ;
      RECT 56.88 6.32 57.275 6.485 ;
      RECT 57.5 5.92 57.79 6.15 ;
      RECT 57.5 5.95 57.96 6.12 ;
      RECT 56.51 2.73 56.8 2.96 ;
      RECT 56.51 2.76 56.97 2.93 ;
      RECT 56.575 1.655 56.74 2.96 ;
      RECT 55.09 1.625 55.38 1.855 ;
      RECT 55.09 1.655 56.74 1.825 ;
      RECT 55.15 0.885 55.32 1.855 ;
      RECT 55.09 0.885 55.38 1.115 ;
      RECT 55.09 7.765 55.38 7.995 ;
      RECT 55.15 7.025 55.32 7.995 ;
      RECT 55.15 7.12 56.74 7.29 ;
      RECT 56.57 5.92 56.74 7.29 ;
      RECT 55.09 7.025 55.38 7.255 ;
      RECT 56.51 5.92 56.8 6.15 ;
      RECT 56.51 5.95 56.97 6.12 ;
      RECT 53.14 3.15 53.48 3.5 ;
      RECT 53.23 2.025 53.4 3.5 ;
      RECT 55.52 1.965 55.87 2.315 ;
      RECT 53.23 2.025 55.87 2.195 ;
      RECT 55.545 6.655 55.87 6.98 ;
      RECT 50.105 6.615 50.455 6.965 ;
      RECT 55.52 6.655 55.87 6.885 ;
      RECT 49.905 6.655 50.455 6.885 ;
      RECT 49.735 6.685 55.87 6.855 ;
      RECT 54.745 2.365 55.065 2.685 ;
      RECT 54.715 2.365 55.065 2.595 ;
      RECT 54.545 2.395 55.065 2.565 ;
      RECT 54.745 6.255 55.065 6.545 ;
      RECT 54.715 6.285 55.065 6.515 ;
      RECT 54.545 6.315 55.065 6.485 ;
      RECT 50.195 3.57 50.515 3.83 ;
      RECT 51.485 2.745 51.625 3.605 ;
      RECT 50.285 3.465 51.625 3.605 ;
      RECT 50.285 3.025 50.425 3.83 ;
      RECT 50.21 3.025 50.5 3.255 ;
      RECT 51.41 2.745 51.7 2.975 ;
      RECT 50.93 3.025 51.22 3.255 ;
      RECT 51.125 1.95 51.265 3.21 ;
      RECT 51.155 1.89 51.475 2.15 ;
      RECT 47.755 2.45 48.075 2.71 ;
      RECT 50.45 2.465 50.74 2.695 ;
      RECT 47.845 2.37 50.665 2.51 ;
      RECT 49.715 1.89 50.035 2.15 ;
      RECT 50.21 1.905 50.5 2.135 ;
      RECT 49.715 1.95 50.5 2.09 ;
      RECT 49.715 3.01 50.035 3.27 ;
      RECT 49.715 2.79 49.945 3.27 ;
      RECT 49.21 2.745 49.5 2.975 ;
      RECT 49.21 2.79 49.945 2.93 ;
      RECT 49.475 7.765 49.765 7.995 ;
      RECT 49.535 7.025 49.705 7.995 ;
      RECT 49.435 7.055 49.815 7.425 ;
      RECT 49.475 7.025 49.765 7.425 ;
      RECT 48.235 3.57 48.555 3.83 ;
      RECT 47.77 3.585 48.06 3.815 ;
      RECT 47.77 3.63 48.555 3.77 ;
      RECT 46.53 2.465 46.82 2.695 ;
      RECT 46.53 2.51 47.465 2.65 ;
      RECT 47.325 1.95 47.465 2.65 ;
      RECT 47.995 1.89 48.315 2.15 ;
      RECT 47.77 1.905 48.315 2.135 ;
      RECT 47.325 1.95 48.315 2.09 ;
      RECT 45.675 3.57 45.995 3.83 ;
      RECT 45.675 3.63 46.745 3.77 ;
      RECT 46.605 3.07 46.745 3.77 ;
      RECT 47.77 3.025 48.06 3.255 ;
      RECT 46.605 3.07 48.06 3.21 ;
      RECT 46.035 1.89 46.355 2.15 ;
      RECT 45.81 1.905 46.355 2.135 ;
      RECT 45.055 2.45 45.375 2.71 ;
      RECT 46.05 2.465 46.34 2.695 ;
      RECT 44.81 2.465 45.375 2.695 ;
      RECT 44.81 2.51 46.34 2.65 ;
      RECT 44.33 3.025 44.62 3.255 ;
      RECT 44.525 1.95 44.665 3.21 ;
      RECT 45.315 1.89 45.635 2.15 ;
      RECT 44.33 1.905 44.62 2.135 ;
      RECT 44.33 1.95 45.635 2.09 ;
      RECT 43.925 3.465 45.025 3.605 ;
      RECT 44.81 3.305 45.1 3.535 ;
      RECT 43.85 3.305 44.14 3.535 ;
      RECT 43.835 1.89 44.155 2.15 ;
      RECT 41.875 1.89 42.195 2.15 ;
      RECT 41.875 1.95 44.155 2.09 ;
      RECT 42.995 3.01 43.315 3.27 ;
      RECT 42.995 3.01 43.825 3.15 ;
      RECT 43.61 2.745 43.825 3.15 ;
      RECT 43.61 2.745 43.9 2.975 ;
      RECT 41.395 2.45 41.715 2.71 ;
      RECT 42.805 2.465 43.095 2.695 ;
      RECT 41.395 2.465 41.94 2.695 ;
      RECT 41.395 2.55 42.345 2.69 ;
      RECT 42.205 2.37 42.345 2.69 ;
      RECT 42.705 2.465 43.095 2.65 ;
      RECT 42.205 2.37 42.845 2.51 ;
      RECT 40.915 3.26 41.235 3.675 ;
      RECT 40.995 1.905 41.15 3.675 ;
      RECT 40.93 1.905 41.22 2.135 ;
      RECT 39.31 7.77 39.6 8 ;
      RECT 39.37 6.29 39.54 8 ;
      RECT 39.36 6.66 39.715 7.015 ;
      RECT 39.31 6.29 39.6 6.52 ;
      RECT 38.905 2.395 39.01 2.965 ;
      RECT 38.905 2.73 39.23 2.96 ;
      RECT 38.905 2.76 39.4 2.93 ;
      RECT 38.905 2.395 39.095 2.96 ;
      RECT 38.32 2.36 38.61 2.59 ;
      RECT 38.32 2.395 39.095 2.565 ;
      RECT 38.38 0.88 38.55 2.59 ;
      RECT 38.32 0.88 38.61 1.11 ;
      RECT 38.32 7.77 38.61 8 ;
      RECT 38.38 6.29 38.55 8 ;
      RECT 38.32 6.29 38.61 6.52 ;
      RECT 38.32 6.325 39.175 6.485 ;
      RECT 39.005 5.92 39.175 6.485 ;
      RECT 38.32 6.32 38.715 6.485 ;
      RECT 38.94 5.92 39.23 6.15 ;
      RECT 38.94 5.95 39.4 6.12 ;
      RECT 37.95 2.73 38.24 2.96 ;
      RECT 37.95 2.76 38.41 2.93 ;
      RECT 38.015 1.655 38.18 2.96 ;
      RECT 36.53 1.625 36.82 1.855 ;
      RECT 36.53 1.655 38.18 1.825 ;
      RECT 36.59 0.885 36.76 1.855 ;
      RECT 36.53 0.885 36.82 1.115 ;
      RECT 36.53 7.765 36.82 7.995 ;
      RECT 36.59 7.025 36.76 7.995 ;
      RECT 36.59 7.12 38.18 7.29 ;
      RECT 38.01 5.92 38.18 7.29 ;
      RECT 36.53 7.025 36.82 7.255 ;
      RECT 37.95 5.92 38.24 6.15 ;
      RECT 37.95 5.95 38.41 6.12 ;
      RECT 34.58 3.15 34.92 3.5 ;
      RECT 34.67 2.025 34.84 3.5 ;
      RECT 36.96 1.965 37.31 2.315 ;
      RECT 34.67 2.025 37.31 2.195 ;
      RECT 36.985 6.655 37.31 6.98 ;
      RECT 31.55 6.61 31.9 6.96 ;
      RECT 36.96 6.655 37.31 6.885 ;
      RECT 31.345 6.655 31.9 6.885 ;
      RECT 31.175 6.685 37.31 6.855 ;
      RECT 36.185 2.365 36.505 2.685 ;
      RECT 36.155 2.365 36.505 2.595 ;
      RECT 35.985 2.395 36.505 2.565 ;
      RECT 36.185 6.255 36.505 6.545 ;
      RECT 36.155 6.285 36.505 6.515 ;
      RECT 35.985 6.315 36.505 6.485 ;
      RECT 31.635 3.57 31.955 3.83 ;
      RECT 32.925 2.745 33.065 3.605 ;
      RECT 31.725 3.465 33.065 3.605 ;
      RECT 31.725 3.025 31.865 3.83 ;
      RECT 31.65 3.025 31.94 3.255 ;
      RECT 32.85 2.745 33.14 2.975 ;
      RECT 32.37 3.025 32.66 3.255 ;
      RECT 32.565 1.95 32.705 3.21 ;
      RECT 32.595 1.89 32.915 2.15 ;
      RECT 29.195 2.45 29.515 2.71 ;
      RECT 31.89 2.465 32.18 2.695 ;
      RECT 29.285 2.37 32.105 2.51 ;
      RECT 31.155 1.89 31.475 2.15 ;
      RECT 31.65 1.905 31.94 2.135 ;
      RECT 31.155 1.95 31.94 2.09 ;
      RECT 31.155 3.01 31.475 3.27 ;
      RECT 31.155 2.79 31.385 3.27 ;
      RECT 30.65 2.745 30.94 2.975 ;
      RECT 30.65 2.79 31.385 2.93 ;
      RECT 30.915 7.765 31.205 7.995 ;
      RECT 30.975 7.025 31.145 7.995 ;
      RECT 30.875 7.055 31.255 7.425 ;
      RECT 30.915 7.025 31.205 7.425 ;
      RECT 29.675 3.57 29.995 3.83 ;
      RECT 29.21 3.585 29.5 3.815 ;
      RECT 29.21 3.63 29.995 3.77 ;
      RECT 27.97 2.465 28.26 2.695 ;
      RECT 27.97 2.51 28.905 2.65 ;
      RECT 28.765 1.95 28.905 2.65 ;
      RECT 29.435 1.89 29.755 2.15 ;
      RECT 29.21 1.905 29.755 2.135 ;
      RECT 28.765 1.95 29.755 2.09 ;
      RECT 27.115 3.57 27.435 3.83 ;
      RECT 27.115 3.63 28.185 3.77 ;
      RECT 28.045 3.07 28.185 3.77 ;
      RECT 29.21 3.025 29.5 3.255 ;
      RECT 28.045 3.07 29.5 3.21 ;
      RECT 27.475 1.89 27.795 2.15 ;
      RECT 27.25 1.905 27.795 2.135 ;
      RECT 26.495 2.45 26.815 2.71 ;
      RECT 27.49 2.465 27.78 2.695 ;
      RECT 26.25 2.465 26.815 2.695 ;
      RECT 26.25 2.51 27.78 2.65 ;
      RECT 25.77 3.025 26.06 3.255 ;
      RECT 25.965 1.95 26.105 3.21 ;
      RECT 26.755 1.89 27.075 2.15 ;
      RECT 25.77 1.905 26.06 2.135 ;
      RECT 25.77 1.95 27.075 2.09 ;
      RECT 25.365 3.465 26.465 3.605 ;
      RECT 26.25 3.305 26.54 3.535 ;
      RECT 25.29 3.305 25.58 3.535 ;
      RECT 25.275 1.89 25.595 2.15 ;
      RECT 23.315 1.89 23.635 2.15 ;
      RECT 23.315 1.95 25.595 2.09 ;
      RECT 24.435 3.01 24.755 3.27 ;
      RECT 24.435 3.01 25.265 3.15 ;
      RECT 25.05 2.745 25.265 3.15 ;
      RECT 25.05 2.745 25.34 2.975 ;
      RECT 22.835 2.45 23.155 2.71 ;
      RECT 24.245 2.465 24.535 2.695 ;
      RECT 22.835 2.465 23.38 2.695 ;
      RECT 22.835 2.55 23.785 2.69 ;
      RECT 23.645 2.37 23.785 2.69 ;
      RECT 24.145 2.465 24.535 2.65 ;
      RECT 23.645 2.37 24.285 2.51 ;
      RECT 22.355 3.26 22.675 3.675 ;
      RECT 22.435 1.905 22.59 3.675 ;
      RECT 22.37 1.905 22.66 2.135 ;
      RECT 20.75 7.77 21.04 8 ;
      RECT 20.81 6.29 20.98 8 ;
      RECT 20.805 6.655 21.155 7.005 ;
      RECT 20.75 6.29 21.04 6.52 ;
      RECT 20.345 2.395 20.45 2.965 ;
      RECT 20.345 2.73 20.67 2.96 ;
      RECT 20.345 2.76 20.84 2.93 ;
      RECT 20.345 2.395 20.535 2.96 ;
      RECT 19.76 2.36 20.05 2.59 ;
      RECT 19.76 2.395 20.535 2.565 ;
      RECT 19.82 0.88 19.99 2.59 ;
      RECT 19.76 0.88 20.05 1.11 ;
      RECT 19.76 7.77 20.05 8 ;
      RECT 19.82 6.29 19.99 8 ;
      RECT 19.76 6.29 20.05 6.52 ;
      RECT 19.76 6.325 20.615 6.485 ;
      RECT 20.445 5.92 20.615 6.485 ;
      RECT 19.76 6.32 20.155 6.485 ;
      RECT 20.38 5.92 20.67 6.15 ;
      RECT 20.38 5.95 20.84 6.12 ;
      RECT 19.39 2.73 19.68 2.96 ;
      RECT 19.39 2.76 19.85 2.93 ;
      RECT 19.455 1.655 19.62 2.96 ;
      RECT 17.97 1.625 18.26 1.855 ;
      RECT 17.97 1.655 19.62 1.825 ;
      RECT 18.03 0.885 18.2 1.855 ;
      RECT 17.97 0.885 18.26 1.115 ;
      RECT 17.97 7.765 18.26 7.995 ;
      RECT 18.03 7.025 18.2 7.995 ;
      RECT 18.03 7.12 19.62 7.29 ;
      RECT 19.45 5.92 19.62 7.29 ;
      RECT 17.97 7.025 18.26 7.255 ;
      RECT 19.39 5.92 19.68 6.15 ;
      RECT 19.39 5.95 19.85 6.12 ;
      RECT 16.02 3.15 16.36 3.5 ;
      RECT 16.11 2.025 16.28 3.5 ;
      RECT 18.4 1.965 18.75 2.315 ;
      RECT 16.11 2.025 18.75 2.195 ;
      RECT 18.425 6.655 18.75 6.98 ;
      RECT 12.99 6.605 13.34 6.955 ;
      RECT 18.4 6.655 18.75 6.885 ;
      RECT 12.785 6.655 13.34 6.885 ;
      RECT 12.615 6.685 18.75 6.855 ;
      RECT 17.625 2.365 17.945 2.685 ;
      RECT 17.595 2.365 17.945 2.595 ;
      RECT 17.425 2.395 17.945 2.565 ;
      RECT 17.625 6.255 17.945 6.545 ;
      RECT 17.595 6.285 17.945 6.515 ;
      RECT 17.425 6.315 17.945 6.485 ;
      RECT 13.075 3.57 13.395 3.83 ;
      RECT 14.365 2.745 14.505 3.605 ;
      RECT 13.165 3.465 14.505 3.605 ;
      RECT 13.165 3.025 13.305 3.83 ;
      RECT 13.09 3.025 13.38 3.255 ;
      RECT 14.29 2.745 14.58 2.975 ;
      RECT 13.81 3.025 14.1 3.255 ;
      RECT 14.005 1.95 14.145 3.21 ;
      RECT 14.035 1.89 14.355 2.15 ;
      RECT 10.635 2.45 10.955 2.71 ;
      RECT 13.33 2.465 13.62 2.695 ;
      RECT 10.725 2.37 13.545 2.51 ;
      RECT 12.595 1.89 12.915 2.15 ;
      RECT 13.09 1.905 13.38 2.135 ;
      RECT 12.595 1.95 13.38 2.09 ;
      RECT 12.595 3.01 12.915 3.27 ;
      RECT 12.595 2.79 12.825 3.27 ;
      RECT 12.09 2.745 12.38 2.975 ;
      RECT 12.09 2.79 12.825 2.93 ;
      RECT 12.355 7.765 12.645 7.995 ;
      RECT 12.415 7.025 12.585 7.995 ;
      RECT 12.315 7.055 12.695 7.425 ;
      RECT 12.355 7.025 12.645 7.425 ;
      RECT 11.115 3.57 11.435 3.83 ;
      RECT 10.65 3.585 10.94 3.815 ;
      RECT 10.65 3.63 11.435 3.77 ;
      RECT 9.41 2.465 9.7 2.695 ;
      RECT 9.41 2.51 10.345 2.65 ;
      RECT 10.205 1.95 10.345 2.65 ;
      RECT 10.875 1.89 11.195 2.15 ;
      RECT 10.65 1.905 11.195 2.135 ;
      RECT 10.205 1.95 11.195 2.09 ;
      RECT 8.555 3.57 8.875 3.83 ;
      RECT 8.555 3.63 9.625 3.77 ;
      RECT 9.485 3.07 9.625 3.77 ;
      RECT 10.65 3.025 10.94 3.255 ;
      RECT 9.485 3.07 10.94 3.21 ;
      RECT 8.915 1.89 9.235 2.15 ;
      RECT 8.69 1.905 9.235 2.135 ;
      RECT 7.935 2.45 8.255 2.71 ;
      RECT 8.93 2.465 9.22 2.695 ;
      RECT 7.69 2.465 8.255 2.695 ;
      RECT 7.69 2.51 9.22 2.65 ;
      RECT 7.21 3.025 7.5 3.255 ;
      RECT 7.405 1.95 7.545 3.21 ;
      RECT 8.195 1.89 8.515 2.15 ;
      RECT 7.21 1.905 7.5 2.135 ;
      RECT 7.21 1.95 8.515 2.09 ;
      RECT 6.805 3.465 7.905 3.605 ;
      RECT 7.69 3.305 7.98 3.535 ;
      RECT 6.73 3.305 7.02 3.535 ;
      RECT 6.715 1.89 7.035 2.15 ;
      RECT 4.755 1.89 5.075 2.15 ;
      RECT 4.755 1.95 7.035 2.09 ;
      RECT 5.875 3.01 6.195 3.27 ;
      RECT 5.875 3.01 6.705 3.15 ;
      RECT 6.49 2.745 6.705 3.15 ;
      RECT 6.49 2.745 6.78 2.975 ;
      RECT 4.275 2.45 4.595 2.71 ;
      RECT 5.685 2.465 5.975 2.695 ;
      RECT 4.275 2.465 4.82 2.695 ;
      RECT 4.275 2.55 5.225 2.69 ;
      RECT 5.085 2.37 5.225 2.69 ;
      RECT 5.585 2.465 5.975 2.65 ;
      RECT 5.085 2.37 5.725 2.51 ;
      RECT 3.795 3.26 4.115 3.675 ;
      RECT 3.875 1.905 4.03 3.675 ;
      RECT 3.81 1.905 4.1 2.135 ;
      RECT 1.54 7.765 1.83 7.995 ;
      RECT 1.6 7.025 1.77 7.995 ;
      RECT 1.51 7.025 1.86 7.315 ;
      RECT 1.135 6.285 1.485 6.575 ;
      RECT 0.995 6.315 1.485 6.485 ;
      RECT 86.315 3.57 86.635 3.83 ;
      RECT 85.715 1.89 86.395 2.15 ;
      RECT 85.835 3.57 86.155 3.83 ;
      RECT 84.355 3.57 84.675 3.83 ;
      RECT 83.875 1.89 84.195 2.15 ;
      RECT 83.155 3.01 83.475 3.27 ;
      RECT 82.435 3.01 82.755 3.27 ;
      RECT 78.995 3.01 79.315 3.27 ;
      RECT 67.755 3.57 68.075 3.83 ;
      RECT 67.155 1.89 67.835 2.15 ;
      RECT 67.275 3.57 67.595 3.83 ;
      RECT 65.795 3.57 66.115 3.83 ;
      RECT 65.315 1.89 65.635 2.15 ;
      RECT 64.595 3.01 64.915 3.27 ;
      RECT 63.875 3.01 64.195 3.27 ;
      RECT 60.435 3.01 60.755 3.27 ;
      RECT 49.195 3.57 49.515 3.83 ;
      RECT 48.595 1.89 49.275 2.15 ;
      RECT 48.715 3.57 49.035 3.83 ;
      RECT 47.235 3.57 47.555 3.83 ;
      RECT 46.755 1.89 47.075 2.15 ;
      RECT 46.035 3.01 46.355 3.27 ;
      RECT 45.315 3.01 45.635 3.27 ;
      RECT 41.875 3.01 42.195 3.27 ;
      RECT 30.635 3.57 30.955 3.83 ;
      RECT 30.035 1.89 30.715 2.15 ;
      RECT 30.155 3.57 30.475 3.83 ;
      RECT 28.675 3.57 28.995 3.83 ;
      RECT 28.195 1.89 28.515 2.15 ;
      RECT 27.475 3.01 27.795 3.27 ;
      RECT 26.755 3.01 27.075 3.27 ;
      RECT 23.315 3.01 23.635 3.27 ;
      RECT 12.075 3.57 12.395 3.83 ;
      RECT 11.475 1.89 12.155 2.15 ;
      RECT 11.595 3.57 11.915 3.83 ;
      RECT 10.115 3.57 10.435 3.83 ;
      RECT 9.635 1.89 9.955 2.15 ;
      RECT 8.915 3.01 9.235 3.27 ;
      RECT 8.195 3.01 8.515 3.27 ;
      RECT 4.755 3.01 5.075 3.27 ;
    LAYER mcon ;
      RECT 95.05 6.32 95.22 6.49 ;
      RECT 95.055 6.315 95.225 6.485 ;
      RECT 76.49 6.32 76.66 6.49 ;
      RECT 76.495 6.315 76.665 6.485 ;
      RECT 57.93 6.32 58.1 6.49 ;
      RECT 57.935 6.315 58.105 6.485 ;
      RECT 39.37 6.32 39.54 6.49 ;
      RECT 39.375 6.315 39.545 6.485 ;
      RECT 20.81 6.32 20.98 6.49 ;
      RECT 20.815 6.315 20.985 6.485 ;
      RECT 95.05 7.8 95.22 7.97 ;
      RECT 94.68 2.76 94.85 2.93 ;
      RECT 94.68 5.95 94.85 6.12 ;
      RECT 94.06 0.91 94.23 1.08 ;
      RECT 94.06 2.39 94.23 2.56 ;
      RECT 94.06 6.32 94.23 6.49 ;
      RECT 94.06 7.8 94.23 7.97 ;
      RECT 93.69 2.76 93.86 2.93 ;
      RECT 93.69 5.95 93.86 6.12 ;
      RECT 92.7 2.025 92.87 2.195 ;
      RECT 92.7 6.685 92.87 6.855 ;
      RECT 92.27 0.915 92.44 1.085 ;
      RECT 92.27 1.655 92.44 1.825 ;
      RECT 92.27 7.055 92.44 7.225 ;
      RECT 92.27 7.795 92.44 7.965 ;
      RECT 91.895 2.395 92.065 2.565 ;
      RECT 91.895 6.315 92.065 6.485 ;
      RECT 88.59 2.775 88.76 2.945 ;
      RECT 88.35 1.935 88.52 2.105 ;
      RECT 88.11 3.055 88.28 3.225 ;
      RECT 87.63 2.495 87.8 2.665 ;
      RECT 87.39 1.935 87.56 2.105 ;
      RECT 87.39 3.055 87.56 3.225 ;
      RECT 87.39 3.615 87.56 3.785 ;
      RECT 87.085 6.685 87.255 6.855 ;
      RECT 86.91 3.055 87.08 3.225 ;
      RECT 86.655 7.055 86.825 7.225 ;
      RECT 86.655 7.795 86.825 7.965 ;
      RECT 86.39 2.775 86.56 2.945 ;
      RECT 86.39 3.615 86.56 3.785 ;
      RECT 85.91 1.935 86.08 2.105 ;
      RECT 85.91 3.615 86.08 3.785 ;
      RECT 84.95 1.935 85.12 2.105 ;
      RECT 84.95 2.495 85.12 2.665 ;
      RECT 84.95 3.055 85.12 3.225 ;
      RECT 84.95 3.615 85.12 3.785 ;
      RECT 84.43 3.615 84.6 3.785 ;
      RECT 83.95 1.935 84.12 2.105 ;
      RECT 83.71 2.495 83.88 2.665 ;
      RECT 83.23 2.495 83.4 2.665 ;
      RECT 83.23 3.055 83.4 3.225 ;
      RECT 82.99 1.935 83.16 2.105 ;
      RECT 82.51 3.055 82.68 3.225 ;
      RECT 81.99 2.495 82.16 2.665 ;
      RECT 81.99 3.335 82.16 3.505 ;
      RECT 81.51 1.935 81.68 2.105 ;
      RECT 81.51 3.055 81.68 3.225 ;
      RECT 81.03 3.335 81.2 3.505 ;
      RECT 80.79 2.775 80.96 2.945 ;
      RECT 79.985 2.495 80.155 2.665 ;
      RECT 79.07 1.935 79.24 2.105 ;
      RECT 79.07 3.055 79.24 3.225 ;
      RECT 78.83 2.495 79 2.665 ;
      RECT 78.11 1.935 78.28 2.105 ;
      RECT 78.11 3.475 78.28 3.645 ;
      RECT 76.49 7.8 76.66 7.97 ;
      RECT 76.12 2.76 76.29 2.93 ;
      RECT 76.12 5.95 76.29 6.12 ;
      RECT 75.5 0.91 75.67 1.08 ;
      RECT 75.5 2.39 75.67 2.56 ;
      RECT 75.5 6.32 75.67 6.49 ;
      RECT 75.5 7.8 75.67 7.97 ;
      RECT 75.13 2.76 75.3 2.93 ;
      RECT 75.13 5.95 75.3 6.12 ;
      RECT 74.14 2.025 74.31 2.195 ;
      RECT 74.14 6.685 74.31 6.855 ;
      RECT 73.71 0.915 73.88 1.085 ;
      RECT 73.71 1.655 73.88 1.825 ;
      RECT 73.71 7.055 73.88 7.225 ;
      RECT 73.71 7.795 73.88 7.965 ;
      RECT 73.335 2.395 73.505 2.565 ;
      RECT 73.335 6.315 73.505 6.485 ;
      RECT 70.03 2.775 70.2 2.945 ;
      RECT 69.79 1.935 69.96 2.105 ;
      RECT 69.55 3.055 69.72 3.225 ;
      RECT 69.07 2.495 69.24 2.665 ;
      RECT 68.83 1.935 69 2.105 ;
      RECT 68.83 3.055 69 3.225 ;
      RECT 68.83 3.615 69 3.785 ;
      RECT 68.525 6.685 68.695 6.855 ;
      RECT 68.35 3.055 68.52 3.225 ;
      RECT 68.095 7.055 68.265 7.225 ;
      RECT 68.095 7.795 68.265 7.965 ;
      RECT 67.83 2.775 68 2.945 ;
      RECT 67.83 3.615 68 3.785 ;
      RECT 67.35 1.935 67.52 2.105 ;
      RECT 67.35 3.615 67.52 3.785 ;
      RECT 66.39 1.935 66.56 2.105 ;
      RECT 66.39 2.495 66.56 2.665 ;
      RECT 66.39 3.055 66.56 3.225 ;
      RECT 66.39 3.615 66.56 3.785 ;
      RECT 65.87 3.615 66.04 3.785 ;
      RECT 65.39 1.935 65.56 2.105 ;
      RECT 65.15 2.495 65.32 2.665 ;
      RECT 64.67 2.495 64.84 2.665 ;
      RECT 64.67 3.055 64.84 3.225 ;
      RECT 64.43 1.935 64.6 2.105 ;
      RECT 63.95 3.055 64.12 3.225 ;
      RECT 63.43 2.495 63.6 2.665 ;
      RECT 63.43 3.335 63.6 3.505 ;
      RECT 62.95 1.935 63.12 2.105 ;
      RECT 62.95 3.055 63.12 3.225 ;
      RECT 62.47 3.335 62.64 3.505 ;
      RECT 62.23 2.775 62.4 2.945 ;
      RECT 61.425 2.495 61.595 2.665 ;
      RECT 60.51 1.935 60.68 2.105 ;
      RECT 60.51 3.055 60.68 3.225 ;
      RECT 60.27 2.495 60.44 2.665 ;
      RECT 59.55 1.935 59.72 2.105 ;
      RECT 59.55 3.475 59.72 3.645 ;
      RECT 57.93 7.8 58.1 7.97 ;
      RECT 57.56 2.76 57.73 2.93 ;
      RECT 57.56 5.95 57.73 6.12 ;
      RECT 56.94 0.91 57.11 1.08 ;
      RECT 56.94 2.39 57.11 2.56 ;
      RECT 56.94 6.32 57.11 6.49 ;
      RECT 56.94 7.8 57.11 7.97 ;
      RECT 56.57 2.76 56.74 2.93 ;
      RECT 56.57 5.95 56.74 6.12 ;
      RECT 55.58 2.025 55.75 2.195 ;
      RECT 55.58 6.685 55.75 6.855 ;
      RECT 55.15 0.915 55.32 1.085 ;
      RECT 55.15 1.655 55.32 1.825 ;
      RECT 55.15 7.055 55.32 7.225 ;
      RECT 55.15 7.795 55.32 7.965 ;
      RECT 54.775 2.395 54.945 2.565 ;
      RECT 54.775 6.315 54.945 6.485 ;
      RECT 51.47 2.775 51.64 2.945 ;
      RECT 51.23 1.935 51.4 2.105 ;
      RECT 50.99 3.055 51.16 3.225 ;
      RECT 50.51 2.495 50.68 2.665 ;
      RECT 50.27 1.935 50.44 2.105 ;
      RECT 50.27 3.055 50.44 3.225 ;
      RECT 50.27 3.615 50.44 3.785 ;
      RECT 49.965 6.685 50.135 6.855 ;
      RECT 49.79 3.055 49.96 3.225 ;
      RECT 49.535 7.055 49.705 7.225 ;
      RECT 49.535 7.795 49.705 7.965 ;
      RECT 49.27 2.775 49.44 2.945 ;
      RECT 49.27 3.615 49.44 3.785 ;
      RECT 48.79 1.935 48.96 2.105 ;
      RECT 48.79 3.615 48.96 3.785 ;
      RECT 47.83 1.935 48 2.105 ;
      RECT 47.83 2.495 48 2.665 ;
      RECT 47.83 3.055 48 3.225 ;
      RECT 47.83 3.615 48 3.785 ;
      RECT 47.31 3.615 47.48 3.785 ;
      RECT 46.83 1.935 47 2.105 ;
      RECT 46.59 2.495 46.76 2.665 ;
      RECT 46.11 2.495 46.28 2.665 ;
      RECT 46.11 3.055 46.28 3.225 ;
      RECT 45.87 1.935 46.04 2.105 ;
      RECT 45.39 3.055 45.56 3.225 ;
      RECT 44.87 2.495 45.04 2.665 ;
      RECT 44.87 3.335 45.04 3.505 ;
      RECT 44.39 1.935 44.56 2.105 ;
      RECT 44.39 3.055 44.56 3.225 ;
      RECT 43.91 3.335 44.08 3.505 ;
      RECT 43.67 2.775 43.84 2.945 ;
      RECT 42.865 2.495 43.035 2.665 ;
      RECT 41.95 1.935 42.12 2.105 ;
      RECT 41.95 3.055 42.12 3.225 ;
      RECT 41.71 2.495 41.88 2.665 ;
      RECT 40.99 1.935 41.16 2.105 ;
      RECT 40.99 3.475 41.16 3.645 ;
      RECT 39.37 7.8 39.54 7.97 ;
      RECT 39 2.76 39.17 2.93 ;
      RECT 39 5.95 39.17 6.12 ;
      RECT 38.38 0.91 38.55 1.08 ;
      RECT 38.38 2.39 38.55 2.56 ;
      RECT 38.38 6.32 38.55 6.49 ;
      RECT 38.38 7.8 38.55 7.97 ;
      RECT 38.01 2.76 38.18 2.93 ;
      RECT 38.01 5.95 38.18 6.12 ;
      RECT 37.02 2.025 37.19 2.195 ;
      RECT 37.02 6.685 37.19 6.855 ;
      RECT 36.59 0.915 36.76 1.085 ;
      RECT 36.59 1.655 36.76 1.825 ;
      RECT 36.59 7.055 36.76 7.225 ;
      RECT 36.59 7.795 36.76 7.965 ;
      RECT 36.215 2.395 36.385 2.565 ;
      RECT 36.215 6.315 36.385 6.485 ;
      RECT 32.91 2.775 33.08 2.945 ;
      RECT 32.67 1.935 32.84 2.105 ;
      RECT 32.43 3.055 32.6 3.225 ;
      RECT 31.95 2.495 32.12 2.665 ;
      RECT 31.71 1.935 31.88 2.105 ;
      RECT 31.71 3.055 31.88 3.225 ;
      RECT 31.71 3.615 31.88 3.785 ;
      RECT 31.405 6.685 31.575 6.855 ;
      RECT 31.23 3.055 31.4 3.225 ;
      RECT 30.975 7.055 31.145 7.225 ;
      RECT 30.975 7.795 31.145 7.965 ;
      RECT 30.71 2.775 30.88 2.945 ;
      RECT 30.71 3.615 30.88 3.785 ;
      RECT 30.23 1.935 30.4 2.105 ;
      RECT 30.23 3.615 30.4 3.785 ;
      RECT 29.27 1.935 29.44 2.105 ;
      RECT 29.27 2.495 29.44 2.665 ;
      RECT 29.27 3.055 29.44 3.225 ;
      RECT 29.27 3.615 29.44 3.785 ;
      RECT 28.75 3.615 28.92 3.785 ;
      RECT 28.27 1.935 28.44 2.105 ;
      RECT 28.03 2.495 28.2 2.665 ;
      RECT 27.55 2.495 27.72 2.665 ;
      RECT 27.55 3.055 27.72 3.225 ;
      RECT 27.31 1.935 27.48 2.105 ;
      RECT 26.83 3.055 27 3.225 ;
      RECT 26.31 2.495 26.48 2.665 ;
      RECT 26.31 3.335 26.48 3.505 ;
      RECT 25.83 1.935 26 2.105 ;
      RECT 25.83 3.055 26 3.225 ;
      RECT 25.35 3.335 25.52 3.505 ;
      RECT 25.11 2.775 25.28 2.945 ;
      RECT 24.305 2.495 24.475 2.665 ;
      RECT 23.39 1.935 23.56 2.105 ;
      RECT 23.39 3.055 23.56 3.225 ;
      RECT 23.15 2.495 23.32 2.665 ;
      RECT 22.43 1.935 22.6 2.105 ;
      RECT 22.43 3.475 22.6 3.645 ;
      RECT 20.81 7.8 20.98 7.97 ;
      RECT 20.44 2.76 20.61 2.93 ;
      RECT 20.44 5.95 20.61 6.12 ;
      RECT 19.82 0.91 19.99 1.08 ;
      RECT 19.82 2.39 19.99 2.56 ;
      RECT 19.82 6.32 19.99 6.49 ;
      RECT 19.82 7.8 19.99 7.97 ;
      RECT 19.45 2.76 19.62 2.93 ;
      RECT 19.45 5.95 19.62 6.12 ;
      RECT 18.46 2.025 18.63 2.195 ;
      RECT 18.46 6.685 18.63 6.855 ;
      RECT 18.03 0.915 18.2 1.085 ;
      RECT 18.03 1.655 18.2 1.825 ;
      RECT 18.03 7.055 18.2 7.225 ;
      RECT 18.03 7.795 18.2 7.965 ;
      RECT 17.655 2.395 17.825 2.565 ;
      RECT 17.655 6.315 17.825 6.485 ;
      RECT 14.35 2.775 14.52 2.945 ;
      RECT 14.11 1.935 14.28 2.105 ;
      RECT 13.87 3.055 14.04 3.225 ;
      RECT 13.39 2.495 13.56 2.665 ;
      RECT 13.15 1.935 13.32 2.105 ;
      RECT 13.15 3.055 13.32 3.225 ;
      RECT 13.15 3.615 13.32 3.785 ;
      RECT 12.845 6.685 13.015 6.855 ;
      RECT 12.67 3.055 12.84 3.225 ;
      RECT 12.415 7.055 12.585 7.225 ;
      RECT 12.415 7.795 12.585 7.965 ;
      RECT 12.15 2.775 12.32 2.945 ;
      RECT 12.15 3.615 12.32 3.785 ;
      RECT 11.67 1.935 11.84 2.105 ;
      RECT 11.67 3.615 11.84 3.785 ;
      RECT 10.71 1.935 10.88 2.105 ;
      RECT 10.71 2.495 10.88 2.665 ;
      RECT 10.71 3.055 10.88 3.225 ;
      RECT 10.71 3.615 10.88 3.785 ;
      RECT 10.19 3.615 10.36 3.785 ;
      RECT 9.71 1.935 9.88 2.105 ;
      RECT 9.47 2.495 9.64 2.665 ;
      RECT 8.99 2.495 9.16 2.665 ;
      RECT 8.99 3.055 9.16 3.225 ;
      RECT 8.75 1.935 8.92 2.105 ;
      RECT 8.27 3.055 8.44 3.225 ;
      RECT 7.75 2.495 7.92 2.665 ;
      RECT 7.75 3.335 7.92 3.505 ;
      RECT 7.27 1.935 7.44 2.105 ;
      RECT 7.27 3.055 7.44 3.225 ;
      RECT 6.79 3.335 6.96 3.505 ;
      RECT 6.55 2.775 6.72 2.945 ;
      RECT 5.745 2.495 5.915 2.665 ;
      RECT 4.83 1.935 5 2.105 ;
      RECT 4.83 3.055 5 3.225 ;
      RECT 4.59 2.495 4.76 2.665 ;
      RECT 3.87 1.935 4.04 2.105 ;
      RECT 3.87 3.475 4.04 3.645 ;
      RECT 1.6 7.055 1.77 7.225 ;
      RECT 1.6 7.795 1.77 7.965 ;
      RECT 1.225 6.315 1.395 6.485 ;
    LAYER li1 ;
      RECT 95.05 5.02 95.22 6.49 ;
      RECT 95.05 6.315 95.225 6.485 ;
      RECT 94.68 1.74 94.85 2.93 ;
      RECT 94.68 1.74 95.15 1.91 ;
      RECT 94.68 6.97 95.15 7.14 ;
      RECT 94.68 5.95 94.85 7.14 ;
      RECT 93.69 1.74 93.86 2.93 ;
      RECT 93.69 1.74 94.16 1.91 ;
      RECT 93.69 6.97 94.16 7.14 ;
      RECT 93.69 5.95 93.86 7.14 ;
      RECT 91.84 2.635 92.01 3.865 ;
      RECT 91.895 0.855 92.065 2.805 ;
      RECT 91.84 0.575 92.01 1.025 ;
      RECT 91.84 7.855 92.01 8.305 ;
      RECT 91.895 6.075 92.065 8.025 ;
      RECT 91.84 5.015 92.01 6.245 ;
      RECT 91.32 0.575 91.49 3.865 ;
      RECT 91.32 2.075 91.725 2.405 ;
      RECT 91.32 1.235 91.725 1.565 ;
      RECT 91.32 5.015 91.49 8.305 ;
      RECT 91.32 7.315 91.725 7.645 ;
      RECT 91.32 6.475 91.725 6.805 ;
      RECT 88.11 3.225 89.08 3.395 ;
      RECT 88.11 3.055 88.28 3.395 ;
      RECT 87.63 2.495 87.8 2.825 ;
      RECT 87.63 2.575 88.36 2.745 ;
      RECT 87.27 3.615 87.56 3.785 ;
      RECT 87.27 2.575 87.44 3.785 ;
      RECT 87.27 3.055 87.56 3.225 ;
      RECT 87.07 2.575 87.44 2.745 ;
      RECT 86.39 2.675 86.56 2.945 ;
      RECT 86.15 2.675 86.56 2.845 ;
      RECT 86.07 2.575 86.4 2.745 ;
      RECT 85.91 3.615 86.56 3.785 ;
      RECT 86.39 3.145 86.56 3.785 ;
      RECT 86.27 3.225 86.56 3.785 ;
      RECT 85.705 5.015 85.875 8.305 ;
      RECT 85.705 7.315 86.11 7.645 ;
      RECT 85.705 6.475 86.11 6.805 ;
      RECT 84.95 2.915 85.12 3.225 ;
      RECT 84.95 2.915 85.84 3.085 ;
      RECT 85.67 2.495 85.84 3.085 ;
      RECT 84.95 2.575 85.44 2.745 ;
      RECT 84.95 2.495 85.12 2.745 ;
      RECT 82.91 3.225 83.4 3.395 ;
      RECT 84.07 2.575 84.24 3.225 ;
      RECT 83.23 3.055 84.24 3.225 ;
      RECT 84.19 2.495 84.36 2.825 ;
      RECT 82.99 1.835 83.16 2.105 ;
      RECT 82.43 1.835 83.16 2.005 ;
      RECT 82.51 2.575 82.68 3.225 ;
      RECT 82.51 2.575 83 2.745 ;
      RECT 81.67 2.575 82.16 2.745 ;
      RECT 81.99 2.495 82.16 2.745 ;
      RECT 81.51 1.835 81.68 2.105 ;
      RECT 80.95 1.835 81.68 2.005 ;
      RECT 81.03 3.225 81.2 3.505 ;
      RECT 79.99 3.225 81.28 3.395 ;
      RECT 79.985 2.575 80.56 2.745 ;
      RECT 79.985 2.495 80.155 2.745 ;
      RECT 79.07 1.835 79.24 2.105 ;
      RECT 79.07 1.835 79.8 2.005 ;
      RECT 79.07 3.055 79.24 3.475 ;
      RECT 78.45 3.14 79.24 3.31 ;
      RECT 78.45 2.915 78.62 3.31 ;
      RECT 78.35 2.495 78.52 3.085 ;
      RECT 78.11 2.575 78.52 2.845 ;
      RECT 76.49 5.02 76.66 6.49 ;
      RECT 76.49 6.315 76.665 6.485 ;
      RECT 76.12 1.74 76.29 2.93 ;
      RECT 76.12 1.74 76.59 1.91 ;
      RECT 76.12 6.97 76.59 7.14 ;
      RECT 76.12 5.95 76.29 7.14 ;
      RECT 75.13 1.74 75.3 2.93 ;
      RECT 75.13 1.74 75.6 1.91 ;
      RECT 75.13 6.97 75.6 7.14 ;
      RECT 75.13 5.95 75.3 7.14 ;
      RECT 73.28 2.635 73.45 3.865 ;
      RECT 73.335 0.855 73.505 2.805 ;
      RECT 73.28 0.575 73.45 1.025 ;
      RECT 73.28 7.855 73.45 8.305 ;
      RECT 73.335 6.075 73.505 8.025 ;
      RECT 73.28 5.015 73.45 6.245 ;
      RECT 72.76 0.575 72.93 3.865 ;
      RECT 72.76 2.075 73.165 2.405 ;
      RECT 72.76 1.235 73.165 1.565 ;
      RECT 72.76 5.015 72.93 8.305 ;
      RECT 72.76 7.315 73.165 7.645 ;
      RECT 72.76 6.475 73.165 6.805 ;
      RECT 69.55 3.225 70.52 3.395 ;
      RECT 69.55 3.055 69.72 3.395 ;
      RECT 69.07 2.495 69.24 2.825 ;
      RECT 69.07 2.575 69.8 2.745 ;
      RECT 68.71 3.615 69 3.785 ;
      RECT 68.71 2.575 68.88 3.785 ;
      RECT 68.71 3.055 69 3.225 ;
      RECT 68.51 2.575 68.88 2.745 ;
      RECT 67.83 2.675 68 2.945 ;
      RECT 67.59 2.675 68 2.845 ;
      RECT 67.51 2.575 67.84 2.745 ;
      RECT 67.35 3.615 68 3.785 ;
      RECT 67.83 3.145 68 3.785 ;
      RECT 67.71 3.225 68 3.785 ;
      RECT 67.145 5.015 67.315 8.305 ;
      RECT 67.145 7.315 67.55 7.645 ;
      RECT 67.145 6.475 67.55 6.805 ;
      RECT 66.39 2.915 66.56 3.225 ;
      RECT 66.39 2.915 67.28 3.085 ;
      RECT 67.11 2.495 67.28 3.085 ;
      RECT 66.39 2.575 66.88 2.745 ;
      RECT 66.39 2.495 66.56 2.745 ;
      RECT 64.35 3.225 64.84 3.395 ;
      RECT 65.51 2.575 65.68 3.225 ;
      RECT 64.67 3.055 65.68 3.225 ;
      RECT 65.63 2.495 65.8 2.825 ;
      RECT 64.43 1.835 64.6 2.105 ;
      RECT 63.87 1.835 64.6 2.005 ;
      RECT 63.95 2.575 64.12 3.225 ;
      RECT 63.95 2.575 64.44 2.745 ;
      RECT 63.11 2.575 63.6 2.745 ;
      RECT 63.43 2.495 63.6 2.745 ;
      RECT 62.95 1.835 63.12 2.105 ;
      RECT 62.39 1.835 63.12 2.005 ;
      RECT 62.47 3.225 62.64 3.505 ;
      RECT 61.43 3.225 62.72 3.395 ;
      RECT 61.425 2.575 62 2.745 ;
      RECT 61.425 2.495 61.595 2.745 ;
      RECT 60.51 1.835 60.68 2.105 ;
      RECT 60.51 1.835 61.24 2.005 ;
      RECT 60.51 3.055 60.68 3.475 ;
      RECT 59.89 3.14 60.68 3.31 ;
      RECT 59.89 2.915 60.06 3.31 ;
      RECT 59.79 2.495 59.96 3.085 ;
      RECT 59.55 2.575 59.96 2.845 ;
      RECT 57.93 5.02 58.1 6.49 ;
      RECT 57.93 6.315 58.105 6.485 ;
      RECT 57.56 1.74 57.73 2.93 ;
      RECT 57.56 1.74 58.03 1.91 ;
      RECT 57.56 6.97 58.03 7.14 ;
      RECT 57.56 5.95 57.73 7.14 ;
      RECT 56.57 1.74 56.74 2.93 ;
      RECT 56.57 1.74 57.04 1.91 ;
      RECT 56.57 6.97 57.04 7.14 ;
      RECT 56.57 5.95 56.74 7.14 ;
      RECT 54.72 2.635 54.89 3.865 ;
      RECT 54.775 0.855 54.945 2.805 ;
      RECT 54.72 0.575 54.89 1.025 ;
      RECT 54.72 7.855 54.89 8.305 ;
      RECT 54.775 6.075 54.945 8.025 ;
      RECT 54.72 5.015 54.89 6.245 ;
      RECT 54.2 0.575 54.37 3.865 ;
      RECT 54.2 2.075 54.605 2.405 ;
      RECT 54.2 1.235 54.605 1.565 ;
      RECT 54.2 5.015 54.37 8.305 ;
      RECT 54.2 7.315 54.605 7.645 ;
      RECT 54.2 6.475 54.605 6.805 ;
      RECT 50.99 3.225 51.96 3.395 ;
      RECT 50.99 3.055 51.16 3.395 ;
      RECT 50.51 2.495 50.68 2.825 ;
      RECT 50.51 2.575 51.24 2.745 ;
      RECT 50.15 3.615 50.44 3.785 ;
      RECT 50.15 2.575 50.32 3.785 ;
      RECT 50.15 3.055 50.44 3.225 ;
      RECT 49.95 2.575 50.32 2.745 ;
      RECT 49.27 2.675 49.44 2.945 ;
      RECT 49.03 2.675 49.44 2.845 ;
      RECT 48.95 2.575 49.28 2.745 ;
      RECT 48.79 3.615 49.44 3.785 ;
      RECT 49.27 3.145 49.44 3.785 ;
      RECT 49.15 3.225 49.44 3.785 ;
      RECT 48.585 5.015 48.755 8.305 ;
      RECT 48.585 7.315 48.99 7.645 ;
      RECT 48.585 6.475 48.99 6.805 ;
      RECT 47.83 2.915 48 3.225 ;
      RECT 47.83 2.915 48.72 3.085 ;
      RECT 48.55 2.495 48.72 3.085 ;
      RECT 47.83 2.575 48.32 2.745 ;
      RECT 47.83 2.495 48 2.745 ;
      RECT 45.79 3.225 46.28 3.395 ;
      RECT 46.95 2.575 47.12 3.225 ;
      RECT 46.11 3.055 47.12 3.225 ;
      RECT 47.07 2.495 47.24 2.825 ;
      RECT 45.87 1.835 46.04 2.105 ;
      RECT 45.31 1.835 46.04 2.005 ;
      RECT 45.39 2.575 45.56 3.225 ;
      RECT 45.39 2.575 45.88 2.745 ;
      RECT 44.55 2.575 45.04 2.745 ;
      RECT 44.87 2.495 45.04 2.745 ;
      RECT 44.39 1.835 44.56 2.105 ;
      RECT 43.83 1.835 44.56 2.005 ;
      RECT 43.91 3.225 44.08 3.505 ;
      RECT 42.87 3.225 44.16 3.395 ;
      RECT 42.865 2.575 43.44 2.745 ;
      RECT 42.865 2.495 43.035 2.745 ;
      RECT 41.95 1.835 42.12 2.105 ;
      RECT 41.95 1.835 42.68 2.005 ;
      RECT 41.95 3.055 42.12 3.475 ;
      RECT 41.33 3.14 42.12 3.31 ;
      RECT 41.33 2.915 41.5 3.31 ;
      RECT 41.23 2.495 41.4 3.085 ;
      RECT 40.99 2.575 41.4 2.845 ;
      RECT 39.37 5.02 39.54 6.49 ;
      RECT 39.37 6.315 39.545 6.485 ;
      RECT 39 1.74 39.17 2.93 ;
      RECT 39 1.74 39.47 1.91 ;
      RECT 39 6.97 39.47 7.14 ;
      RECT 39 5.95 39.17 7.14 ;
      RECT 38.01 1.74 38.18 2.93 ;
      RECT 38.01 1.74 38.48 1.91 ;
      RECT 38.01 6.97 38.48 7.14 ;
      RECT 38.01 5.95 38.18 7.14 ;
      RECT 36.16 2.635 36.33 3.865 ;
      RECT 36.215 0.855 36.385 2.805 ;
      RECT 36.16 0.575 36.33 1.025 ;
      RECT 36.16 7.855 36.33 8.305 ;
      RECT 36.215 6.075 36.385 8.025 ;
      RECT 36.16 5.015 36.33 6.245 ;
      RECT 35.64 0.575 35.81 3.865 ;
      RECT 35.64 2.075 36.045 2.405 ;
      RECT 35.64 1.235 36.045 1.565 ;
      RECT 35.64 5.015 35.81 8.305 ;
      RECT 35.64 7.315 36.045 7.645 ;
      RECT 35.64 6.475 36.045 6.805 ;
      RECT 32.43 3.225 33.4 3.395 ;
      RECT 32.43 3.055 32.6 3.395 ;
      RECT 31.95 2.495 32.12 2.825 ;
      RECT 31.95 2.575 32.68 2.745 ;
      RECT 31.59 3.615 31.88 3.785 ;
      RECT 31.59 2.575 31.76 3.785 ;
      RECT 31.59 3.055 31.88 3.225 ;
      RECT 31.39 2.575 31.76 2.745 ;
      RECT 30.71 2.675 30.88 2.945 ;
      RECT 30.47 2.675 30.88 2.845 ;
      RECT 30.39 2.575 30.72 2.745 ;
      RECT 30.23 3.615 30.88 3.785 ;
      RECT 30.71 3.145 30.88 3.785 ;
      RECT 30.59 3.225 30.88 3.785 ;
      RECT 30.025 5.015 30.195 8.305 ;
      RECT 30.025 7.315 30.43 7.645 ;
      RECT 30.025 6.475 30.43 6.805 ;
      RECT 29.27 2.915 29.44 3.225 ;
      RECT 29.27 2.915 30.16 3.085 ;
      RECT 29.99 2.495 30.16 3.085 ;
      RECT 29.27 2.575 29.76 2.745 ;
      RECT 29.27 2.495 29.44 2.745 ;
      RECT 27.23 3.225 27.72 3.395 ;
      RECT 28.39 2.575 28.56 3.225 ;
      RECT 27.55 3.055 28.56 3.225 ;
      RECT 28.51 2.495 28.68 2.825 ;
      RECT 27.31 1.835 27.48 2.105 ;
      RECT 26.75 1.835 27.48 2.005 ;
      RECT 26.83 2.575 27 3.225 ;
      RECT 26.83 2.575 27.32 2.745 ;
      RECT 25.99 2.575 26.48 2.745 ;
      RECT 26.31 2.495 26.48 2.745 ;
      RECT 25.83 1.835 26 2.105 ;
      RECT 25.27 1.835 26 2.005 ;
      RECT 25.35 3.225 25.52 3.505 ;
      RECT 24.31 3.225 25.6 3.395 ;
      RECT 24.305 2.575 24.88 2.745 ;
      RECT 24.305 2.495 24.475 2.745 ;
      RECT 23.39 1.835 23.56 2.105 ;
      RECT 23.39 1.835 24.12 2.005 ;
      RECT 23.39 3.055 23.56 3.475 ;
      RECT 22.77 3.14 23.56 3.31 ;
      RECT 22.77 2.915 22.94 3.31 ;
      RECT 22.67 2.495 22.84 3.085 ;
      RECT 22.43 2.575 22.84 2.845 ;
      RECT 20.81 5.02 20.98 6.49 ;
      RECT 20.81 6.315 20.985 6.485 ;
      RECT 20.44 1.74 20.61 2.93 ;
      RECT 20.44 1.74 20.91 1.91 ;
      RECT 20.44 6.97 20.91 7.14 ;
      RECT 20.44 5.95 20.61 7.14 ;
      RECT 19.45 1.74 19.62 2.93 ;
      RECT 19.45 1.74 19.92 1.91 ;
      RECT 19.45 6.97 19.92 7.14 ;
      RECT 19.45 5.95 19.62 7.14 ;
      RECT 17.6 2.635 17.77 3.865 ;
      RECT 17.655 0.855 17.825 2.805 ;
      RECT 17.6 0.575 17.77 1.025 ;
      RECT 17.6 7.855 17.77 8.305 ;
      RECT 17.655 6.075 17.825 8.025 ;
      RECT 17.6 5.015 17.77 6.245 ;
      RECT 17.08 0.575 17.25 3.865 ;
      RECT 17.08 2.075 17.485 2.405 ;
      RECT 17.08 1.235 17.485 1.565 ;
      RECT 17.08 5.015 17.25 8.305 ;
      RECT 17.08 7.315 17.485 7.645 ;
      RECT 17.08 6.475 17.485 6.805 ;
      RECT 13.87 3.225 14.84 3.395 ;
      RECT 13.87 3.055 14.04 3.395 ;
      RECT 13.39 2.495 13.56 2.825 ;
      RECT 13.39 2.575 14.12 2.745 ;
      RECT 13.03 3.615 13.32 3.785 ;
      RECT 13.03 2.575 13.2 3.785 ;
      RECT 13.03 3.055 13.32 3.225 ;
      RECT 12.83 2.575 13.2 2.745 ;
      RECT 12.15 2.675 12.32 2.945 ;
      RECT 11.91 2.675 12.32 2.845 ;
      RECT 11.83 2.575 12.16 2.745 ;
      RECT 11.67 3.615 12.32 3.785 ;
      RECT 12.15 3.145 12.32 3.785 ;
      RECT 12.03 3.225 12.32 3.785 ;
      RECT 11.465 5.015 11.635 8.305 ;
      RECT 11.465 7.315 11.87 7.645 ;
      RECT 11.465 6.475 11.87 6.805 ;
      RECT 10.71 2.915 10.88 3.225 ;
      RECT 10.71 2.915 11.6 3.085 ;
      RECT 11.43 2.495 11.6 3.085 ;
      RECT 10.71 2.575 11.2 2.745 ;
      RECT 10.71 2.495 10.88 2.745 ;
      RECT 8.67 3.225 9.16 3.395 ;
      RECT 9.83 2.575 10 3.225 ;
      RECT 8.99 3.055 10 3.225 ;
      RECT 9.95 2.495 10.12 2.825 ;
      RECT 8.75 1.835 8.92 2.105 ;
      RECT 8.19 1.835 8.92 2.005 ;
      RECT 8.27 2.575 8.44 3.225 ;
      RECT 8.27 2.575 8.76 2.745 ;
      RECT 7.43 2.575 7.92 2.745 ;
      RECT 7.75 2.495 7.92 2.745 ;
      RECT 7.27 1.835 7.44 2.105 ;
      RECT 6.71 1.835 7.44 2.005 ;
      RECT 6.79 3.225 6.96 3.505 ;
      RECT 5.75 3.225 7.04 3.395 ;
      RECT 5.745 2.575 6.32 2.745 ;
      RECT 5.745 2.495 5.915 2.745 ;
      RECT 4.83 1.835 5 2.105 ;
      RECT 4.83 1.835 5.56 2.005 ;
      RECT 4.83 3.055 5 3.475 ;
      RECT 4.21 3.14 5 3.31 ;
      RECT 4.21 2.915 4.38 3.31 ;
      RECT 4.11 2.495 4.28 3.085 ;
      RECT 3.87 2.575 4.28 2.845 ;
      RECT 1.17 7.855 1.34 8.305 ;
      RECT 1.225 6.075 1.395 8.025 ;
      RECT 1.17 5.015 1.34 6.245 ;
      RECT 0.65 5.015 0.82 8.305 ;
      RECT 0.65 7.315 1.055 7.645 ;
      RECT 0.65 6.475 1.055 6.805 ;
      RECT 95.05 7.8 95.22 8.31 ;
      RECT 94.06 0.57 94.23 1.08 ;
      RECT 94.06 2.39 94.23 3.86 ;
      RECT 94.06 5.02 94.23 6.49 ;
      RECT 94.06 7.8 94.23 8.31 ;
      RECT 92.7 0.575 92.87 3.865 ;
      RECT 92.7 5.015 92.87 8.305 ;
      RECT 92.27 0.575 92.44 1.085 ;
      RECT 92.27 1.655 92.44 3.865 ;
      RECT 92.27 5.015 92.44 7.225 ;
      RECT 92.27 7.795 92.44 8.305 ;
      RECT 88.59 2.495 88.76 2.945 ;
      RECT 88.35 1.755 88.52 2.105 ;
      RECT 87.39 1.755 87.56 2.105 ;
      RECT 87.085 5.015 87.255 8.305 ;
      RECT 86.91 3.055 87.08 3.475 ;
      RECT 86.655 5.015 86.825 7.225 ;
      RECT 86.655 7.795 86.825 8.305 ;
      RECT 85.91 1.755 86.08 2.105 ;
      RECT 84.95 1.755 85.12 2.105 ;
      RECT 84.95 3.485 85.12 3.815 ;
      RECT 84.43 3.145 84.6 3.785 ;
      RECT 83.95 1.755 84.12 2.105 ;
      RECT 83.71 2.495 83.88 2.825 ;
      RECT 83.23 2.495 83.4 2.825 ;
      RECT 81.99 3.145 82.16 3.505 ;
      RECT 81.51 3.055 81.68 3.475 ;
      RECT 80.79 2.495 80.96 2.945 ;
      RECT 78.83 2.495 79 2.825 ;
      RECT 78.11 1.755 78.28 2.105 ;
      RECT 78.11 3.285 78.28 3.645 ;
      RECT 76.49 7.8 76.66 8.31 ;
      RECT 75.5 0.57 75.67 1.08 ;
      RECT 75.5 2.39 75.67 3.86 ;
      RECT 75.5 5.02 75.67 6.49 ;
      RECT 75.5 7.8 75.67 8.31 ;
      RECT 74.14 0.575 74.31 3.865 ;
      RECT 74.14 5.015 74.31 8.305 ;
      RECT 73.71 0.575 73.88 1.085 ;
      RECT 73.71 1.655 73.88 3.865 ;
      RECT 73.71 5.015 73.88 7.225 ;
      RECT 73.71 7.795 73.88 8.305 ;
      RECT 70.03 2.495 70.2 2.945 ;
      RECT 69.79 1.755 69.96 2.105 ;
      RECT 68.83 1.755 69 2.105 ;
      RECT 68.525 5.015 68.695 8.305 ;
      RECT 68.35 3.055 68.52 3.475 ;
      RECT 68.095 5.015 68.265 7.225 ;
      RECT 68.095 7.795 68.265 8.305 ;
      RECT 67.35 1.755 67.52 2.105 ;
      RECT 66.39 1.755 66.56 2.105 ;
      RECT 66.39 3.485 66.56 3.815 ;
      RECT 65.87 3.145 66.04 3.785 ;
      RECT 65.39 1.755 65.56 2.105 ;
      RECT 65.15 2.495 65.32 2.825 ;
      RECT 64.67 2.495 64.84 2.825 ;
      RECT 63.43 3.145 63.6 3.505 ;
      RECT 62.95 3.055 63.12 3.475 ;
      RECT 62.23 2.495 62.4 2.945 ;
      RECT 60.27 2.495 60.44 2.825 ;
      RECT 59.55 1.755 59.72 2.105 ;
      RECT 59.55 3.285 59.72 3.645 ;
      RECT 57.93 7.8 58.1 8.31 ;
      RECT 56.94 0.57 57.11 1.08 ;
      RECT 56.94 2.39 57.11 3.86 ;
      RECT 56.94 5.02 57.11 6.49 ;
      RECT 56.94 7.8 57.11 8.31 ;
      RECT 55.58 0.575 55.75 3.865 ;
      RECT 55.58 5.015 55.75 8.305 ;
      RECT 55.15 0.575 55.32 1.085 ;
      RECT 55.15 1.655 55.32 3.865 ;
      RECT 55.15 5.015 55.32 7.225 ;
      RECT 55.15 7.795 55.32 8.305 ;
      RECT 51.47 2.495 51.64 2.945 ;
      RECT 51.23 1.755 51.4 2.105 ;
      RECT 50.27 1.755 50.44 2.105 ;
      RECT 49.965 5.015 50.135 8.305 ;
      RECT 49.79 3.055 49.96 3.475 ;
      RECT 49.535 5.015 49.705 7.225 ;
      RECT 49.535 7.795 49.705 8.305 ;
      RECT 48.79 1.755 48.96 2.105 ;
      RECT 47.83 1.755 48 2.105 ;
      RECT 47.83 3.485 48 3.815 ;
      RECT 47.31 3.145 47.48 3.785 ;
      RECT 46.83 1.755 47 2.105 ;
      RECT 46.59 2.495 46.76 2.825 ;
      RECT 46.11 2.495 46.28 2.825 ;
      RECT 44.87 3.145 45.04 3.505 ;
      RECT 44.39 3.055 44.56 3.475 ;
      RECT 43.67 2.495 43.84 2.945 ;
      RECT 41.71 2.495 41.88 2.825 ;
      RECT 40.99 1.755 41.16 2.105 ;
      RECT 40.99 3.285 41.16 3.645 ;
      RECT 39.37 7.8 39.54 8.31 ;
      RECT 38.38 0.57 38.55 1.08 ;
      RECT 38.38 2.39 38.55 3.86 ;
      RECT 38.38 5.02 38.55 6.49 ;
      RECT 38.38 7.8 38.55 8.31 ;
      RECT 37.02 0.575 37.19 3.865 ;
      RECT 37.02 5.015 37.19 8.305 ;
      RECT 36.59 0.575 36.76 1.085 ;
      RECT 36.59 1.655 36.76 3.865 ;
      RECT 36.59 5.015 36.76 7.225 ;
      RECT 36.59 7.795 36.76 8.305 ;
      RECT 32.91 2.495 33.08 2.945 ;
      RECT 32.67 1.755 32.84 2.105 ;
      RECT 31.71 1.755 31.88 2.105 ;
      RECT 31.405 5.015 31.575 8.305 ;
      RECT 31.23 3.055 31.4 3.475 ;
      RECT 30.975 5.015 31.145 7.225 ;
      RECT 30.975 7.795 31.145 8.305 ;
      RECT 30.23 1.755 30.4 2.105 ;
      RECT 29.27 1.755 29.44 2.105 ;
      RECT 29.27 3.485 29.44 3.815 ;
      RECT 28.75 3.145 28.92 3.785 ;
      RECT 28.27 1.755 28.44 2.105 ;
      RECT 28.03 2.495 28.2 2.825 ;
      RECT 27.55 2.495 27.72 2.825 ;
      RECT 26.31 3.145 26.48 3.505 ;
      RECT 25.83 3.055 26 3.475 ;
      RECT 25.11 2.495 25.28 2.945 ;
      RECT 23.15 2.495 23.32 2.825 ;
      RECT 22.43 1.755 22.6 2.105 ;
      RECT 22.43 3.285 22.6 3.645 ;
      RECT 20.81 7.8 20.98 8.31 ;
      RECT 19.82 0.57 19.99 1.08 ;
      RECT 19.82 2.39 19.99 3.86 ;
      RECT 19.82 5.02 19.99 6.49 ;
      RECT 19.82 7.8 19.99 8.31 ;
      RECT 18.46 0.575 18.63 3.865 ;
      RECT 18.46 5.015 18.63 8.305 ;
      RECT 18.03 0.575 18.2 1.085 ;
      RECT 18.03 1.655 18.2 3.865 ;
      RECT 18.03 5.015 18.2 7.225 ;
      RECT 18.03 7.795 18.2 8.305 ;
      RECT 14.35 2.495 14.52 2.945 ;
      RECT 14.11 1.755 14.28 2.105 ;
      RECT 13.15 1.755 13.32 2.105 ;
      RECT 12.845 5.015 13.015 8.305 ;
      RECT 12.67 3.055 12.84 3.475 ;
      RECT 12.415 5.015 12.585 7.225 ;
      RECT 12.415 7.795 12.585 8.305 ;
      RECT 11.67 1.755 11.84 2.105 ;
      RECT 10.71 1.755 10.88 2.105 ;
      RECT 10.71 3.485 10.88 3.815 ;
      RECT 10.19 3.145 10.36 3.785 ;
      RECT 9.71 1.755 9.88 2.105 ;
      RECT 9.47 2.495 9.64 2.825 ;
      RECT 8.99 2.495 9.16 2.825 ;
      RECT 7.75 3.145 7.92 3.505 ;
      RECT 7.27 3.055 7.44 3.475 ;
      RECT 6.55 2.495 6.72 2.945 ;
      RECT 4.59 2.495 4.76 2.825 ;
      RECT 3.87 1.755 4.04 2.105 ;
      RECT 3.87 3.285 4.04 3.645 ;
      RECT 1.6 5.015 1.77 7.225 ;
      RECT 1.6 7.795 1.77 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r1 ;
  SIZE 79.1 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 17.52 0.915 17.69 1.085 ;
        RECT 17.515 0.91 17.685 1.08 ;
        RECT 17.515 2.39 17.685 2.56 ;
      LAYER li1 ;
        RECT 17.52 0.915 17.69 1.085 ;
        RECT 17.515 0.57 17.685 1.08 ;
        RECT 17.515 2.39 17.685 3.86 ;
      LAYER met1 ;
        RECT 17.455 2.36 17.745 2.59 ;
        RECT 17.455 0.88 17.745 1.11 ;
        RECT 17.515 0.88 17.685 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 32.78 0.915 32.95 1.085 ;
        RECT 32.775 0.91 32.945 1.08 ;
        RECT 32.775 2.39 32.945 2.56 ;
      LAYER li1 ;
        RECT 32.78 0.915 32.95 1.085 ;
        RECT 32.775 0.57 32.945 1.08 ;
        RECT 32.775 2.39 32.945 3.86 ;
      LAYER met1 ;
        RECT 32.715 2.36 33.005 2.59 ;
        RECT 32.715 0.88 33.005 1.11 ;
        RECT 32.775 0.88 32.945 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 48.04 0.915 48.21 1.085 ;
        RECT 48.035 0.91 48.205 1.08 ;
        RECT 48.035 2.39 48.205 2.56 ;
      LAYER li1 ;
        RECT 48.04 0.915 48.21 1.085 ;
        RECT 48.035 0.57 48.205 1.08 ;
        RECT 48.035 2.39 48.205 3.86 ;
      LAYER met1 ;
        RECT 47.975 2.36 48.265 2.59 ;
        RECT 47.975 0.88 48.265 1.11 ;
        RECT 48.035 0.88 48.205 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 63.3 0.915 63.47 1.085 ;
        RECT 63.295 0.91 63.465 1.08 ;
        RECT 63.295 2.39 63.465 2.56 ;
      LAYER li1 ;
        RECT 63.3 0.915 63.47 1.085 ;
        RECT 63.295 0.57 63.465 1.08 ;
        RECT 63.295 2.39 63.465 3.86 ;
      LAYER met1 ;
        RECT 63.235 2.36 63.525 2.59 ;
        RECT 63.235 0.88 63.525 1.11 ;
        RECT 63.295 0.88 63.465 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 78.56 0.915 78.73 1.085 ;
        RECT 78.555 0.91 78.725 1.08 ;
        RECT 78.555 2.39 78.725 2.56 ;
      LAYER li1 ;
        RECT 78.56 0.915 78.73 1.085 ;
        RECT 78.555 0.57 78.725 1.08 ;
        RECT 78.555 2.39 78.725 3.86 ;
      LAYER met1 ;
        RECT 78.495 2.36 78.785 2.59 ;
        RECT 78.495 0.88 78.785 1.11 ;
        RECT 78.555 0.88 78.725 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 13.285 5.86 13.625 6.21 ;
        RECT 13.285 2.705 13.625 3.055 ;
        RECT 13.365 2.705 13.535 6.21 ;
      LAYER li1 ;
        RECT 13.365 1.66 13.535 2.935 ;
        RECT 13.365 5.945 13.535 7.22 ;
        RECT 7.75 5.945 7.92 7.22 ;
      LAYER met1 ;
        RECT 13.285 2.765 13.765 2.935 ;
        RECT 13.285 2.705 13.625 3.055 ;
        RECT 7.69 5.945 13.765 6.115 ;
        RECT 13.285 5.86 13.625 6.21 ;
        RECT 7.69 5.915 7.98 6.145 ;
      LAYER mcon ;
        RECT 7.75 5.945 7.92 6.115 ;
        RECT 13.365 5.945 13.535 6.115 ;
        RECT 13.365 2.765 13.535 2.935 ;
      LAYER via1 ;
        RECT 13.385 5.96 13.535 6.11 ;
        RECT 13.385 2.805 13.535 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 28.545 5.86 28.885 6.21 ;
        RECT 28.545 2.705 28.885 3.055 ;
        RECT 28.625 2.705 28.795 6.21 ;
      LAYER li1 ;
        RECT 28.625 1.66 28.795 2.935 ;
        RECT 28.625 5.945 28.795 7.22 ;
        RECT 23.01 5.945 23.18 7.22 ;
      LAYER met1 ;
        RECT 28.545 2.765 29.025 2.935 ;
        RECT 28.545 2.705 28.885 3.055 ;
        RECT 22.95 5.945 29.025 6.115 ;
        RECT 28.545 5.86 28.885 6.21 ;
        RECT 22.95 5.915 23.24 6.145 ;
      LAYER mcon ;
        RECT 23.01 5.945 23.18 6.115 ;
        RECT 28.625 5.945 28.795 6.115 ;
        RECT 28.625 2.765 28.795 2.935 ;
      LAYER via1 ;
        RECT 28.645 5.96 28.795 6.11 ;
        RECT 28.645 2.805 28.795 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 43.805 5.86 44.145 6.21 ;
        RECT 43.805 2.705 44.145 3.055 ;
        RECT 43.885 2.705 44.055 6.21 ;
      LAYER li1 ;
        RECT 43.885 1.66 44.055 2.935 ;
        RECT 43.885 5.945 44.055 7.22 ;
        RECT 38.27 5.945 38.44 7.22 ;
      LAYER met1 ;
        RECT 43.805 2.765 44.285 2.935 ;
        RECT 43.805 2.705 44.145 3.055 ;
        RECT 38.21 5.945 44.285 6.115 ;
        RECT 43.805 5.86 44.145 6.21 ;
        RECT 38.21 5.915 38.5 6.145 ;
      LAYER mcon ;
        RECT 38.27 5.945 38.44 6.115 ;
        RECT 43.885 5.945 44.055 6.115 ;
        RECT 43.885 2.765 44.055 2.935 ;
      LAYER via1 ;
        RECT 43.905 5.96 44.055 6.11 ;
        RECT 43.905 2.805 44.055 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 59.065 5.86 59.405 6.21 ;
        RECT 59.065 2.705 59.405 3.055 ;
        RECT 59.145 2.705 59.315 6.21 ;
      LAYER li1 ;
        RECT 59.145 1.66 59.315 2.935 ;
        RECT 59.145 5.945 59.315 7.22 ;
        RECT 53.53 5.945 53.7 7.22 ;
      LAYER met1 ;
        RECT 59.065 2.765 59.545 2.935 ;
        RECT 59.065 2.705 59.405 3.055 ;
        RECT 53.47 5.945 59.545 6.115 ;
        RECT 59.065 5.86 59.405 6.21 ;
        RECT 53.47 5.915 53.76 6.145 ;
      LAYER mcon ;
        RECT 53.53 5.945 53.7 6.115 ;
        RECT 59.145 5.945 59.315 6.115 ;
        RECT 59.145 2.765 59.315 2.935 ;
      LAYER via1 ;
        RECT 59.165 5.96 59.315 6.11 ;
        RECT 59.165 2.805 59.315 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 74.325 5.86 74.665 6.21 ;
        RECT 74.325 2.705 74.665 3.055 ;
        RECT 74.405 2.705 74.575 6.21 ;
      LAYER li1 ;
        RECT 74.405 1.66 74.575 2.935 ;
        RECT 74.405 5.945 74.575 7.22 ;
        RECT 68.79 5.945 68.96 7.22 ;
      LAYER met1 ;
        RECT 74.325 2.765 74.805 2.935 ;
        RECT 74.325 2.705 74.665 3.055 ;
        RECT 68.73 5.945 74.805 6.115 ;
        RECT 74.325 5.86 74.665 6.21 ;
        RECT 68.73 5.915 69.02 6.145 ;
      LAYER mcon ;
        RECT 68.79 5.945 68.96 6.115 ;
        RECT 74.405 5.945 74.575 6.115 ;
        RECT 74.405 2.765 74.575 2.935 ;
      LAYER via1 ;
        RECT 74.425 5.96 74.575 6.11 ;
        RECT 74.425 2.805 74.575 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.235 5.945 0.405 7.22 ;
      LAYER met1 ;
        RECT 0.175 5.945 0.635 6.115 ;
        RECT 0.175 5.915 0.465 6.145 ;
      LAYER mcon ;
        RECT 0.235 5.945 0.405 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.67 4.265 2.475 4.645 ;
      LAYER met2 ;
        RECT 1.86 4.265 2.24 4.645 ;
      LAYER li1 ;
        RECT 0.05 4.44 79.1 4.745 ;
        RECT 72.16 4.135 79.1 4.745 ;
        RECT 76.965 4.13 78.945 4.75 ;
        RECT 78.125 3.4 78.295 5.48 ;
        RECT 77.135 3.4 77.305 5.48 ;
        RECT 74.395 3.405 74.565 5.475 ;
        RECT 64.59 4.13 73.33 4.3 ;
        RECT 2.135 4.305 79.1 4.745 ;
        RECT 71.62 3.63 71.79 4.3 ;
        RECT 69.7 3.63 69.87 4.3 ;
        RECT 68.78 4.305 68.95 5.475 ;
        RECT 68.76 3.63 68.93 4.3 ;
        RECT 67.3 3.63 67.47 4.3 ;
        RECT 65.38 3.63 65.55 4.3 ;
        RECT 56.9 4.14 64.595 4.745 ;
        RECT 49.33 4.135 63.84 4.3 ;
        RECT 61.705 4.13 63.685 4.75 ;
        RECT 62.865 3.4 63.035 5.48 ;
        RECT 61.875 3.4 62.045 5.48 ;
        RECT 59.135 3.405 59.305 5.475 ;
        RECT 49.33 4.13 58.07 4.3 ;
        RECT 56.36 3.63 56.53 4.3 ;
        RECT 54.44 3.63 54.61 4.3 ;
        RECT 53.52 4.305 53.69 5.475 ;
        RECT 53.5 3.63 53.67 4.3 ;
        RECT 52.04 3.63 52.21 4.3 ;
        RECT 50.12 3.63 50.29 4.3 ;
        RECT 41.64 4.14 49.335 4.745 ;
        RECT 34.07 4.135 48.58 4.3 ;
        RECT 46.445 4.13 48.425 4.75 ;
        RECT 47.605 3.4 47.775 5.48 ;
        RECT 46.615 3.4 46.785 5.48 ;
        RECT 43.875 3.405 44.045 5.475 ;
        RECT 34.07 4.13 42.81 4.3 ;
        RECT 41.1 3.63 41.27 4.3 ;
        RECT 39.18 3.63 39.35 4.3 ;
        RECT 38.26 4.305 38.43 5.475 ;
        RECT 38.24 3.63 38.41 4.3 ;
        RECT 36.78 3.63 36.95 4.3 ;
        RECT 34.86 3.63 35.03 4.3 ;
        RECT 26.38 4.14 34.075 4.745 ;
        RECT 18.81 4.135 33.32 4.3 ;
        RECT 31.185 4.13 33.165 4.75 ;
        RECT 32.345 3.4 32.515 5.48 ;
        RECT 31.355 3.4 31.525 5.48 ;
        RECT 28.615 3.405 28.785 5.475 ;
        RECT 18.81 4.13 27.55 4.3 ;
        RECT 25.84 3.63 26.01 4.3 ;
        RECT 23.92 3.63 24.09 4.3 ;
        RECT 23 4.305 23.17 5.475 ;
        RECT 22.98 3.63 23.15 4.3 ;
        RECT 21.52 3.63 21.69 4.3 ;
        RECT 19.6 3.63 19.77 4.3 ;
        RECT 11.12 4.14 18.815 4.745 ;
        RECT 3.55 4.135 18.06 4.3 ;
        RECT 15.925 4.13 17.905 4.75 ;
        RECT 17.085 3.4 17.255 5.48 ;
        RECT 16.095 3.4 16.265 5.48 ;
        RECT 13.355 3.405 13.525 5.475 ;
        RECT 3.55 4.13 12.29 4.3 ;
        RECT 10.58 3.63 10.75 4.3 ;
        RECT 8.66 3.63 8.83 4.3 ;
        RECT 7.74 4.305 7.91 5.475 ;
        RECT 7.72 3.63 7.89 4.3 ;
        RECT 6.26 3.63 6.43 4.3 ;
        RECT 4.34 3.63 4.51 4.3 ;
        RECT 0.05 4.14 3.695 4.34 ;
        RECT 2.035 4.44 2.205 8.305 ;
        RECT 0.05 4.14 1.965 4.745 ;
        RECT 0.225 4.14 0.395 5.475 ;
      LAYER met1 ;
        RECT 0.05 4.14 79.1 4.745 ;
        RECT 64.59 4.135 79.1 4.745 ;
        RECT 76.965 4.13 78.945 4.75 ;
        RECT 64.59 3.98 73.33 4.745 ;
        RECT 49.33 4.135 63.84 4.745 ;
        RECT 61.705 4.13 63.685 4.75 ;
        RECT 49.33 3.98 58.07 4.745 ;
        RECT 34.07 4.135 48.58 4.745 ;
        RECT 46.445 4.13 48.425 4.75 ;
        RECT 34.07 3.98 42.81 4.745 ;
        RECT 18.81 4.135 33.32 4.745 ;
        RECT 31.185 4.13 33.165 4.75 ;
        RECT 18.81 3.98 27.55 4.745 ;
        RECT 3.55 4.135 18.06 4.745 ;
        RECT 15.925 4.13 17.905 4.75 ;
        RECT 3.55 3.98 12.29 4.745 ;
        RECT 1.975 6.655 2.265 6.885 ;
        RECT 1.805 6.685 2.265 6.855 ;
      LAYER via2 ;
        RECT 1.95 4.355 2.15 4.555 ;
      LAYER mcon ;
        RECT 2.035 6.685 2.205 6.855 ;
        RECT 2.345 4.545 2.515 4.715 ;
        RECT 3.69 4.13 3.86 4.3 ;
        RECT 4.15 4.13 4.32 4.3 ;
        RECT 4.61 4.13 4.78 4.3 ;
        RECT 5.07 4.13 5.24 4.3 ;
        RECT 5.53 4.13 5.7 4.3 ;
        RECT 5.99 4.13 6.16 4.3 ;
        RECT 6.45 4.13 6.62 4.3 ;
        RECT 6.91 4.13 7.08 4.3 ;
        RECT 7.37 4.13 7.54 4.3 ;
        RECT 7.83 4.13 8 4.3 ;
        RECT 8.29 4.13 8.46 4.3 ;
        RECT 8.75 4.13 8.92 4.3 ;
        RECT 9.21 4.13 9.38 4.3 ;
        RECT 9.67 4.13 9.84 4.3 ;
        RECT 9.86 4.545 10.03 4.715 ;
        RECT 10.13 4.13 10.3 4.3 ;
        RECT 10.59 4.13 10.76 4.3 ;
        RECT 11.05 4.13 11.22 4.3 ;
        RECT 11.51 4.13 11.68 4.3 ;
        RECT 11.97 4.13 12.14 4.3 ;
        RECT 15.475 4.545 15.645 4.715 ;
        RECT 15.475 4.165 15.645 4.335 ;
        RECT 16.175 4.55 16.345 4.72 ;
        RECT 16.175 4.16 16.345 4.33 ;
        RECT 17.165 4.55 17.335 4.72 ;
        RECT 17.165 4.16 17.335 4.33 ;
        RECT 18.95 4.13 19.12 4.3 ;
        RECT 19.41 4.13 19.58 4.3 ;
        RECT 19.87 4.13 20.04 4.3 ;
        RECT 20.33 4.13 20.5 4.3 ;
        RECT 20.79 4.13 20.96 4.3 ;
        RECT 21.25 4.13 21.42 4.3 ;
        RECT 21.71 4.13 21.88 4.3 ;
        RECT 22.17 4.13 22.34 4.3 ;
        RECT 22.63 4.13 22.8 4.3 ;
        RECT 23.09 4.13 23.26 4.3 ;
        RECT 23.55 4.13 23.72 4.3 ;
        RECT 24.01 4.13 24.18 4.3 ;
        RECT 24.47 4.13 24.64 4.3 ;
        RECT 24.93 4.13 25.1 4.3 ;
        RECT 25.12 4.545 25.29 4.715 ;
        RECT 25.39 4.13 25.56 4.3 ;
        RECT 25.85 4.13 26.02 4.3 ;
        RECT 26.31 4.13 26.48 4.3 ;
        RECT 26.77 4.13 26.94 4.3 ;
        RECT 27.23 4.13 27.4 4.3 ;
        RECT 30.735 4.545 30.905 4.715 ;
        RECT 30.735 4.165 30.905 4.335 ;
        RECT 31.435 4.55 31.605 4.72 ;
        RECT 31.435 4.16 31.605 4.33 ;
        RECT 32.425 4.55 32.595 4.72 ;
        RECT 32.425 4.16 32.595 4.33 ;
        RECT 34.21 4.13 34.38 4.3 ;
        RECT 34.67 4.13 34.84 4.3 ;
        RECT 35.13 4.13 35.3 4.3 ;
        RECT 35.59 4.13 35.76 4.3 ;
        RECT 36.05 4.13 36.22 4.3 ;
        RECT 36.51 4.13 36.68 4.3 ;
        RECT 36.97 4.13 37.14 4.3 ;
        RECT 37.43 4.13 37.6 4.3 ;
        RECT 37.89 4.13 38.06 4.3 ;
        RECT 38.35 4.13 38.52 4.3 ;
        RECT 38.81 4.13 38.98 4.3 ;
        RECT 39.27 4.13 39.44 4.3 ;
        RECT 39.73 4.13 39.9 4.3 ;
        RECT 40.19 4.13 40.36 4.3 ;
        RECT 40.38 4.545 40.55 4.715 ;
        RECT 40.65 4.13 40.82 4.3 ;
        RECT 41.11 4.13 41.28 4.3 ;
        RECT 41.57 4.13 41.74 4.3 ;
        RECT 42.03 4.13 42.2 4.3 ;
        RECT 42.49 4.13 42.66 4.3 ;
        RECT 45.995 4.545 46.165 4.715 ;
        RECT 45.995 4.165 46.165 4.335 ;
        RECT 46.695 4.55 46.865 4.72 ;
        RECT 46.695 4.16 46.865 4.33 ;
        RECT 47.685 4.55 47.855 4.72 ;
        RECT 47.685 4.16 47.855 4.33 ;
        RECT 49.47 4.13 49.64 4.3 ;
        RECT 49.93 4.13 50.1 4.3 ;
        RECT 50.39 4.13 50.56 4.3 ;
        RECT 50.85 4.13 51.02 4.3 ;
        RECT 51.31 4.13 51.48 4.3 ;
        RECT 51.77 4.13 51.94 4.3 ;
        RECT 52.23 4.13 52.4 4.3 ;
        RECT 52.69 4.13 52.86 4.3 ;
        RECT 53.15 4.13 53.32 4.3 ;
        RECT 53.61 4.13 53.78 4.3 ;
        RECT 54.07 4.13 54.24 4.3 ;
        RECT 54.53 4.13 54.7 4.3 ;
        RECT 54.99 4.13 55.16 4.3 ;
        RECT 55.45 4.13 55.62 4.3 ;
        RECT 55.64 4.545 55.81 4.715 ;
        RECT 55.91 4.13 56.08 4.3 ;
        RECT 56.37 4.13 56.54 4.3 ;
        RECT 56.83 4.13 57 4.3 ;
        RECT 57.29 4.13 57.46 4.3 ;
        RECT 57.75 4.13 57.92 4.3 ;
        RECT 61.255 4.545 61.425 4.715 ;
        RECT 61.255 4.165 61.425 4.335 ;
        RECT 61.955 4.55 62.125 4.72 ;
        RECT 61.955 4.16 62.125 4.33 ;
        RECT 62.945 4.55 63.115 4.72 ;
        RECT 62.945 4.16 63.115 4.33 ;
        RECT 64.73 4.13 64.9 4.3 ;
        RECT 65.19 4.13 65.36 4.3 ;
        RECT 65.65 4.13 65.82 4.3 ;
        RECT 66.11 4.13 66.28 4.3 ;
        RECT 66.57 4.13 66.74 4.3 ;
        RECT 67.03 4.13 67.2 4.3 ;
        RECT 67.49 4.13 67.66 4.3 ;
        RECT 67.95 4.13 68.12 4.3 ;
        RECT 68.41 4.13 68.58 4.3 ;
        RECT 68.87 4.13 69.04 4.3 ;
        RECT 69.33 4.13 69.5 4.3 ;
        RECT 69.79 4.13 69.96 4.3 ;
        RECT 70.25 4.13 70.42 4.3 ;
        RECT 70.71 4.13 70.88 4.3 ;
        RECT 70.9 4.545 71.07 4.715 ;
        RECT 71.17 4.13 71.34 4.3 ;
        RECT 71.63 4.13 71.8 4.3 ;
        RECT 72.09 4.13 72.26 4.3 ;
        RECT 72.55 4.13 72.72 4.3 ;
        RECT 73.01 4.13 73.18 4.3 ;
        RECT 76.515 4.545 76.685 4.715 ;
        RECT 76.515 4.165 76.685 4.335 ;
        RECT 77.215 4.55 77.385 4.72 ;
        RECT 77.215 4.16 77.385 4.33 ;
        RECT 78.205 4.55 78.375 4.72 ;
        RECT 78.205 4.16 78.375 4.33 ;
      LAYER via1 ;
        RECT 1.975 4.38 2.125 4.53 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 65.42 1.85 66.15 2.18 ;
        RECT 50.16 1.85 50.89 2.18 ;
        RECT 34.9 1.85 35.63 2.18 ;
        RECT 19.64 1.85 20.37 2.18 ;
        RECT 4.38 1.85 5.11 2.18 ;
        RECT 0.05 0 0.855 0.38 ;
        RECT 0.01 8.5 0.815 8.88 ;
      LAYER met2 ;
        RECT 65.56 1.86 65.95 2.18 ;
        RECT 65.56 1.83 65.84 2.2 ;
        RECT 50.3 1.86 50.69 2.18 ;
        RECT 50.3 1.83 50.58 2.2 ;
        RECT 35.04 1.86 35.43 2.18 ;
        RECT 35.04 1.83 35.32 2.2 ;
        RECT 19.78 1.86 20.17 2.18 ;
        RECT 19.78 1.83 20.06 2.2 ;
        RECT 4.52 1.86 4.91 2.18 ;
        RECT 4.52 1.83 4.8 2.2 ;
        RECT 0.24 0 0.62 0.38 ;
        RECT 0.2 8.5 0.58 8.88 ;
        RECT 0.285 0 0.44 8.88 ;
      LAYER li1 ;
        RECT 78.92 0 79.1 0.305 ;
        RECT 0.515 0 79.1 0.3 ;
        RECT 78.125 0 78.295 0.93 ;
        RECT 77.135 0 77.305 0.93 ;
        RECT 63.66 0 76.97 0.305 ;
        RECT 74.395 0 74.565 0.935 ;
        RECT 73.135 0 73.33 1.585 ;
        RECT 64.59 0 73.33 1.58 ;
        RECT 72.56 0 72.73 2.08 ;
        RECT 71.62 0 71.79 2.08 ;
        RECT 71.465 0 71.79 1.585 ;
        RECT 70.66 0 70.83 2.08 ;
        RECT 69.615 0 69.81 1.595 ;
        RECT 68.74 0 68.91 2.08 ;
        RECT 67.78 0 67.95 2.08 ;
        RECT 65.86 0 66.135 1.595 ;
        RECT 65.86 0 66.03 2.08 ;
        RECT 62.865 0 63.035 0.93 ;
        RECT 61.875 0 62.045 0.93 ;
        RECT 48.4 0 61.71 0.305 ;
        RECT 59.135 0 59.305 0.935 ;
        RECT 57.875 0 58.07 1.585 ;
        RECT 49.33 0 58.07 1.58 ;
        RECT 57.3 0 57.47 2.08 ;
        RECT 56.36 0 56.53 2.08 ;
        RECT 56.205 0 56.53 1.585 ;
        RECT 55.4 0 55.57 2.08 ;
        RECT 54.355 0 54.55 1.595 ;
        RECT 53.48 0 53.65 2.08 ;
        RECT 52.52 0 52.69 2.08 ;
        RECT 50.6 0 50.875 1.595 ;
        RECT 50.6 0 50.77 2.08 ;
        RECT 47.605 0 47.775 0.93 ;
        RECT 46.615 0 46.785 0.93 ;
        RECT 33.14 0 46.45 0.305 ;
        RECT 43.875 0 44.045 0.935 ;
        RECT 42.615 0 42.81 1.585 ;
        RECT 34.07 0 42.81 1.58 ;
        RECT 42.04 0 42.21 2.08 ;
        RECT 41.1 0 41.27 2.08 ;
        RECT 40.945 0 41.27 1.585 ;
        RECT 40.14 0 40.31 2.08 ;
        RECT 39.095 0 39.29 1.595 ;
        RECT 38.22 0 38.39 2.08 ;
        RECT 37.26 0 37.43 2.08 ;
        RECT 35.34 0 35.615 1.595 ;
        RECT 35.34 0 35.51 2.08 ;
        RECT 32.345 0 32.515 0.93 ;
        RECT 31.355 0 31.525 0.93 ;
        RECT 17.88 0 31.19 0.305 ;
        RECT 28.615 0 28.785 0.935 ;
        RECT 27.355 0 27.55 1.585 ;
        RECT 18.81 0 27.55 1.58 ;
        RECT 26.78 0 26.95 2.08 ;
        RECT 25.84 0 26.01 2.08 ;
        RECT 25.685 0 26.01 1.585 ;
        RECT 24.88 0 25.05 2.08 ;
        RECT 23.835 0 24.03 1.595 ;
        RECT 22.96 0 23.13 2.08 ;
        RECT 22 0 22.17 2.08 ;
        RECT 20.08 0 20.355 1.595 ;
        RECT 20.08 0 20.25 2.08 ;
        RECT 17.085 0 17.255 0.93 ;
        RECT 16.095 0 16.265 0.93 ;
        RECT 0.05 0.245 15.93 0.305 ;
        RECT 13.355 0 13.525 0.935 ;
        RECT 12.095 0 12.29 1.585 ;
        RECT 3.55 0 12.29 1.58 ;
        RECT 11.52 0 11.69 2.08 ;
        RECT 10.58 0 10.75 2.08 ;
        RECT 10.425 0 10.75 1.585 ;
        RECT 9.62 0 9.79 2.08 ;
        RECT 8.575 0 8.77 1.595 ;
        RECT 7.7 0 7.87 2.08 ;
        RECT 6.74 0 6.91 2.08 ;
        RECT 4.82 0 5.095 1.595 ;
        RECT 4.82 0 4.99 2.08 ;
        RECT 0.05 0.245 0.855 0.315 ;
        RECT 0.345 0.245 0.515 0.335 ;
        RECT 0.05 0 79.1 0.075 ;
        RECT 0.05 0 0.345 0.315 ;
        RECT 0.01 8.58 79.1 8.88 ;
        RECT 78.92 8.575 79.1 8.88 ;
        RECT 78.125 7.95 78.295 8.88 ;
        RECT 77.135 7.95 77.305 8.88 ;
        RECT 63.66 8.575 76.97 8.88 ;
        RECT 74.395 7.945 74.565 8.88 ;
        RECT 68.78 7.945 68.95 8.88 ;
        RECT 62.865 7.95 63.035 8.88 ;
        RECT 61.875 7.95 62.045 8.88 ;
        RECT 48.4 8.575 61.71 8.88 ;
        RECT 59.135 7.945 59.305 8.88 ;
        RECT 53.52 7.945 53.69 8.88 ;
        RECT 47.605 7.95 47.775 8.88 ;
        RECT 46.615 7.95 46.785 8.88 ;
        RECT 33.14 8.575 46.45 8.88 ;
        RECT 43.875 7.945 44.045 8.88 ;
        RECT 38.26 7.945 38.43 8.88 ;
        RECT 32.345 7.95 32.515 8.88 ;
        RECT 31.355 7.95 31.525 8.88 ;
        RECT 17.88 8.575 31.19 8.88 ;
        RECT 28.615 7.945 28.785 8.88 ;
        RECT 23 7.945 23.17 8.88 ;
        RECT 17.085 7.95 17.255 8.88 ;
        RECT 16.095 7.95 16.265 8.88 ;
        RECT 0.01 8.575 15.93 8.88 ;
        RECT 13.355 7.945 13.525 8.88 ;
        RECT 7.74 7.945 7.91 8.88 ;
        RECT 0.01 8.565 0.815 8.88 ;
        RECT 0.225 8.545 0.475 8.88 ;
        RECT 0.225 7.945 0.395 8.88 ;
        RECT 69.785 6.075 69.955 8.025 ;
        RECT 69.73 7.855 69.9 8.305 ;
        RECT 69.73 5.015 69.9 6.245 ;
        RECT 66.46 2.57 66.83 2.74 ;
        RECT 66.46 1.93 66.63 2.74 ;
        RECT 66.34 1.93 66.63 2.1 ;
        RECT 65.14 2.49 65.31 2.94 ;
        RECT 54.525 6.075 54.695 8.025 ;
        RECT 54.47 7.855 54.64 8.305 ;
        RECT 54.47 5.015 54.64 6.245 ;
        RECT 51.2 2.57 51.57 2.74 ;
        RECT 51.2 1.93 51.37 2.74 ;
        RECT 51.08 1.93 51.37 2.1 ;
        RECT 49.88 2.49 50.05 2.94 ;
        RECT 39.265 6.075 39.435 8.025 ;
        RECT 39.21 7.855 39.38 8.305 ;
        RECT 39.21 5.015 39.38 6.245 ;
        RECT 35.94 2.57 36.31 2.74 ;
        RECT 35.94 1.93 36.11 2.74 ;
        RECT 35.82 1.93 36.11 2.1 ;
        RECT 34.62 2.49 34.79 2.94 ;
        RECT 24.005 6.075 24.175 8.025 ;
        RECT 23.95 7.855 24.12 8.305 ;
        RECT 23.95 5.015 24.12 6.245 ;
        RECT 20.68 2.57 21.05 2.74 ;
        RECT 20.68 1.93 20.85 2.74 ;
        RECT 20.56 1.93 20.85 2.1 ;
        RECT 19.36 2.49 19.53 2.94 ;
        RECT 8.745 6.075 8.915 8.025 ;
        RECT 8.69 7.855 8.86 8.305 ;
        RECT 8.69 5.015 8.86 6.245 ;
        RECT 5.42 2.57 5.79 2.74 ;
        RECT 5.42 1.93 5.59 2.74 ;
        RECT 5.3 1.93 5.59 2.1 ;
        RECT 4.1 2.49 4.27 2.94 ;
      LAYER met1 ;
        RECT 78.92 0 79.1 0.305 ;
        RECT 0.05 0 79.1 0.3 ;
        RECT 63.66 0 76.97 0.305 ;
        RECT 64.59 0 73.33 1.74 ;
        RECT 66.28 1.9 66.57 2.13 ;
        RECT 65.39 1.95 66.57 2.09 ;
        RECT 65.575 1.89 65.98 2.15 ;
        RECT 65.575 0 65.865 2.15 ;
        RECT 65.15 2.37 65.77 2.51 ;
        RECT 65.63 0 65.77 2.51 ;
        RECT 65.39 1.95 65.77 2.21 ;
        RECT 65.08 2.74 65.37 2.97 ;
        RECT 65.15 2.37 65.29 2.97 ;
        RECT 48.4 0 61.71 0.305 ;
        RECT 49.33 0 58.07 1.74 ;
        RECT 51.02 1.9 51.31 2.13 ;
        RECT 50.13 1.95 51.31 2.09 ;
        RECT 50.315 1.89 50.72 2.15 ;
        RECT 50.315 0 50.605 2.15 ;
        RECT 49.89 2.37 50.51 2.51 ;
        RECT 50.37 0 50.51 2.51 ;
        RECT 50.13 1.95 50.51 2.21 ;
        RECT 49.82 2.74 50.11 2.97 ;
        RECT 49.89 2.37 50.03 2.97 ;
        RECT 33.14 0 46.45 0.305 ;
        RECT 34.07 0 42.81 1.74 ;
        RECT 35.76 1.9 36.05 2.13 ;
        RECT 34.87 1.95 36.05 2.09 ;
        RECT 35.055 1.89 35.46 2.15 ;
        RECT 35.055 0 35.345 2.15 ;
        RECT 34.63 2.37 35.25 2.51 ;
        RECT 35.11 0 35.25 2.51 ;
        RECT 34.87 1.95 35.25 2.21 ;
        RECT 34.56 2.74 34.85 2.97 ;
        RECT 34.63 2.37 34.77 2.97 ;
        RECT 17.88 0 31.19 0.305 ;
        RECT 18.81 0 27.55 1.74 ;
        RECT 20.5 1.9 20.79 2.13 ;
        RECT 19.61 1.95 20.79 2.09 ;
        RECT 19.795 1.89 20.2 2.15 ;
        RECT 19.795 0 20.085 2.15 ;
        RECT 19.37 2.37 19.99 2.51 ;
        RECT 19.85 0 19.99 2.51 ;
        RECT 19.61 1.95 19.99 2.21 ;
        RECT 19.3 2.74 19.59 2.97 ;
        RECT 19.37 2.37 19.51 2.97 ;
        RECT 0.05 0 15.93 0.305 ;
        RECT 3.55 0 12.29 1.74 ;
        RECT 5.24 1.9 5.53 2.13 ;
        RECT 4.35 1.95 5.53 2.09 ;
        RECT 4.535 1.89 4.94 2.15 ;
        RECT 4.535 0 4.825 2.15 ;
        RECT 4.11 2.37 4.73 2.51 ;
        RECT 4.59 0 4.73 2.51 ;
        RECT 4.35 1.95 4.73 2.21 ;
        RECT 4.04 2.74 4.33 2.97 ;
        RECT 4.11 2.37 4.25 2.97 ;
        RECT 0.05 0 0.855 0.315 ;
        RECT 0.255 0 0.605 0.335 ;
        RECT 0.01 8.58 79.1 8.88 ;
        RECT 78.92 8.575 79.1 8.88 ;
        RECT 63.66 8.575 76.97 8.88 ;
        RECT 69.725 6.285 70.015 6.515 ;
        RECT 69.56 6.315 69.73 8.88 ;
        RECT 69.555 6.315 70.015 6.485 ;
        RECT 48.4 8.575 61.71 8.88 ;
        RECT 54.465 6.285 54.755 6.515 ;
        RECT 54.3 6.315 54.47 8.88 ;
        RECT 54.295 6.315 54.755 6.485 ;
        RECT 33.14 8.575 46.45 8.88 ;
        RECT 39.205 6.285 39.495 6.515 ;
        RECT 39.04 6.315 39.21 8.88 ;
        RECT 39.035 6.315 39.495 6.485 ;
        RECT 17.88 8.575 31.19 8.88 ;
        RECT 23.945 6.285 24.235 6.515 ;
        RECT 23.78 6.315 23.95 8.88 ;
        RECT 23.775 6.315 24.235 6.485 ;
        RECT 0.01 8.575 15.93 8.88 ;
        RECT 8.685 6.285 8.975 6.515 ;
        RECT 8.52 6.315 8.69 8.88 ;
        RECT 8.515 6.315 8.975 6.485 ;
        RECT 0.01 8.565 0.815 8.88 ;
        RECT 0.215 8.545 0.565 8.88 ;
      LAYER via2 ;
        RECT 0.29 8.59 0.49 8.79 ;
        RECT 0.33 0.09 0.53 0.29 ;
        RECT 4.56 1.92 4.76 2.12 ;
        RECT 19.82 1.92 20.02 2.12 ;
        RECT 35.08 1.92 35.28 2.12 ;
        RECT 50.34 1.92 50.54 2.12 ;
        RECT 65.6 1.92 65.8 2.12 ;
      LAYER mcon ;
        RECT 0.305 8.605 0.475 8.775 ;
        RECT 0.985 8.605 1.155 8.775 ;
        RECT 1.665 8.605 1.835 8.775 ;
        RECT 2.345 8.605 2.515 8.775 ;
        RECT 4.1 2.77 4.27 2.94 ;
        RECT 5.3 1.93 5.47 2.1 ;
        RECT 7.82 8.605 7.99 8.775 ;
        RECT 8.5 8.605 8.67 8.775 ;
        RECT 8.745 6.315 8.915 6.485 ;
        RECT 9.18 8.605 9.35 8.775 ;
        RECT 9.86 8.605 10.03 8.775 ;
        RECT 13.435 8.605 13.605 8.775 ;
        RECT 13.435 0.105 13.605 0.275 ;
        RECT 14.115 8.605 14.285 8.775 ;
        RECT 14.115 0.105 14.285 0.275 ;
        RECT 14.795 8.605 14.965 8.775 ;
        RECT 14.795 0.105 14.965 0.275 ;
        RECT 15.475 8.605 15.645 8.775 ;
        RECT 15.475 0.105 15.645 0.275 ;
        RECT 16.175 8.61 16.345 8.78 ;
        RECT 16.175 0.1 16.345 0.27 ;
        RECT 17.165 8.61 17.335 8.78 ;
        RECT 17.165 0.1 17.335 0.27 ;
        RECT 19.36 2.77 19.53 2.94 ;
        RECT 20.56 1.93 20.73 2.1 ;
        RECT 23.08 8.605 23.25 8.775 ;
        RECT 23.76 8.605 23.93 8.775 ;
        RECT 24.005 6.315 24.175 6.485 ;
        RECT 24.44 8.605 24.61 8.775 ;
        RECT 25.12 8.605 25.29 8.775 ;
        RECT 28.695 8.605 28.865 8.775 ;
        RECT 28.695 0.105 28.865 0.275 ;
        RECT 29.375 8.605 29.545 8.775 ;
        RECT 29.375 0.105 29.545 0.275 ;
        RECT 30.055 8.605 30.225 8.775 ;
        RECT 30.055 0.105 30.225 0.275 ;
        RECT 30.735 8.605 30.905 8.775 ;
        RECT 30.735 0.105 30.905 0.275 ;
        RECT 31.435 8.61 31.605 8.78 ;
        RECT 31.435 0.1 31.605 0.27 ;
        RECT 32.425 8.61 32.595 8.78 ;
        RECT 32.425 0.1 32.595 0.27 ;
        RECT 34.62 2.77 34.79 2.94 ;
        RECT 35.82 1.93 35.99 2.1 ;
        RECT 38.34 8.605 38.51 8.775 ;
        RECT 39.02 8.605 39.19 8.775 ;
        RECT 39.265 6.315 39.435 6.485 ;
        RECT 39.7 8.605 39.87 8.775 ;
        RECT 40.38 8.605 40.55 8.775 ;
        RECT 43.955 8.605 44.125 8.775 ;
        RECT 43.955 0.105 44.125 0.275 ;
        RECT 44.635 8.605 44.805 8.775 ;
        RECT 44.635 0.105 44.805 0.275 ;
        RECT 45.315 8.605 45.485 8.775 ;
        RECT 45.315 0.105 45.485 0.275 ;
        RECT 45.995 8.605 46.165 8.775 ;
        RECT 45.995 0.105 46.165 0.275 ;
        RECT 46.695 8.61 46.865 8.78 ;
        RECT 46.695 0.1 46.865 0.27 ;
        RECT 47.685 8.61 47.855 8.78 ;
        RECT 47.685 0.1 47.855 0.27 ;
        RECT 49.88 2.77 50.05 2.94 ;
        RECT 51.08 1.93 51.25 2.1 ;
        RECT 53.6 8.605 53.77 8.775 ;
        RECT 54.28 8.605 54.45 8.775 ;
        RECT 54.525 6.315 54.695 6.485 ;
        RECT 54.96 8.605 55.13 8.775 ;
        RECT 55.64 8.605 55.81 8.775 ;
        RECT 59.215 8.605 59.385 8.775 ;
        RECT 59.215 0.105 59.385 0.275 ;
        RECT 59.895 8.605 60.065 8.775 ;
        RECT 59.895 0.105 60.065 0.275 ;
        RECT 60.575 8.605 60.745 8.775 ;
        RECT 60.575 0.105 60.745 0.275 ;
        RECT 61.255 8.605 61.425 8.775 ;
        RECT 61.255 0.105 61.425 0.275 ;
        RECT 61.955 8.61 62.125 8.78 ;
        RECT 61.955 0.1 62.125 0.27 ;
        RECT 62.945 8.61 63.115 8.78 ;
        RECT 62.945 0.1 63.115 0.27 ;
        RECT 65.14 2.77 65.31 2.94 ;
        RECT 66.34 1.93 66.51 2.1 ;
        RECT 68.86 8.605 69.03 8.775 ;
        RECT 69.54 8.605 69.71 8.775 ;
        RECT 69.785 6.315 69.955 6.485 ;
        RECT 70.22 8.605 70.39 8.775 ;
        RECT 70.9 8.605 71.07 8.775 ;
        RECT 74.475 8.605 74.645 8.775 ;
        RECT 74.475 0.105 74.645 0.275 ;
        RECT 75.155 8.605 75.325 8.775 ;
        RECT 75.155 0.105 75.325 0.275 ;
        RECT 75.835 8.605 76.005 8.775 ;
        RECT 75.835 0.105 76.005 0.275 ;
        RECT 76.515 8.605 76.685 8.775 ;
        RECT 76.515 0.105 76.685 0.275 ;
        RECT 77.215 8.61 77.385 8.78 ;
        RECT 77.215 0.1 77.385 0.27 ;
        RECT 78.205 8.61 78.375 8.78 ;
        RECT 78.205 0.1 78.375 0.27 ;
      LAYER via1 ;
        RECT 0.315 8.615 0.465 8.765 ;
        RECT 0.355 0.115 0.505 0.265 ;
        RECT 4.705 1.945 4.855 2.095 ;
        RECT 19.965 1.945 20.115 2.095 ;
        RECT 35.225 1.945 35.375 2.095 ;
        RECT 50.485 1.945 50.635 2.095 ;
        RECT 65.745 1.945 65.895 2.095 ;
    END
  END vssd1
  OBS
    LAYER met4 ;
      RECT 66.74 2.97 67.07 3.3 ;
      RECT 66.75 2.5 67.07 3.3 ;
      RECT 68.9 2.48 69.23 2.84 ;
      RECT 66.75 2.5 69.23 2.8 ;
      RECT 51.48 2.97 51.81 3.3 ;
      RECT 51.49 2.5 51.81 3.3 ;
      RECT 53.64 2.48 53.97 2.84 ;
      RECT 51.49 2.5 53.97 2.8 ;
      RECT 36.22 2.97 36.55 3.3 ;
      RECT 36.23 2.5 36.55 3.3 ;
      RECT 38.38 2.48 38.71 2.84 ;
      RECT 36.23 2.5 38.71 2.8 ;
      RECT 20.96 2.97 21.29 3.3 ;
      RECT 20.97 2.5 21.29 3.3 ;
      RECT 23.12 2.48 23.45 2.84 ;
      RECT 20.97 2.5 23.45 2.8 ;
      RECT 5.7 2.97 6.03 3.3 ;
      RECT 5.71 2.5 6.03 3.3 ;
      RECT 7.86 2.48 8.19 2.84 ;
      RECT 5.71 2.5 8.19 2.8 ;
    LAYER via3 ;
      RECT 68.96 2.57 69.16 2.77 ;
      RECT 66.8 3.04 67 3.24 ;
      RECT 53.7 2.57 53.9 2.77 ;
      RECT 51.54 3.04 51.74 3.24 ;
      RECT 38.44 2.57 38.64 2.77 ;
      RECT 36.28 3.04 36.48 3.24 ;
      RECT 23.18 2.57 23.38 2.77 ;
      RECT 21.02 3.04 21.22 3.24 ;
      RECT 7.92 2.57 8.12 2.77 ;
      RECT 5.76 3.04 5.96 3.24 ;
    LAYER met3 ;
      RECT 70.06 7.055 70.43 7.425 ;
      RECT 70.095 4.475 70.395 7.425 ;
      RECT 68.655 4.475 70.395 4.775 ;
      RECT 65.86 4.255 68.955 4.555 ;
      RECT 68.655 2.515 68.955 4.775 ;
      RECT 65.86 2.97 66.16 4.555 ;
      RECT 69.38 3.51 69.71 3.86 ;
      RECT 67.47 3.55 69.71 3.85 ;
      RECT 67.47 2.41 67.77 3.85 ;
      RECT 65.55 2.97 66.28 3.3 ;
      RECT 68.45 2.52 69.23 2.86 ;
      RECT 68.92 2.48 69.23 2.86 ;
      RECT 67.46 2.41 67.79 2.74 ;
      RECT 68.9 2.51 69.23 2.86 ;
      RECT 66.74 2.41 67.06 3.33 ;
      RECT 66.74 2.41 67.07 2.95 ;
      RECT 54.8 7.055 55.17 7.425 ;
      RECT 54.835 4.475 55.135 7.425 ;
      RECT 53.395 4.475 55.135 4.775 ;
      RECT 50.6 4.255 53.695 4.555 ;
      RECT 53.395 2.515 53.695 4.775 ;
      RECT 50.6 2.97 50.9 4.555 ;
      RECT 54.12 3.51 54.45 3.86 ;
      RECT 52.21 3.55 54.45 3.85 ;
      RECT 52.21 2.41 52.51 3.85 ;
      RECT 50.29 2.97 51.02 3.3 ;
      RECT 53.19 2.52 53.97 2.86 ;
      RECT 53.66 2.48 53.97 2.86 ;
      RECT 52.2 2.41 52.53 2.74 ;
      RECT 53.64 2.51 53.97 2.86 ;
      RECT 51.48 2.41 51.8 3.33 ;
      RECT 51.48 2.41 51.81 2.95 ;
      RECT 39.54 7.055 39.91 7.425 ;
      RECT 39.575 4.475 39.875 7.425 ;
      RECT 38.135 4.475 39.875 4.775 ;
      RECT 35.34 4.255 38.435 4.555 ;
      RECT 38.135 2.515 38.435 4.775 ;
      RECT 35.34 2.97 35.64 4.555 ;
      RECT 38.86 3.51 39.19 3.86 ;
      RECT 36.95 3.55 39.19 3.85 ;
      RECT 36.95 2.41 37.25 3.85 ;
      RECT 35.03 2.97 35.76 3.3 ;
      RECT 37.93 2.52 38.71 2.86 ;
      RECT 38.4 2.48 38.71 2.86 ;
      RECT 36.94 2.41 37.27 2.74 ;
      RECT 38.38 2.51 38.71 2.86 ;
      RECT 36.22 2.41 36.54 3.33 ;
      RECT 36.22 2.41 36.55 2.95 ;
      RECT 24.28 7.055 24.65 7.425 ;
      RECT 24.315 4.475 24.615 7.425 ;
      RECT 22.875 4.475 24.615 4.775 ;
      RECT 20.08 4.255 23.175 4.555 ;
      RECT 22.875 2.515 23.175 4.775 ;
      RECT 20.08 2.97 20.38 4.555 ;
      RECT 23.6 3.51 23.93 3.86 ;
      RECT 21.69 3.55 23.93 3.85 ;
      RECT 21.69 2.41 21.99 3.85 ;
      RECT 19.77 2.97 20.5 3.3 ;
      RECT 22.67 2.52 23.45 2.86 ;
      RECT 23.14 2.48 23.45 2.86 ;
      RECT 21.68 2.41 22.01 2.74 ;
      RECT 23.12 2.51 23.45 2.86 ;
      RECT 20.96 2.41 21.28 3.33 ;
      RECT 20.96 2.41 21.29 2.95 ;
      RECT 9.02 7.055 9.39 7.425 ;
      RECT 9.055 4.475 9.355 7.425 ;
      RECT 7.615 4.475 9.355 4.775 ;
      RECT 4.82 4.255 7.915 4.555 ;
      RECT 7.615 2.515 7.915 4.775 ;
      RECT 4.82 2.97 5.12 4.555 ;
      RECT 8.34 3.51 8.67 3.86 ;
      RECT 6.43 3.55 8.67 3.85 ;
      RECT 6.43 2.41 6.73 3.85 ;
      RECT 4.51 2.97 5.24 3.3 ;
      RECT 7.41 2.52 8.19 2.86 ;
      RECT 7.88 2.48 8.19 2.86 ;
      RECT 6.42 2.41 6.75 2.74 ;
      RECT 7.86 2.51 8.19 2.86 ;
      RECT 5.7 2.41 6.02 3.33 ;
      RECT 5.7 2.41 6.03 2.95 ;
      RECT 72.3 1.85 73.03 2.18 ;
      RECT 70.61 1.87 71.34 2.2 ;
      RECT 69.57 1.85 70.3 2.2 ;
      RECT 68.02 1.88 68.75 2.21 ;
      RECT 57.04 1.85 57.77 2.18 ;
      RECT 55.35 1.87 56.08 2.2 ;
      RECT 54.31 1.85 55.04 2.2 ;
      RECT 52.76 1.88 53.49 2.21 ;
      RECT 41.78 1.85 42.51 2.18 ;
      RECT 40.09 1.87 40.82 2.2 ;
      RECT 39.05 1.85 39.78 2.2 ;
      RECT 37.5 1.88 38.23 2.21 ;
      RECT 26.52 1.85 27.25 2.18 ;
      RECT 24.83 1.87 25.56 2.2 ;
      RECT 23.79 1.85 24.52 2.2 ;
      RECT 22.24 1.88 22.97 2.21 ;
      RECT 11.26 1.85 11.99 2.18 ;
      RECT 9.57 1.87 10.3 2.2 ;
      RECT 8.53 1.85 9.26 2.2 ;
      RECT 6.98 1.88 7.71 2.21 ;
    LAYER via2 ;
      RECT 72.53 1.92 72.73 2.12 ;
      RECT 70.67 1.93 70.87 2.13 ;
      RECT 70.145 7.14 70.345 7.34 ;
      RECT 69.65 1.94 69.85 2.14 ;
      RECT 69.44 3.57 69.64 3.77 ;
      RECT 68.96 2.57 69.16 2.77 ;
      RECT 68.21 1.94 68.41 2.14 ;
      RECT 67.52 2.48 67.72 2.68 ;
      RECT 66.81 2.48 67.01 2.68 ;
      RECT 65.84 3.04 66.04 3.24 ;
      RECT 57.27 1.92 57.47 2.12 ;
      RECT 55.41 1.93 55.61 2.13 ;
      RECT 54.885 7.14 55.085 7.34 ;
      RECT 54.39 1.94 54.59 2.14 ;
      RECT 54.18 3.57 54.38 3.77 ;
      RECT 53.7 2.57 53.9 2.77 ;
      RECT 52.95 1.94 53.15 2.14 ;
      RECT 52.26 2.48 52.46 2.68 ;
      RECT 51.55 2.48 51.75 2.68 ;
      RECT 50.58 3.04 50.78 3.24 ;
      RECT 42.01 1.92 42.21 2.12 ;
      RECT 40.15 1.93 40.35 2.13 ;
      RECT 39.625 7.14 39.825 7.34 ;
      RECT 39.13 1.94 39.33 2.14 ;
      RECT 38.92 3.57 39.12 3.77 ;
      RECT 38.44 2.57 38.64 2.77 ;
      RECT 37.69 1.94 37.89 2.14 ;
      RECT 37 2.48 37.2 2.68 ;
      RECT 36.29 2.48 36.49 2.68 ;
      RECT 35.32 3.04 35.52 3.24 ;
      RECT 26.75 1.92 26.95 2.12 ;
      RECT 24.89 1.93 25.09 2.13 ;
      RECT 24.365 7.14 24.565 7.34 ;
      RECT 23.87 1.94 24.07 2.14 ;
      RECT 23.66 3.57 23.86 3.77 ;
      RECT 23.18 2.57 23.38 2.77 ;
      RECT 22.43 1.94 22.63 2.14 ;
      RECT 21.74 2.48 21.94 2.68 ;
      RECT 21.03 2.48 21.23 2.68 ;
      RECT 20.06 3.04 20.26 3.24 ;
      RECT 11.49 1.92 11.69 2.12 ;
      RECT 9.63 1.93 9.83 2.13 ;
      RECT 9.105 7.14 9.305 7.34 ;
      RECT 8.61 1.94 8.81 2.14 ;
      RECT 8.4 3.57 8.6 3.77 ;
      RECT 7.92 2.57 8.12 2.77 ;
      RECT 7.17 1.94 7.37 2.14 ;
      RECT 6.48 2.48 6.68 2.68 ;
      RECT 5.77 2.48 5.97 2.68 ;
      RECT 4.8 3.04 5 3.24 ;
    LAYER met2 ;
      RECT 1.23 8.4 78.73 8.57 ;
      RECT 78.56 7.275 78.73 8.57 ;
      RECT 1.23 6.255 1.4 8.57 ;
      RECT 78.53 7.275 78.88 7.625 ;
      RECT 1.17 6.255 1.46 6.605 ;
      RECT 75.37 6.22 75.69 6.545 ;
      RECT 75.4 5.695 75.57 6.545 ;
      RECT 75.4 5.695 75.575 6.045 ;
      RECT 75.4 5.695 76.375 5.87 ;
      RECT 76.2 1.965 76.375 5.87 ;
      RECT 76.145 1.965 76.495 2.315 ;
      RECT 76.17 6.655 76.495 6.98 ;
      RECT 75.055 6.745 76.495 6.915 ;
      RECT 75.055 2.395 75.215 6.915 ;
      RECT 75.37 2.365 75.69 2.685 ;
      RECT 75.055 2.395 75.69 2.565 ;
      RECT 72.5 3.54 72.76 3.86 ;
      RECT 72.56 1.83 72.7 3.86 ;
      RECT 73.765 2.7 74.105 3.05 ;
      RECT 73.14 2.77 74.105 2.97 ;
      RECT 73.14 1.94 73.34 2.97 ;
      RECT 72.39 2.39 72.7 2.76 ;
      RECT 73.855 2.695 74.025 3.05 ;
      RECT 72.46 1.95 72.7 2.76 ;
      RECT 72.49 1.83 72.77 2.2 ;
      RECT 72.49 1.94 73.34 2.14 ;
      RECT 71.81 2.42 72.07 2.74 ;
      RECT 71.15 2.51 72.07 2.65 ;
      RECT 71.15 1.57 71.29 2.65 ;
      RECT 67.61 1.86 67.87 2.18 ;
      RECT 67.79 1.57 67.93 2.09 ;
      RECT 67.79 1.57 71.29 1.71 ;
      RECT 63.245 6.655 63.595 7.005 ;
      RECT 70.73 6.61 71.08 6.96 ;
      RECT 63.245 6.685 71.08 6.885 ;
      RECT 70.64 3.26 70.9 3.58 ;
      RECT 70.7 1.85 70.84 3.58 ;
      RECT 70.63 1.85 70.91 2.22 ;
      RECT 68.03 4.01 70.47 4.15 ;
      RECT 70.33 2.7 70.47 4.15 ;
      RECT 68.03 3.63 68.17 4.15 ;
      RECT 67.73 3.63 68.17 3.86 ;
      RECT 65.39 3.63 68.17 3.77 ;
      RECT 67.73 3.54 67.99 3.86 ;
      RECT 65.39 3.35 65.53 3.77 ;
      RECT 64.88 3.26 65.14 3.58 ;
      RECT 64.88 3.35 65.53 3.49 ;
      RECT 64.94 1.86 65.08 3.58 ;
      RECT 70.27 2.7 70.53 3.02 ;
      RECT 64.88 1.86 65.14 2.18 ;
      RECT 69.89 3.54 70.15 3.86 ;
      RECT 69.95 1.95 70.09 3.86 ;
      RECT 69.61 1.95 70.09 2.22 ;
      RECT 69.41 1.85 69.89 2.2 ;
      RECT 69.4 3.49 69.68 3.86 ;
      RECT 69.47 2.39 69.61 3.86 ;
      RECT 69.41 2.39 69.67 3.02 ;
      RECT 69.4 2.39 69.68 2.76 ;
      RECT 68.33 3.54 68.59 3.86 ;
      RECT 68.33 3.35 68.53 3.86 ;
      RECT 68.14 3.35 68.53 3.49 ;
      RECT 68.14 1.86 68.28 3.49 ;
      RECT 68.14 1.86 68.45 2.23 ;
      RECT 68.08 1.86 68.45 2.18 ;
      RECT 65.8 2.95 66.08 3.32 ;
      RECT 67.25 2.98 67.51 3.3 ;
      RECT 65.63 3.07 67.51 3.21 ;
      RECT 65.63 2.95 66.08 3.21 ;
      RECT 65.57 2.39 65.83 3.02 ;
      RECT 65.56 2.39 65.84 2.76 ;
      RECT 66.64 2.39 67.05 2.76 ;
      RECT 66.05 2.42 66.31 2.74 ;
      RECT 66.05 2.51 67.05 2.65 ;
      RECT 60.11 6.22 60.43 6.545 ;
      RECT 60.14 5.695 60.31 6.545 ;
      RECT 60.14 5.695 60.315 6.045 ;
      RECT 60.14 5.695 61.115 5.87 ;
      RECT 60.94 1.965 61.115 5.87 ;
      RECT 60.885 1.965 61.235 2.315 ;
      RECT 60.91 6.655 61.235 6.98 ;
      RECT 59.795 6.745 61.235 6.915 ;
      RECT 59.795 2.395 59.955 6.915 ;
      RECT 60.11 2.365 60.43 2.685 ;
      RECT 59.795 2.395 60.43 2.565 ;
      RECT 57.24 3.54 57.5 3.86 ;
      RECT 57.3 1.83 57.44 3.86 ;
      RECT 58.505 2.7 58.845 3.05 ;
      RECT 57.88 2.77 58.845 2.97 ;
      RECT 57.88 1.94 58.08 2.97 ;
      RECT 57.13 2.39 57.44 2.76 ;
      RECT 58.595 2.695 58.765 3.05 ;
      RECT 57.2 1.95 57.44 2.76 ;
      RECT 57.23 1.83 57.51 2.2 ;
      RECT 57.23 1.94 58.08 2.14 ;
      RECT 56.55 2.42 56.81 2.74 ;
      RECT 55.89 2.51 56.81 2.65 ;
      RECT 55.89 1.57 56.03 2.65 ;
      RECT 52.35 1.86 52.61 2.18 ;
      RECT 52.53 1.57 52.67 2.09 ;
      RECT 52.53 1.57 56.03 1.71 ;
      RECT 47.985 6.655 48.335 7.005 ;
      RECT 55.475 6.61 55.825 6.96 ;
      RECT 47.985 6.685 55.825 6.885 ;
      RECT 55.38 3.26 55.64 3.58 ;
      RECT 55.44 1.85 55.58 3.58 ;
      RECT 55.37 1.85 55.65 2.22 ;
      RECT 52.77 4.01 55.21 4.15 ;
      RECT 55.07 2.7 55.21 4.15 ;
      RECT 52.77 3.63 52.91 4.15 ;
      RECT 52.47 3.63 52.91 3.86 ;
      RECT 50.13 3.63 52.91 3.77 ;
      RECT 52.47 3.54 52.73 3.86 ;
      RECT 50.13 3.35 50.27 3.77 ;
      RECT 49.62 3.26 49.88 3.58 ;
      RECT 49.62 3.35 50.27 3.49 ;
      RECT 49.68 1.86 49.82 3.58 ;
      RECT 55.01 2.7 55.27 3.02 ;
      RECT 49.62 1.86 49.88 2.18 ;
      RECT 54.63 3.54 54.89 3.86 ;
      RECT 54.69 1.95 54.83 3.86 ;
      RECT 54.35 1.95 54.83 2.22 ;
      RECT 54.15 1.85 54.63 2.2 ;
      RECT 54.14 3.49 54.42 3.86 ;
      RECT 54.21 2.39 54.35 3.86 ;
      RECT 54.15 2.39 54.41 3.02 ;
      RECT 54.14 2.39 54.42 2.76 ;
      RECT 53.07 3.54 53.33 3.86 ;
      RECT 53.07 3.35 53.27 3.86 ;
      RECT 52.88 3.35 53.27 3.49 ;
      RECT 52.88 1.86 53.02 3.49 ;
      RECT 52.88 1.86 53.19 2.23 ;
      RECT 52.82 1.86 53.19 2.18 ;
      RECT 50.54 2.95 50.82 3.32 ;
      RECT 51.99 2.98 52.25 3.3 ;
      RECT 50.37 3.07 52.25 3.21 ;
      RECT 50.37 2.95 50.82 3.21 ;
      RECT 50.31 2.39 50.57 3.02 ;
      RECT 50.3 2.39 50.58 2.76 ;
      RECT 51.38 2.39 51.79 2.76 ;
      RECT 50.79 2.42 51.05 2.74 ;
      RECT 50.79 2.51 51.79 2.65 ;
      RECT 44.85 6.22 45.17 6.545 ;
      RECT 44.88 5.695 45.05 6.545 ;
      RECT 44.88 5.695 45.055 6.045 ;
      RECT 44.88 5.695 45.855 5.87 ;
      RECT 45.68 1.965 45.855 5.87 ;
      RECT 45.625 1.965 45.975 2.315 ;
      RECT 45.65 6.655 45.975 6.98 ;
      RECT 44.535 6.745 45.975 6.915 ;
      RECT 44.535 2.395 44.695 6.915 ;
      RECT 44.85 2.365 45.17 2.685 ;
      RECT 44.535 2.395 45.17 2.565 ;
      RECT 41.98 3.54 42.24 3.86 ;
      RECT 42.04 1.83 42.18 3.86 ;
      RECT 43.245 2.7 43.585 3.05 ;
      RECT 42.62 2.77 43.585 2.97 ;
      RECT 42.62 1.94 42.82 2.97 ;
      RECT 41.87 2.39 42.18 2.76 ;
      RECT 43.335 2.695 43.505 3.05 ;
      RECT 41.94 1.95 42.18 2.76 ;
      RECT 41.97 1.83 42.25 2.2 ;
      RECT 41.97 1.94 42.82 2.14 ;
      RECT 41.29 2.42 41.55 2.74 ;
      RECT 40.63 2.51 41.55 2.65 ;
      RECT 40.63 1.57 40.77 2.65 ;
      RECT 37.09 1.86 37.35 2.18 ;
      RECT 37.27 1.57 37.41 2.09 ;
      RECT 37.27 1.57 40.77 1.71 ;
      RECT 32.77 6.66 33.12 7.01 ;
      RECT 40.21 6.615 40.56 6.965 ;
      RECT 32.77 6.69 40.56 6.89 ;
      RECT 40.12 3.26 40.38 3.58 ;
      RECT 40.18 1.85 40.32 3.58 ;
      RECT 40.11 1.85 40.39 2.22 ;
      RECT 37.51 4.01 39.95 4.15 ;
      RECT 39.81 2.7 39.95 4.15 ;
      RECT 37.51 3.63 37.65 4.15 ;
      RECT 37.21 3.63 37.65 3.86 ;
      RECT 34.87 3.63 37.65 3.77 ;
      RECT 37.21 3.54 37.47 3.86 ;
      RECT 34.87 3.35 35.01 3.77 ;
      RECT 34.36 3.26 34.62 3.58 ;
      RECT 34.36 3.35 35.01 3.49 ;
      RECT 34.42 1.86 34.56 3.58 ;
      RECT 39.75 2.7 40.01 3.02 ;
      RECT 34.36 1.86 34.62 2.18 ;
      RECT 39.37 3.54 39.63 3.86 ;
      RECT 39.43 1.95 39.57 3.86 ;
      RECT 39.09 1.95 39.57 2.22 ;
      RECT 38.89 1.85 39.37 2.2 ;
      RECT 38.88 3.49 39.16 3.86 ;
      RECT 38.95 2.39 39.09 3.86 ;
      RECT 38.89 2.39 39.15 3.02 ;
      RECT 38.88 2.39 39.16 2.76 ;
      RECT 37.81 3.54 38.07 3.86 ;
      RECT 37.81 3.35 38.01 3.86 ;
      RECT 37.62 3.35 38.01 3.49 ;
      RECT 37.62 1.86 37.76 3.49 ;
      RECT 37.62 1.86 37.93 2.23 ;
      RECT 37.56 1.86 37.93 2.18 ;
      RECT 35.28 2.95 35.56 3.32 ;
      RECT 36.73 2.98 36.99 3.3 ;
      RECT 35.11 3.07 36.99 3.21 ;
      RECT 35.11 2.95 35.56 3.21 ;
      RECT 35.05 2.39 35.31 3.02 ;
      RECT 35.04 2.39 35.32 2.76 ;
      RECT 36.12 2.39 36.53 2.76 ;
      RECT 35.53 2.42 35.79 2.74 ;
      RECT 35.53 2.51 36.53 2.65 ;
      RECT 29.59 6.22 29.91 6.545 ;
      RECT 29.62 5.695 29.79 6.545 ;
      RECT 29.62 5.695 29.795 6.045 ;
      RECT 29.62 5.695 30.595 5.87 ;
      RECT 30.42 1.965 30.595 5.87 ;
      RECT 30.365 1.965 30.715 2.315 ;
      RECT 30.39 6.655 30.715 6.98 ;
      RECT 29.275 6.745 30.715 6.915 ;
      RECT 29.275 2.395 29.435 6.915 ;
      RECT 29.59 2.365 29.91 2.685 ;
      RECT 29.275 2.395 29.91 2.565 ;
      RECT 26.72 3.54 26.98 3.86 ;
      RECT 26.78 1.83 26.92 3.86 ;
      RECT 27.985 2.7 28.325 3.05 ;
      RECT 27.36 2.77 28.325 2.97 ;
      RECT 27.36 1.94 27.56 2.97 ;
      RECT 26.61 2.39 26.92 2.76 ;
      RECT 28.075 2.695 28.245 3.05 ;
      RECT 26.68 1.95 26.92 2.76 ;
      RECT 26.71 1.83 26.99 2.2 ;
      RECT 26.71 1.94 27.56 2.14 ;
      RECT 26.03 2.42 26.29 2.74 ;
      RECT 25.37 2.51 26.29 2.65 ;
      RECT 25.37 1.57 25.51 2.65 ;
      RECT 21.83 1.86 22.09 2.18 ;
      RECT 22.01 1.57 22.15 2.09 ;
      RECT 22.01 1.57 25.51 1.71 ;
      RECT 17.51 6.655 17.86 7.005 ;
      RECT 24.95 6.61 25.3 6.96 ;
      RECT 17.51 6.685 25.3 6.885 ;
      RECT 24.86 3.26 25.12 3.58 ;
      RECT 24.92 1.85 25.06 3.58 ;
      RECT 24.85 1.85 25.13 2.22 ;
      RECT 22.25 4.01 24.69 4.15 ;
      RECT 24.55 2.7 24.69 4.15 ;
      RECT 22.25 3.63 22.39 4.15 ;
      RECT 21.95 3.63 22.39 3.86 ;
      RECT 19.61 3.63 22.39 3.77 ;
      RECT 21.95 3.54 22.21 3.86 ;
      RECT 19.61 3.35 19.75 3.77 ;
      RECT 19.1 3.26 19.36 3.58 ;
      RECT 19.1 3.35 19.75 3.49 ;
      RECT 19.16 1.86 19.3 3.58 ;
      RECT 24.49 2.7 24.75 3.02 ;
      RECT 19.1 1.86 19.36 2.18 ;
      RECT 24.11 3.54 24.37 3.86 ;
      RECT 24.17 1.95 24.31 3.86 ;
      RECT 23.83 1.95 24.31 2.22 ;
      RECT 23.63 1.85 24.11 2.2 ;
      RECT 23.62 3.49 23.9 3.86 ;
      RECT 23.69 2.39 23.83 3.86 ;
      RECT 23.63 2.39 23.89 3.02 ;
      RECT 23.62 2.39 23.9 2.76 ;
      RECT 22.55 3.54 22.81 3.86 ;
      RECT 22.55 3.35 22.75 3.86 ;
      RECT 22.36 3.35 22.75 3.49 ;
      RECT 22.36 1.86 22.5 3.49 ;
      RECT 22.36 1.86 22.67 2.23 ;
      RECT 22.3 1.86 22.67 2.18 ;
      RECT 20.02 2.95 20.3 3.32 ;
      RECT 21.47 2.98 21.73 3.3 ;
      RECT 19.85 3.07 21.73 3.21 ;
      RECT 19.85 2.95 20.3 3.21 ;
      RECT 19.79 2.39 20.05 3.02 ;
      RECT 19.78 2.39 20.06 2.76 ;
      RECT 20.86 2.39 21.27 2.76 ;
      RECT 20.27 2.42 20.53 2.74 ;
      RECT 20.27 2.51 21.27 2.65 ;
      RECT 14.33 6.22 14.65 6.545 ;
      RECT 14.36 5.695 14.53 6.545 ;
      RECT 14.36 5.695 14.535 6.045 ;
      RECT 14.36 5.695 15.335 5.87 ;
      RECT 15.16 1.965 15.335 5.87 ;
      RECT 15.105 1.965 15.455 2.315 ;
      RECT 15.13 6.655 15.455 6.98 ;
      RECT 14.015 6.745 15.455 6.915 ;
      RECT 14.015 2.395 14.175 6.915 ;
      RECT 14.33 2.365 14.65 2.685 ;
      RECT 14.015 2.395 14.65 2.565 ;
      RECT 11.46 3.54 11.72 3.86 ;
      RECT 11.52 1.83 11.66 3.86 ;
      RECT 12.725 2.7 13.065 3.05 ;
      RECT 12.1 2.77 13.065 2.97 ;
      RECT 12.1 1.94 12.3 2.97 ;
      RECT 11.35 2.39 11.66 2.76 ;
      RECT 12.815 2.695 12.985 3.05 ;
      RECT 11.42 1.95 11.66 2.76 ;
      RECT 11.45 1.83 11.73 2.2 ;
      RECT 11.45 1.94 12.3 2.14 ;
      RECT 10.77 2.42 11.03 2.74 ;
      RECT 10.11 2.51 11.03 2.65 ;
      RECT 10.11 1.57 10.25 2.65 ;
      RECT 6.57 1.86 6.83 2.18 ;
      RECT 6.75 1.57 6.89 2.09 ;
      RECT 6.75 1.57 10.25 1.71 ;
      RECT 1.545 6.995 1.835 7.345 ;
      RECT 1.545 7.065 2.765 7.235 ;
      RECT 2.595 6.685 2.765 7.235 ;
      RECT 9.69 6.605 10.04 6.955 ;
      RECT 2.595 6.685 10.04 6.855 ;
      RECT 9.6 3.26 9.86 3.58 ;
      RECT 9.66 1.85 9.8 3.58 ;
      RECT 9.59 1.85 9.87 2.22 ;
      RECT 6.99 4.01 9.43 4.15 ;
      RECT 9.29 2.7 9.43 4.15 ;
      RECT 6.99 3.63 7.13 4.15 ;
      RECT 6.69 3.63 7.13 3.86 ;
      RECT 4.35 3.63 7.13 3.77 ;
      RECT 6.69 3.54 6.95 3.86 ;
      RECT 4.35 3.35 4.49 3.77 ;
      RECT 3.84 3.26 4.1 3.58 ;
      RECT 3.84 3.35 4.49 3.49 ;
      RECT 3.9 1.86 4.04 3.58 ;
      RECT 9.23 2.7 9.49 3.02 ;
      RECT 3.84 1.86 4.1 2.18 ;
      RECT 8.85 3.54 9.11 3.86 ;
      RECT 8.91 1.95 9.05 3.86 ;
      RECT 8.57 1.95 9.05 2.22 ;
      RECT 8.37 1.85 8.85 2.2 ;
      RECT 8.36 3.49 8.64 3.86 ;
      RECT 8.43 2.39 8.57 3.86 ;
      RECT 8.37 2.39 8.63 3.02 ;
      RECT 8.36 2.39 8.64 2.76 ;
      RECT 7.29 3.54 7.55 3.86 ;
      RECT 7.29 3.35 7.49 3.86 ;
      RECT 7.1 3.35 7.49 3.49 ;
      RECT 7.1 1.86 7.24 3.49 ;
      RECT 7.1 1.86 7.41 2.23 ;
      RECT 7.04 1.86 7.41 2.18 ;
      RECT 4.76 2.95 5.04 3.32 ;
      RECT 6.21 2.98 6.47 3.3 ;
      RECT 4.59 3.07 6.47 3.21 ;
      RECT 4.59 2.95 5.04 3.21 ;
      RECT 4.53 2.39 4.79 3.02 ;
      RECT 4.52 2.39 4.8 2.76 ;
      RECT 5.6 2.39 6.01 2.76 ;
      RECT 5.01 2.42 5.27 2.74 ;
      RECT 5.01 2.51 6.01 2.65 ;
      RECT 70.06 7.055 70.43 7.425 ;
      RECT 68.92 2.39 69.2 2.86 ;
      RECT 68.68 1.86 68.96 2.2 ;
      RECT 67.48 2.39 67.76 2.76 ;
      RECT 64.925 1.215 65.295 1.22 ;
      RECT 54.8 7.055 55.17 7.425 ;
      RECT 53.66 2.39 53.94 2.86 ;
      RECT 53.42 1.86 53.7 2.2 ;
      RECT 52.22 2.39 52.5 2.76 ;
      RECT 49.665 1.215 50.035 1.22 ;
      RECT 39.54 7.055 39.91 7.425 ;
      RECT 38.4 2.39 38.68 2.86 ;
      RECT 38.16 1.86 38.44 2.2 ;
      RECT 36.96 2.39 37.24 2.76 ;
      RECT 34.405 1.215 34.775 1.22 ;
      RECT 24.28 7.055 24.65 7.425 ;
      RECT 23.14 2.39 23.42 2.86 ;
      RECT 22.9 1.86 23.18 2.2 ;
      RECT 21.7 2.39 21.98 2.76 ;
      RECT 19.145 1.215 19.515 1.22 ;
      RECT 9.02 7.055 9.39 7.425 ;
      RECT 7.88 2.39 8.16 2.86 ;
      RECT 7.64 1.86 7.92 2.2 ;
      RECT 6.44 2.39 6.72 2.76 ;
      RECT 3.885 1.215 4.255 1.22 ;
    LAYER via1 ;
      RECT 78.63 7.375 78.78 7.525 ;
      RECT 76.26 6.74 76.41 6.89 ;
      RECT 76.245 2.065 76.395 2.215 ;
      RECT 75.455 2.45 75.605 2.6 ;
      RECT 75.455 6.325 75.605 6.475 ;
      RECT 73.865 2.8 74.015 2.95 ;
      RECT 72.555 1.945 72.705 2.095 ;
      RECT 72.555 3.625 72.705 3.775 ;
      RECT 71.865 2.505 72.015 2.655 ;
      RECT 70.83 6.71 70.98 6.86 ;
      RECT 70.695 1.945 70.845 2.095 ;
      RECT 70.695 3.345 70.845 3.495 ;
      RECT 70.325 2.785 70.475 2.935 ;
      RECT 70.17 7.165 70.32 7.315 ;
      RECT 69.945 3.625 70.095 3.775 ;
      RECT 69.465 1.945 69.615 2.095 ;
      RECT 69.465 2.785 69.615 2.935 ;
      RECT 68.985 2.505 69.135 2.655 ;
      RECT 68.745 1.945 68.895 2.095 ;
      RECT 68.385 3.625 68.535 3.775 ;
      RECT 68.135 1.945 68.285 2.095 ;
      RECT 67.785 3.625 67.935 3.775 ;
      RECT 67.665 1.945 67.815 2.095 ;
      RECT 67.545 2.505 67.695 2.655 ;
      RECT 67.305 3.065 67.455 3.215 ;
      RECT 66.105 2.505 66.255 2.655 ;
      RECT 65.625 2.785 65.775 2.935 ;
      RECT 64.935 1.945 65.085 2.095 ;
      RECT 64.935 3.345 65.085 3.495 ;
      RECT 63.345 6.755 63.495 6.905 ;
      RECT 61 6.74 61.15 6.89 ;
      RECT 60.985 2.065 61.135 2.215 ;
      RECT 60.195 2.45 60.345 2.6 ;
      RECT 60.195 6.325 60.345 6.475 ;
      RECT 58.605 2.8 58.755 2.95 ;
      RECT 57.295 1.945 57.445 2.095 ;
      RECT 57.295 3.625 57.445 3.775 ;
      RECT 56.605 2.505 56.755 2.655 ;
      RECT 55.575 6.71 55.725 6.86 ;
      RECT 55.435 1.945 55.585 2.095 ;
      RECT 55.435 3.345 55.585 3.495 ;
      RECT 55.065 2.785 55.215 2.935 ;
      RECT 54.91 7.165 55.06 7.315 ;
      RECT 54.685 3.625 54.835 3.775 ;
      RECT 54.205 1.945 54.355 2.095 ;
      RECT 54.205 2.785 54.355 2.935 ;
      RECT 53.725 2.505 53.875 2.655 ;
      RECT 53.485 1.945 53.635 2.095 ;
      RECT 53.125 3.625 53.275 3.775 ;
      RECT 52.875 1.945 53.025 2.095 ;
      RECT 52.525 3.625 52.675 3.775 ;
      RECT 52.405 1.945 52.555 2.095 ;
      RECT 52.285 2.505 52.435 2.655 ;
      RECT 52.045 3.065 52.195 3.215 ;
      RECT 50.845 2.505 50.995 2.655 ;
      RECT 50.365 2.785 50.515 2.935 ;
      RECT 49.675 1.945 49.825 2.095 ;
      RECT 49.675 3.345 49.825 3.495 ;
      RECT 48.085 6.755 48.235 6.905 ;
      RECT 45.74 6.74 45.89 6.89 ;
      RECT 45.725 2.065 45.875 2.215 ;
      RECT 44.935 2.45 45.085 2.6 ;
      RECT 44.935 6.325 45.085 6.475 ;
      RECT 43.345 2.8 43.495 2.95 ;
      RECT 42.035 1.945 42.185 2.095 ;
      RECT 42.035 3.625 42.185 3.775 ;
      RECT 41.345 2.505 41.495 2.655 ;
      RECT 40.31 6.715 40.46 6.865 ;
      RECT 40.175 1.945 40.325 2.095 ;
      RECT 40.175 3.345 40.325 3.495 ;
      RECT 39.805 2.785 39.955 2.935 ;
      RECT 39.65 7.165 39.8 7.315 ;
      RECT 39.425 3.625 39.575 3.775 ;
      RECT 38.945 1.945 39.095 2.095 ;
      RECT 38.945 2.785 39.095 2.935 ;
      RECT 38.465 2.505 38.615 2.655 ;
      RECT 38.225 1.945 38.375 2.095 ;
      RECT 37.865 3.625 38.015 3.775 ;
      RECT 37.615 1.945 37.765 2.095 ;
      RECT 37.265 3.625 37.415 3.775 ;
      RECT 37.145 1.945 37.295 2.095 ;
      RECT 37.025 2.505 37.175 2.655 ;
      RECT 36.785 3.065 36.935 3.215 ;
      RECT 35.585 2.505 35.735 2.655 ;
      RECT 35.105 2.785 35.255 2.935 ;
      RECT 34.415 1.945 34.565 2.095 ;
      RECT 34.415 3.345 34.565 3.495 ;
      RECT 32.87 6.76 33.02 6.91 ;
      RECT 30.48 6.74 30.63 6.89 ;
      RECT 30.465 2.065 30.615 2.215 ;
      RECT 29.675 2.45 29.825 2.6 ;
      RECT 29.675 6.325 29.825 6.475 ;
      RECT 28.085 2.8 28.235 2.95 ;
      RECT 26.775 1.945 26.925 2.095 ;
      RECT 26.775 3.625 26.925 3.775 ;
      RECT 26.085 2.505 26.235 2.655 ;
      RECT 25.05 6.71 25.2 6.86 ;
      RECT 24.915 1.945 25.065 2.095 ;
      RECT 24.915 3.345 25.065 3.495 ;
      RECT 24.545 2.785 24.695 2.935 ;
      RECT 24.39 7.165 24.54 7.315 ;
      RECT 24.165 3.625 24.315 3.775 ;
      RECT 23.685 1.945 23.835 2.095 ;
      RECT 23.685 2.785 23.835 2.935 ;
      RECT 23.205 2.505 23.355 2.655 ;
      RECT 22.965 1.945 23.115 2.095 ;
      RECT 22.605 3.625 22.755 3.775 ;
      RECT 22.355 1.945 22.505 2.095 ;
      RECT 22.005 3.625 22.155 3.775 ;
      RECT 21.885 1.945 22.035 2.095 ;
      RECT 21.765 2.505 21.915 2.655 ;
      RECT 21.525 3.065 21.675 3.215 ;
      RECT 20.325 2.505 20.475 2.655 ;
      RECT 19.845 2.785 19.995 2.935 ;
      RECT 19.155 1.945 19.305 2.095 ;
      RECT 19.155 3.345 19.305 3.495 ;
      RECT 17.61 6.755 17.76 6.905 ;
      RECT 15.22 6.74 15.37 6.89 ;
      RECT 15.205 2.065 15.355 2.215 ;
      RECT 14.415 2.45 14.565 2.6 ;
      RECT 14.415 6.325 14.565 6.475 ;
      RECT 12.825 2.8 12.975 2.95 ;
      RECT 11.515 1.945 11.665 2.095 ;
      RECT 11.515 3.625 11.665 3.775 ;
      RECT 10.825 2.505 10.975 2.655 ;
      RECT 9.79 6.705 9.94 6.855 ;
      RECT 9.655 1.945 9.805 2.095 ;
      RECT 9.655 3.345 9.805 3.495 ;
      RECT 9.285 2.785 9.435 2.935 ;
      RECT 9.13 7.165 9.28 7.315 ;
      RECT 8.905 3.625 9.055 3.775 ;
      RECT 8.425 1.945 8.575 2.095 ;
      RECT 8.425 2.785 8.575 2.935 ;
      RECT 7.945 2.505 8.095 2.655 ;
      RECT 7.705 1.945 7.855 2.095 ;
      RECT 7.345 3.625 7.495 3.775 ;
      RECT 7.095 1.945 7.245 2.095 ;
      RECT 6.745 3.625 6.895 3.775 ;
      RECT 6.625 1.945 6.775 2.095 ;
      RECT 6.505 2.505 6.655 2.655 ;
      RECT 6.265 3.065 6.415 3.215 ;
      RECT 5.065 2.505 5.215 2.655 ;
      RECT 4.585 2.785 4.735 2.935 ;
      RECT 3.895 1.945 4.045 2.095 ;
      RECT 3.895 3.345 4.045 3.495 ;
      RECT 1.615 7.095 1.765 7.245 ;
      RECT 1.24 6.355 1.39 6.505 ;
    LAYER met1 ;
      RECT 78.495 7.77 78.785 8 ;
      RECT 78.555 6.29 78.725 8 ;
      RECT 78.53 7.275 78.88 7.625 ;
      RECT 78.495 6.29 78.785 6.52 ;
      RECT 78.09 2.395 78.195 2.965 ;
      RECT 78.09 2.73 78.415 2.96 ;
      RECT 78.09 2.76 78.585 2.93 ;
      RECT 78.09 2.395 78.28 2.96 ;
      RECT 77.505 2.36 77.795 2.59 ;
      RECT 77.505 2.395 78.28 2.565 ;
      RECT 77.565 0.88 77.735 2.59 ;
      RECT 77.505 0.88 77.795 1.11 ;
      RECT 77.505 7.77 77.795 8 ;
      RECT 77.565 6.29 77.735 8 ;
      RECT 77.505 6.29 77.795 6.52 ;
      RECT 77.505 6.325 78.36 6.485 ;
      RECT 78.19 5.92 78.36 6.485 ;
      RECT 77.505 6.32 77.9 6.485 ;
      RECT 78.125 5.92 78.415 6.15 ;
      RECT 78.125 5.95 78.585 6.12 ;
      RECT 77.135 2.73 77.425 2.96 ;
      RECT 77.135 2.76 77.595 2.93 ;
      RECT 77.2 1.655 77.365 2.96 ;
      RECT 75.715 1.625 76.005 1.855 ;
      RECT 75.715 1.655 77.365 1.825 ;
      RECT 75.775 0.885 75.945 1.855 ;
      RECT 75.715 0.885 76.005 1.115 ;
      RECT 75.715 7.765 76.005 7.995 ;
      RECT 75.775 7.025 75.945 7.995 ;
      RECT 75.775 7.12 77.365 7.29 ;
      RECT 77.195 5.92 77.365 7.29 ;
      RECT 75.715 7.025 76.005 7.255 ;
      RECT 77.135 5.92 77.425 6.15 ;
      RECT 77.135 5.95 77.595 6.12 ;
      RECT 73.765 2.7 74.105 3.05 ;
      RECT 73.855 2.025 74.025 3.05 ;
      RECT 76.145 1.965 76.495 2.315 ;
      RECT 73.855 2.025 76.495 2.195 ;
      RECT 76.17 6.655 76.495 6.98 ;
      RECT 70.73 6.61 71.08 6.96 ;
      RECT 76.145 6.655 76.495 6.885 ;
      RECT 70.53 6.655 71.08 6.885 ;
      RECT 70.36 6.685 76.495 6.855 ;
      RECT 75.37 2.365 75.69 2.685 ;
      RECT 75.34 2.365 75.69 2.595 ;
      RECT 75.17 2.395 75.69 2.565 ;
      RECT 75.37 6.255 75.69 6.545 ;
      RECT 75.34 6.285 75.69 6.515 ;
      RECT 75.17 6.315 75.69 6.485 ;
      RECT 72.47 1.89 72.79 2.15 ;
      RECT 72.04 1.9 72.33 2.13 ;
      RECT 72.04 1.95 72.79 2.09 ;
      RECT 72.47 3.57 72.79 3.83 ;
      RECT 72.04 3.58 72.33 3.81 ;
      RECT 72.04 3.63 72.79 3.77 ;
      RECT 71.8 3.02 72.09 3.25 ;
      RECT 71.8 3.07 72.37 3.21 ;
      RECT 72.23 2.93 72.49 3.07 ;
      RECT 72.28 2.74 72.57 2.97 ;
      RECT 70.43 2.93 71.53 3.07 ;
      RECT 70.24 2.73 70.56 2.99 ;
      RECT 71.32 2.74 71.61 2.97 ;
      RECT 70.24 2.74 70.65 2.99 ;
      RECT 70.61 1.89 70.93 2.15 ;
      RECT 71.08 1.9 71.37 2.13 ;
      RECT 70.61 1.95 71.37 2.09 ;
      RECT 67.91 3.15 70.09 3.29 ;
      RECT 69.95 2.16 70.09 3.29 ;
      RECT 67.91 3.07 69.21 3.29 ;
      RECT 68.92 3.02 69.21 3.29 ;
      RECT 67.91 2.79 68.25 3.29 ;
      RECT 67.96 2.74 68.25 3.29 ;
      RECT 70.84 2.46 71.13 2.69 ;
      RECT 69.95 2.37 71.05 2.51 ;
      RECT 69.88 2.16 70.17 2.41 ;
      RECT 70.1 7.765 70.39 7.995 ;
      RECT 70.16 7.025 70.33 7.995 ;
      RECT 70.06 7.055 70.43 7.425 ;
      RECT 70.1 7.025 70.39 7.425 ;
      RECT 69.86 3.57 70.18 3.83 ;
      RECT 69.86 3.58 70.38 3.81 ;
      RECT 68.44 2.46 68.73 2.69 ;
      RECT 68.59 2.07 68.73 2.69 ;
      RECT 68.59 2.07 68.89 2.21 ;
      RECT 69.38 1.89 69.7 2.15 ;
      RECT 68.66 1.89 68.98 2.15 ;
      RECT 69.16 1.9 69.7 2.13 ;
      RECT 68.66 1.95 69.7 2.09 ;
      RECT 68.3 3.57 68.62 3.83 ;
      RECT 68.2 3.58 68.62 3.81 ;
      RECT 66.28 3.02 66.57 3.25 ;
      RECT 66.28 3.02 66.73 3.21 ;
      RECT 66.59 2.55 66.73 3.21 ;
      RECT 66.71 1.95 66.85 2.69 ;
      RECT 67.58 1.89 67.9 2.15 ;
      RECT 66.76 1.9 67.05 2.13 ;
      RECT 66.71 1.95 67.9 2.09 ;
      RECT 67.46 2.45 67.78 2.71 ;
      RECT 67 2.46 67.29 2.69 ;
      RECT 67 2.51 67.78 2.65 ;
      RECT 67.22 3.01 67.54 3.27 ;
      RECT 67.22 3.02 67.77 3.25 ;
      RECT 66.76 3.58 67.05 3.81 ;
      RECT 65.87 3.46 66.97 3.6 ;
      RECT 65.8 3.3 66.09 3.53 ;
      RECT 63.235 7.77 63.525 8 ;
      RECT 63.295 6.29 63.465 8 ;
      RECT 63.245 6.655 63.595 7.005 ;
      RECT 63.235 6.29 63.525 6.52 ;
      RECT 62.83 2.395 62.935 2.965 ;
      RECT 62.83 2.73 63.155 2.96 ;
      RECT 62.83 2.76 63.325 2.93 ;
      RECT 62.83 2.395 63.02 2.96 ;
      RECT 62.245 2.36 62.535 2.59 ;
      RECT 62.245 2.395 63.02 2.565 ;
      RECT 62.305 0.88 62.475 2.59 ;
      RECT 62.245 0.88 62.535 1.11 ;
      RECT 62.245 7.77 62.535 8 ;
      RECT 62.305 6.29 62.475 8 ;
      RECT 62.245 6.29 62.535 6.52 ;
      RECT 62.245 6.325 63.1 6.485 ;
      RECT 62.93 5.92 63.1 6.485 ;
      RECT 62.245 6.32 62.64 6.485 ;
      RECT 62.865 5.92 63.155 6.15 ;
      RECT 62.865 5.95 63.325 6.12 ;
      RECT 61.875 2.73 62.165 2.96 ;
      RECT 61.875 2.76 62.335 2.93 ;
      RECT 61.94 1.655 62.105 2.96 ;
      RECT 60.455 1.625 60.745 1.855 ;
      RECT 60.455 1.655 62.105 1.825 ;
      RECT 60.515 0.885 60.685 1.855 ;
      RECT 60.455 0.885 60.745 1.115 ;
      RECT 60.455 7.765 60.745 7.995 ;
      RECT 60.515 7.025 60.685 7.995 ;
      RECT 60.515 7.12 62.105 7.29 ;
      RECT 61.935 5.92 62.105 7.29 ;
      RECT 60.455 7.025 60.745 7.255 ;
      RECT 61.875 5.92 62.165 6.15 ;
      RECT 61.875 5.95 62.335 6.12 ;
      RECT 58.505 2.7 58.845 3.05 ;
      RECT 58.595 2.025 58.765 3.05 ;
      RECT 60.885 1.965 61.235 2.315 ;
      RECT 58.595 2.025 61.235 2.195 ;
      RECT 60.91 6.655 61.235 6.98 ;
      RECT 55.475 6.61 55.825 6.96 ;
      RECT 60.885 6.655 61.235 6.885 ;
      RECT 55.27 6.655 55.825 6.885 ;
      RECT 55.1 6.685 61.235 6.855 ;
      RECT 60.11 2.365 60.43 2.685 ;
      RECT 60.08 2.365 60.43 2.595 ;
      RECT 59.91 2.395 60.43 2.565 ;
      RECT 60.11 6.255 60.43 6.545 ;
      RECT 60.08 6.285 60.43 6.515 ;
      RECT 59.91 6.315 60.43 6.485 ;
      RECT 57.21 1.89 57.53 2.15 ;
      RECT 56.78 1.9 57.07 2.13 ;
      RECT 56.78 1.95 57.53 2.09 ;
      RECT 57.21 3.57 57.53 3.83 ;
      RECT 56.78 3.58 57.07 3.81 ;
      RECT 56.78 3.63 57.53 3.77 ;
      RECT 56.54 3.02 56.83 3.25 ;
      RECT 56.54 3.07 57.11 3.21 ;
      RECT 56.97 2.93 57.23 3.07 ;
      RECT 57.02 2.74 57.31 2.97 ;
      RECT 55.17 2.93 56.27 3.07 ;
      RECT 54.98 2.73 55.3 2.99 ;
      RECT 56.06 2.74 56.35 2.97 ;
      RECT 54.98 2.74 55.39 2.99 ;
      RECT 55.35 1.89 55.67 2.15 ;
      RECT 55.82 1.9 56.11 2.13 ;
      RECT 55.35 1.95 56.11 2.09 ;
      RECT 52.65 3.15 54.83 3.29 ;
      RECT 54.69 2.16 54.83 3.29 ;
      RECT 52.65 3.07 53.95 3.29 ;
      RECT 53.66 3.02 53.95 3.29 ;
      RECT 52.65 2.79 52.99 3.29 ;
      RECT 52.7 2.74 52.99 3.29 ;
      RECT 55.58 2.46 55.87 2.69 ;
      RECT 54.69 2.37 55.79 2.51 ;
      RECT 54.62 2.16 54.91 2.41 ;
      RECT 54.84 7.765 55.13 7.995 ;
      RECT 54.9 7.025 55.07 7.995 ;
      RECT 54.8 7.055 55.17 7.425 ;
      RECT 54.84 7.025 55.13 7.425 ;
      RECT 54.6 3.57 54.92 3.83 ;
      RECT 54.6 3.58 55.12 3.81 ;
      RECT 53.18 2.46 53.47 2.69 ;
      RECT 53.33 2.07 53.47 2.69 ;
      RECT 53.33 2.07 53.63 2.21 ;
      RECT 54.12 1.89 54.44 2.15 ;
      RECT 53.4 1.89 53.72 2.15 ;
      RECT 53.9 1.9 54.44 2.13 ;
      RECT 53.4 1.95 54.44 2.09 ;
      RECT 53.04 3.57 53.36 3.83 ;
      RECT 52.94 3.58 53.36 3.81 ;
      RECT 51.02 3.02 51.31 3.25 ;
      RECT 51.02 3.02 51.47 3.21 ;
      RECT 51.33 2.55 51.47 3.21 ;
      RECT 51.45 1.95 51.59 2.69 ;
      RECT 52.32 1.89 52.64 2.15 ;
      RECT 51.5 1.9 51.79 2.13 ;
      RECT 51.45 1.95 52.64 2.09 ;
      RECT 52.2 2.45 52.52 2.71 ;
      RECT 51.74 2.46 52.03 2.69 ;
      RECT 51.74 2.51 52.52 2.65 ;
      RECT 51.96 3.01 52.28 3.27 ;
      RECT 51.96 3.02 52.51 3.25 ;
      RECT 51.5 3.58 51.79 3.81 ;
      RECT 50.61 3.46 51.71 3.6 ;
      RECT 50.54 3.3 50.83 3.53 ;
      RECT 47.975 7.77 48.265 8 ;
      RECT 48.035 6.29 48.205 8 ;
      RECT 47.985 6.655 48.335 7.005 ;
      RECT 47.975 6.29 48.265 6.52 ;
      RECT 47.57 2.395 47.675 2.965 ;
      RECT 47.57 2.73 47.895 2.96 ;
      RECT 47.57 2.76 48.065 2.93 ;
      RECT 47.57 2.395 47.76 2.96 ;
      RECT 46.985 2.36 47.275 2.59 ;
      RECT 46.985 2.395 47.76 2.565 ;
      RECT 47.045 0.88 47.215 2.59 ;
      RECT 46.985 0.88 47.275 1.11 ;
      RECT 46.985 7.77 47.275 8 ;
      RECT 47.045 6.29 47.215 8 ;
      RECT 46.985 6.29 47.275 6.52 ;
      RECT 46.985 6.325 47.84 6.485 ;
      RECT 47.67 5.92 47.84 6.485 ;
      RECT 46.985 6.32 47.38 6.485 ;
      RECT 47.605 5.92 47.895 6.15 ;
      RECT 47.605 5.95 48.065 6.12 ;
      RECT 46.615 2.73 46.905 2.96 ;
      RECT 46.615 2.76 47.075 2.93 ;
      RECT 46.68 1.655 46.845 2.96 ;
      RECT 45.195 1.625 45.485 1.855 ;
      RECT 45.195 1.655 46.845 1.825 ;
      RECT 45.255 0.885 45.425 1.855 ;
      RECT 45.195 0.885 45.485 1.115 ;
      RECT 45.195 7.765 45.485 7.995 ;
      RECT 45.255 7.025 45.425 7.995 ;
      RECT 45.255 7.12 46.845 7.29 ;
      RECT 46.675 5.92 46.845 7.29 ;
      RECT 45.195 7.025 45.485 7.255 ;
      RECT 46.615 5.92 46.905 6.15 ;
      RECT 46.615 5.95 47.075 6.12 ;
      RECT 43.245 2.7 43.585 3.05 ;
      RECT 43.335 2.025 43.505 3.05 ;
      RECT 45.625 1.965 45.975 2.315 ;
      RECT 43.335 2.025 45.975 2.195 ;
      RECT 45.65 6.655 45.975 6.98 ;
      RECT 40.21 6.615 40.56 6.965 ;
      RECT 45.625 6.655 45.975 6.885 ;
      RECT 40.01 6.655 40.56 6.885 ;
      RECT 39.84 6.685 45.975 6.855 ;
      RECT 44.85 2.365 45.17 2.685 ;
      RECT 44.82 2.365 45.17 2.595 ;
      RECT 44.65 2.395 45.17 2.565 ;
      RECT 44.85 6.255 45.17 6.545 ;
      RECT 44.82 6.285 45.17 6.515 ;
      RECT 44.65 6.315 45.17 6.485 ;
      RECT 41.95 1.89 42.27 2.15 ;
      RECT 41.52 1.9 41.81 2.13 ;
      RECT 41.52 1.95 42.27 2.09 ;
      RECT 41.95 3.57 42.27 3.83 ;
      RECT 41.52 3.58 41.81 3.81 ;
      RECT 41.52 3.63 42.27 3.77 ;
      RECT 41.28 3.02 41.57 3.25 ;
      RECT 41.28 3.07 41.85 3.21 ;
      RECT 41.71 2.93 41.97 3.07 ;
      RECT 41.76 2.74 42.05 2.97 ;
      RECT 39.91 2.93 41.01 3.07 ;
      RECT 39.72 2.73 40.04 2.99 ;
      RECT 40.8 2.74 41.09 2.97 ;
      RECT 39.72 2.74 40.13 2.99 ;
      RECT 40.09 1.89 40.41 2.15 ;
      RECT 40.56 1.9 40.85 2.13 ;
      RECT 40.09 1.95 40.85 2.09 ;
      RECT 37.39 3.15 39.57 3.29 ;
      RECT 39.43 2.16 39.57 3.29 ;
      RECT 37.39 3.07 38.69 3.29 ;
      RECT 38.4 3.02 38.69 3.29 ;
      RECT 37.39 2.79 37.73 3.29 ;
      RECT 37.44 2.74 37.73 3.29 ;
      RECT 40.32 2.46 40.61 2.69 ;
      RECT 39.43 2.37 40.53 2.51 ;
      RECT 39.36 2.16 39.65 2.41 ;
      RECT 39.58 7.765 39.87 7.995 ;
      RECT 39.64 7.025 39.81 7.995 ;
      RECT 39.54 7.055 39.91 7.425 ;
      RECT 39.58 7.025 39.87 7.425 ;
      RECT 39.34 3.57 39.66 3.83 ;
      RECT 39.34 3.58 39.86 3.81 ;
      RECT 37.92 2.46 38.21 2.69 ;
      RECT 38.07 2.07 38.21 2.69 ;
      RECT 38.07 2.07 38.37 2.21 ;
      RECT 38.86 1.89 39.18 2.15 ;
      RECT 38.14 1.89 38.46 2.15 ;
      RECT 38.64 1.9 39.18 2.13 ;
      RECT 38.14 1.95 39.18 2.09 ;
      RECT 37.78 3.57 38.1 3.83 ;
      RECT 37.68 3.58 38.1 3.81 ;
      RECT 35.76 3.02 36.05 3.25 ;
      RECT 35.76 3.02 36.21 3.21 ;
      RECT 36.07 2.55 36.21 3.21 ;
      RECT 36.19 1.95 36.33 2.69 ;
      RECT 37.06 1.89 37.38 2.15 ;
      RECT 36.24 1.9 36.53 2.13 ;
      RECT 36.19 1.95 37.38 2.09 ;
      RECT 36.94 2.45 37.26 2.71 ;
      RECT 36.48 2.46 36.77 2.69 ;
      RECT 36.48 2.51 37.26 2.65 ;
      RECT 36.7 3.01 37.02 3.27 ;
      RECT 36.7 3.02 37.25 3.25 ;
      RECT 36.24 3.58 36.53 3.81 ;
      RECT 35.35 3.46 36.45 3.6 ;
      RECT 35.28 3.3 35.57 3.53 ;
      RECT 32.715 7.77 33.005 8 ;
      RECT 32.775 6.29 32.945 8 ;
      RECT 32.765 6.66 33.12 7.015 ;
      RECT 32.715 6.29 33.005 6.52 ;
      RECT 32.31 2.395 32.415 2.965 ;
      RECT 32.31 2.73 32.635 2.96 ;
      RECT 32.31 2.76 32.805 2.93 ;
      RECT 32.31 2.395 32.5 2.96 ;
      RECT 31.725 2.36 32.015 2.59 ;
      RECT 31.725 2.395 32.5 2.565 ;
      RECT 31.785 0.88 31.955 2.59 ;
      RECT 31.725 0.88 32.015 1.11 ;
      RECT 31.725 7.77 32.015 8 ;
      RECT 31.785 6.29 31.955 8 ;
      RECT 31.725 6.29 32.015 6.52 ;
      RECT 31.725 6.325 32.58 6.485 ;
      RECT 32.41 5.92 32.58 6.485 ;
      RECT 31.725 6.32 32.12 6.485 ;
      RECT 32.345 5.92 32.635 6.15 ;
      RECT 32.345 5.95 32.805 6.12 ;
      RECT 31.355 2.73 31.645 2.96 ;
      RECT 31.355 2.76 31.815 2.93 ;
      RECT 31.42 1.655 31.585 2.96 ;
      RECT 29.935 1.625 30.225 1.855 ;
      RECT 29.935 1.655 31.585 1.825 ;
      RECT 29.995 0.885 30.165 1.855 ;
      RECT 29.935 0.885 30.225 1.115 ;
      RECT 29.935 7.765 30.225 7.995 ;
      RECT 29.995 7.025 30.165 7.995 ;
      RECT 29.995 7.12 31.585 7.29 ;
      RECT 31.415 5.92 31.585 7.29 ;
      RECT 29.935 7.025 30.225 7.255 ;
      RECT 31.355 5.92 31.645 6.15 ;
      RECT 31.355 5.95 31.815 6.12 ;
      RECT 27.985 2.7 28.325 3.05 ;
      RECT 28.075 2.025 28.245 3.05 ;
      RECT 30.365 1.965 30.715 2.315 ;
      RECT 28.075 2.025 30.715 2.195 ;
      RECT 30.39 6.655 30.715 6.98 ;
      RECT 24.95 6.61 25.3 6.96 ;
      RECT 30.365 6.655 30.715 6.885 ;
      RECT 24.75 6.655 25.3 6.885 ;
      RECT 24.58 6.685 30.715 6.855 ;
      RECT 29.59 2.365 29.91 2.685 ;
      RECT 29.56 2.365 29.91 2.595 ;
      RECT 29.39 2.395 29.91 2.565 ;
      RECT 29.59 6.255 29.91 6.545 ;
      RECT 29.56 6.285 29.91 6.515 ;
      RECT 29.39 6.315 29.91 6.485 ;
      RECT 26.69 1.89 27.01 2.15 ;
      RECT 26.26 1.9 26.55 2.13 ;
      RECT 26.26 1.95 27.01 2.09 ;
      RECT 26.69 3.57 27.01 3.83 ;
      RECT 26.26 3.58 26.55 3.81 ;
      RECT 26.26 3.63 27.01 3.77 ;
      RECT 26.02 3.02 26.31 3.25 ;
      RECT 26.02 3.07 26.59 3.21 ;
      RECT 26.45 2.93 26.71 3.07 ;
      RECT 26.5 2.74 26.79 2.97 ;
      RECT 24.65 2.93 25.75 3.07 ;
      RECT 24.46 2.73 24.78 2.99 ;
      RECT 25.54 2.74 25.83 2.97 ;
      RECT 24.46 2.74 24.87 2.99 ;
      RECT 24.83 1.89 25.15 2.15 ;
      RECT 25.3 1.9 25.59 2.13 ;
      RECT 24.83 1.95 25.59 2.09 ;
      RECT 22.13 3.15 24.31 3.29 ;
      RECT 24.17 2.16 24.31 3.29 ;
      RECT 22.13 3.07 23.43 3.29 ;
      RECT 23.14 3.02 23.43 3.29 ;
      RECT 22.13 2.79 22.47 3.29 ;
      RECT 22.18 2.74 22.47 3.29 ;
      RECT 25.06 2.46 25.35 2.69 ;
      RECT 24.17 2.37 25.27 2.51 ;
      RECT 24.1 2.16 24.39 2.41 ;
      RECT 24.32 7.765 24.61 7.995 ;
      RECT 24.38 7.025 24.55 7.995 ;
      RECT 24.28 7.055 24.65 7.425 ;
      RECT 24.32 7.025 24.61 7.425 ;
      RECT 24.08 3.57 24.4 3.83 ;
      RECT 24.08 3.58 24.6 3.81 ;
      RECT 22.66 2.46 22.95 2.69 ;
      RECT 22.81 2.07 22.95 2.69 ;
      RECT 22.81 2.07 23.11 2.21 ;
      RECT 23.6 1.89 23.92 2.15 ;
      RECT 22.88 1.89 23.2 2.15 ;
      RECT 23.38 1.9 23.92 2.13 ;
      RECT 22.88 1.95 23.92 2.09 ;
      RECT 22.52 3.57 22.84 3.83 ;
      RECT 22.42 3.58 22.84 3.81 ;
      RECT 20.5 3.02 20.79 3.25 ;
      RECT 20.5 3.02 20.95 3.21 ;
      RECT 20.81 2.55 20.95 3.21 ;
      RECT 20.93 1.95 21.07 2.69 ;
      RECT 21.8 1.89 22.12 2.15 ;
      RECT 20.98 1.9 21.27 2.13 ;
      RECT 20.93 1.95 22.12 2.09 ;
      RECT 21.68 2.45 22 2.71 ;
      RECT 21.22 2.46 21.51 2.69 ;
      RECT 21.22 2.51 22 2.65 ;
      RECT 21.44 3.01 21.76 3.27 ;
      RECT 21.44 3.02 21.99 3.25 ;
      RECT 20.98 3.58 21.27 3.81 ;
      RECT 20.09 3.46 21.19 3.6 ;
      RECT 20.02 3.3 20.31 3.53 ;
      RECT 17.455 7.77 17.745 8 ;
      RECT 17.515 6.29 17.685 8 ;
      RECT 17.51 6.655 17.86 7.005 ;
      RECT 17.455 6.29 17.745 6.52 ;
      RECT 17.05 2.395 17.155 2.965 ;
      RECT 17.05 2.73 17.375 2.96 ;
      RECT 17.05 2.76 17.545 2.93 ;
      RECT 17.05 2.395 17.24 2.96 ;
      RECT 16.465 2.36 16.755 2.59 ;
      RECT 16.465 2.395 17.24 2.565 ;
      RECT 16.525 0.88 16.695 2.59 ;
      RECT 16.465 0.88 16.755 1.11 ;
      RECT 16.465 7.77 16.755 8 ;
      RECT 16.525 6.29 16.695 8 ;
      RECT 16.465 6.29 16.755 6.52 ;
      RECT 16.465 6.325 17.32 6.485 ;
      RECT 17.15 5.92 17.32 6.485 ;
      RECT 16.465 6.32 16.86 6.485 ;
      RECT 17.085 5.92 17.375 6.15 ;
      RECT 17.085 5.95 17.545 6.12 ;
      RECT 16.095 2.73 16.385 2.96 ;
      RECT 16.095 2.76 16.555 2.93 ;
      RECT 16.16 1.655 16.325 2.96 ;
      RECT 14.675 1.625 14.965 1.855 ;
      RECT 14.675 1.655 16.325 1.825 ;
      RECT 14.735 0.885 14.905 1.855 ;
      RECT 14.675 0.885 14.965 1.115 ;
      RECT 14.675 7.765 14.965 7.995 ;
      RECT 14.735 7.025 14.905 7.995 ;
      RECT 14.735 7.12 16.325 7.29 ;
      RECT 16.155 5.92 16.325 7.29 ;
      RECT 14.675 7.025 14.965 7.255 ;
      RECT 16.095 5.92 16.385 6.15 ;
      RECT 16.095 5.95 16.555 6.12 ;
      RECT 12.725 2.7 13.065 3.05 ;
      RECT 12.815 2.025 12.985 3.05 ;
      RECT 15.105 1.965 15.455 2.315 ;
      RECT 12.815 2.025 15.455 2.195 ;
      RECT 15.13 6.655 15.455 6.98 ;
      RECT 9.69 6.605 10.04 6.955 ;
      RECT 15.105 6.655 15.455 6.885 ;
      RECT 9.49 6.655 10.04 6.885 ;
      RECT 9.32 6.685 15.455 6.855 ;
      RECT 14.33 2.365 14.65 2.685 ;
      RECT 14.3 2.365 14.65 2.595 ;
      RECT 14.13 2.395 14.65 2.565 ;
      RECT 14.33 6.255 14.65 6.545 ;
      RECT 14.3 6.285 14.65 6.515 ;
      RECT 14.13 6.315 14.65 6.485 ;
      RECT 11.43 1.89 11.75 2.15 ;
      RECT 11 1.9 11.29 2.13 ;
      RECT 11 1.95 11.75 2.09 ;
      RECT 11.43 3.57 11.75 3.83 ;
      RECT 11 3.58 11.29 3.81 ;
      RECT 11 3.63 11.75 3.77 ;
      RECT 10.76 3.02 11.05 3.25 ;
      RECT 10.76 3.07 11.33 3.21 ;
      RECT 11.19 2.93 11.45 3.07 ;
      RECT 11.24 2.74 11.53 2.97 ;
      RECT 9.39 2.93 10.49 3.07 ;
      RECT 9.2 2.73 9.52 2.99 ;
      RECT 10.28 2.74 10.57 2.97 ;
      RECT 9.2 2.74 9.61 2.99 ;
      RECT 9.57 1.89 9.89 2.15 ;
      RECT 10.04 1.9 10.33 2.13 ;
      RECT 9.57 1.95 10.33 2.09 ;
      RECT 6.87 3.15 9.05 3.29 ;
      RECT 8.91 2.16 9.05 3.29 ;
      RECT 6.87 3.07 8.17 3.29 ;
      RECT 7.88 3.02 8.17 3.29 ;
      RECT 6.87 2.79 7.21 3.29 ;
      RECT 6.92 2.74 7.21 3.29 ;
      RECT 9.8 2.46 10.09 2.69 ;
      RECT 8.91 2.37 10.01 2.51 ;
      RECT 8.84 2.16 9.13 2.41 ;
      RECT 9.06 7.765 9.35 7.995 ;
      RECT 9.12 7.025 9.29 7.995 ;
      RECT 9.02 7.055 9.39 7.425 ;
      RECT 9.06 7.025 9.35 7.425 ;
      RECT 8.82 3.57 9.14 3.83 ;
      RECT 8.82 3.58 9.34 3.81 ;
      RECT 7.4 2.46 7.69 2.69 ;
      RECT 7.55 2.07 7.69 2.69 ;
      RECT 7.55 2.07 7.85 2.21 ;
      RECT 8.34 1.89 8.66 2.15 ;
      RECT 7.62 1.89 7.94 2.15 ;
      RECT 8.12 1.9 8.66 2.13 ;
      RECT 7.62 1.95 8.66 2.09 ;
      RECT 7.26 3.57 7.58 3.83 ;
      RECT 7.16 3.58 7.58 3.81 ;
      RECT 5.24 3.02 5.53 3.25 ;
      RECT 5.24 3.02 5.69 3.21 ;
      RECT 5.55 2.55 5.69 3.21 ;
      RECT 5.67 1.95 5.81 2.69 ;
      RECT 6.54 1.89 6.86 2.15 ;
      RECT 5.72 1.9 6.01 2.13 ;
      RECT 5.67 1.95 6.86 2.09 ;
      RECT 6.42 2.45 6.74 2.71 ;
      RECT 5.96 2.46 6.25 2.69 ;
      RECT 5.96 2.51 6.74 2.65 ;
      RECT 6.18 3.01 6.5 3.27 ;
      RECT 6.18 3.02 6.73 3.25 ;
      RECT 5.72 3.58 6.01 3.81 ;
      RECT 4.83 3.46 5.93 3.6 ;
      RECT 4.76 3.3 5.05 3.53 ;
      RECT 1.545 7.765 1.835 7.995 ;
      RECT 1.605 7.025 1.775 7.995 ;
      RECT 1.515 7.025 1.865 7.315 ;
      RECT 1.14 6.285 1.49 6.575 ;
      RECT 1 6.315 1.49 6.485 ;
      RECT 71.78 2.45 72.1 2.71 ;
      RECT 70.61 3.29 70.93 3.55 ;
      RECT 69.38 2.73 69.7 2.99 ;
      RECT 68.9 2.45 69.22 2.71 ;
      RECT 68.05 1.89 68.45 2.15 ;
      RECT 67.7 3.57 68.02 3.83 ;
      RECT 66.02 2.45 66.34 2.71 ;
      RECT 65.54 2.73 65.86 2.99 ;
      RECT 64.85 1.89 65.17 2.15 ;
      RECT 64.85 3.29 65.17 3.55 ;
      RECT 56.52 2.45 56.84 2.71 ;
      RECT 55.35 3.29 55.67 3.55 ;
      RECT 54.12 2.73 54.44 2.99 ;
      RECT 53.64 2.45 53.96 2.71 ;
      RECT 52.79 1.89 53.19 2.15 ;
      RECT 52.44 3.57 52.76 3.83 ;
      RECT 50.76 2.45 51.08 2.71 ;
      RECT 50.28 2.73 50.6 2.99 ;
      RECT 49.59 1.89 49.91 2.15 ;
      RECT 49.59 3.29 49.91 3.55 ;
      RECT 41.26 2.45 41.58 2.71 ;
      RECT 40.09 3.29 40.41 3.55 ;
      RECT 38.86 2.73 39.18 2.99 ;
      RECT 38.38 2.45 38.7 2.71 ;
      RECT 37.53 1.89 37.93 2.15 ;
      RECT 37.18 3.57 37.5 3.83 ;
      RECT 35.5 2.45 35.82 2.71 ;
      RECT 35.02 2.73 35.34 2.99 ;
      RECT 34.33 1.89 34.65 2.15 ;
      RECT 34.33 3.29 34.65 3.55 ;
      RECT 26 2.45 26.32 2.71 ;
      RECT 24.83 3.29 25.15 3.55 ;
      RECT 23.6 2.73 23.92 2.99 ;
      RECT 23.12 2.45 23.44 2.71 ;
      RECT 22.27 1.89 22.67 2.15 ;
      RECT 21.92 3.57 22.24 3.83 ;
      RECT 20.24 2.45 20.56 2.71 ;
      RECT 19.76 2.73 20.08 2.99 ;
      RECT 19.07 1.89 19.39 2.15 ;
      RECT 19.07 3.29 19.39 3.55 ;
      RECT 10.74 2.45 11.06 2.71 ;
      RECT 9.57 3.29 9.89 3.55 ;
      RECT 8.34 2.73 8.66 2.99 ;
      RECT 7.86 2.45 8.18 2.71 ;
      RECT 7.01 1.89 7.41 2.15 ;
      RECT 6.66 3.57 6.98 3.83 ;
      RECT 4.98 2.45 5.3 2.71 ;
      RECT 4.5 2.73 4.82 2.99 ;
      RECT 3.81 1.89 4.13 2.15 ;
      RECT 3.81 3.29 4.13 3.55 ;
    LAYER mcon ;
      RECT 78.555 6.32 78.725 6.49 ;
      RECT 78.56 6.315 78.73 6.485 ;
      RECT 63.295 6.32 63.465 6.49 ;
      RECT 63.3 6.315 63.47 6.485 ;
      RECT 48.035 6.32 48.205 6.49 ;
      RECT 48.04 6.315 48.21 6.485 ;
      RECT 32.775 6.32 32.945 6.49 ;
      RECT 32.78 6.315 32.95 6.485 ;
      RECT 17.515 6.32 17.685 6.49 ;
      RECT 17.52 6.315 17.69 6.485 ;
      RECT 78.555 7.8 78.725 7.97 ;
      RECT 78.185 2.76 78.355 2.93 ;
      RECT 78.185 5.95 78.355 6.12 ;
      RECT 77.565 0.91 77.735 1.08 ;
      RECT 77.565 2.39 77.735 2.56 ;
      RECT 77.565 6.32 77.735 6.49 ;
      RECT 77.565 7.8 77.735 7.97 ;
      RECT 77.195 2.76 77.365 2.93 ;
      RECT 77.195 5.95 77.365 6.12 ;
      RECT 76.205 2.025 76.375 2.195 ;
      RECT 76.205 6.685 76.375 6.855 ;
      RECT 75.775 0.915 75.945 1.085 ;
      RECT 75.775 1.655 75.945 1.825 ;
      RECT 75.775 7.055 75.945 7.225 ;
      RECT 75.775 7.795 75.945 7.965 ;
      RECT 75.4 2.395 75.57 2.565 ;
      RECT 75.4 6.315 75.57 6.485 ;
      RECT 72.34 2.77 72.51 2.94 ;
      RECT 72.1 1.93 72.27 2.1 ;
      RECT 72.1 3.61 72.27 3.78 ;
      RECT 71.86 2.49 72.03 2.66 ;
      RECT 71.86 3.05 72.03 3.22 ;
      RECT 71.38 2.77 71.55 2.94 ;
      RECT 71.14 1.93 71.31 2.1 ;
      RECT 70.9 2.49 71.07 2.66 ;
      RECT 70.69 3.33 70.86 3.5 ;
      RECT 70.59 6.685 70.76 6.855 ;
      RECT 70.42 2.77 70.59 2.94 ;
      RECT 70.16 7.055 70.33 7.225 ;
      RECT 70.16 7.795 70.33 7.965 ;
      RECT 70.15 3.61 70.32 3.78 ;
      RECT 69.94 2.19 70.11 2.36 ;
      RECT 69.46 2.77 69.63 2.94 ;
      RECT 69.22 1.93 69.39 2.1 ;
      RECT 68.98 2.49 69.15 2.66 ;
      RECT 68.98 3.05 69.15 3.22 ;
      RECT 68.5 2.49 68.67 2.66 ;
      RECT 68.26 3.61 68.43 3.78 ;
      RECT 68.22 1.93 68.39 2.1 ;
      RECT 68.02 2.77 68.19 2.94 ;
      RECT 67.78 3.61 67.95 3.78 ;
      RECT 67.54 3.05 67.71 3.22 ;
      RECT 67.06 2.49 67.23 2.66 ;
      RECT 66.82 1.93 66.99 2.1 ;
      RECT 66.82 3.61 66.99 3.78 ;
      RECT 66.34 3.05 66.51 3.22 ;
      RECT 66.1 2.49 66.27 2.66 ;
      RECT 65.86 3.33 66.03 3.5 ;
      RECT 65.62 2.77 65.79 2.94 ;
      RECT 64.93 1.93 65.1 2.1 ;
      RECT 64.93 3.33 65.1 3.5 ;
      RECT 63.295 7.8 63.465 7.97 ;
      RECT 62.925 2.76 63.095 2.93 ;
      RECT 62.925 5.95 63.095 6.12 ;
      RECT 62.305 0.91 62.475 1.08 ;
      RECT 62.305 2.39 62.475 2.56 ;
      RECT 62.305 6.32 62.475 6.49 ;
      RECT 62.305 7.8 62.475 7.97 ;
      RECT 61.935 2.76 62.105 2.93 ;
      RECT 61.935 5.95 62.105 6.12 ;
      RECT 60.945 2.025 61.115 2.195 ;
      RECT 60.945 6.685 61.115 6.855 ;
      RECT 60.515 0.915 60.685 1.085 ;
      RECT 60.515 1.655 60.685 1.825 ;
      RECT 60.515 7.055 60.685 7.225 ;
      RECT 60.515 7.795 60.685 7.965 ;
      RECT 60.14 2.395 60.31 2.565 ;
      RECT 60.14 6.315 60.31 6.485 ;
      RECT 57.08 2.77 57.25 2.94 ;
      RECT 56.84 1.93 57.01 2.1 ;
      RECT 56.84 3.61 57.01 3.78 ;
      RECT 56.6 2.49 56.77 2.66 ;
      RECT 56.6 3.05 56.77 3.22 ;
      RECT 56.12 2.77 56.29 2.94 ;
      RECT 55.88 1.93 56.05 2.1 ;
      RECT 55.64 2.49 55.81 2.66 ;
      RECT 55.43 3.33 55.6 3.5 ;
      RECT 55.33 6.685 55.5 6.855 ;
      RECT 55.16 2.77 55.33 2.94 ;
      RECT 54.9 7.055 55.07 7.225 ;
      RECT 54.9 7.795 55.07 7.965 ;
      RECT 54.89 3.61 55.06 3.78 ;
      RECT 54.68 2.19 54.85 2.36 ;
      RECT 54.2 2.77 54.37 2.94 ;
      RECT 53.96 1.93 54.13 2.1 ;
      RECT 53.72 2.49 53.89 2.66 ;
      RECT 53.72 3.05 53.89 3.22 ;
      RECT 53.24 2.49 53.41 2.66 ;
      RECT 53 3.61 53.17 3.78 ;
      RECT 52.96 1.93 53.13 2.1 ;
      RECT 52.76 2.77 52.93 2.94 ;
      RECT 52.52 3.61 52.69 3.78 ;
      RECT 52.28 3.05 52.45 3.22 ;
      RECT 51.8 2.49 51.97 2.66 ;
      RECT 51.56 1.93 51.73 2.1 ;
      RECT 51.56 3.61 51.73 3.78 ;
      RECT 51.08 3.05 51.25 3.22 ;
      RECT 50.84 2.49 51.01 2.66 ;
      RECT 50.6 3.33 50.77 3.5 ;
      RECT 50.36 2.77 50.53 2.94 ;
      RECT 49.67 1.93 49.84 2.1 ;
      RECT 49.67 3.33 49.84 3.5 ;
      RECT 48.035 7.8 48.205 7.97 ;
      RECT 47.665 2.76 47.835 2.93 ;
      RECT 47.665 5.95 47.835 6.12 ;
      RECT 47.045 0.91 47.215 1.08 ;
      RECT 47.045 2.39 47.215 2.56 ;
      RECT 47.045 6.32 47.215 6.49 ;
      RECT 47.045 7.8 47.215 7.97 ;
      RECT 46.675 2.76 46.845 2.93 ;
      RECT 46.675 5.95 46.845 6.12 ;
      RECT 45.685 2.025 45.855 2.195 ;
      RECT 45.685 6.685 45.855 6.855 ;
      RECT 45.255 0.915 45.425 1.085 ;
      RECT 45.255 1.655 45.425 1.825 ;
      RECT 45.255 7.055 45.425 7.225 ;
      RECT 45.255 7.795 45.425 7.965 ;
      RECT 44.88 2.395 45.05 2.565 ;
      RECT 44.88 6.315 45.05 6.485 ;
      RECT 41.82 2.77 41.99 2.94 ;
      RECT 41.58 1.93 41.75 2.1 ;
      RECT 41.58 3.61 41.75 3.78 ;
      RECT 41.34 2.49 41.51 2.66 ;
      RECT 41.34 3.05 41.51 3.22 ;
      RECT 40.86 2.77 41.03 2.94 ;
      RECT 40.62 1.93 40.79 2.1 ;
      RECT 40.38 2.49 40.55 2.66 ;
      RECT 40.17 3.33 40.34 3.5 ;
      RECT 40.07 6.685 40.24 6.855 ;
      RECT 39.9 2.77 40.07 2.94 ;
      RECT 39.64 7.055 39.81 7.225 ;
      RECT 39.64 7.795 39.81 7.965 ;
      RECT 39.63 3.61 39.8 3.78 ;
      RECT 39.42 2.19 39.59 2.36 ;
      RECT 38.94 2.77 39.11 2.94 ;
      RECT 38.7 1.93 38.87 2.1 ;
      RECT 38.46 2.49 38.63 2.66 ;
      RECT 38.46 3.05 38.63 3.22 ;
      RECT 37.98 2.49 38.15 2.66 ;
      RECT 37.74 3.61 37.91 3.78 ;
      RECT 37.7 1.93 37.87 2.1 ;
      RECT 37.5 2.77 37.67 2.94 ;
      RECT 37.26 3.61 37.43 3.78 ;
      RECT 37.02 3.05 37.19 3.22 ;
      RECT 36.54 2.49 36.71 2.66 ;
      RECT 36.3 1.93 36.47 2.1 ;
      RECT 36.3 3.61 36.47 3.78 ;
      RECT 35.82 3.05 35.99 3.22 ;
      RECT 35.58 2.49 35.75 2.66 ;
      RECT 35.34 3.33 35.51 3.5 ;
      RECT 35.1 2.77 35.27 2.94 ;
      RECT 34.41 1.93 34.58 2.1 ;
      RECT 34.41 3.33 34.58 3.5 ;
      RECT 32.775 7.8 32.945 7.97 ;
      RECT 32.405 2.76 32.575 2.93 ;
      RECT 32.405 5.95 32.575 6.12 ;
      RECT 31.785 0.91 31.955 1.08 ;
      RECT 31.785 2.39 31.955 2.56 ;
      RECT 31.785 6.32 31.955 6.49 ;
      RECT 31.785 7.8 31.955 7.97 ;
      RECT 31.415 2.76 31.585 2.93 ;
      RECT 31.415 5.95 31.585 6.12 ;
      RECT 30.425 2.025 30.595 2.195 ;
      RECT 30.425 6.685 30.595 6.855 ;
      RECT 29.995 0.915 30.165 1.085 ;
      RECT 29.995 1.655 30.165 1.825 ;
      RECT 29.995 7.055 30.165 7.225 ;
      RECT 29.995 7.795 30.165 7.965 ;
      RECT 29.62 2.395 29.79 2.565 ;
      RECT 29.62 6.315 29.79 6.485 ;
      RECT 26.56 2.77 26.73 2.94 ;
      RECT 26.32 1.93 26.49 2.1 ;
      RECT 26.32 3.61 26.49 3.78 ;
      RECT 26.08 2.49 26.25 2.66 ;
      RECT 26.08 3.05 26.25 3.22 ;
      RECT 25.6 2.77 25.77 2.94 ;
      RECT 25.36 1.93 25.53 2.1 ;
      RECT 25.12 2.49 25.29 2.66 ;
      RECT 24.91 3.33 25.08 3.5 ;
      RECT 24.81 6.685 24.98 6.855 ;
      RECT 24.64 2.77 24.81 2.94 ;
      RECT 24.38 7.055 24.55 7.225 ;
      RECT 24.38 7.795 24.55 7.965 ;
      RECT 24.37 3.61 24.54 3.78 ;
      RECT 24.16 2.19 24.33 2.36 ;
      RECT 23.68 2.77 23.85 2.94 ;
      RECT 23.44 1.93 23.61 2.1 ;
      RECT 23.2 2.49 23.37 2.66 ;
      RECT 23.2 3.05 23.37 3.22 ;
      RECT 22.72 2.49 22.89 2.66 ;
      RECT 22.48 3.61 22.65 3.78 ;
      RECT 22.44 1.93 22.61 2.1 ;
      RECT 22.24 2.77 22.41 2.94 ;
      RECT 22 3.61 22.17 3.78 ;
      RECT 21.76 3.05 21.93 3.22 ;
      RECT 21.28 2.49 21.45 2.66 ;
      RECT 21.04 1.93 21.21 2.1 ;
      RECT 21.04 3.61 21.21 3.78 ;
      RECT 20.56 3.05 20.73 3.22 ;
      RECT 20.32 2.49 20.49 2.66 ;
      RECT 20.08 3.33 20.25 3.5 ;
      RECT 19.84 2.77 20.01 2.94 ;
      RECT 19.15 1.93 19.32 2.1 ;
      RECT 19.15 3.33 19.32 3.5 ;
      RECT 17.515 7.8 17.685 7.97 ;
      RECT 17.145 2.76 17.315 2.93 ;
      RECT 17.145 5.95 17.315 6.12 ;
      RECT 16.525 0.91 16.695 1.08 ;
      RECT 16.525 2.39 16.695 2.56 ;
      RECT 16.525 6.32 16.695 6.49 ;
      RECT 16.525 7.8 16.695 7.97 ;
      RECT 16.155 2.76 16.325 2.93 ;
      RECT 16.155 5.95 16.325 6.12 ;
      RECT 15.165 2.025 15.335 2.195 ;
      RECT 15.165 6.685 15.335 6.855 ;
      RECT 14.735 0.915 14.905 1.085 ;
      RECT 14.735 1.655 14.905 1.825 ;
      RECT 14.735 7.055 14.905 7.225 ;
      RECT 14.735 7.795 14.905 7.965 ;
      RECT 14.36 2.395 14.53 2.565 ;
      RECT 14.36 6.315 14.53 6.485 ;
      RECT 11.3 2.77 11.47 2.94 ;
      RECT 11.06 1.93 11.23 2.1 ;
      RECT 11.06 3.61 11.23 3.78 ;
      RECT 10.82 2.49 10.99 2.66 ;
      RECT 10.82 3.05 10.99 3.22 ;
      RECT 10.34 2.77 10.51 2.94 ;
      RECT 10.1 1.93 10.27 2.1 ;
      RECT 9.86 2.49 10.03 2.66 ;
      RECT 9.65 3.33 9.82 3.5 ;
      RECT 9.55 6.685 9.72 6.855 ;
      RECT 9.38 2.77 9.55 2.94 ;
      RECT 9.12 7.055 9.29 7.225 ;
      RECT 9.12 7.795 9.29 7.965 ;
      RECT 9.11 3.61 9.28 3.78 ;
      RECT 8.9 2.19 9.07 2.36 ;
      RECT 8.42 2.77 8.59 2.94 ;
      RECT 8.18 1.93 8.35 2.1 ;
      RECT 7.94 2.49 8.11 2.66 ;
      RECT 7.94 3.05 8.11 3.22 ;
      RECT 7.46 2.49 7.63 2.66 ;
      RECT 7.22 3.61 7.39 3.78 ;
      RECT 7.18 1.93 7.35 2.1 ;
      RECT 6.98 2.77 7.15 2.94 ;
      RECT 6.74 3.61 6.91 3.78 ;
      RECT 6.5 3.05 6.67 3.22 ;
      RECT 6.02 2.49 6.19 2.66 ;
      RECT 5.78 1.93 5.95 2.1 ;
      RECT 5.78 3.61 5.95 3.78 ;
      RECT 5.3 3.05 5.47 3.22 ;
      RECT 5.06 2.49 5.23 2.66 ;
      RECT 4.82 3.33 4.99 3.5 ;
      RECT 4.58 2.77 4.75 2.94 ;
      RECT 3.89 1.93 4.06 2.1 ;
      RECT 3.89 3.33 4.06 3.5 ;
      RECT 1.605 7.055 1.775 7.225 ;
      RECT 1.605 7.795 1.775 7.965 ;
      RECT 1.23 6.315 1.4 6.485 ;
    LAYER li1 ;
      RECT 78.555 5.02 78.725 6.49 ;
      RECT 78.555 6.315 78.73 6.485 ;
      RECT 78.185 1.74 78.355 2.93 ;
      RECT 78.185 1.74 78.655 1.91 ;
      RECT 78.185 6.97 78.655 7.14 ;
      RECT 78.185 5.95 78.355 7.14 ;
      RECT 77.195 1.74 77.365 2.93 ;
      RECT 77.195 1.74 77.665 1.91 ;
      RECT 77.195 6.97 77.665 7.14 ;
      RECT 77.195 5.95 77.365 7.14 ;
      RECT 75.345 2.635 75.515 3.865 ;
      RECT 75.4 0.855 75.57 2.805 ;
      RECT 75.345 0.575 75.515 1.025 ;
      RECT 75.345 7.855 75.515 8.305 ;
      RECT 75.4 6.075 75.57 8.025 ;
      RECT 75.345 5.015 75.515 6.245 ;
      RECT 74.825 0.575 74.995 3.865 ;
      RECT 74.825 2.075 75.23 2.405 ;
      RECT 74.825 1.235 75.23 1.565 ;
      RECT 74.825 5.015 74.995 8.305 ;
      RECT 74.825 7.315 75.23 7.645 ;
      RECT 74.825 6.475 75.23 6.805 ;
      RECT 72.1 3.61 72.61 3.78 ;
      RECT 72.44 3.22 72.61 3.78 ;
      RECT 72.55 3.14 72.72 3.47 ;
      RECT 72.34 2.53 72.61 2.94 ;
      RECT 72.22 2.53 72.61 2.74 ;
      RECT 70.69 3.14 70.86 3.5 ;
      RECT 70.69 3.22 72.03 3.39 ;
      RECT 71.86 3.05 72.03 3.39 ;
      RECT 70.42 2.57 70.59 2.94 ;
      RECT 69.94 2.57 70.59 2.84 ;
      RECT 69.86 2.57 70.67 2.74 ;
      RECT 69.22 1.81 69.39 2.1 ;
      RECT 69.22 1.81 70.46 1.98 ;
      RECT 69.94 2.15 70.11 2.36 ;
      RECT 69.58 2.15 70.11 2.32 ;
      RECT 69.21 5.015 69.38 8.305 ;
      RECT 69.21 7.315 69.615 7.645 ;
      RECT 69.21 6.475 69.615 6.805 ;
      RECT 68.98 3.22 69.47 3.39 ;
      RECT 68.98 3.05 69.15 3.39 ;
      RECT 68.26 3.22 68.43 3.78 ;
      RECT 68.15 3.22 68.48 3.39 ;
      RECT 68.22 1.83 68.39 2.1 ;
      RECT 68.26 1.75 68.43 2.08 ;
      RECT 68.12 1.83 68.43 2.05 ;
      RECT 66.7 3.22 66.99 3.78 ;
      RECT 66.82 3.14 66.99 3.78 ;
      RECT 63.295 5.02 63.465 6.49 ;
      RECT 63.295 6.315 63.47 6.485 ;
      RECT 62.925 1.74 63.095 2.93 ;
      RECT 62.925 1.74 63.395 1.91 ;
      RECT 62.925 6.97 63.395 7.14 ;
      RECT 62.925 5.95 63.095 7.14 ;
      RECT 61.935 1.74 62.105 2.93 ;
      RECT 61.935 1.74 62.405 1.91 ;
      RECT 61.935 6.97 62.405 7.14 ;
      RECT 61.935 5.95 62.105 7.14 ;
      RECT 60.085 2.635 60.255 3.865 ;
      RECT 60.14 0.855 60.31 2.805 ;
      RECT 60.085 0.575 60.255 1.025 ;
      RECT 60.085 7.855 60.255 8.305 ;
      RECT 60.14 6.075 60.31 8.025 ;
      RECT 60.085 5.015 60.255 6.245 ;
      RECT 59.565 0.575 59.735 3.865 ;
      RECT 59.565 2.075 59.97 2.405 ;
      RECT 59.565 1.235 59.97 1.565 ;
      RECT 59.565 5.015 59.735 8.305 ;
      RECT 59.565 7.315 59.97 7.645 ;
      RECT 59.565 6.475 59.97 6.805 ;
      RECT 56.84 3.61 57.35 3.78 ;
      RECT 57.18 3.22 57.35 3.78 ;
      RECT 57.29 3.14 57.46 3.47 ;
      RECT 57.08 2.53 57.35 2.94 ;
      RECT 56.96 2.53 57.35 2.74 ;
      RECT 55.43 3.14 55.6 3.5 ;
      RECT 55.43 3.22 56.77 3.39 ;
      RECT 56.6 3.05 56.77 3.39 ;
      RECT 55.16 2.57 55.33 2.94 ;
      RECT 54.68 2.57 55.33 2.84 ;
      RECT 54.6 2.57 55.41 2.74 ;
      RECT 53.96 1.81 54.13 2.1 ;
      RECT 53.96 1.81 55.2 1.98 ;
      RECT 54.68 2.15 54.85 2.36 ;
      RECT 54.32 2.15 54.85 2.32 ;
      RECT 53.95 5.015 54.12 8.305 ;
      RECT 53.95 7.315 54.355 7.645 ;
      RECT 53.95 6.475 54.355 6.805 ;
      RECT 53.72 3.22 54.21 3.39 ;
      RECT 53.72 3.05 53.89 3.39 ;
      RECT 53 3.22 53.17 3.78 ;
      RECT 52.89 3.22 53.22 3.39 ;
      RECT 52.96 1.83 53.13 2.1 ;
      RECT 53 1.75 53.17 2.08 ;
      RECT 52.86 1.83 53.17 2.05 ;
      RECT 51.44 3.22 51.73 3.78 ;
      RECT 51.56 3.14 51.73 3.78 ;
      RECT 48.035 5.02 48.205 6.49 ;
      RECT 48.035 6.315 48.21 6.485 ;
      RECT 47.665 1.74 47.835 2.93 ;
      RECT 47.665 1.74 48.135 1.91 ;
      RECT 47.665 6.97 48.135 7.14 ;
      RECT 47.665 5.95 47.835 7.14 ;
      RECT 46.675 1.74 46.845 2.93 ;
      RECT 46.675 1.74 47.145 1.91 ;
      RECT 46.675 6.97 47.145 7.14 ;
      RECT 46.675 5.95 46.845 7.14 ;
      RECT 44.825 2.635 44.995 3.865 ;
      RECT 44.88 0.855 45.05 2.805 ;
      RECT 44.825 0.575 44.995 1.025 ;
      RECT 44.825 7.855 44.995 8.305 ;
      RECT 44.88 6.075 45.05 8.025 ;
      RECT 44.825 5.015 44.995 6.245 ;
      RECT 44.305 0.575 44.475 3.865 ;
      RECT 44.305 2.075 44.71 2.405 ;
      RECT 44.305 1.235 44.71 1.565 ;
      RECT 44.305 5.015 44.475 8.305 ;
      RECT 44.305 7.315 44.71 7.645 ;
      RECT 44.305 6.475 44.71 6.805 ;
      RECT 41.58 3.61 42.09 3.78 ;
      RECT 41.92 3.22 42.09 3.78 ;
      RECT 42.03 3.14 42.2 3.47 ;
      RECT 41.82 2.53 42.09 2.94 ;
      RECT 41.7 2.53 42.09 2.74 ;
      RECT 40.17 3.14 40.34 3.5 ;
      RECT 40.17 3.22 41.51 3.39 ;
      RECT 41.34 3.05 41.51 3.39 ;
      RECT 39.9 2.57 40.07 2.94 ;
      RECT 39.42 2.57 40.07 2.84 ;
      RECT 39.34 2.57 40.15 2.74 ;
      RECT 38.7 1.81 38.87 2.1 ;
      RECT 38.7 1.81 39.94 1.98 ;
      RECT 39.42 2.15 39.59 2.36 ;
      RECT 39.06 2.15 39.59 2.32 ;
      RECT 38.69 5.015 38.86 8.305 ;
      RECT 38.69 7.315 39.095 7.645 ;
      RECT 38.69 6.475 39.095 6.805 ;
      RECT 38.46 3.22 38.95 3.39 ;
      RECT 38.46 3.05 38.63 3.39 ;
      RECT 37.74 3.22 37.91 3.78 ;
      RECT 37.63 3.22 37.96 3.39 ;
      RECT 37.7 1.83 37.87 2.1 ;
      RECT 37.74 1.75 37.91 2.08 ;
      RECT 37.6 1.83 37.91 2.05 ;
      RECT 36.18 3.22 36.47 3.78 ;
      RECT 36.3 3.14 36.47 3.78 ;
      RECT 32.775 5.02 32.945 6.49 ;
      RECT 32.775 6.315 32.95 6.485 ;
      RECT 32.405 1.74 32.575 2.93 ;
      RECT 32.405 1.74 32.875 1.91 ;
      RECT 32.405 6.97 32.875 7.14 ;
      RECT 32.405 5.95 32.575 7.14 ;
      RECT 31.415 1.74 31.585 2.93 ;
      RECT 31.415 1.74 31.885 1.91 ;
      RECT 31.415 6.97 31.885 7.14 ;
      RECT 31.415 5.95 31.585 7.14 ;
      RECT 29.565 2.635 29.735 3.865 ;
      RECT 29.62 0.855 29.79 2.805 ;
      RECT 29.565 0.575 29.735 1.025 ;
      RECT 29.565 7.855 29.735 8.305 ;
      RECT 29.62 6.075 29.79 8.025 ;
      RECT 29.565 5.015 29.735 6.245 ;
      RECT 29.045 0.575 29.215 3.865 ;
      RECT 29.045 2.075 29.45 2.405 ;
      RECT 29.045 1.235 29.45 1.565 ;
      RECT 29.045 5.015 29.215 8.305 ;
      RECT 29.045 7.315 29.45 7.645 ;
      RECT 29.045 6.475 29.45 6.805 ;
      RECT 26.32 3.61 26.83 3.78 ;
      RECT 26.66 3.22 26.83 3.78 ;
      RECT 26.77 3.14 26.94 3.47 ;
      RECT 26.56 2.53 26.83 2.94 ;
      RECT 26.44 2.53 26.83 2.74 ;
      RECT 24.91 3.14 25.08 3.5 ;
      RECT 24.91 3.22 26.25 3.39 ;
      RECT 26.08 3.05 26.25 3.39 ;
      RECT 24.64 2.57 24.81 2.94 ;
      RECT 24.16 2.57 24.81 2.84 ;
      RECT 24.08 2.57 24.89 2.74 ;
      RECT 23.44 1.81 23.61 2.1 ;
      RECT 23.44 1.81 24.68 1.98 ;
      RECT 24.16 2.15 24.33 2.36 ;
      RECT 23.8 2.15 24.33 2.32 ;
      RECT 23.43 5.015 23.6 8.305 ;
      RECT 23.43 7.315 23.835 7.645 ;
      RECT 23.43 6.475 23.835 6.805 ;
      RECT 23.2 3.22 23.69 3.39 ;
      RECT 23.2 3.05 23.37 3.39 ;
      RECT 22.48 3.22 22.65 3.78 ;
      RECT 22.37 3.22 22.7 3.39 ;
      RECT 22.44 1.83 22.61 2.1 ;
      RECT 22.48 1.75 22.65 2.08 ;
      RECT 22.34 1.83 22.65 2.05 ;
      RECT 20.92 3.22 21.21 3.78 ;
      RECT 21.04 3.14 21.21 3.78 ;
      RECT 17.515 5.02 17.685 6.49 ;
      RECT 17.515 6.315 17.69 6.485 ;
      RECT 17.145 1.74 17.315 2.93 ;
      RECT 17.145 1.74 17.615 1.91 ;
      RECT 17.145 6.97 17.615 7.14 ;
      RECT 17.145 5.95 17.315 7.14 ;
      RECT 16.155 1.74 16.325 2.93 ;
      RECT 16.155 1.74 16.625 1.91 ;
      RECT 16.155 6.97 16.625 7.14 ;
      RECT 16.155 5.95 16.325 7.14 ;
      RECT 14.305 2.635 14.475 3.865 ;
      RECT 14.36 0.855 14.53 2.805 ;
      RECT 14.305 0.575 14.475 1.025 ;
      RECT 14.305 7.855 14.475 8.305 ;
      RECT 14.36 6.075 14.53 8.025 ;
      RECT 14.305 5.015 14.475 6.245 ;
      RECT 13.785 0.575 13.955 3.865 ;
      RECT 13.785 2.075 14.19 2.405 ;
      RECT 13.785 1.235 14.19 1.565 ;
      RECT 13.785 5.015 13.955 8.305 ;
      RECT 13.785 7.315 14.19 7.645 ;
      RECT 13.785 6.475 14.19 6.805 ;
      RECT 11.06 3.61 11.57 3.78 ;
      RECT 11.4 3.22 11.57 3.78 ;
      RECT 11.51 3.14 11.68 3.47 ;
      RECT 11.3 2.53 11.57 2.94 ;
      RECT 11.18 2.53 11.57 2.74 ;
      RECT 9.65 3.14 9.82 3.5 ;
      RECT 9.65 3.22 10.99 3.39 ;
      RECT 10.82 3.05 10.99 3.39 ;
      RECT 9.38 2.57 9.55 2.94 ;
      RECT 8.9 2.57 9.55 2.84 ;
      RECT 8.82 2.57 9.63 2.74 ;
      RECT 8.18 1.81 8.35 2.1 ;
      RECT 8.18 1.81 9.42 1.98 ;
      RECT 8.9 2.15 9.07 2.36 ;
      RECT 8.54 2.15 9.07 2.32 ;
      RECT 8.17 5.015 8.34 8.305 ;
      RECT 8.17 7.315 8.575 7.645 ;
      RECT 8.17 6.475 8.575 6.805 ;
      RECT 7.94 3.22 8.43 3.39 ;
      RECT 7.94 3.05 8.11 3.39 ;
      RECT 7.22 3.22 7.39 3.78 ;
      RECT 7.11 3.22 7.44 3.39 ;
      RECT 7.18 1.83 7.35 2.1 ;
      RECT 7.22 1.75 7.39 2.08 ;
      RECT 7.08 1.83 7.39 2.05 ;
      RECT 5.66 3.22 5.95 3.78 ;
      RECT 5.78 3.14 5.95 3.78 ;
      RECT 1.175 7.855 1.345 8.305 ;
      RECT 1.23 6.075 1.4 8.025 ;
      RECT 1.175 5.015 1.345 6.245 ;
      RECT 0.655 5.015 0.825 8.305 ;
      RECT 0.655 7.315 1.06 7.645 ;
      RECT 0.655 6.475 1.06 6.805 ;
      RECT 78.555 7.8 78.725 8.31 ;
      RECT 77.565 0.57 77.735 1.08 ;
      RECT 77.565 2.39 77.735 3.86 ;
      RECT 77.565 5.02 77.735 6.49 ;
      RECT 77.565 7.8 77.735 8.31 ;
      RECT 76.205 0.575 76.375 3.865 ;
      RECT 76.205 5.015 76.375 8.305 ;
      RECT 75.775 0.575 75.945 1.085 ;
      RECT 75.775 1.655 75.945 3.865 ;
      RECT 75.775 5.015 75.945 7.225 ;
      RECT 75.775 7.795 75.945 8.305 ;
      RECT 72.1 1.75 72.27 2.1 ;
      RECT 71.86 2.49 72.03 2.82 ;
      RECT 71.38 2.49 71.55 2.94 ;
      RECT 71.14 1.75 71.31 2.1 ;
      RECT 70.9 2.49 71.07 2.82 ;
      RECT 70.59 5.015 70.76 8.305 ;
      RECT 70.16 5.015 70.33 7.225 ;
      RECT 70.16 7.795 70.33 8.305 ;
      RECT 70.15 3.48 70.32 3.81 ;
      RECT 69.46 2.49 69.63 2.94 ;
      RECT 68.98 2.49 69.15 2.82 ;
      RECT 68.5 2.49 68.67 2.82 ;
      RECT 68.02 2.49 68.19 2.94 ;
      RECT 67.78 3.48 67.95 3.81 ;
      RECT 67.54 2.49 67.71 3.22 ;
      RECT 67.06 2.49 67.23 2.82 ;
      RECT 66.82 1.75 66.99 2.1 ;
      RECT 66.34 3.05 66.51 3.47 ;
      RECT 66.1 2.49 66.27 2.82 ;
      RECT 65.86 3.14 66.03 3.5 ;
      RECT 65.62 2.49 65.79 2.94 ;
      RECT 64.93 1.75 65.1 2.1 ;
      RECT 64.93 3.14 65.1 3.5 ;
      RECT 63.295 7.8 63.465 8.31 ;
      RECT 62.305 0.57 62.475 1.08 ;
      RECT 62.305 2.39 62.475 3.86 ;
      RECT 62.305 5.02 62.475 6.49 ;
      RECT 62.305 7.8 62.475 8.31 ;
      RECT 60.945 0.575 61.115 3.865 ;
      RECT 60.945 5.015 61.115 8.305 ;
      RECT 60.515 0.575 60.685 1.085 ;
      RECT 60.515 1.655 60.685 3.865 ;
      RECT 60.515 5.015 60.685 7.225 ;
      RECT 60.515 7.795 60.685 8.305 ;
      RECT 56.84 1.75 57.01 2.1 ;
      RECT 56.6 2.49 56.77 2.82 ;
      RECT 56.12 2.49 56.29 2.94 ;
      RECT 55.88 1.75 56.05 2.1 ;
      RECT 55.64 2.49 55.81 2.82 ;
      RECT 55.33 5.015 55.5 8.305 ;
      RECT 54.9 5.015 55.07 7.225 ;
      RECT 54.9 7.795 55.07 8.305 ;
      RECT 54.89 3.48 55.06 3.81 ;
      RECT 54.2 2.49 54.37 2.94 ;
      RECT 53.72 2.49 53.89 2.82 ;
      RECT 53.24 2.49 53.41 2.82 ;
      RECT 52.76 2.49 52.93 2.94 ;
      RECT 52.52 3.48 52.69 3.81 ;
      RECT 52.28 2.49 52.45 3.22 ;
      RECT 51.8 2.49 51.97 2.82 ;
      RECT 51.56 1.75 51.73 2.1 ;
      RECT 51.08 3.05 51.25 3.47 ;
      RECT 50.84 2.49 51.01 2.82 ;
      RECT 50.6 3.14 50.77 3.5 ;
      RECT 50.36 2.49 50.53 2.94 ;
      RECT 49.67 1.75 49.84 2.1 ;
      RECT 49.67 3.14 49.84 3.5 ;
      RECT 48.035 7.8 48.205 8.31 ;
      RECT 47.045 0.57 47.215 1.08 ;
      RECT 47.045 2.39 47.215 3.86 ;
      RECT 47.045 5.02 47.215 6.49 ;
      RECT 47.045 7.8 47.215 8.31 ;
      RECT 45.685 0.575 45.855 3.865 ;
      RECT 45.685 5.015 45.855 8.305 ;
      RECT 45.255 0.575 45.425 1.085 ;
      RECT 45.255 1.655 45.425 3.865 ;
      RECT 45.255 5.015 45.425 7.225 ;
      RECT 45.255 7.795 45.425 8.305 ;
      RECT 41.58 1.75 41.75 2.1 ;
      RECT 41.34 2.49 41.51 2.82 ;
      RECT 40.86 2.49 41.03 2.94 ;
      RECT 40.62 1.75 40.79 2.1 ;
      RECT 40.38 2.49 40.55 2.82 ;
      RECT 40.07 5.015 40.24 8.305 ;
      RECT 39.64 5.015 39.81 7.225 ;
      RECT 39.64 7.795 39.81 8.305 ;
      RECT 39.63 3.48 39.8 3.81 ;
      RECT 38.94 2.49 39.11 2.94 ;
      RECT 38.46 2.49 38.63 2.82 ;
      RECT 37.98 2.49 38.15 2.82 ;
      RECT 37.5 2.49 37.67 2.94 ;
      RECT 37.26 3.48 37.43 3.81 ;
      RECT 37.02 2.49 37.19 3.22 ;
      RECT 36.54 2.49 36.71 2.82 ;
      RECT 36.3 1.75 36.47 2.1 ;
      RECT 35.82 3.05 35.99 3.47 ;
      RECT 35.58 2.49 35.75 2.82 ;
      RECT 35.34 3.14 35.51 3.5 ;
      RECT 35.1 2.49 35.27 2.94 ;
      RECT 34.41 1.75 34.58 2.1 ;
      RECT 34.41 3.14 34.58 3.5 ;
      RECT 32.775 7.8 32.945 8.31 ;
      RECT 31.785 0.57 31.955 1.08 ;
      RECT 31.785 2.39 31.955 3.86 ;
      RECT 31.785 5.02 31.955 6.49 ;
      RECT 31.785 7.8 31.955 8.31 ;
      RECT 30.425 0.575 30.595 3.865 ;
      RECT 30.425 5.015 30.595 8.305 ;
      RECT 29.995 0.575 30.165 1.085 ;
      RECT 29.995 1.655 30.165 3.865 ;
      RECT 29.995 5.015 30.165 7.225 ;
      RECT 29.995 7.795 30.165 8.305 ;
      RECT 26.32 1.75 26.49 2.1 ;
      RECT 26.08 2.49 26.25 2.82 ;
      RECT 25.6 2.49 25.77 2.94 ;
      RECT 25.36 1.75 25.53 2.1 ;
      RECT 25.12 2.49 25.29 2.82 ;
      RECT 24.81 5.015 24.98 8.305 ;
      RECT 24.38 5.015 24.55 7.225 ;
      RECT 24.38 7.795 24.55 8.305 ;
      RECT 24.37 3.48 24.54 3.81 ;
      RECT 23.68 2.49 23.85 2.94 ;
      RECT 23.2 2.49 23.37 2.82 ;
      RECT 22.72 2.49 22.89 2.82 ;
      RECT 22.24 2.49 22.41 2.94 ;
      RECT 22 3.48 22.17 3.81 ;
      RECT 21.76 2.49 21.93 3.22 ;
      RECT 21.28 2.49 21.45 2.82 ;
      RECT 21.04 1.75 21.21 2.1 ;
      RECT 20.56 3.05 20.73 3.47 ;
      RECT 20.32 2.49 20.49 2.82 ;
      RECT 20.08 3.14 20.25 3.5 ;
      RECT 19.84 2.49 20.01 2.94 ;
      RECT 19.15 1.75 19.32 2.1 ;
      RECT 19.15 3.14 19.32 3.5 ;
      RECT 17.515 7.8 17.685 8.31 ;
      RECT 16.525 0.57 16.695 1.08 ;
      RECT 16.525 2.39 16.695 3.86 ;
      RECT 16.525 5.02 16.695 6.49 ;
      RECT 16.525 7.8 16.695 8.31 ;
      RECT 15.165 0.575 15.335 3.865 ;
      RECT 15.165 5.015 15.335 8.305 ;
      RECT 14.735 0.575 14.905 1.085 ;
      RECT 14.735 1.655 14.905 3.865 ;
      RECT 14.735 5.015 14.905 7.225 ;
      RECT 14.735 7.795 14.905 8.305 ;
      RECT 11.06 1.75 11.23 2.1 ;
      RECT 10.82 2.49 10.99 2.82 ;
      RECT 10.34 2.49 10.51 2.94 ;
      RECT 10.1 1.75 10.27 2.1 ;
      RECT 9.86 2.49 10.03 2.82 ;
      RECT 9.55 5.015 9.72 8.305 ;
      RECT 9.12 5.015 9.29 7.225 ;
      RECT 9.12 7.795 9.29 8.305 ;
      RECT 9.11 3.48 9.28 3.81 ;
      RECT 8.42 2.49 8.59 2.94 ;
      RECT 7.94 2.49 8.11 2.82 ;
      RECT 7.46 2.49 7.63 2.82 ;
      RECT 6.98 2.49 7.15 2.94 ;
      RECT 6.74 3.48 6.91 3.81 ;
      RECT 6.5 2.49 6.67 3.22 ;
      RECT 6.02 2.49 6.19 2.82 ;
      RECT 5.78 1.75 5.95 2.1 ;
      RECT 5.3 3.05 5.47 3.47 ;
      RECT 5.06 2.49 5.23 2.82 ;
      RECT 4.82 3.14 4.99 3.5 ;
      RECT 4.58 2.49 4.75 2.94 ;
      RECT 3.89 1.75 4.06 2.1 ;
      RECT 3.89 3.14 4.06 3.5 ;
      RECT 1.605 5.015 1.775 7.225 ;
      RECT 1.605 7.795 1.775 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r2 ;
  SIZE 79.095 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 17.515 0.915 17.685 1.085 ;
        RECT 17.51 0.91 17.68 1.08 ;
        RECT 17.51 2.39 17.68 2.56 ;
      LAYER li1 ;
        RECT 17.515 0.915 17.685 1.085 ;
        RECT 17.51 0.57 17.68 1.08 ;
        RECT 17.51 2.39 17.68 3.86 ;
      LAYER met1 ;
        RECT 17.45 2.36 17.74 2.59 ;
        RECT 17.45 0.88 17.74 1.11 ;
        RECT 17.51 0.88 17.68 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 32.775 0.915 32.945 1.085 ;
        RECT 32.77 0.91 32.94 1.08 ;
        RECT 32.77 2.39 32.94 2.56 ;
      LAYER li1 ;
        RECT 32.775 0.915 32.945 1.085 ;
        RECT 32.77 0.57 32.94 1.08 ;
        RECT 32.77 2.39 32.94 3.86 ;
      LAYER met1 ;
        RECT 32.71 2.36 33 2.59 ;
        RECT 32.71 0.88 33 1.11 ;
        RECT 32.77 0.88 32.94 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 48.035 0.915 48.205 1.085 ;
        RECT 48.03 0.91 48.2 1.08 ;
        RECT 48.03 2.39 48.2 2.56 ;
      LAYER li1 ;
        RECT 48.035 0.915 48.205 1.085 ;
        RECT 48.03 0.57 48.2 1.08 ;
        RECT 48.03 2.39 48.2 3.86 ;
      LAYER met1 ;
        RECT 47.97 2.36 48.26 2.59 ;
        RECT 47.97 0.88 48.26 1.11 ;
        RECT 48.03 0.88 48.2 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 63.295 0.915 63.465 1.085 ;
        RECT 63.29 0.91 63.46 1.08 ;
        RECT 63.29 2.39 63.46 2.56 ;
      LAYER li1 ;
        RECT 63.295 0.915 63.465 1.085 ;
        RECT 63.29 0.57 63.46 1.08 ;
        RECT 63.29 2.39 63.46 3.86 ;
      LAYER met1 ;
        RECT 63.23 2.36 63.52 2.59 ;
        RECT 63.23 0.88 63.52 1.11 ;
        RECT 63.29 0.88 63.46 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 78.555 0.915 78.725 1.085 ;
        RECT 78.55 0.91 78.72 1.08 ;
        RECT 78.55 2.39 78.72 2.56 ;
      LAYER li1 ;
        RECT 78.555 0.915 78.725 1.085 ;
        RECT 78.55 0.57 78.72 1.08 ;
        RECT 78.55 2.39 78.72 3.86 ;
      LAYER met1 ;
        RECT 78.49 2.36 78.78 2.59 ;
        RECT 78.49 0.88 78.78 1.11 ;
        RECT 78.55 0.88 78.72 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 13.28 5.86 13.62 6.21 ;
        RECT 13.28 2.705 13.62 3.055 ;
        RECT 13.36 2.705 13.53 6.21 ;
      LAYER li1 ;
        RECT 13.36 1.66 13.53 2.935 ;
        RECT 13.36 5.945 13.53 7.22 ;
        RECT 7.745 5.945 7.915 7.22 ;
      LAYER met1 ;
        RECT 13.28 2.765 13.76 2.935 ;
        RECT 13.28 2.705 13.62 3.055 ;
        RECT 7.685 5.945 13.76 6.115 ;
        RECT 13.28 5.86 13.62 6.21 ;
        RECT 7.685 5.915 7.975 6.145 ;
      LAYER mcon ;
        RECT 7.745 5.945 7.915 6.115 ;
        RECT 13.36 5.945 13.53 6.115 ;
        RECT 13.36 2.765 13.53 2.935 ;
      LAYER via1 ;
        RECT 13.38 5.96 13.53 6.11 ;
        RECT 13.38 2.805 13.53 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 28.54 5.86 28.88 6.21 ;
        RECT 28.54 2.705 28.88 3.055 ;
        RECT 28.62 2.705 28.79 6.21 ;
      LAYER li1 ;
        RECT 28.62 1.66 28.79 2.935 ;
        RECT 28.62 5.945 28.79 7.22 ;
        RECT 23.005 5.945 23.175 7.22 ;
      LAYER met1 ;
        RECT 28.54 2.765 29.02 2.935 ;
        RECT 28.54 2.705 28.88 3.055 ;
        RECT 22.945 5.945 29.02 6.115 ;
        RECT 28.54 5.86 28.88 6.21 ;
        RECT 22.945 5.915 23.235 6.145 ;
      LAYER mcon ;
        RECT 23.005 5.945 23.175 6.115 ;
        RECT 28.62 5.945 28.79 6.115 ;
        RECT 28.62 2.765 28.79 2.935 ;
      LAYER via1 ;
        RECT 28.64 5.96 28.79 6.11 ;
        RECT 28.64 2.805 28.79 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 43.8 5.86 44.14 6.21 ;
        RECT 43.8 2.705 44.14 3.055 ;
        RECT 43.88 2.705 44.05 6.21 ;
      LAYER li1 ;
        RECT 43.88 1.66 44.05 2.935 ;
        RECT 43.88 5.945 44.05 7.22 ;
        RECT 38.265 5.945 38.435 7.22 ;
      LAYER met1 ;
        RECT 43.8 2.765 44.28 2.935 ;
        RECT 43.8 2.705 44.14 3.055 ;
        RECT 38.205 5.945 44.28 6.115 ;
        RECT 43.8 5.86 44.14 6.21 ;
        RECT 38.205 5.915 38.495 6.145 ;
      LAYER mcon ;
        RECT 38.265 5.945 38.435 6.115 ;
        RECT 43.88 5.945 44.05 6.115 ;
        RECT 43.88 2.765 44.05 2.935 ;
      LAYER via1 ;
        RECT 43.9 5.96 44.05 6.11 ;
        RECT 43.9 2.805 44.05 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 59.06 5.86 59.4 6.21 ;
        RECT 59.06 2.705 59.4 3.055 ;
        RECT 59.14 2.705 59.31 6.21 ;
      LAYER li1 ;
        RECT 59.14 1.66 59.31 2.935 ;
        RECT 59.14 5.945 59.31 7.22 ;
        RECT 53.525 5.945 53.695 7.22 ;
      LAYER met1 ;
        RECT 59.06 2.765 59.54 2.935 ;
        RECT 59.06 2.705 59.4 3.055 ;
        RECT 53.465 5.945 59.54 6.115 ;
        RECT 59.06 5.86 59.4 6.21 ;
        RECT 53.465 5.915 53.755 6.145 ;
      LAYER mcon ;
        RECT 53.525 5.945 53.695 6.115 ;
        RECT 59.14 5.945 59.31 6.115 ;
        RECT 59.14 2.765 59.31 2.935 ;
      LAYER via1 ;
        RECT 59.16 5.96 59.31 6.11 ;
        RECT 59.16 2.805 59.31 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 74.32 5.86 74.66 6.21 ;
        RECT 74.32 2.705 74.66 3.055 ;
        RECT 74.4 2.705 74.57 6.21 ;
      LAYER li1 ;
        RECT 74.4 1.66 74.57 2.935 ;
        RECT 74.4 5.945 74.57 7.22 ;
        RECT 68.785 5.945 68.955 7.22 ;
      LAYER met1 ;
        RECT 74.32 2.765 74.8 2.935 ;
        RECT 74.32 2.705 74.66 3.055 ;
        RECT 68.725 5.945 74.8 6.115 ;
        RECT 74.32 5.86 74.66 6.21 ;
        RECT 68.725 5.915 69.015 6.145 ;
      LAYER mcon ;
        RECT 68.785 5.945 68.955 6.115 ;
        RECT 74.4 5.945 74.57 6.115 ;
        RECT 74.4 2.765 74.57 2.935 ;
      LAYER via1 ;
        RECT 74.42 5.96 74.57 6.11 ;
        RECT 74.42 2.805 74.57 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 5.945 0.4 7.22 ;
      LAYER met1 ;
        RECT 0.17 5.945 0.63 6.115 ;
        RECT 0.17 5.915 0.46 6.145 ;
      LAYER mcon ;
        RECT 0.23 5.945 0.4 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.48 4.275 2.285 4.655 ;
      LAYER met2 ;
        RECT 1.67 4.275 2.05 4.655 ;
      LAYER li1 ;
        RECT 0 4.44 79.095 4.745 ;
        RECT 72.155 4.135 79.095 4.745 ;
        RECT 76.96 4.13 78.94 4.75 ;
        RECT 78.12 3.4 78.29 5.48 ;
        RECT 77.13 3.4 77.3 5.48 ;
        RECT 74.39 3.405 74.56 5.475 ;
        RECT 64.585 4.13 73.325 4.3 ;
        RECT 1.945 4.305 79.095 4.745 ;
        RECT 71.615 3.63 71.785 4.3 ;
        RECT 69.695 3.63 69.865 4.3 ;
        RECT 68.775 4.305 68.945 5.475 ;
        RECT 68.755 3.63 68.925 4.3 ;
        RECT 67.295 3.63 67.465 4.3 ;
        RECT 65.375 3.63 65.545 4.3 ;
        RECT 56.895 4.14 64.59 4.745 ;
        RECT 49.325 4.135 63.835 4.3 ;
        RECT 61.7 4.13 63.68 4.75 ;
        RECT 62.86 3.4 63.03 5.48 ;
        RECT 61.87 3.4 62.04 5.48 ;
        RECT 59.13 3.405 59.3 5.475 ;
        RECT 49.325 4.13 58.065 4.3 ;
        RECT 56.355 3.63 56.525 4.3 ;
        RECT 54.435 3.63 54.605 4.3 ;
        RECT 53.515 4.305 53.685 5.475 ;
        RECT 53.495 3.63 53.665 4.3 ;
        RECT 52.035 3.63 52.205 4.3 ;
        RECT 50.115 3.63 50.285 4.3 ;
        RECT 41.635 4.14 49.33 4.745 ;
        RECT 34.065 4.135 48.575 4.3 ;
        RECT 46.44 4.13 48.42 4.75 ;
        RECT 47.6 3.4 47.77 5.48 ;
        RECT 46.61 3.4 46.78 5.48 ;
        RECT 43.87 3.405 44.04 5.475 ;
        RECT 34.065 4.13 42.805 4.3 ;
        RECT 41.095 3.63 41.265 4.3 ;
        RECT 39.175 3.63 39.345 4.3 ;
        RECT 38.255 4.305 38.425 5.475 ;
        RECT 38.235 3.63 38.405 4.3 ;
        RECT 36.775 3.63 36.945 4.3 ;
        RECT 34.855 3.63 35.025 4.3 ;
        RECT 26.375 4.14 34.07 4.745 ;
        RECT 18.805 4.135 33.315 4.3 ;
        RECT 31.18 4.13 33.16 4.75 ;
        RECT 32.34 3.4 32.51 5.48 ;
        RECT 31.35 3.4 31.52 5.48 ;
        RECT 28.61 3.405 28.78 5.475 ;
        RECT 18.805 4.13 27.545 4.3 ;
        RECT 25.835 3.63 26.005 4.3 ;
        RECT 23.915 3.63 24.085 4.3 ;
        RECT 22.995 4.305 23.165 5.475 ;
        RECT 22.975 3.63 23.145 4.3 ;
        RECT 21.515 3.63 21.685 4.3 ;
        RECT 19.595 3.63 19.765 4.3 ;
        RECT 11.115 4.14 18.81 4.745 ;
        RECT 3.545 4.135 18.055 4.3 ;
        RECT 15.92 4.13 17.9 4.75 ;
        RECT 17.08 3.4 17.25 5.48 ;
        RECT 16.09 3.4 16.26 5.48 ;
        RECT 13.35 3.405 13.52 5.475 ;
        RECT 3.545 4.13 12.285 4.3 ;
        RECT 10.575 3.63 10.745 4.3 ;
        RECT 8.655 3.63 8.825 4.3 ;
        RECT 7.735 4.305 7.905 5.475 ;
        RECT 7.715 3.63 7.885 4.3 ;
        RECT 6.255 3.63 6.425 4.3 ;
        RECT 4.335 3.63 4.505 4.3 ;
        RECT 0 4.14 3.69 4.35 ;
        RECT 2.03 4.14 2.2 8.305 ;
        RECT 0 4.14 1.775 4.745 ;
        RECT 0.22 4.14 0.39 5.475 ;
      LAYER met1 ;
        RECT 0 4.14 79.095 4.745 ;
        RECT 64.585 4.135 79.095 4.745 ;
        RECT 76.96 4.13 78.94 4.75 ;
        RECT 64.585 3.98 73.325 4.745 ;
        RECT 49.325 4.135 63.835 4.745 ;
        RECT 61.7 4.13 63.68 4.75 ;
        RECT 49.325 3.98 58.065 4.745 ;
        RECT 34.065 4.135 48.575 4.745 ;
        RECT 46.44 4.13 48.42 4.75 ;
        RECT 34.065 3.98 42.805 4.745 ;
        RECT 18.805 4.135 33.315 4.745 ;
        RECT 31.18 4.13 33.16 4.75 ;
        RECT 18.805 3.98 27.545 4.745 ;
        RECT 3.545 4.135 18.055 4.745 ;
        RECT 15.92 4.13 17.9 4.75 ;
        RECT 3.545 3.98 12.285 4.745 ;
        RECT 1.97 6.655 2.26 6.885 ;
        RECT 1.8 6.685 2.26 6.855 ;
      LAYER via2 ;
        RECT 1.76 4.365 1.96 4.565 ;
      LAYER mcon ;
        RECT 2.03 6.685 2.2 6.855 ;
        RECT 2.34 4.545 2.51 4.715 ;
        RECT 3.685 4.13 3.855 4.3 ;
        RECT 4.145 4.13 4.315 4.3 ;
        RECT 4.605 4.13 4.775 4.3 ;
        RECT 5.065 4.13 5.235 4.3 ;
        RECT 5.525 4.13 5.695 4.3 ;
        RECT 5.985 4.13 6.155 4.3 ;
        RECT 6.445 4.13 6.615 4.3 ;
        RECT 6.905 4.13 7.075 4.3 ;
        RECT 7.365 4.13 7.535 4.3 ;
        RECT 7.825 4.13 7.995 4.3 ;
        RECT 8.285 4.13 8.455 4.3 ;
        RECT 8.745 4.13 8.915 4.3 ;
        RECT 9.205 4.13 9.375 4.3 ;
        RECT 9.665 4.13 9.835 4.3 ;
        RECT 9.855 4.545 10.025 4.715 ;
        RECT 10.125 4.13 10.295 4.3 ;
        RECT 10.585 4.13 10.755 4.3 ;
        RECT 11.045 4.13 11.215 4.3 ;
        RECT 11.505 4.13 11.675 4.3 ;
        RECT 11.965 4.13 12.135 4.3 ;
        RECT 15.47 4.545 15.64 4.715 ;
        RECT 15.47 4.165 15.64 4.335 ;
        RECT 16.17 4.55 16.34 4.72 ;
        RECT 16.17 4.16 16.34 4.33 ;
        RECT 17.16 4.55 17.33 4.72 ;
        RECT 17.16 4.16 17.33 4.33 ;
        RECT 18.945 4.13 19.115 4.3 ;
        RECT 19.405 4.13 19.575 4.3 ;
        RECT 19.865 4.13 20.035 4.3 ;
        RECT 20.325 4.13 20.495 4.3 ;
        RECT 20.785 4.13 20.955 4.3 ;
        RECT 21.245 4.13 21.415 4.3 ;
        RECT 21.705 4.13 21.875 4.3 ;
        RECT 22.165 4.13 22.335 4.3 ;
        RECT 22.625 4.13 22.795 4.3 ;
        RECT 23.085 4.13 23.255 4.3 ;
        RECT 23.545 4.13 23.715 4.3 ;
        RECT 24.005 4.13 24.175 4.3 ;
        RECT 24.465 4.13 24.635 4.3 ;
        RECT 24.925 4.13 25.095 4.3 ;
        RECT 25.115 4.545 25.285 4.715 ;
        RECT 25.385 4.13 25.555 4.3 ;
        RECT 25.845 4.13 26.015 4.3 ;
        RECT 26.305 4.13 26.475 4.3 ;
        RECT 26.765 4.13 26.935 4.3 ;
        RECT 27.225 4.13 27.395 4.3 ;
        RECT 30.73 4.545 30.9 4.715 ;
        RECT 30.73 4.165 30.9 4.335 ;
        RECT 31.43 4.55 31.6 4.72 ;
        RECT 31.43 4.16 31.6 4.33 ;
        RECT 32.42 4.55 32.59 4.72 ;
        RECT 32.42 4.16 32.59 4.33 ;
        RECT 34.205 4.13 34.375 4.3 ;
        RECT 34.665 4.13 34.835 4.3 ;
        RECT 35.125 4.13 35.295 4.3 ;
        RECT 35.585 4.13 35.755 4.3 ;
        RECT 36.045 4.13 36.215 4.3 ;
        RECT 36.505 4.13 36.675 4.3 ;
        RECT 36.965 4.13 37.135 4.3 ;
        RECT 37.425 4.13 37.595 4.3 ;
        RECT 37.885 4.13 38.055 4.3 ;
        RECT 38.345 4.13 38.515 4.3 ;
        RECT 38.805 4.13 38.975 4.3 ;
        RECT 39.265 4.13 39.435 4.3 ;
        RECT 39.725 4.13 39.895 4.3 ;
        RECT 40.185 4.13 40.355 4.3 ;
        RECT 40.375 4.545 40.545 4.715 ;
        RECT 40.645 4.13 40.815 4.3 ;
        RECT 41.105 4.13 41.275 4.3 ;
        RECT 41.565 4.13 41.735 4.3 ;
        RECT 42.025 4.13 42.195 4.3 ;
        RECT 42.485 4.13 42.655 4.3 ;
        RECT 45.99 4.545 46.16 4.715 ;
        RECT 45.99 4.165 46.16 4.335 ;
        RECT 46.69 4.55 46.86 4.72 ;
        RECT 46.69 4.16 46.86 4.33 ;
        RECT 47.68 4.55 47.85 4.72 ;
        RECT 47.68 4.16 47.85 4.33 ;
        RECT 49.465 4.13 49.635 4.3 ;
        RECT 49.925 4.13 50.095 4.3 ;
        RECT 50.385 4.13 50.555 4.3 ;
        RECT 50.845 4.13 51.015 4.3 ;
        RECT 51.305 4.13 51.475 4.3 ;
        RECT 51.765 4.13 51.935 4.3 ;
        RECT 52.225 4.13 52.395 4.3 ;
        RECT 52.685 4.13 52.855 4.3 ;
        RECT 53.145 4.13 53.315 4.3 ;
        RECT 53.605 4.13 53.775 4.3 ;
        RECT 54.065 4.13 54.235 4.3 ;
        RECT 54.525 4.13 54.695 4.3 ;
        RECT 54.985 4.13 55.155 4.3 ;
        RECT 55.445 4.13 55.615 4.3 ;
        RECT 55.635 4.545 55.805 4.715 ;
        RECT 55.905 4.13 56.075 4.3 ;
        RECT 56.365 4.13 56.535 4.3 ;
        RECT 56.825 4.13 56.995 4.3 ;
        RECT 57.285 4.13 57.455 4.3 ;
        RECT 57.745 4.13 57.915 4.3 ;
        RECT 61.25 4.545 61.42 4.715 ;
        RECT 61.25 4.165 61.42 4.335 ;
        RECT 61.95 4.55 62.12 4.72 ;
        RECT 61.95 4.16 62.12 4.33 ;
        RECT 62.94 4.55 63.11 4.72 ;
        RECT 62.94 4.16 63.11 4.33 ;
        RECT 64.725 4.13 64.895 4.3 ;
        RECT 65.185 4.13 65.355 4.3 ;
        RECT 65.645 4.13 65.815 4.3 ;
        RECT 66.105 4.13 66.275 4.3 ;
        RECT 66.565 4.13 66.735 4.3 ;
        RECT 67.025 4.13 67.195 4.3 ;
        RECT 67.485 4.13 67.655 4.3 ;
        RECT 67.945 4.13 68.115 4.3 ;
        RECT 68.405 4.13 68.575 4.3 ;
        RECT 68.865 4.13 69.035 4.3 ;
        RECT 69.325 4.13 69.495 4.3 ;
        RECT 69.785 4.13 69.955 4.3 ;
        RECT 70.245 4.13 70.415 4.3 ;
        RECT 70.705 4.13 70.875 4.3 ;
        RECT 70.895 4.545 71.065 4.715 ;
        RECT 71.165 4.13 71.335 4.3 ;
        RECT 71.625 4.13 71.795 4.3 ;
        RECT 72.085 4.13 72.255 4.3 ;
        RECT 72.545 4.13 72.715 4.3 ;
        RECT 73.005 4.13 73.175 4.3 ;
        RECT 76.51 4.545 76.68 4.715 ;
        RECT 76.51 4.165 76.68 4.335 ;
        RECT 77.21 4.55 77.38 4.72 ;
        RECT 77.21 4.16 77.38 4.33 ;
        RECT 78.2 4.55 78.37 4.72 ;
        RECT 78.2 4.16 78.37 4.33 ;
      LAYER via1 ;
        RECT 1.785 4.39 1.935 4.54 ;
    END
  END vccd1
  OBS
    LAYER met4 ;
      RECT 66.735 2.97 67.065 3.3 ;
      RECT 66.745 2.5 67.065 3.3 ;
      RECT 68.895 2.48 69.225 2.84 ;
      RECT 66.745 2.5 69.225 2.8 ;
      RECT 51.475 2.97 51.805 3.3 ;
      RECT 51.485 2.5 51.805 3.3 ;
      RECT 53.635 2.48 53.965 2.84 ;
      RECT 51.485 2.5 53.965 2.8 ;
      RECT 36.215 2.97 36.545 3.3 ;
      RECT 36.225 2.5 36.545 3.3 ;
      RECT 38.375 2.48 38.705 2.84 ;
      RECT 36.225 2.5 38.705 2.8 ;
      RECT 20.955 2.97 21.285 3.3 ;
      RECT 20.965 2.5 21.285 3.3 ;
      RECT 23.115 2.48 23.445 2.84 ;
      RECT 20.965 2.5 23.445 2.8 ;
      RECT 5.695 2.97 6.025 3.3 ;
      RECT 5.705 2.5 6.025 3.3 ;
      RECT 7.855 2.48 8.185 2.84 ;
      RECT 5.705 2.5 8.185 2.8 ;
    LAYER via3 ;
      RECT 68.955 2.57 69.155 2.77 ;
      RECT 66.795 3.04 66.995 3.24 ;
      RECT 53.695 2.57 53.895 2.77 ;
      RECT 51.535 3.04 51.735 3.24 ;
      RECT 38.435 2.57 38.635 2.77 ;
      RECT 36.275 3.04 36.475 3.24 ;
      RECT 23.175 2.57 23.375 2.77 ;
      RECT 21.015 3.04 21.215 3.24 ;
      RECT 7.915 2.57 8.115 2.77 ;
      RECT 5.755 3.04 5.955 3.24 ;
    LAYER met3 ;
      RECT 73.76 1.105 74.1 3.065 ;
      RECT 68.015 1.88 68.745 2.21 ;
      RECT 68.17 1.105 68.47 2.21 ;
      RECT 68.17 1.105 74.1 1.405 ;
      RECT 70.055 7.055 70.425 7.425 ;
      RECT 70.09 4.475 70.39 7.425 ;
      RECT 68.65 4.475 70.39 4.775 ;
      RECT 65.855 4.255 68.95 4.555 ;
      RECT 68.65 2.515 68.95 4.775 ;
      RECT 65.855 2.97 66.155 4.555 ;
      RECT 69.375 3.51 69.705 3.86 ;
      RECT 67.465 3.55 69.705 3.85 ;
      RECT 67.465 2.41 67.765 3.85 ;
      RECT 65.545 2.97 66.275 3.3 ;
      RECT 68.445 2.52 69.225 2.86 ;
      RECT 68.915 2.48 69.225 2.86 ;
      RECT 67.455 2.41 67.785 2.74 ;
      RECT 68.895 2.51 69.225 2.86 ;
      RECT 66.735 2.41 67.055 3.33 ;
      RECT 66.735 2.41 67.065 2.95 ;
      RECT 58.5 1.105 58.84 3.065 ;
      RECT 52.755 1.88 53.485 2.21 ;
      RECT 52.91 1.105 53.21 2.21 ;
      RECT 52.91 1.105 58.84 1.405 ;
      RECT 54.795 7.055 55.165 7.425 ;
      RECT 54.83 4.475 55.13 7.425 ;
      RECT 53.39 4.475 55.13 4.775 ;
      RECT 50.595 4.255 53.69 4.555 ;
      RECT 53.39 2.515 53.69 4.775 ;
      RECT 50.595 2.97 50.895 4.555 ;
      RECT 54.115 3.51 54.445 3.86 ;
      RECT 52.205 3.55 54.445 3.85 ;
      RECT 52.205 2.41 52.505 3.85 ;
      RECT 50.285 2.97 51.015 3.3 ;
      RECT 53.185 2.52 53.965 2.86 ;
      RECT 53.655 2.48 53.965 2.86 ;
      RECT 52.195 2.41 52.525 2.74 ;
      RECT 53.635 2.51 53.965 2.86 ;
      RECT 51.475 2.41 51.795 3.33 ;
      RECT 51.475 2.41 51.805 2.95 ;
      RECT 43.24 1.105 43.58 3.065 ;
      RECT 37.495 1.88 38.225 2.21 ;
      RECT 37.65 1.105 37.95 2.21 ;
      RECT 37.65 1.105 43.58 1.405 ;
      RECT 39.535 7.055 39.905 7.425 ;
      RECT 39.57 4.475 39.87 7.425 ;
      RECT 38.13 4.475 39.87 4.775 ;
      RECT 35.335 4.255 38.43 4.555 ;
      RECT 38.13 2.515 38.43 4.775 ;
      RECT 35.335 2.97 35.635 4.555 ;
      RECT 38.855 3.51 39.185 3.86 ;
      RECT 36.945 3.55 39.185 3.85 ;
      RECT 36.945 2.41 37.245 3.85 ;
      RECT 35.025 2.97 35.755 3.3 ;
      RECT 37.925 2.52 38.705 2.86 ;
      RECT 38.395 2.48 38.705 2.86 ;
      RECT 36.935 2.41 37.265 2.74 ;
      RECT 38.375 2.51 38.705 2.86 ;
      RECT 36.215 2.41 36.535 3.33 ;
      RECT 36.215 2.41 36.545 2.95 ;
      RECT 27.98 1.105 28.32 3.065 ;
      RECT 22.235 1.88 22.965 2.21 ;
      RECT 22.39 1.105 22.69 2.21 ;
      RECT 22.39 1.105 28.32 1.405 ;
      RECT 24.275 7.055 24.645 7.425 ;
      RECT 24.31 4.475 24.61 7.425 ;
      RECT 22.87 4.475 24.61 4.775 ;
      RECT 20.075 4.255 23.17 4.555 ;
      RECT 22.87 2.515 23.17 4.775 ;
      RECT 20.075 2.97 20.375 4.555 ;
      RECT 23.595 3.51 23.925 3.86 ;
      RECT 21.685 3.55 23.925 3.85 ;
      RECT 21.685 2.41 21.985 3.85 ;
      RECT 19.765 2.97 20.495 3.3 ;
      RECT 22.665 2.52 23.445 2.86 ;
      RECT 23.135 2.48 23.445 2.86 ;
      RECT 21.675 2.41 22.005 2.74 ;
      RECT 23.115 2.51 23.445 2.86 ;
      RECT 20.955 2.41 21.275 3.33 ;
      RECT 20.955 2.41 21.285 2.95 ;
      RECT 12.72 1.105 13.06 3.065 ;
      RECT 6.975 1.88 7.705 2.21 ;
      RECT 7.13 1.105 7.43 2.21 ;
      RECT 7.13 1.105 13.06 1.405 ;
      RECT 9.015 7.055 9.385 7.425 ;
      RECT 9.05 4.475 9.35 7.425 ;
      RECT 7.61 4.475 9.35 4.775 ;
      RECT 4.815 4.255 7.91 4.555 ;
      RECT 7.61 2.515 7.91 4.775 ;
      RECT 4.815 2.97 5.115 4.555 ;
      RECT 8.335 3.51 8.665 3.86 ;
      RECT 6.425 3.55 8.665 3.85 ;
      RECT 6.425 2.41 6.725 3.85 ;
      RECT 4.505 2.97 5.235 3.3 ;
      RECT 7.405 2.52 8.185 2.86 ;
      RECT 7.875 2.48 8.185 2.86 ;
      RECT 6.415 2.41 6.745 2.74 ;
      RECT 7.855 2.51 8.185 2.86 ;
      RECT 5.695 2.41 6.015 3.33 ;
      RECT 5.695 2.41 6.025 2.95 ;
      RECT 72.295 1.85 73.025 2.18 ;
      RECT 70.605 1.87 71.335 2.2 ;
      RECT 69.565 1.85 70.295 2.2 ;
      RECT 65.415 1.85 66.145 2.18 ;
      RECT 57.035 1.85 57.765 2.18 ;
      RECT 55.345 1.87 56.075 2.2 ;
      RECT 54.305 1.85 55.035 2.2 ;
      RECT 50.155 1.85 50.885 2.18 ;
      RECT 41.775 1.85 42.505 2.18 ;
      RECT 40.085 1.87 40.815 2.2 ;
      RECT 39.045 1.85 39.775 2.2 ;
      RECT 34.895 1.85 35.625 2.18 ;
      RECT 26.515 1.85 27.245 2.18 ;
      RECT 24.825 1.87 25.555 2.2 ;
      RECT 23.785 1.85 24.515 2.2 ;
      RECT 19.635 1.85 20.365 2.18 ;
      RECT 11.255 1.85 11.985 2.18 ;
      RECT 9.565 1.87 10.295 2.2 ;
      RECT 8.525 1.85 9.255 2.2 ;
      RECT 4.375 1.85 5.105 2.18 ;
      RECT 0.005 8.5 0.81 8.88 ;
      RECT 0 0 0.805 0.38 ;
    LAYER via2 ;
      RECT 73.835 2.775 74.035 2.975 ;
      RECT 72.525 1.92 72.725 2.12 ;
      RECT 70.665 1.93 70.865 2.13 ;
      RECT 70.14 7.14 70.34 7.34 ;
      RECT 69.645 1.94 69.845 2.14 ;
      RECT 69.435 3.57 69.635 3.77 ;
      RECT 68.955 2.57 69.155 2.77 ;
      RECT 68.205 1.94 68.405 2.14 ;
      RECT 67.515 2.48 67.715 2.68 ;
      RECT 66.805 2.48 67.005 2.68 ;
      RECT 65.835 3.04 66.035 3.24 ;
      RECT 65.595 1.92 65.795 2.12 ;
      RECT 58.575 2.775 58.775 2.975 ;
      RECT 57.265 1.92 57.465 2.12 ;
      RECT 55.405 1.93 55.605 2.13 ;
      RECT 54.88 7.14 55.08 7.34 ;
      RECT 54.385 1.94 54.585 2.14 ;
      RECT 54.175 3.57 54.375 3.77 ;
      RECT 53.695 2.57 53.895 2.77 ;
      RECT 52.945 1.94 53.145 2.14 ;
      RECT 52.255 2.48 52.455 2.68 ;
      RECT 51.545 2.48 51.745 2.68 ;
      RECT 50.575 3.04 50.775 3.24 ;
      RECT 50.335 1.92 50.535 2.12 ;
      RECT 43.315 2.775 43.515 2.975 ;
      RECT 42.005 1.92 42.205 2.12 ;
      RECT 40.145 1.93 40.345 2.13 ;
      RECT 39.62 7.14 39.82 7.34 ;
      RECT 39.125 1.94 39.325 2.14 ;
      RECT 38.915 3.57 39.115 3.77 ;
      RECT 38.435 2.57 38.635 2.77 ;
      RECT 37.685 1.94 37.885 2.14 ;
      RECT 36.995 2.48 37.195 2.68 ;
      RECT 36.285 2.48 36.485 2.68 ;
      RECT 35.315 3.04 35.515 3.24 ;
      RECT 35.075 1.92 35.275 2.12 ;
      RECT 28.055 2.775 28.255 2.975 ;
      RECT 26.745 1.92 26.945 2.12 ;
      RECT 24.885 1.93 25.085 2.13 ;
      RECT 24.36 7.14 24.56 7.34 ;
      RECT 23.865 1.94 24.065 2.14 ;
      RECT 23.655 3.57 23.855 3.77 ;
      RECT 23.175 2.57 23.375 2.77 ;
      RECT 22.425 1.94 22.625 2.14 ;
      RECT 21.735 2.48 21.935 2.68 ;
      RECT 21.025 2.48 21.225 2.68 ;
      RECT 20.055 3.04 20.255 3.24 ;
      RECT 19.815 1.92 20.015 2.12 ;
      RECT 12.795 2.775 12.995 2.975 ;
      RECT 11.485 1.92 11.685 2.12 ;
      RECT 9.625 1.93 9.825 2.13 ;
      RECT 9.1 7.14 9.3 7.34 ;
      RECT 8.605 1.94 8.805 2.14 ;
      RECT 8.395 3.57 8.595 3.77 ;
      RECT 7.915 2.57 8.115 2.77 ;
      RECT 7.165 1.94 7.365 2.14 ;
      RECT 6.475 2.48 6.675 2.68 ;
      RECT 5.765 2.48 5.965 2.68 ;
      RECT 4.795 3.04 4.995 3.24 ;
      RECT 4.555 1.92 4.755 2.12 ;
      RECT 0.285 8.59 0.485 8.79 ;
      RECT 0.28 0.09 0.48 0.29 ;
    LAYER met2 ;
      RECT 1.23 8.4 78.725 8.57 ;
      RECT 78.555 7.275 78.725 8.57 ;
      RECT 1.23 6.255 1.4 8.57 ;
      RECT 78.525 7.275 78.875 7.625 ;
      RECT 1.165 6.255 1.455 6.605 ;
      RECT 75.365 6.22 75.685 6.545 ;
      RECT 75.395 5.695 75.565 6.545 ;
      RECT 75.395 5.695 75.57 6.045 ;
      RECT 75.395 5.695 76.37 5.87 ;
      RECT 76.195 1.965 76.37 5.87 ;
      RECT 76.14 1.965 76.49 2.315 ;
      RECT 76.165 6.655 76.49 6.98 ;
      RECT 75.05 6.745 76.49 6.915 ;
      RECT 75.05 2.395 75.21 6.915 ;
      RECT 75.365 2.365 75.685 2.685 ;
      RECT 75.05 2.395 75.685 2.565 ;
      RECT 73.79 2.685 74.08 3.065 ;
      RECT 73.76 2.7 74.1 3.05 ;
      RECT 72.495 3.54 72.755 3.86 ;
      RECT 72.555 1.83 72.695 3.86 ;
      RECT 72.385 2.39 72.695 2.76 ;
      RECT 72.455 1.95 72.695 2.76 ;
      RECT 72.485 1.83 72.765 2.2 ;
      RECT 72.485 1.94 72.77 2.14 ;
      RECT 71.805 2.42 72.065 2.74 ;
      RECT 71.145 2.51 72.065 2.65 ;
      RECT 71.145 1.57 71.285 2.65 ;
      RECT 67.605 1.86 67.865 2.18 ;
      RECT 67.785 1.57 67.925 2.09 ;
      RECT 67.785 1.57 71.285 1.71 ;
      RECT 63.24 6.655 63.59 7.005 ;
      RECT 70.725 6.61 71.075 6.96 ;
      RECT 63.24 6.685 71.075 6.885 ;
      RECT 70.635 3.26 70.895 3.58 ;
      RECT 70.695 1.85 70.835 3.58 ;
      RECT 70.625 1.85 70.905 2.22 ;
      RECT 68.025 4.01 70.465 4.15 ;
      RECT 70.325 2.7 70.465 4.15 ;
      RECT 68.025 3.63 68.165 4.15 ;
      RECT 67.725 3.63 68.165 3.86 ;
      RECT 65.385 3.63 68.165 3.77 ;
      RECT 67.725 3.54 67.985 3.86 ;
      RECT 65.385 3.35 65.525 3.77 ;
      RECT 64.875 3.26 65.135 3.58 ;
      RECT 64.875 3.35 65.525 3.49 ;
      RECT 64.935 1.86 65.075 3.58 ;
      RECT 70.265 2.7 70.525 3.02 ;
      RECT 64.875 1.86 65.135 2.18 ;
      RECT 69.885 3.54 70.145 3.86 ;
      RECT 69.945 1.95 70.085 3.86 ;
      RECT 69.605 1.95 70.085 2.22 ;
      RECT 69.405 1.85 69.885 2.2 ;
      RECT 69.395 3.49 69.675 3.86 ;
      RECT 69.465 2.39 69.605 3.86 ;
      RECT 69.405 2.39 69.665 3.02 ;
      RECT 69.395 2.39 69.675 2.76 ;
      RECT 68.325 3.54 68.585 3.86 ;
      RECT 68.325 3.35 68.525 3.86 ;
      RECT 68.135 3.35 68.525 3.49 ;
      RECT 68.135 1.86 68.275 3.49 ;
      RECT 68.135 1.86 68.445 2.23 ;
      RECT 68.075 1.86 68.445 2.18 ;
      RECT 65.795 2.95 66.075 3.32 ;
      RECT 67.245 2.98 67.505 3.3 ;
      RECT 65.625 3.07 67.505 3.21 ;
      RECT 65.625 2.95 66.075 3.21 ;
      RECT 65.565 2.39 65.825 3.02 ;
      RECT 65.555 2.39 65.835 2.76 ;
      RECT 66.635 2.39 67.045 2.76 ;
      RECT 66.045 2.42 66.305 2.74 ;
      RECT 66.045 2.51 67.045 2.65 ;
      RECT 65.555 1.83 65.835 2.2 ;
      RECT 65.555 1.86 65.945 2.18 ;
      RECT 60.105 6.22 60.425 6.545 ;
      RECT 60.135 5.695 60.305 6.545 ;
      RECT 60.135 5.695 60.31 6.045 ;
      RECT 60.135 5.695 61.11 5.87 ;
      RECT 60.935 1.965 61.11 5.87 ;
      RECT 60.88 1.965 61.23 2.315 ;
      RECT 60.905 6.655 61.23 6.98 ;
      RECT 59.79 6.745 61.23 6.915 ;
      RECT 59.79 2.395 59.95 6.915 ;
      RECT 60.105 2.365 60.425 2.685 ;
      RECT 59.79 2.395 60.425 2.565 ;
      RECT 58.53 2.685 58.82 3.065 ;
      RECT 58.5 2.7 58.84 3.05 ;
      RECT 57.235 3.54 57.495 3.86 ;
      RECT 57.295 1.83 57.435 3.86 ;
      RECT 57.125 2.39 57.435 2.76 ;
      RECT 57.195 1.95 57.435 2.76 ;
      RECT 57.225 1.83 57.505 2.2 ;
      RECT 57.225 1.94 57.51 2.14 ;
      RECT 56.545 2.42 56.805 2.74 ;
      RECT 55.885 2.51 56.805 2.65 ;
      RECT 55.885 1.57 56.025 2.65 ;
      RECT 52.345 1.86 52.605 2.18 ;
      RECT 52.525 1.57 52.665 2.09 ;
      RECT 52.525 1.57 56.025 1.71 ;
      RECT 47.98 6.655 48.33 7.005 ;
      RECT 55.47 6.61 55.82 6.96 ;
      RECT 47.98 6.685 55.82 6.885 ;
      RECT 55.375 3.26 55.635 3.58 ;
      RECT 55.435 1.85 55.575 3.58 ;
      RECT 55.365 1.85 55.645 2.22 ;
      RECT 52.765 4.01 55.205 4.15 ;
      RECT 55.065 2.7 55.205 4.15 ;
      RECT 52.765 3.63 52.905 4.15 ;
      RECT 52.465 3.63 52.905 3.86 ;
      RECT 50.125 3.63 52.905 3.77 ;
      RECT 52.465 3.54 52.725 3.86 ;
      RECT 50.125 3.35 50.265 3.77 ;
      RECT 49.615 3.26 49.875 3.58 ;
      RECT 49.615 3.35 50.265 3.49 ;
      RECT 49.675 1.86 49.815 3.58 ;
      RECT 55.005 2.7 55.265 3.02 ;
      RECT 49.615 1.86 49.875 2.18 ;
      RECT 54.625 3.54 54.885 3.86 ;
      RECT 54.685 1.95 54.825 3.86 ;
      RECT 54.345 1.95 54.825 2.22 ;
      RECT 54.145 1.85 54.625 2.2 ;
      RECT 54.135 3.49 54.415 3.86 ;
      RECT 54.205 2.39 54.345 3.86 ;
      RECT 54.145 2.39 54.405 3.02 ;
      RECT 54.135 2.39 54.415 2.76 ;
      RECT 53.065 3.54 53.325 3.86 ;
      RECT 53.065 3.35 53.265 3.86 ;
      RECT 52.875 3.35 53.265 3.49 ;
      RECT 52.875 1.86 53.015 3.49 ;
      RECT 52.875 1.86 53.185 2.23 ;
      RECT 52.815 1.86 53.185 2.18 ;
      RECT 50.535 2.95 50.815 3.32 ;
      RECT 51.985 2.98 52.245 3.3 ;
      RECT 50.365 3.07 52.245 3.21 ;
      RECT 50.365 2.95 50.815 3.21 ;
      RECT 50.305 2.39 50.565 3.02 ;
      RECT 50.295 2.39 50.575 2.76 ;
      RECT 51.375 2.39 51.785 2.76 ;
      RECT 50.785 2.42 51.045 2.74 ;
      RECT 50.785 2.51 51.785 2.65 ;
      RECT 50.295 1.83 50.575 2.2 ;
      RECT 50.295 1.86 50.685 2.18 ;
      RECT 44.845 6.22 45.165 6.545 ;
      RECT 44.875 5.695 45.045 6.545 ;
      RECT 44.875 5.695 45.05 6.045 ;
      RECT 44.875 5.695 45.85 5.87 ;
      RECT 45.675 1.965 45.85 5.87 ;
      RECT 45.62 1.965 45.97 2.315 ;
      RECT 45.645 6.655 45.97 6.98 ;
      RECT 44.53 6.745 45.97 6.915 ;
      RECT 44.53 2.395 44.69 6.915 ;
      RECT 44.845 2.365 45.165 2.685 ;
      RECT 44.53 2.395 45.165 2.565 ;
      RECT 43.27 2.685 43.56 3.065 ;
      RECT 43.24 2.7 43.58 3.05 ;
      RECT 41.975 3.54 42.235 3.86 ;
      RECT 42.035 1.83 42.175 3.86 ;
      RECT 41.865 2.39 42.175 2.76 ;
      RECT 41.935 1.95 42.175 2.76 ;
      RECT 41.965 1.83 42.245 2.2 ;
      RECT 41.965 1.94 42.25 2.14 ;
      RECT 41.285 2.42 41.545 2.74 ;
      RECT 40.625 2.51 41.545 2.65 ;
      RECT 40.625 1.57 40.765 2.65 ;
      RECT 37.085 1.86 37.345 2.18 ;
      RECT 37.265 1.57 37.405 2.09 ;
      RECT 37.265 1.57 40.765 1.71 ;
      RECT 32.765 6.66 33.115 7.01 ;
      RECT 40.205 6.615 40.555 6.965 ;
      RECT 32.765 6.69 40.555 6.89 ;
      RECT 40.115 3.26 40.375 3.58 ;
      RECT 40.175 1.85 40.315 3.58 ;
      RECT 40.105 1.85 40.385 2.22 ;
      RECT 37.505 4.01 39.945 4.15 ;
      RECT 39.805 2.7 39.945 4.15 ;
      RECT 37.505 3.63 37.645 4.15 ;
      RECT 37.205 3.63 37.645 3.86 ;
      RECT 34.865 3.63 37.645 3.77 ;
      RECT 37.205 3.54 37.465 3.86 ;
      RECT 34.865 3.35 35.005 3.77 ;
      RECT 34.355 3.26 34.615 3.58 ;
      RECT 34.355 3.35 35.005 3.49 ;
      RECT 34.415 1.86 34.555 3.58 ;
      RECT 39.745 2.7 40.005 3.02 ;
      RECT 34.355 1.86 34.615 2.18 ;
      RECT 39.365 3.54 39.625 3.86 ;
      RECT 39.425 1.95 39.565 3.86 ;
      RECT 39.085 1.95 39.565 2.22 ;
      RECT 38.885 1.85 39.365 2.2 ;
      RECT 38.875 3.49 39.155 3.86 ;
      RECT 38.945 2.39 39.085 3.86 ;
      RECT 38.885 2.39 39.145 3.02 ;
      RECT 38.875 2.39 39.155 2.76 ;
      RECT 37.805 3.54 38.065 3.86 ;
      RECT 37.805 3.35 38.005 3.86 ;
      RECT 37.615 3.35 38.005 3.49 ;
      RECT 37.615 1.86 37.755 3.49 ;
      RECT 37.615 1.86 37.925 2.23 ;
      RECT 37.555 1.86 37.925 2.18 ;
      RECT 35.275 2.95 35.555 3.32 ;
      RECT 36.725 2.98 36.985 3.3 ;
      RECT 35.105 3.07 36.985 3.21 ;
      RECT 35.105 2.95 35.555 3.21 ;
      RECT 35.045 2.39 35.305 3.02 ;
      RECT 35.035 2.39 35.315 2.76 ;
      RECT 36.115 2.39 36.525 2.76 ;
      RECT 35.525 2.42 35.785 2.74 ;
      RECT 35.525 2.51 36.525 2.65 ;
      RECT 35.035 1.83 35.315 2.2 ;
      RECT 35.035 1.86 35.425 2.18 ;
      RECT 29.585 6.22 29.905 6.545 ;
      RECT 29.615 5.695 29.785 6.545 ;
      RECT 29.615 5.695 29.79 6.045 ;
      RECT 29.615 5.695 30.59 5.87 ;
      RECT 30.415 1.965 30.59 5.87 ;
      RECT 30.36 1.965 30.71 2.315 ;
      RECT 30.385 6.655 30.71 6.98 ;
      RECT 29.27 6.745 30.71 6.915 ;
      RECT 29.27 2.395 29.43 6.915 ;
      RECT 29.585 2.365 29.905 2.685 ;
      RECT 29.27 2.395 29.905 2.565 ;
      RECT 28.01 2.685 28.3 3.065 ;
      RECT 27.98 2.7 28.32 3.05 ;
      RECT 26.715 3.54 26.975 3.86 ;
      RECT 26.775 1.83 26.915 3.86 ;
      RECT 26.605 2.39 26.915 2.76 ;
      RECT 26.675 1.95 26.915 2.76 ;
      RECT 26.705 1.83 26.985 2.2 ;
      RECT 26.705 1.94 26.99 2.14 ;
      RECT 26.025 2.42 26.285 2.74 ;
      RECT 25.365 2.51 26.285 2.65 ;
      RECT 25.365 1.57 25.505 2.65 ;
      RECT 21.825 1.86 22.085 2.18 ;
      RECT 22.005 1.57 22.145 2.09 ;
      RECT 22.005 1.57 25.505 1.71 ;
      RECT 17.505 6.655 17.855 7.005 ;
      RECT 24.945 6.61 25.295 6.96 ;
      RECT 17.505 6.685 25.295 6.885 ;
      RECT 24.855 3.26 25.115 3.58 ;
      RECT 24.915 1.85 25.055 3.58 ;
      RECT 24.845 1.85 25.125 2.22 ;
      RECT 22.245 4.01 24.685 4.15 ;
      RECT 24.545 2.7 24.685 4.15 ;
      RECT 22.245 3.63 22.385 4.15 ;
      RECT 21.945 3.63 22.385 3.86 ;
      RECT 19.605 3.63 22.385 3.77 ;
      RECT 21.945 3.54 22.205 3.86 ;
      RECT 19.605 3.35 19.745 3.77 ;
      RECT 19.095 3.26 19.355 3.58 ;
      RECT 19.095 3.35 19.745 3.49 ;
      RECT 19.155 1.86 19.295 3.58 ;
      RECT 24.485 2.7 24.745 3.02 ;
      RECT 19.095 1.86 19.355 2.18 ;
      RECT 24.105 3.54 24.365 3.86 ;
      RECT 24.165 1.95 24.305 3.86 ;
      RECT 23.825 1.95 24.305 2.22 ;
      RECT 23.625 1.85 24.105 2.2 ;
      RECT 23.615 3.49 23.895 3.86 ;
      RECT 23.685 2.39 23.825 3.86 ;
      RECT 23.625 2.39 23.885 3.02 ;
      RECT 23.615 2.39 23.895 2.76 ;
      RECT 22.545 3.54 22.805 3.86 ;
      RECT 22.545 3.35 22.745 3.86 ;
      RECT 22.355 3.35 22.745 3.49 ;
      RECT 22.355 1.86 22.495 3.49 ;
      RECT 22.355 1.86 22.665 2.23 ;
      RECT 22.295 1.86 22.665 2.18 ;
      RECT 20.015 2.95 20.295 3.32 ;
      RECT 21.465 2.98 21.725 3.3 ;
      RECT 19.845 3.07 21.725 3.21 ;
      RECT 19.845 2.95 20.295 3.21 ;
      RECT 19.785 2.39 20.045 3.02 ;
      RECT 19.775 2.39 20.055 2.76 ;
      RECT 20.855 2.39 21.265 2.76 ;
      RECT 20.265 2.42 20.525 2.74 ;
      RECT 20.265 2.51 21.265 2.65 ;
      RECT 19.775 1.83 20.055 2.2 ;
      RECT 19.775 1.86 20.165 2.18 ;
      RECT 14.325 6.22 14.645 6.545 ;
      RECT 14.355 5.695 14.525 6.545 ;
      RECT 14.355 5.695 14.53 6.045 ;
      RECT 14.355 5.695 15.33 5.87 ;
      RECT 15.155 1.965 15.33 5.87 ;
      RECT 15.1 1.965 15.45 2.315 ;
      RECT 15.125 6.655 15.45 6.98 ;
      RECT 14.01 6.745 15.45 6.915 ;
      RECT 14.01 2.395 14.17 6.915 ;
      RECT 14.325 2.365 14.645 2.685 ;
      RECT 14.01 2.395 14.645 2.565 ;
      RECT 12.75 2.685 13.04 3.065 ;
      RECT 12.72 2.7 13.06 3.05 ;
      RECT 11.455 3.54 11.715 3.86 ;
      RECT 11.515 1.83 11.655 3.86 ;
      RECT 11.345 2.39 11.655 2.76 ;
      RECT 11.415 1.95 11.655 2.76 ;
      RECT 11.445 1.83 11.725 2.2 ;
      RECT 11.445 1.94 11.73 2.14 ;
      RECT 10.765 2.42 11.025 2.74 ;
      RECT 10.105 2.51 11.025 2.65 ;
      RECT 10.105 1.57 10.245 2.65 ;
      RECT 6.565 1.86 6.825 2.18 ;
      RECT 6.745 1.57 6.885 2.09 ;
      RECT 6.745 1.57 10.245 1.71 ;
      RECT 1.54 6.995 1.83 7.345 ;
      RECT 1.54 7.05 2.795 7.22 ;
      RECT 2.625 6.685 2.795 7.22 ;
      RECT 9.685 6.605 10.035 6.955 ;
      RECT 2.625 6.685 10.035 6.855 ;
      RECT 9.595 3.26 9.855 3.58 ;
      RECT 9.655 1.85 9.795 3.58 ;
      RECT 9.585 1.85 9.865 2.22 ;
      RECT 6.985 4.01 9.425 4.15 ;
      RECT 9.285 2.7 9.425 4.15 ;
      RECT 6.985 3.63 7.125 4.15 ;
      RECT 6.685 3.63 7.125 3.86 ;
      RECT 4.345 3.63 7.125 3.77 ;
      RECT 6.685 3.54 6.945 3.86 ;
      RECT 4.345 3.35 4.485 3.77 ;
      RECT 3.835 3.26 4.095 3.58 ;
      RECT 3.835 3.35 4.485 3.49 ;
      RECT 3.895 1.86 4.035 3.58 ;
      RECT 9.225 2.7 9.485 3.02 ;
      RECT 3.835 1.86 4.095 2.18 ;
      RECT 8.845 3.54 9.105 3.86 ;
      RECT 8.905 1.95 9.045 3.86 ;
      RECT 8.565 1.95 9.045 2.22 ;
      RECT 8.365 1.85 8.845 2.2 ;
      RECT 8.355 3.49 8.635 3.86 ;
      RECT 8.425 2.39 8.565 3.86 ;
      RECT 8.365 2.39 8.625 3.02 ;
      RECT 8.355 2.39 8.635 2.76 ;
      RECT 7.285 3.54 7.545 3.86 ;
      RECT 7.285 3.35 7.485 3.86 ;
      RECT 7.095 3.35 7.485 3.49 ;
      RECT 7.095 1.86 7.235 3.49 ;
      RECT 7.095 1.86 7.405 2.23 ;
      RECT 7.035 1.86 7.405 2.18 ;
      RECT 4.755 2.95 5.035 3.32 ;
      RECT 6.205 2.98 6.465 3.3 ;
      RECT 4.585 3.07 6.465 3.21 ;
      RECT 4.585 2.95 5.035 3.21 ;
      RECT 4.525 2.39 4.785 3.02 ;
      RECT 4.515 2.39 4.795 2.76 ;
      RECT 5.595 2.39 6.005 2.76 ;
      RECT 5.005 2.42 5.265 2.74 ;
      RECT 5.005 2.51 6.005 2.65 ;
      RECT 4.515 1.83 4.795 2.2 ;
      RECT 4.515 1.86 4.905 2.18 ;
      RECT 0.195 8.5 0.575 8.88 ;
      RECT 0.235 0 0.4 8.88 ;
      RECT 0.19 0 0.57 0.38 ;
      RECT 70.055 7.055 70.425 7.425 ;
      RECT 68.915 2.39 69.195 2.86 ;
      RECT 68.675 1.86 68.955 2.2 ;
      RECT 67.475 2.39 67.755 2.76 ;
      RECT 64.92 1.215 65.29 1.22 ;
      RECT 54.795 7.055 55.165 7.425 ;
      RECT 53.655 2.39 53.935 2.86 ;
      RECT 53.415 1.86 53.695 2.2 ;
      RECT 52.215 2.39 52.495 2.76 ;
      RECT 49.66 1.215 50.03 1.22 ;
      RECT 39.535 7.055 39.905 7.425 ;
      RECT 38.395 2.39 38.675 2.86 ;
      RECT 38.155 1.86 38.435 2.2 ;
      RECT 36.955 2.39 37.235 2.76 ;
      RECT 34.4 1.215 34.77 1.22 ;
      RECT 24.275 7.055 24.645 7.425 ;
      RECT 23.135 2.39 23.415 2.86 ;
      RECT 22.895 1.86 23.175 2.2 ;
      RECT 21.695 2.39 21.975 2.76 ;
      RECT 19.14 1.215 19.51 1.22 ;
      RECT 9.015 7.055 9.385 7.425 ;
      RECT 7.875 2.39 8.155 2.86 ;
      RECT 7.635 1.86 7.915 2.2 ;
      RECT 6.435 2.39 6.715 2.76 ;
      RECT 3.88 1.215 4.25 1.22 ;
    LAYER via1 ;
      RECT 78.625 7.375 78.775 7.525 ;
      RECT 76.255 6.74 76.405 6.89 ;
      RECT 76.24 2.065 76.39 2.215 ;
      RECT 75.45 2.45 75.6 2.6 ;
      RECT 75.45 6.325 75.6 6.475 ;
      RECT 73.86 2.8 74.01 2.95 ;
      RECT 72.55 1.945 72.7 2.095 ;
      RECT 72.55 3.625 72.7 3.775 ;
      RECT 71.86 2.505 72.01 2.655 ;
      RECT 70.825 6.71 70.975 6.86 ;
      RECT 70.69 1.945 70.84 2.095 ;
      RECT 70.69 3.345 70.84 3.495 ;
      RECT 70.32 2.785 70.47 2.935 ;
      RECT 70.165 7.165 70.315 7.315 ;
      RECT 69.94 3.625 70.09 3.775 ;
      RECT 69.46 1.945 69.61 2.095 ;
      RECT 69.46 2.785 69.61 2.935 ;
      RECT 68.98 2.505 69.13 2.655 ;
      RECT 68.74 1.945 68.89 2.095 ;
      RECT 68.38 3.625 68.53 3.775 ;
      RECT 68.13 1.945 68.28 2.095 ;
      RECT 67.78 3.625 67.93 3.775 ;
      RECT 67.66 1.945 67.81 2.095 ;
      RECT 67.54 2.505 67.69 2.655 ;
      RECT 67.3 3.065 67.45 3.215 ;
      RECT 66.1 2.505 66.25 2.655 ;
      RECT 65.74 1.945 65.89 2.095 ;
      RECT 65.62 2.785 65.77 2.935 ;
      RECT 64.93 1.945 65.08 2.095 ;
      RECT 64.93 3.345 65.08 3.495 ;
      RECT 63.34 6.755 63.49 6.905 ;
      RECT 60.995 6.74 61.145 6.89 ;
      RECT 60.98 2.065 61.13 2.215 ;
      RECT 60.19 2.45 60.34 2.6 ;
      RECT 60.19 6.325 60.34 6.475 ;
      RECT 58.6 2.8 58.75 2.95 ;
      RECT 57.29 1.945 57.44 2.095 ;
      RECT 57.29 3.625 57.44 3.775 ;
      RECT 56.6 2.505 56.75 2.655 ;
      RECT 55.57 6.71 55.72 6.86 ;
      RECT 55.43 1.945 55.58 2.095 ;
      RECT 55.43 3.345 55.58 3.495 ;
      RECT 55.06 2.785 55.21 2.935 ;
      RECT 54.905 7.165 55.055 7.315 ;
      RECT 54.68 3.625 54.83 3.775 ;
      RECT 54.2 1.945 54.35 2.095 ;
      RECT 54.2 2.785 54.35 2.935 ;
      RECT 53.72 2.505 53.87 2.655 ;
      RECT 53.48 1.945 53.63 2.095 ;
      RECT 53.12 3.625 53.27 3.775 ;
      RECT 52.87 1.945 53.02 2.095 ;
      RECT 52.52 3.625 52.67 3.775 ;
      RECT 52.4 1.945 52.55 2.095 ;
      RECT 52.28 2.505 52.43 2.655 ;
      RECT 52.04 3.065 52.19 3.215 ;
      RECT 50.84 2.505 50.99 2.655 ;
      RECT 50.48 1.945 50.63 2.095 ;
      RECT 50.36 2.785 50.51 2.935 ;
      RECT 49.67 1.945 49.82 2.095 ;
      RECT 49.67 3.345 49.82 3.495 ;
      RECT 48.08 6.755 48.23 6.905 ;
      RECT 45.735 6.74 45.885 6.89 ;
      RECT 45.72 2.065 45.87 2.215 ;
      RECT 44.93 2.45 45.08 2.6 ;
      RECT 44.93 6.325 45.08 6.475 ;
      RECT 43.34 2.8 43.49 2.95 ;
      RECT 42.03 1.945 42.18 2.095 ;
      RECT 42.03 3.625 42.18 3.775 ;
      RECT 41.34 2.505 41.49 2.655 ;
      RECT 40.305 6.715 40.455 6.865 ;
      RECT 40.17 1.945 40.32 2.095 ;
      RECT 40.17 3.345 40.32 3.495 ;
      RECT 39.8 2.785 39.95 2.935 ;
      RECT 39.645 7.165 39.795 7.315 ;
      RECT 39.42 3.625 39.57 3.775 ;
      RECT 38.94 1.945 39.09 2.095 ;
      RECT 38.94 2.785 39.09 2.935 ;
      RECT 38.46 2.505 38.61 2.655 ;
      RECT 38.22 1.945 38.37 2.095 ;
      RECT 37.86 3.625 38.01 3.775 ;
      RECT 37.61 1.945 37.76 2.095 ;
      RECT 37.26 3.625 37.41 3.775 ;
      RECT 37.14 1.945 37.29 2.095 ;
      RECT 37.02 2.505 37.17 2.655 ;
      RECT 36.78 3.065 36.93 3.215 ;
      RECT 35.58 2.505 35.73 2.655 ;
      RECT 35.22 1.945 35.37 2.095 ;
      RECT 35.1 2.785 35.25 2.935 ;
      RECT 34.41 1.945 34.56 2.095 ;
      RECT 34.41 3.345 34.56 3.495 ;
      RECT 32.865 6.76 33.015 6.91 ;
      RECT 30.475 6.74 30.625 6.89 ;
      RECT 30.46 2.065 30.61 2.215 ;
      RECT 29.67 2.45 29.82 2.6 ;
      RECT 29.67 6.325 29.82 6.475 ;
      RECT 28.08 2.8 28.23 2.95 ;
      RECT 26.77 1.945 26.92 2.095 ;
      RECT 26.77 3.625 26.92 3.775 ;
      RECT 26.08 2.505 26.23 2.655 ;
      RECT 25.045 6.71 25.195 6.86 ;
      RECT 24.91 1.945 25.06 2.095 ;
      RECT 24.91 3.345 25.06 3.495 ;
      RECT 24.54 2.785 24.69 2.935 ;
      RECT 24.385 7.165 24.535 7.315 ;
      RECT 24.16 3.625 24.31 3.775 ;
      RECT 23.68 1.945 23.83 2.095 ;
      RECT 23.68 2.785 23.83 2.935 ;
      RECT 23.2 2.505 23.35 2.655 ;
      RECT 22.96 1.945 23.11 2.095 ;
      RECT 22.6 3.625 22.75 3.775 ;
      RECT 22.35 1.945 22.5 2.095 ;
      RECT 22 3.625 22.15 3.775 ;
      RECT 21.88 1.945 22.03 2.095 ;
      RECT 21.76 2.505 21.91 2.655 ;
      RECT 21.52 3.065 21.67 3.215 ;
      RECT 20.32 2.505 20.47 2.655 ;
      RECT 19.96 1.945 20.11 2.095 ;
      RECT 19.84 2.785 19.99 2.935 ;
      RECT 19.15 1.945 19.3 2.095 ;
      RECT 19.15 3.345 19.3 3.495 ;
      RECT 17.605 6.755 17.755 6.905 ;
      RECT 15.215 6.74 15.365 6.89 ;
      RECT 15.2 2.065 15.35 2.215 ;
      RECT 14.41 2.45 14.56 2.6 ;
      RECT 14.41 6.325 14.56 6.475 ;
      RECT 12.82 2.8 12.97 2.95 ;
      RECT 11.51 1.945 11.66 2.095 ;
      RECT 11.51 3.625 11.66 3.775 ;
      RECT 10.82 2.505 10.97 2.655 ;
      RECT 9.785 6.705 9.935 6.855 ;
      RECT 9.65 1.945 9.8 2.095 ;
      RECT 9.65 3.345 9.8 3.495 ;
      RECT 9.28 2.785 9.43 2.935 ;
      RECT 9.125 7.165 9.275 7.315 ;
      RECT 8.9 3.625 9.05 3.775 ;
      RECT 8.42 1.945 8.57 2.095 ;
      RECT 8.42 2.785 8.57 2.935 ;
      RECT 7.94 2.505 8.09 2.655 ;
      RECT 7.7 1.945 7.85 2.095 ;
      RECT 7.34 3.625 7.49 3.775 ;
      RECT 7.09 1.945 7.24 2.095 ;
      RECT 6.74 3.625 6.89 3.775 ;
      RECT 6.62 1.945 6.77 2.095 ;
      RECT 6.5 2.505 6.65 2.655 ;
      RECT 6.26 3.065 6.41 3.215 ;
      RECT 5.06 2.505 5.21 2.655 ;
      RECT 4.7 1.945 4.85 2.095 ;
      RECT 4.58 2.785 4.73 2.935 ;
      RECT 3.89 1.945 4.04 2.095 ;
      RECT 3.89 3.345 4.04 3.495 ;
      RECT 1.61 7.095 1.76 7.245 ;
      RECT 1.235 6.355 1.385 6.505 ;
      RECT 0.31 8.615 0.46 8.765 ;
      RECT 0.305 0.115 0.455 0.265 ;
    LAYER met1 ;
      RECT 65.075 2.74 65.365 2.97 ;
      RECT 49.815 2.74 50.105 2.97 ;
      RECT 34.555 2.74 34.845 2.97 ;
      RECT 19.295 2.74 19.585 2.97 ;
      RECT 4.035 2.74 4.325 2.97 ;
      RECT 65.145 2.37 65.285 2.97 ;
      RECT 49.885 2.37 50.025 2.97 ;
      RECT 34.625 2.37 34.765 2.97 ;
      RECT 19.365 2.37 19.505 2.97 ;
      RECT 4.105 2.37 4.245 2.97 ;
      RECT 65.145 2.37 65.765 2.51 ;
      RECT 65.625 0 65.765 2.51 ;
      RECT 49.885 2.37 50.505 2.51 ;
      RECT 50.365 0 50.505 2.51 ;
      RECT 34.625 2.37 35.245 2.51 ;
      RECT 35.105 0 35.245 2.51 ;
      RECT 19.365 2.37 19.985 2.51 ;
      RECT 19.845 0 19.985 2.51 ;
      RECT 4.105 2.37 4.725 2.51 ;
      RECT 4.585 0 4.725 2.51 ;
      RECT 65.385 1.95 65.765 2.21 ;
      RECT 50.125 1.95 50.505 2.21 ;
      RECT 34.865 1.95 35.245 2.21 ;
      RECT 19.605 1.95 19.985 2.21 ;
      RECT 4.345 1.95 4.725 2.21 ;
      RECT 65.57 1.89 65.975 2.15 ;
      RECT 50.31 1.89 50.715 2.15 ;
      RECT 35.05 1.89 35.455 2.15 ;
      RECT 19.79 1.89 20.195 2.15 ;
      RECT 4.53 1.89 4.935 2.15 ;
      RECT 66.275 1.9 66.565 2.13 ;
      RECT 51.015 1.9 51.305 2.13 ;
      RECT 35.755 1.9 36.045 2.13 ;
      RECT 20.495 1.9 20.785 2.13 ;
      RECT 5.235 1.9 5.525 2.13 ;
      RECT 65.385 1.95 66.565 2.09 ;
      RECT 50.125 1.95 51.305 2.09 ;
      RECT 34.865 1.95 36.045 2.09 ;
      RECT 19.605 1.95 20.785 2.09 ;
      RECT 4.345 1.95 5.525 2.09 ;
      RECT 65.57 0 65.86 2.15 ;
      RECT 50.31 0 50.6 2.15 ;
      RECT 35.05 0 35.34 2.15 ;
      RECT 19.79 0 20.08 2.15 ;
      RECT 4.53 0 4.82 2.15 ;
      RECT 64.585 0 73.325 1.74 ;
      RECT 49.325 0 58.065 1.74 ;
      RECT 34.065 0 42.805 1.74 ;
      RECT 18.805 0 27.545 1.74 ;
      RECT 3.545 0 12.285 1.74 ;
      RECT 0.205 0 0.555 0.335 ;
      RECT 0 0 0.805 0.315 ;
      RECT 78.915 0 79.095 0.305 ;
      RECT 63.655 0 76.965 0.305 ;
      RECT 48.395 0 61.705 0.305 ;
      RECT 33.135 0 46.445 0.305 ;
      RECT 17.875 0 31.185 0.305 ;
      RECT 0 0 15.925 0.305 ;
      RECT 0 0 79.095 0.3 ;
      RECT 0 8.58 79.095 8.88 ;
      RECT 78.915 8.575 79.095 8.88 ;
      RECT 63.655 8.575 76.965 8.88 ;
      RECT 48.395 8.575 61.705 8.88 ;
      RECT 33.135 8.575 46.445 8.88 ;
      RECT 17.875 8.575 31.185 8.88 ;
      RECT 0 8.575 15.925 8.88 ;
      RECT 69.555 6.315 69.725 8.88 ;
      RECT 54.295 6.315 54.465 8.88 ;
      RECT 39.035 6.315 39.205 8.88 ;
      RECT 23.775 6.315 23.945 8.88 ;
      RECT 8.515 6.315 8.685 8.88 ;
      RECT 0.005 8.565 0.81 8.88 ;
      RECT 0.21 8.545 0.56 8.88 ;
      RECT 69.72 6.285 70.01 6.515 ;
      RECT 54.46 6.285 54.75 6.515 ;
      RECT 39.2 6.285 39.49 6.515 ;
      RECT 23.94 6.285 24.23 6.515 ;
      RECT 8.68 6.285 8.97 6.515 ;
      RECT 69.55 6.315 70.01 6.485 ;
      RECT 54.29 6.315 54.75 6.485 ;
      RECT 39.03 6.315 39.49 6.485 ;
      RECT 23.77 6.315 24.23 6.485 ;
      RECT 8.51 6.315 8.97 6.485 ;
      RECT 78.49 7.77 78.78 8 ;
      RECT 78.55 6.29 78.72 8 ;
      RECT 78.525 7.275 78.875 7.625 ;
      RECT 78.49 6.29 78.78 6.52 ;
      RECT 78.085 2.395 78.19 2.965 ;
      RECT 78.085 2.73 78.41 2.96 ;
      RECT 78.085 2.76 78.58 2.93 ;
      RECT 78.085 2.395 78.275 2.96 ;
      RECT 77.5 2.36 77.79 2.59 ;
      RECT 77.5 2.395 78.275 2.565 ;
      RECT 77.56 0.88 77.73 2.59 ;
      RECT 77.5 0.88 77.79 1.11 ;
      RECT 77.5 7.77 77.79 8 ;
      RECT 77.56 6.29 77.73 8 ;
      RECT 77.5 6.29 77.79 6.52 ;
      RECT 77.5 6.325 78.355 6.485 ;
      RECT 78.185 5.92 78.355 6.485 ;
      RECT 77.5 6.32 77.895 6.485 ;
      RECT 78.12 5.92 78.41 6.15 ;
      RECT 78.12 5.95 78.58 6.12 ;
      RECT 77.13 2.73 77.42 2.96 ;
      RECT 77.13 2.76 77.59 2.93 ;
      RECT 77.195 1.655 77.36 2.96 ;
      RECT 75.71 1.625 76 1.855 ;
      RECT 75.71 1.655 77.36 1.825 ;
      RECT 75.77 0.885 75.94 1.855 ;
      RECT 75.71 0.885 76 1.115 ;
      RECT 75.71 7.765 76 7.995 ;
      RECT 75.77 7.025 75.94 7.995 ;
      RECT 75.77 7.12 77.36 7.29 ;
      RECT 77.19 5.92 77.36 7.29 ;
      RECT 75.71 7.025 76 7.255 ;
      RECT 77.13 5.92 77.42 6.15 ;
      RECT 77.13 5.95 77.59 6.12 ;
      RECT 73.76 2.7 74.1 3.05 ;
      RECT 73.85 2.025 74.02 3.05 ;
      RECT 76.14 1.965 76.49 2.315 ;
      RECT 73.85 2.025 76.49 2.195 ;
      RECT 76.165 6.655 76.49 6.98 ;
      RECT 70.725 6.61 71.075 6.96 ;
      RECT 76.14 6.655 76.49 6.885 ;
      RECT 70.525 6.655 71.075 6.885 ;
      RECT 70.355 6.685 76.49 6.855 ;
      RECT 75.365 2.365 75.685 2.685 ;
      RECT 75.335 2.365 75.685 2.595 ;
      RECT 75.165 2.395 75.685 2.565 ;
      RECT 75.365 6.255 75.685 6.545 ;
      RECT 75.335 6.285 75.685 6.515 ;
      RECT 75.165 6.315 75.685 6.485 ;
      RECT 72.465 1.89 72.785 2.15 ;
      RECT 72.035 1.9 72.325 2.13 ;
      RECT 72.035 1.95 72.785 2.09 ;
      RECT 72.465 3.57 72.785 3.83 ;
      RECT 72.035 3.58 72.325 3.81 ;
      RECT 72.035 3.63 72.785 3.77 ;
      RECT 71.795 3.02 72.085 3.25 ;
      RECT 71.795 3.07 72.365 3.21 ;
      RECT 72.225 2.93 72.485 3.07 ;
      RECT 72.275 2.74 72.565 2.97 ;
      RECT 70.425 2.93 71.525 3.07 ;
      RECT 70.235 2.73 70.555 2.99 ;
      RECT 71.315 2.74 71.605 2.97 ;
      RECT 70.235 2.74 70.645 2.99 ;
      RECT 70.605 1.89 70.925 2.15 ;
      RECT 71.075 1.9 71.365 2.13 ;
      RECT 70.605 1.95 71.365 2.09 ;
      RECT 67.905 3.15 70.085 3.29 ;
      RECT 69.945 2.16 70.085 3.29 ;
      RECT 67.905 3.07 69.205 3.29 ;
      RECT 68.915 3.02 69.205 3.29 ;
      RECT 67.905 2.79 68.245 3.29 ;
      RECT 67.955 2.74 68.245 3.29 ;
      RECT 70.835 2.46 71.125 2.69 ;
      RECT 69.945 2.37 71.045 2.51 ;
      RECT 69.875 2.16 70.165 2.41 ;
      RECT 70.095 7.765 70.385 7.995 ;
      RECT 70.155 7.025 70.325 7.995 ;
      RECT 70.055 7.055 70.425 7.425 ;
      RECT 70.095 7.025 70.385 7.425 ;
      RECT 69.855 3.57 70.175 3.83 ;
      RECT 69.855 3.58 70.375 3.81 ;
      RECT 68.435 2.46 68.725 2.69 ;
      RECT 68.585 2.07 68.725 2.69 ;
      RECT 68.585 2.07 68.885 2.21 ;
      RECT 69.375 1.89 69.695 2.15 ;
      RECT 68.655 1.89 68.975 2.15 ;
      RECT 69.155 1.9 69.695 2.13 ;
      RECT 68.655 1.95 69.695 2.09 ;
      RECT 68.295 3.57 68.615 3.83 ;
      RECT 68.195 3.58 68.615 3.81 ;
      RECT 66.275 3.02 66.565 3.25 ;
      RECT 66.275 3.02 66.725 3.21 ;
      RECT 66.585 2.55 66.725 3.21 ;
      RECT 66.705 1.95 66.845 2.69 ;
      RECT 67.575 1.89 67.895 2.15 ;
      RECT 66.755 1.9 67.045 2.13 ;
      RECT 66.705 1.95 67.895 2.09 ;
      RECT 67.455 2.45 67.775 2.71 ;
      RECT 66.995 2.46 67.285 2.69 ;
      RECT 66.995 2.51 67.775 2.65 ;
      RECT 67.215 3.01 67.535 3.27 ;
      RECT 67.215 3.02 67.765 3.25 ;
      RECT 66.755 3.58 67.045 3.81 ;
      RECT 65.865 3.46 66.965 3.6 ;
      RECT 65.795 3.3 66.085 3.53 ;
      RECT 63.23 7.77 63.52 8 ;
      RECT 63.29 6.29 63.46 8 ;
      RECT 63.24 6.655 63.59 7.005 ;
      RECT 63.23 6.29 63.52 6.52 ;
      RECT 62.825 2.395 62.93 2.965 ;
      RECT 62.825 2.73 63.15 2.96 ;
      RECT 62.825 2.76 63.32 2.93 ;
      RECT 62.825 2.395 63.015 2.96 ;
      RECT 62.24 2.36 62.53 2.59 ;
      RECT 62.24 2.395 63.015 2.565 ;
      RECT 62.3 0.88 62.47 2.59 ;
      RECT 62.24 0.88 62.53 1.11 ;
      RECT 62.24 7.77 62.53 8 ;
      RECT 62.3 6.29 62.47 8 ;
      RECT 62.24 6.29 62.53 6.52 ;
      RECT 62.24 6.325 63.095 6.485 ;
      RECT 62.925 5.92 63.095 6.485 ;
      RECT 62.24 6.32 62.635 6.485 ;
      RECT 62.86 5.92 63.15 6.15 ;
      RECT 62.86 5.95 63.32 6.12 ;
      RECT 61.87 2.73 62.16 2.96 ;
      RECT 61.87 2.76 62.33 2.93 ;
      RECT 61.935 1.655 62.1 2.96 ;
      RECT 60.45 1.625 60.74 1.855 ;
      RECT 60.45 1.655 62.1 1.825 ;
      RECT 60.51 0.885 60.68 1.855 ;
      RECT 60.45 0.885 60.74 1.115 ;
      RECT 60.45 7.765 60.74 7.995 ;
      RECT 60.51 7.025 60.68 7.995 ;
      RECT 60.51 7.12 62.1 7.29 ;
      RECT 61.93 5.92 62.1 7.29 ;
      RECT 60.45 7.025 60.74 7.255 ;
      RECT 61.87 5.92 62.16 6.15 ;
      RECT 61.87 5.95 62.33 6.12 ;
      RECT 58.5 2.7 58.84 3.05 ;
      RECT 58.59 2.025 58.76 3.05 ;
      RECT 60.88 1.965 61.23 2.315 ;
      RECT 58.59 2.025 61.23 2.195 ;
      RECT 60.905 6.655 61.23 6.98 ;
      RECT 55.47 6.61 55.82 6.96 ;
      RECT 60.88 6.655 61.23 6.885 ;
      RECT 55.265 6.655 55.82 6.885 ;
      RECT 55.095 6.685 61.23 6.855 ;
      RECT 60.105 2.365 60.425 2.685 ;
      RECT 60.075 2.365 60.425 2.595 ;
      RECT 59.905 2.395 60.425 2.565 ;
      RECT 60.105 6.255 60.425 6.545 ;
      RECT 60.075 6.285 60.425 6.515 ;
      RECT 59.905 6.315 60.425 6.485 ;
      RECT 57.205 1.89 57.525 2.15 ;
      RECT 56.775 1.9 57.065 2.13 ;
      RECT 56.775 1.95 57.525 2.09 ;
      RECT 57.205 3.57 57.525 3.83 ;
      RECT 56.775 3.58 57.065 3.81 ;
      RECT 56.775 3.63 57.525 3.77 ;
      RECT 56.535 3.02 56.825 3.25 ;
      RECT 56.535 3.07 57.105 3.21 ;
      RECT 56.965 2.93 57.225 3.07 ;
      RECT 57.015 2.74 57.305 2.97 ;
      RECT 55.165 2.93 56.265 3.07 ;
      RECT 54.975 2.73 55.295 2.99 ;
      RECT 56.055 2.74 56.345 2.97 ;
      RECT 54.975 2.74 55.385 2.99 ;
      RECT 55.345 1.89 55.665 2.15 ;
      RECT 55.815 1.9 56.105 2.13 ;
      RECT 55.345 1.95 56.105 2.09 ;
      RECT 52.645 3.15 54.825 3.29 ;
      RECT 54.685 2.16 54.825 3.29 ;
      RECT 52.645 3.07 53.945 3.29 ;
      RECT 53.655 3.02 53.945 3.29 ;
      RECT 52.645 2.79 52.985 3.29 ;
      RECT 52.695 2.74 52.985 3.29 ;
      RECT 55.575 2.46 55.865 2.69 ;
      RECT 54.685 2.37 55.785 2.51 ;
      RECT 54.615 2.16 54.905 2.41 ;
      RECT 54.835 7.765 55.125 7.995 ;
      RECT 54.895 7.025 55.065 7.995 ;
      RECT 54.795 7.055 55.165 7.425 ;
      RECT 54.835 7.025 55.125 7.425 ;
      RECT 54.595 3.57 54.915 3.83 ;
      RECT 54.595 3.58 55.115 3.81 ;
      RECT 53.175 2.46 53.465 2.69 ;
      RECT 53.325 2.07 53.465 2.69 ;
      RECT 53.325 2.07 53.625 2.21 ;
      RECT 54.115 1.89 54.435 2.15 ;
      RECT 53.395 1.89 53.715 2.15 ;
      RECT 53.895 1.9 54.435 2.13 ;
      RECT 53.395 1.95 54.435 2.09 ;
      RECT 53.035 3.57 53.355 3.83 ;
      RECT 52.935 3.58 53.355 3.81 ;
      RECT 51.015 3.02 51.305 3.25 ;
      RECT 51.015 3.02 51.465 3.21 ;
      RECT 51.325 2.55 51.465 3.21 ;
      RECT 51.445 1.95 51.585 2.69 ;
      RECT 52.315 1.89 52.635 2.15 ;
      RECT 51.495 1.9 51.785 2.13 ;
      RECT 51.445 1.95 52.635 2.09 ;
      RECT 52.195 2.45 52.515 2.71 ;
      RECT 51.735 2.46 52.025 2.69 ;
      RECT 51.735 2.51 52.515 2.65 ;
      RECT 51.955 3.01 52.275 3.27 ;
      RECT 51.955 3.02 52.505 3.25 ;
      RECT 51.495 3.58 51.785 3.81 ;
      RECT 50.605 3.46 51.705 3.6 ;
      RECT 50.535 3.3 50.825 3.53 ;
      RECT 47.97 7.77 48.26 8 ;
      RECT 48.03 6.29 48.2 8 ;
      RECT 47.98 6.655 48.33 7.005 ;
      RECT 47.97 6.29 48.26 6.52 ;
      RECT 47.565 2.395 47.67 2.965 ;
      RECT 47.565 2.73 47.89 2.96 ;
      RECT 47.565 2.76 48.06 2.93 ;
      RECT 47.565 2.395 47.755 2.96 ;
      RECT 46.98 2.36 47.27 2.59 ;
      RECT 46.98 2.395 47.755 2.565 ;
      RECT 47.04 0.88 47.21 2.59 ;
      RECT 46.98 0.88 47.27 1.11 ;
      RECT 46.98 7.77 47.27 8 ;
      RECT 47.04 6.29 47.21 8 ;
      RECT 46.98 6.29 47.27 6.52 ;
      RECT 46.98 6.325 47.835 6.485 ;
      RECT 47.665 5.92 47.835 6.485 ;
      RECT 46.98 6.32 47.375 6.485 ;
      RECT 47.6 5.92 47.89 6.15 ;
      RECT 47.6 5.95 48.06 6.12 ;
      RECT 46.61 2.73 46.9 2.96 ;
      RECT 46.61 2.76 47.07 2.93 ;
      RECT 46.675 1.655 46.84 2.96 ;
      RECT 45.19 1.625 45.48 1.855 ;
      RECT 45.19 1.655 46.84 1.825 ;
      RECT 45.25 0.885 45.42 1.855 ;
      RECT 45.19 0.885 45.48 1.115 ;
      RECT 45.19 7.765 45.48 7.995 ;
      RECT 45.25 7.025 45.42 7.995 ;
      RECT 45.25 7.12 46.84 7.29 ;
      RECT 46.67 5.92 46.84 7.29 ;
      RECT 45.19 7.025 45.48 7.255 ;
      RECT 46.61 5.92 46.9 6.15 ;
      RECT 46.61 5.95 47.07 6.12 ;
      RECT 43.24 2.7 43.58 3.05 ;
      RECT 43.33 2.025 43.5 3.05 ;
      RECT 45.62 1.965 45.97 2.315 ;
      RECT 43.33 2.025 45.97 2.195 ;
      RECT 45.645 6.655 45.97 6.98 ;
      RECT 40.205 6.615 40.555 6.965 ;
      RECT 45.62 6.655 45.97 6.885 ;
      RECT 40.005 6.655 40.555 6.885 ;
      RECT 39.835 6.685 45.97 6.855 ;
      RECT 44.845 2.365 45.165 2.685 ;
      RECT 44.815 2.365 45.165 2.595 ;
      RECT 44.645 2.395 45.165 2.565 ;
      RECT 44.845 6.255 45.165 6.545 ;
      RECT 44.815 6.285 45.165 6.515 ;
      RECT 44.645 6.315 45.165 6.485 ;
      RECT 41.945 1.89 42.265 2.15 ;
      RECT 41.515 1.9 41.805 2.13 ;
      RECT 41.515 1.95 42.265 2.09 ;
      RECT 41.945 3.57 42.265 3.83 ;
      RECT 41.515 3.58 41.805 3.81 ;
      RECT 41.515 3.63 42.265 3.77 ;
      RECT 41.275 3.02 41.565 3.25 ;
      RECT 41.275 3.07 41.845 3.21 ;
      RECT 41.705 2.93 41.965 3.07 ;
      RECT 41.755 2.74 42.045 2.97 ;
      RECT 39.905 2.93 41.005 3.07 ;
      RECT 39.715 2.73 40.035 2.99 ;
      RECT 40.795 2.74 41.085 2.97 ;
      RECT 39.715 2.74 40.125 2.99 ;
      RECT 40.085 1.89 40.405 2.15 ;
      RECT 40.555 1.9 40.845 2.13 ;
      RECT 40.085 1.95 40.845 2.09 ;
      RECT 37.385 3.15 39.565 3.29 ;
      RECT 39.425 2.16 39.565 3.29 ;
      RECT 37.385 3.07 38.685 3.29 ;
      RECT 38.395 3.02 38.685 3.29 ;
      RECT 37.385 2.79 37.725 3.29 ;
      RECT 37.435 2.74 37.725 3.29 ;
      RECT 40.315 2.46 40.605 2.69 ;
      RECT 39.425 2.37 40.525 2.51 ;
      RECT 39.355 2.16 39.645 2.41 ;
      RECT 39.575 7.765 39.865 7.995 ;
      RECT 39.635 7.025 39.805 7.995 ;
      RECT 39.535 7.055 39.905 7.425 ;
      RECT 39.575 7.025 39.865 7.425 ;
      RECT 39.335 3.57 39.655 3.83 ;
      RECT 39.335 3.58 39.855 3.81 ;
      RECT 37.915 2.46 38.205 2.69 ;
      RECT 38.065 2.07 38.205 2.69 ;
      RECT 38.065 2.07 38.365 2.21 ;
      RECT 38.855 1.89 39.175 2.15 ;
      RECT 38.135 1.89 38.455 2.15 ;
      RECT 38.635 1.9 39.175 2.13 ;
      RECT 38.135 1.95 39.175 2.09 ;
      RECT 37.775 3.57 38.095 3.83 ;
      RECT 37.675 3.58 38.095 3.81 ;
      RECT 35.755 3.02 36.045 3.25 ;
      RECT 35.755 3.02 36.205 3.21 ;
      RECT 36.065 2.55 36.205 3.21 ;
      RECT 36.185 1.95 36.325 2.69 ;
      RECT 37.055 1.89 37.375 2.15 ;
      RECT 36.235 1.9 36.525 2.13 ;
      RECT 36.185 1.95 37.375 2.09 ;
      RECT 36.935 2.45 37.255 2.71 ;
      RECT 36.475 2.46 36.765 2.69 ;
      RECT 36.475 2.51 37.255 2.65 ;
      RECT 36.695 3.01 37.015 3.27 ;
      RECT 36.695 3.02 37.245 3.25 ;
      RECT 36.235 3.58 36.525 3.81 ;
      RECT 35.345 3.46 36.445 3.6 ;
      RECT 35.275 3.3 35.565 3.53 ;
      RECT 32.71 7.77 33 8 ;
      RECT 32.77 6.29 32.94 8 ;
      RECT 32.76 6.66 33.115 7.015 ;
      RECT 32.71 6.29 33 6.52 ;
      RECT 32.305 2.395 32.41 2.965 ;
      RECT 32.305 2.73 32.63 2.96 ;
      RECT 32.305 2.76 32.8 2.93 ;
      RECT 32.305 2.395 32.495 2.96 ;
      RECT 31.72 2.36 32.01 2.59 ;
      RECT 31.72 2.395 32.495 2.565 ;
      RECT 31.78 0.88 31.95 2.59 ;
      RECT 31.72 0.88 32.01 1.11 ;
      RECT 31.72 7.77 32.01 8 ;
      RECT 31.78 6.29 31.95 8 ;
      RECT 31.72 6.29 32.01 6.52 ;
      RECT 31.72 6.325 32.575 6.485 ;
      RECT 32.405 5.92 32.575 6.485 ;
      RECT 31.72 6.32 32.115 6.485 ;
      RECT 32.34 5.92 32.63 6.15 ;
      RECT 32.34 5.95 32.8 6.12 ;
      RECT 31.35 2.73 31.64 2.96 ;
      RECT 31.35 2.76 31.81 2.93 ;
      RECT 31.415 1.655 31.58 2.96 ;
      RECT 29.93 1.625 30.22 1.855 ;
      RECT 29.93 1.655 31.58 1.825 ;
      RECT 29.99 0.885 30.16 1.855 ;
      RECT 29.93 0.885 30.22 1.115 ;
      RECT 29.93 7.765 30.22 7.995 ;
      RECT 29.99 7.025 30.16 7.995 ;
      RECT 29.99 7.12 31.58 7.29 ;
      RECT 31.41 5.92 31.58 7.29 ;
      RECT 29.93 7.025 30.22 7.255 ;
      RECT 31.35 5.92 31.64 6.15 ;
      RECT 31.35 5.95 31.81 6.12 ;
      RECT 27.98 2.7 28.32 3.05 ;
      RECT 28.07 2.025 28.24 3.05 ;
      RECT 30.36 1.965 30.71 2.315 ;
      RECT 28.07 2.025 30.71 2.195 ;
      RECT 30.385 6.655 30.71 6.98 ;
      RECT 24.945 6.61 25.295 6.96 ;
      RECT 30.36 6.655 30.71 6.885 ;
      RECT 24.745 6.655 25.295 6.885 ;
      RECT 24.575 6.685 30.71 6.855 ;
      RECT 29.585 2.365 29.905 2.685 ;
      RECT 29.555 2.365 29.905 2.595 ;
      RECT 29.385 2.395 29.905 2.565 ;
      RECT 29.585 6.255 29.905 6.545 ;
      RECT 29.555 6.285 29.905 6.515 ;
      RECT 29.385 6.315 29.905 6.485 ;
      RECT 26.685 1.89 27.005 2.15 ;
      RECT 26.255 1.9 26.545 2.13 ;
      RECT 26.255 1.95 27.005 2.09 ;
      RECT 26.685 3.57 27.005 3.83 ;
      RECT 26.255 3.58 26.545 3.81 ;
      RECT 26.255 3.63 27.005 3.77 ;
      RECT 26.015 3.02 26.305 3.25 ;
      RECT 26.015 3.07 26.585 3.21 ;
      RECT 26.445 2.93 26.705 3.07 ;
      RECT 26.495 2.74 26.785 2.97 ;
      RECT 24.645 2.93 25.745 3.07 ;
      RECT 24.455 2.73 24.775 2.99 ;
      RECT 25.535 2.74 25.825 2.97 ;
      RECT 24.455 2.74 24.865 2.99 ;
      RECT 24.825 1.89 25.145 2.15 ;
      RECT 25.295 1.9 25.585 2.13 ;
      RECT 24.825 1.95 25.585 2.09 ;
      RECT 22.125 3.15 24.305 3.29 ;
      RECT 24.165 2.16 24.305 3.29 ;
      RECT 22.125 3.07 23.425 3.29 ;
      RECT 23.135 3.02 23.425 3.29 ;
      RECT 22.125 2.79 22.465 3.29 ;
      RECT 22.175 2.74 22.465 3.29 ;
      RECT 25.055 2.46 25.345 2.69 ;
      RECT 24.165 2.37 25.265 2.51 ;
      RECT 24.095 2.16 24.385 2.41 ;
      RECT 24.315 7.765 24.605 7.995 ;
      RECT 24.375 7.025 24.545 7.995 ;
      RECT 24.275 7.055 24.645 7.425 ;
      RECT 24.315 7.025 24.605 7.425 ;
      RECT 24.075 3.57 24.395 3.83 ;
      RECT 24.075 3.58 24.595 3.81 ;
      RECT 22.655 2.46 22.945 2.69 ;
      RECT 22.805 2.07 22.945 2.69 ;
      RECT 22.805 2.07 23.105 2.21 ;
      RECT 23.595 1.89 23.915 2.15 ;
      RECT 22.875 1.89 23.195 2.15 ;
      RECT 23.375 1.9 23.915 2.13 ;
      RECT 22.875 1.95 23.915 2.09 ;
      RECT 22.515 3.57 22.835 3.83 ;
      RECT 22.415 3.58 22.835 3.81 ;
      RECT 20.495 3.02 20.785 3.25 ;
      RECT 20.495 3.02 20.945 3.21 ;
      RECT 20.805 2.55 20.945 3.21 ;
      RECT 20.925 1.95 21.065 2.69 ;
      RECT 21.795 1.89 22.115 2.15 ;
      RECT 20.975 1.9 21.265 2.13 ;
      RECT 20.925 1.95 22.115 2.09 ;
      RECT 21.675 2.45 21.995 2.71 ;
      RECT 21.215 2.46 21.505 2.69 ;
      RECT 21.215 2.51 21.995 2.65 ;
      RECT 21.435 3.01 21.755 3.27 ;
      RECT 21.435 3.02 21.985 3.25 ;
      RECT 20.975 3.58 21.265 3.81 ;
      RECT 20.085 3.46 21.185 3.6 ;
      RECT 20.015 3.3 20.305 3.53 ;
      RECT 17.45 7.77 17.74 8 ;
      RECT 17.51 6.29 17.68 8 ;
      RECT 17.505 6.655 17.855 7.005 ;
      RECT 17.45 6.29 17.74 6.52 ;
      RECT 17.045 2.395 17.15 2.965 ;
      RECT 17.045 2.73 17.37 2.96 ;
      RECT 17.045 2.76 17.54 2.93 ;
      RECT 17.045 2.395 17.235 2.96 ;
      RECT 16.46 2.36 16.75 2.59 ;
      RECT 16.46 2.395 17.235 2.565 ;
      RECT 16.52 0.88 16.69 2.59 ;
      RECT 16.46 0.88 16.75 1.11 ;
      RECT 16.46 7.77 16.75 8 ;
      RECT 16.52 6.29 16.69 8 ;
      RECT 16.46 6.29 16.75 6.52 ;
      RECT 16.46 6.325 17.315 6.485 ;
      RECT 17.145 5.92 17.315 6.485 ;
      RECT 16.46 6.32 16.855 6.485 ;
      RECT 17.08 5.92 17.37 6.15 ;
      RECT 17.08 5.95 17.54 6.12 ;
      RECT 16.09 2.73 16.38 2.96 ;
      RECT 16.09 2.76 16.55 2.93 ;
      RECT 16.155 1.655 16.32 2.96 ;
      RECT 14.67 1.625 14.96 1.855 ;
      RECT 14.67 1.655 16.32 1.825 ;
      RECT 14.73 0.885 14.9 1.855 ;
      RECT 14.67 0.885 14.96 1.115 ;
      RECT 14.67 7.765 14.96 7.995 ;
      RECT 14.73 7.025 14.9 7.995 ;
      RECT 14.73 7.12 16.32 7.29 ;
      RECT 16.15 5.92 16.32 7.29 ;
      RECT 14.67 7.025 14.96 7.255 ;
      RECT 16.09 5.92 16.38 6.15 ;
      RECT 16.09 5.95 16.55 6.12 ;
      RECT 12.72 2.7 13.06 3.05 ;
      RECT 12.81 2.025 12.98 3.05 ;
      RECT 15.1 1.965 15.45 2.315 ;
      RECT 12.81 2.025 15.45 2.195 ;
      RECT 15.125 6.655 15.45 6.98 ;
      RECT 9.685 6.605 10.035 6.955 ;
      RECT 15.1 6.655 15.45 6.885 ;
      RECT 9.485 6.655 10.035 6.885 ;
      RECT 9.315 6.685 15.45 6.855 ;
      RECT 14.325 2.365 14.645 2.685 ;
      RECT 14.295 2.365 14.645 2.595 ;
      RECT 14.125 2.395 14.645 2.565 ;
      RECT 14.325 6.255 14.645 6.545 ;
      RECT 14.295 6.285 14.645 6.515 ;
      RECT 14.125 6.315 14.645 6.485 ;
      RECT 11.425 1.89 11.745 2.15 ;
      RECT 10.995 1.9 11.285 2.13 ;
      RECT 10.995 1.95 11.745 2.09 ;
      RECT 11.425 3.57 11.745 3.83 ;
      RECT 10.995 3.58 11.285 3.81 ;
      RECT 10.995 3.63 11.745 3.77 ;
      RECT 10.755 3.02 11.045 3.25 ;
      RECT 10.755 3.07 11.325 3.21 ;
      RECT 11.185 2.93 11.445 3.07 ;
      RECT 11.235 2.74 11.525 2.97 ;
      RECT 9.385 2.93 10.485 3.07 ;
      RECT 9.195 2.73 9.515 2.99 ;
      RECT 10.275 2.74 10.565 2.97 ;
      RECT 9.195 2.74 9.605 2.99 ;
      RECT 9.565 1.89 9.885 2.15 ;
      RECT 10.035 1.9 10.325 2.13 ;
      RECT 9.565 1.95 10.325 2.09 ;
      RECT 6.865 3.15 9.045 3.29 ;
      RECT 8.905 2.16 9.045 3.29 ;
      RECT 6.865 3.07 8.165 3.29 ;
      RECT 7.875 3.02 8.165 3.29 ;
      RECT 6.865 2.79 7.205 3.29 ;
      RECT 6.915 2.74 7.205 3.29 ;
      RECT 9.795 2.46 10.085 2.69 ;
      RECT 8.905 2.37 10.005 2.51 ;
      RECT 8.835 2.16 9.125 2.41 ;
      RECT 9.055 7.765 9.345 7.995 ;
      RECT 9.115 7.025 9.285 7.995 ;
      RECT 9.015 7.055 9.385 7.425 ;
      RECT 9.055 7.025 9.345 7.425 ;
      RECT 8.815 3.57 9.135 3.83 ;
      RECT 8.815 3.58 9.335 3.81 ;
      RECT 7.395 2.46 7.685 2.69 ;
      RECT 7.545 2.07 7.685 2.69 ;
      RECT 7.545 2.07 7.845 2.21 ;
      RECT 8.335 1.89 8.655 2.15 ;
      RECT 7.615 1.89 7.935 2.15 ;
      RECT 8.115 1.9 8.655 2.13 ;
      RECT 7.615 1.95 8.655 2.09 ;
      RECT 7.255 3.57 7.575 3.83 ;
      RECT 7.155 3.58 7.575 3.81 ;
      RECT 5.235 3.02 5.525 3.25 ;
      RECT 5.235 3.02 5.685 3.21 ;
      RECT 5.545 2.55 5.685 3.21 ;
      RECT 5.665 1.95 5.805 2.69 ;
      RECT 6.535 1.89 6.855 2.15 ;
      RECT 5.715 1.9 6.005 2.13 ;
      RECT 5.665 1.95 6.855 2.09 ;
      RECT 6.415 2.45 6.735 2.71 ;
      RECT 5.955 2.46 6.245 2.69 ;
      RECT 5.955 2.51 6.735 2.65 ;
      RECT 6.175 3.01 6.495 3.27 ;
      RECT 6.175 3.02 6.725 3.25 ;
      RECT 5.715 3.58 6.005 3.81 ;
      RECT 4.825 3.46 5.925 3.6 ;
      RECT 4.755 3.3 5.045 3.53 ;
      RECT 1.54 7.765 1.83 7.995 ;
      RECT 1.6 7.025 1.77 7.995 ;
      RECT 1.51 7.025 1.86 7.315 ;
      RECT 1.135 6.285 1.485 6.575 ;
      RECT 0.995 6.315 1.485 6.485 ;
      RECT 71.775 2.45 72.095 2.71 ;
      RECT 70.605 3.29 70.925 3.55 ;
      RECT 69.375 2.73 69.695 2.99 ;
      RECT 68.895 2.45 69.215 2.71 ;
      RECT 68.045 1.89 68.445 2.15 ;
      RECT 67.695 3.57 68.015 3.83 ;
      RECT 66.015 2.45 66.335 2.71 ;
      RECT 65.535 2.73 65.855 2.99 ;
      RECT 64.845 1.89 65.165 2.15 ;
      RECT 64.845 3.29 65.165 3.55 ;
      RECT 56.515 2.45 56.835 2.71 ;
      RECT 55.345 3.29 55.665 3.55 ;
      RECT 54.115 2.73 54.435 2.99 ;
      RECT 53.635 2.45 53.955 2.71 ;
      RECT 52.785 1.89 53.185 2.15 ;
      RECT 52.435 3.57 52.755 3.83 ;
      RECT 50.755 2.45 51.075 2.71 ;
      RECT 50.275 2.73 50.595 2.99 ;
      RECT 49.585 1.89 49.905 2.15 ;
      RECT 49.585 3.29 49.905 3.55 ;
      RECT 41.255 2.45 41.575 2.71 ;
      RECT 40.085 3.29 40.405 3.55 ;
      RECT 38.855 2.73 39.175 2.99 ;
      RECT 38.375 2.45 38.695 2.71 ;
      RECT 37.525 1.89 37.925 2.15 ;
      RECT 37.175 3.57 37.495 3.83 ;
      RECT 35.495 2.45 35.815 2.71 ;
      RECT 35.015 2.73 35.335 2.99 ;
      RECT 34.325 1.89 34.645 2.15 ;
      RECT 34.325 3.29 34.645 3.55 ;
      RECT 25.995 2.45 26.315 2.71 ;
      RECT 24.825 3.29 25.145 3.55 ;
      RECT 23.595 2.73 23.915 2.99 ;
      RECT 23.115 2.45 23.435 2.71 ;
      RECT 22.265 1.89 22.665 2.15 ;
      RECT 21.915 3.57 22.235 3.83 ;
      RECT 20.235 2.45 20.555 2.71 ;
      RECT 19.755 2.73 20.075 2.99 ;
      RECT 19.065 1.89 19.385 2.15 ;
      RECT 19.065 3.29 19.385 3.55 ;
      RECT 10.735 2.45 11.055 2.71 ;
      RECT 9.565 3.29 9.885 3.55 ;
      RECT 8.335 2.73 8.655 2.99 ;
      RECT 7.855 2.45 8.175 2.71 ;
      RECT 7.005 1.89 7.405 2.15 ;
      RECT 6.655 3.57 6.975 3.83 ;
      RECT 4.975 2.45 5.295 2.71 ;
      RECT 4.495 2.73 4.815 2.99 ;
      RECT 3.805 1.89 4.125 2.15 ;
      RECT 3.805 3.29 4.125 3.55 ;
    LAYER mcon ;
      RECT 78.55 6.32 78.72 6.49 ;
      RECT 78.555 6.315 78.725 6.485 ;
      RECT 63.29 6.32 63.46 6.49 ;
      RECT 63.295 6.315 63.465 6.485 ;
      RECT 48.03 6.32 48.2 6.49 ;
      RECT 48.035 6.315 48.205 6.485 ;
      RECT 32.77 6.32 32.94 6.49 ;
      RECT 32.775 6.315 32.945 6.485 ;
      RECT 17.51 6.32 17.68 6.49 ;
      RECT 17.515 6.315 17.685 6.485 ;
      RECT 78.55 7.8 78.72 7.97 ;
      RECT 78.2 0.1 78.37 0.27 ;
      RECT 78.2 8.61 78.37 8.78 ;
      RECT 78.18 2.76 78.35 2.93 ;
      RECT 78.18 5.95 78.35 6.12 ;
      RECT 77.56 0.91 77.73 1.08 ;
      RECT 77.56 2.39 77.73 2.56 ;
      RECT 77.56 6.32 77.73 6.49 ;
      RECT 77.56 7.8 77.73 7.97 ;
      RECT 77.21 0.1 77.38 0.27 ;
      RECT 77.21 8.61 77.38 8.78 ;
      RECT 77.19 2.76 77.36 2.93 ;
      RECT 77.19 5.95 77.36 6.12 ;
      RECT 76.51 0.105 76.68 0.275 ;
      RECT 76.51 8.605 76.68 8.775 ;
      RECT 76.2 2.025 76.37 2.195 ;
      RECT 76.2 6.685 76.37 6.855 ;
      RECT 75.83 0.105 76 0.275 ;
      RECT 75.83 8.605 76 8.775 ;
      RECT 75.77 0.915 75.94 1.085 ;
      RECT 75.77 1.655 75.94 1.825 ;
      RECT 75.77 7.055 75.94 7.225 ;
      RECT 75.77 7.795 75.94 7.965 ;
      RECT 75.395 2.395 75.565 2.565 ;
      RECT 75.395 6.315 75.565 6.485 ;
      RECT 75.15 0.105 75.32 0.275 ;
      RECT 75.15 8.605 75.32 8.775 ;
      RECT 74.47 0.105 74.64 0.275 ;
      RECT 74.47 8.605 74.64 8.775 ;
      RECT 72.335 2.77 72.505 2.94 ;
      RECT 72.095 1.93 72.265 2.1 ;
      RECT 72.095 3.61 72.265 3.78 ;
      RECT 71.855 2.49 72.025 2.66 ;
      RECT 71.855 3.05 72.025 3.22 ;
      RECT 71.375 2.77 71.545 2.94 ;
      RECT 71.135 1.93 71.305 2.1 ;
      RECT 70.895 2.49 71.065 2.66 ;
      RECT 70.895 8.605 71.065 8.775 ;
      RECT 70.685 3.33 70.855 3.5 ;
      RECT 70.585 6.685 70.755 6.855 ;
      RECT 70.415 2.77 70.585 2.94 ;
      RECT 70.215 8.605 70.385 8.775 ;
      RECT 70.155 7.055 70.325 7.225 ;
      RECT 70.155 7.795 70.325 7.965 ;
      RECT 70.145 3.61 70.315 3.78 ;
      RECT 69.935 2.19 70.105 2.36 ;
      RECT 69.78 6.315 69.95 6.485 ;
      RECT 69.535 8.605 69.705 8.775 ;
      RECT 69.455 2.77 69.625 2.94 ;
      RECT 69.215 1.93 69.385 2.1 ;
      RECT 68.975 2.49 69.145 2.66 ;
      RECT 68.975 3.05 69.145 3.22 ;
      RECT 68.855 8.605 69.025 8.775 ;
      RECT 68.495 2.49 68.665 2.66 ;
      RECT 68.255 3.61 68.425 3.78 ;
      RECT 68.215 1.93 68.385 2.1 ;
      RECT 68.015 2.77 68.185 2.94 ;
      RECT 67.775 3.61 67.945 3.78 ;
      RECT 67.535 3.05 67.705 3.22 ;
      RECT 67.055 2.49 67.225 2.66 ;
      RECT 66.815 1.93 66.985 2.1 ;
      RECT 66.815 3.61 66.985 3.78 ;
      RECT 66.335 1.93 66.505 2.1 ;
      RECT 66.335 3.05 66.505 3.22 ;
      RECT 66.095 2.49 66.265 2.66 ;
      RECT 65.855 3.33 66.025 3.5 ;
      RECT 65.615 2.77 65.785 2.94 ;
      RECT 65.135 2.77 65.305 2.94 ;
      RECT 64.925 1.93 65.095 2.1 ;
      RECT 64.925 3.33 65.095 3.5 ;
      RECT 63.29 7.8 63.46 7.97 ;
      RECT 62.94 0.1 63.11 0.27 ;
      RECT 62.94 8.61 63.11 8.78 ;
      RECT 62.92 2.76 63.09 2.93 ;
      RECT 62.92 5.95 63.09 6.12 ;
      RECT 62.3 0.91 62.47 1.08 ;
      RECT 62.3 2.39 62.47 2.56 ;
      RECT 62.3 6.32 62.47 6.49 ;
      RECT 62.3 7.8 62.47 7.97 ;
      RECT 61.95 0.1 62.12 0.27 ;
      RECT 61.95 8.61 62.12 8.78 ;
      RECT 61.93 2.76 62.1 2.93 ;
      RECT 61.93 5.95 62.1 6.12 ;
      RECT 61.25 0.105 61.42 0.275 ;
      RECT 61.25 8.605 61.42 8.775 ;
      RECT 60.94 2.025 61.11 2.195 ;
      RECT 60.94 6.685 61.11 6.855 ;
      RECT 60.57 0.105 60.74 0.275 ;
      RECT 60.57 8.605 60.74 8.775 ;
      RECT 60.51 0.915 60.68 1.085 ;
      RECT 60.51 1.655 60.68 1.825 ;
      RECT 60.51 7.055 60.68 7.225 ;
      RECT 60.51 7.795 60.68 7.965 ;
      RECT 60.135 2.395 60.305 2.565 ;
      RECT 60.135 6.315 60.305 6.485 ;
      RECT 59.89 0.105 60.06 0.275 ;
      RECT 59.89 8.605 60.06 8.775 ;
      RECT 59.21 0.105 59.38 0.275 ;
      RECT 59.21 8.605 59.38 8.775 ;
      RECT 57.075 2.77 57.245 2.94 ;
      RECT 56.835 1.93 57.005 2.1 ;
      RECT 56.835 3.61 57.005 3.78 ;
      RECT 56.595 2.49 56.765 2.66 ;
      RECT 56.595 3.05 56.765 3.22 ;
      RECT 56.115 2.77 56.285 2.94 ;
      RECT 55.875 1.93 56.045 2.1 ;
      RECT 55.635 2.49 55.805 2.66 ;
      RECT 55.635 8.605 55.805 8.775 ;
      RECT 55.425 3.33 55.595 3.5 ;
      RECT 55.325 6.685 55.495 6.855 ;
      RECT 55.155 2.77 55.325 2.94 ;
      RECT 54.955 8.605 55.125 8.775 ;
      RECT 54.895 7.055 55.065 7.225 ;
      RECT 54.895 7.795 55.065 7.965 ;
      RECT 54.885 3.61 55.055 3.78 ;
      RECT 54.675 2.19 54.845 2.36 ;
      RECT 54.52 6.315 54.69 6.485 ;
      RECT 54.275 8.605 54.445 8.775 ;
      RECT 54.195 2.77 54.365 2.94 ;
      RECT 53.955 1.93 54.125 2.1 ;
      RECT 53.715 2.49 53.885 2.66 ;
      RECT 53.715 3.05 53.885 3.22 ;
      RECT 53.595 8.605 53.765 8.775 ;
      RECT 53.235 2.49 53.405 2.66 ;
      RECT 52.995 3.61 53.165 3.78 ;
      RECT 52.955 1.93 53.125 2.1 ;
      RECT 52.755 2.77 52.925 2.94 ;
      RECT 52.515 3.61 52.685 3.78 ;
      RECT 52.275 3.05 52.445 3.22 ;
      RECT 51.795 2.49 51.965 2.66 ;
      RECT 51.555 1.93 51.725 2.1 ;
      RECT 51.555 3.61 51.725 3.78 ;
      RECT 51.075 1.93 51.245 2.1 ;
      RECT 51.075 3.05 51.245 3.22 ;
      RECT 50.835 2.49 51.005 2.66 ;
      RECT 50.595 3.33 50.765 3.5 ;
      RECT 50.355 2.77 50.525 2.94 ;
      RECT 49.875 2.77 50.045 2.94 ;
      RECT 49.665 1.93 49.835 2.1 ;
      RECT 49.665 3.33 49.835 3.5 ;
      RECT 48.03 7.8 48.2 7.97 ;
      RECT 47.68 0.1 47.85 0.27 ;
      RECT 47.68 8.61 47.85 8.78 ;
      RECT 47.66 2.76 47.83 2.93 ;
      RECT 47.66 5.95 47.83 6.12 ;
      RECT 47.04 0.91 47.21 1.08 ;
      RECT 47.04 2.39 47.21 2.56 ;
      RECT 47.04 6.32 47.21 6.49 ;
      RECT 47.04 7.8 47.21 7.97 ;
      RECT 46.69 0.1 46.86 0.27 ;
      RECT 46.69 8.61 46.86 8.78 ;
      RECT 46.67 2.76 46.84 2.93 ;
      RECT 46.67 5.95 46.84 6.12 ;
      RECT 45.99 0.105 46.16 0.275 ;
      RECT 45.99 8.605 46.16 8.775 ;
      RECT 45.68 2.025 45.85 2.195 ;
      RECT 45.68 6.685 45.85 6.855 ;
      RECT 45.31 0.105 45.48 0.275 ;
      RECT 45.31 8.605 45.48 8.775 ;
      RECT 45.25 0.915 45.42 1.085 ;
      RECT 45.25 1.655 45.42 1.825 ;
      RECT 45.25 7.055 45.42 7.225 ;
      RECT 45.25 7.795 45.42 7.965 ;
      RECT 44.875 2.395 45.045 2.565 ;
      RECT 44.875 6.315 45.045 6.485 ;
      RECT 44.63 0.105 44.8 0.275 ;
      RECT 44.63 8.605 44.8 8.775 ;
      RECT 43.95 0.105 44.12 0.275 ;
      RECT 43.95 8.605 44.12 8.775 ;
      RECT 41.815 2.77 41.985 2.94 ;
      RECT 41.575 1.93 41.745 2.1 ;
      RECT 41.575 3.61 41.745 3.78 ;
      RECT 41.335 2.49 41.505 2.66 ;
      RECT 41.335 3.05 41.505 3.22 ;
      RECT 40.855 2.77 41.025 2.94 ;
      RECT 40.615 1.93 40.785 2.1 ;
      RECT 40.375 2.49 40.545 2.66 ;
      RECT 40.375 8.605 40.545 8.775 ;
      RECT 40.165 3.33 40.335 3.5 ;
      RECT 40.065 6.685 40.235 6.855 ;
      RECT 39.895 2.77 40.065 2.94 ;
      RECT 39.695 8.605 39.865 8.775 ;
      RECT 39.635 7.055 39.805 7.225 ;
      RECT 39.635 7.795 39.805 7.965 ;
      RECT 39.625 3.61 39.795 3.78 ;
      RECT 39.415 2.19 39.585 2.36 ;
      RECT 39.26 6.315 39.43 6.485 ;
      RECT 39.015 8.605 39.185 8.775 ;
      RECT 38.935 2.77 39.105 2.94 ;
      RECT 38.695 1.93 38.865 2.1 ;
      RECT 38.455 2.49 38.625 2.66 ;
      RECT 38.455 3.05 38.625 3.22 ;
      RECT 38.335 8.605 38.505 8.775 ;
      RECT 37.975 2.49 38.145 2.66 ;
      RECT 37.735 3.61 37.905 3.78 ;
      RECT 37.695 1.93 37.865 2.1 ;
      RECT 37.495 2.77 37.665 2.94 ;
      RECT 37.255 3.61 37.425 3.78 ;
      RECT 37.015 3.05 37.185 3.22 ;
      RECT 36.535 2.49 36.705 2.66 ;
      RECT 36.295 1.93 36.465 2.1 ;
      RECT 36.295 3.61 36.465 3.78 ;
      RECT 35.815 1.93 35.985 2.1 ;
      RECT 35.815 3.05 35.985 3.22 ;
      RECT 35.575 2.49 35.745 2.66 ;
      RECT 35.335 3.33 35.505 3.5 ;
      RECT 35.095 2.77 35.265 2.94 ;
      RECT 34.615 2.77 34.785 2.94 ;
      RECT 34.405 1.93 34.575 2.1 ;
      RECT 34.405 3.33 34.575 3.5 ;
      RECT 32.77 7.8 32.94 7.97 ;
      RECT 32.42 0.1 32.59 0.27 ;
      RECT 32.42 8.61 32.59 8.78 ;
      RECT 32.4 2.76 32.57 2.93 ;
      RECT 32.4 5.95 32.57 6.12 ;
      RECT 31.78 0.91 31.95 1.08 ;
      RECT 31.78 2.39 31.95 2.56 ;
      RECT 31.78 6.32 31.95 6.49 ;
      RECT 31.78 7.8 31.95 7.97 ;
      RECT 31.43 0.1 31.6 0.27 ;
      RECT 31.43 8.61 31.6 8.78 ;
      RECT 31.41 2.76 31.58 2.93 ;
      RECT 31.41 5.95 31.58 6.12 ;
      RECT 30.73 0.105 30.9 0.275 ;
      RECT 30.73 8.605 30.9 8.775 ;
      RECT 30.42 2.025 30.59 2.195 ;
      RECT 30.42 6.685 30.59 6.855 ;
      RECT 30.05 0.105 30.22 0.275 ;
      RECT 30.05 8.605 30.22 8.775 ;
      RECT 29.99 0.915 30.16 1.085 ;
      RECT 29.99 1.655 30.16 1.825 ;
      RECT 29.99 7.055 30.16 7.225 ;
      RECT 29.99 7.795 30.16 7.965 ;
      RECT 29.615 2.395 29.785 2.565 ;
      RECT 29.615 6.315 29.785 6.485 ;
      RECT 29.37 0.105 29.54 0.275 ;
      RECT 29.37 8.605 29.54 8.775 ;
      RECT 28.69 0.105 28.86 0.275 ;
      RECT 28.69 8.605 28.86 8.775 ;
      RECT 26.555 2.77 26.725 2.94 ;
      RECT 26.315 1.93 26.485 2.1 ;
      RECT 26.315 3.61 26.485 3.78 ;
      RECT 26.075 2.49 26.245 2.66 ;
      RECT 26.075 3.05 26.245 3.22 ;
      RECT 25.595 2.77 25.765 2.94 ;
      RECT 25.355 1.93 25.525 2.1 ;
      RECT 25.115 2.49 25.285 2.66 ;
      RECT 25.115 8.605 25.285 8.775 ;
      RECT 24.905 3.33 25.075 3.5 ;
      RECT 24.805 6.685 24.975 6.855 ;
      RECT 24.635 2.77 24.805 2.94 ;
      RECT 24.435 8.605 24.605 8.775 ;
      RECT 24.375 7.055 24.545 7.225 ;
      RECT 24.375 7.795 24.545 7.965 ;
      RECT 24.365 3.61 24.535 3.78 ;
      RECT 24.155 2.19 24.325 2.36 ;
      RECT 24 6.315 24.17 6.485 ;
      RECT 23.755 8.605 23.925 8.775 ;
      RECT 23.675 2.77 23.845 2.94 ;
      RECT 23.435 1.93 23.605 2.1 ;
      RECT 23.195 2.49 23.365 2.66 ;
      RECT 23.195 3.05 23.365 3.22 ;
      RECT 23.075 8.605 23.245 8.775 ;
      RECT 22.715 2.49 22.885 2.66 ;
      RECT 22.475 3.61 22.645 3.78 ;
      RECT 22.435 1.93 22.605 2.1 ;
      RECT 22.235 2.77 22.405 2.94 ;
      RECT 21.995 3.61 22.165 3.78 ;
      RECT 21.755 3.05 21.925 3.22 ;
      RECT 21.275 2.49 21.445 2.66 ;
      RECT 21.035 1.93 21.205 2.1 ;
      RECT 21.035 3.61 21.205 3.78 ;
      RECT 20.555 1.93 20.725 2.1 ;
      RECT 20.555 3.05 20.725 3.22 ;
      RECT 20.315 2.49 20.485 2.66 ;
      RECT 20.075 3.33 20.245 3.5 ;
      RECT 19.835 2.77 20.005 2.94 ;
      RECT 19.355 2.77 19.525 2.94 ;
      RECT 19.145 1.93 19.315 2.1 ;
      RECT 19.145 3.33 19.315 3.5 ;
      RECT 17.51 7.8 17.68 7.97 ;
      RECT 17.16 0.1 17.33 0.27 ;
      RECT 17.16 8.61 17.33 8.78 ;
      RECT 17.14 2.76 17.31 2.93 ;
      RECT 17.14 5.95 17.31 6.12 ;
      RECT 16.52 0.91 16.69 1.08 ;
      RECT 16.52 2.39 16.69 2.56 ;
      RECT 16.52 6.32 16.69 6.49 ;
      RECT 16.52 7.8 16.69 7.97 ;
      RECT 16.17 0.1 16.34 0.27 ;
      RECT 16.17 8.61 16.34 8.78 ;
      RECT 16.15 2.76 16.32 2.93 ;
      RECT 16.15 5.95 16.32 6.12 ;
      RECT 15.47 0.105 15.64 0.275 ;
      RECT 15.47 8.605 15.64 8.775 ;
      RECT 15.16 2.025 15.33 2.195 ;
      RECT 15.16 6.685 15.33 6.855 ;
      RECT 14.79 0.105 14.96 0.275 ;
      RECT 14.79 8.605 14.96 8.775 ;
      RECT 14.73 0.915 14.9 1.085 ;
      RECT 14.73 1.655 14.9 1.825 ;
      RECT 14.73 7.055 14.9 7.225 ;
      RECT 14.73 7.795 14.9 7.965 ;
      RECT 14.355 2.395 14.525 2.565 ;
      RECT 14.355 6.315 14.525 6.485 ;
      RECT 14.11 0.105 14.28 0.275 ;
      RECT 14.11 8.605 14.28 8.775 ;
      RECT 13.43 0.105 13.6 0.275 ;
      RECT 13.43 8.605 13.6 8.775 ;
      RECT 11.295 2.77 11.465 2.94 ;
      RECT 11.055 1.93 11.225 2.1 ;
      RECT 11.055 3.61 11.225 3.78 ;
      RECT 10.815 2.49 10.985 2.66 ;
      RECT 10.815 3.05 10.985 3.22 ;
      RECT 10.335 2.77 10.505 2.94 ;
      RECT 10.095 1.93 10.265 2.1 ;
      RECT 9.855 2.49 10.025 2.66 ;
      RECT 9.855 8.605 10.025 8.775 ;
      RECT 9.645 3.33 9.815 3.5 ;
      RECT 9.545 6.685 9.715 6.855 ;
      RECT 9.375 2.77 9.545 2.94 ;
      RECT 9.175 8.605 9.345 8.775 ;
      RECT 9.115 7.055 9.285 7.225 ;
      RECT 9.115 7.795 9.285 7.965 ;
      RECT 9.105 3.61 9.275 3.78 ;
      RECT 8.895 2.19 9.065 2.36 ;
      RECT 8.74 6.315 8.91 6.485 ;
      RECT 8.495 8.605 8.665 8.775 ;
      RECT 8.415 2.77 8.585 2.94 ;
      RECT 8.175 1.93 8.345 2.1 ;
      RECT 7.935 2.49 8.105 2.66 ;
      RECT 7.935 3.05 8.105 3.22 ;
      RECT 7.815 8.605 7.985 8.775 ;
      RECT 7.455 2.49 7.625 2.66 ;
      RECT 7.215 3.61 7.385 3.78 ;
      RECT 7.175 1.93 7.345 2.1 ;
      RECT 6.975 2.77 7.145 2.94 ;
      RECT 6.735 3.61 6.905 3.78 ;
      RECT 6.495 3.05 6.665 3.22 ;
      RECT 6.015 2.49 6.185 2.66 ;
      RECT 5.775 1.93 5.945 2.1 ;
      RECT 5.775 3.61 5.945 3.78 ;
      RECT 5.295 1.93 5.465 2.1 ;
      RECT 5.295 3.05 5.465 3.22 ;
      RECT 5.055 2.49 5.225 2.66 ;
      RECT 4.815 3.33 4.985 3.5 ;
      RECT 4.575 2.77 4.745 2.94 ;
      RECT 4.095 2.77 4.265 2.94 ;
      RECT 3.885 1.93 4.055 2.1 ;
      RECT 3.885 3.33 4.055 3.5 ;
      RECT 2.34 8.605 2.51 8.775 ;
      RECT 1.66 8.605 1.83 8.775 ;
      RECT 1.6 7.055 1.77 7.225 ;
      RECT 1.6 7.795 1.77 7.965 ;
      RECT 1.225 6.315 1.395 6.485 ;
      RECT 0.98 8.605 1.15 8.775 ;
      RECT 0.3 8.605 0.47 8.775 ;
    LAYER li1 ;
      RECT 72.555 0 72.725 2.08 ;
      RECT 71.615 0 71.785 2.08 ;
      RECT 70.655 0 70.825 2.08 ;
      RECT 68.735 0 68.905 2.08 ;
      RECT 67.775 0 67.945 2.08 ;
      RECT 65.855 0 66.025 2.08 ;
      RECT 57.295 0 57.465 2.08 ;
      RECT 56.355 0 56.525 2.08 ;
      RECT 55.395 0 55.565 2.08 ;
      RECT 53.475 0 53.645 2.08 ;
      RECT 52.515 0 52.685 2.08 ;
      RECT 50.595 0 50.765 2.08 ;
      RECT 42.035 0 42.205 2.08 ;
      RECT 41.095 0 41.265 2.08 ;
      RECT 40.135 0 40.305 2.08 ;
      RECT 38.215 0 38.385 2.08 ;
      RECT 37.255 0 37.425 2.08 ;
      RECT 35.335 0 35.505 2.08 ;
      RECT 26.775 0 26.945 2.08 ;
      RECT 25.835 0 26.005 2.08 ;
      RECT 24.875 0 25.045 2.08 ;
      RECT 22.955 0 23.125 2.08 ;
      RECT 21.995 0 22.165 2.08 ;
      RECT 20.075 0 20.245 2.08 ;
      RECT 11.515 0 11.685 2.08 ;
      RECT 10.575 0 10.745 2.08 ;
      RECT 9.615 0 9.785 2.08 ;
      RECT 7.695 0 7.865 2.08 ;
      RECT 6.735 0 6.905 2.08 ;
      RECT 4.815 0 4.985 2.08 ;
      RECT 69.61 0 69.805 1.595 ;
      RECT 65.855 0 66.13 1.595 ;
      RECT 54.35 0 54.545 1.595 ;
      RECT 50.595 0 50.87 1.595 ;
      RECT 39.09 0 39.285 1.595 ;
      RECT 35.335 0 35.61 1.595 ;
      RECT 23.83 0 24.025 1.595 ;
      RECT 20.075 0 20.35 1.595 ;
      RECT 8.57 0 8.765 1.595 ;
      RECT 4.815 0 5.09 1.595 ;
      RECT 73.13 0 73.325 1.585 ;
      RECT 71.46 0 71.785 1.585 ;
      RECT 57.87 0 58.065 1.585 ;
      RECT 56.2 0 56.525 1.585 ;
      RECT 42.61 0 42.805 1.585 ;
      RECT 40.94 0 41.265 1.585 ;
      RECT 27.35 0 27.545 1.585 ;
      RECT 25.68 0 26.005 1.585 ;
      RECT 12.09 0 12.285 1.585 ;
      RECT 10.42 0 10.745 1.585 ;
      RECT 64.585 0 73.325 1.58 ;
      RECT 49.325 0 58.065 1.58 ;
      RECT 34.065 0 42.805 1.58 ;
      RECT 18.805 0 27.545 1.58 ;
      RECT 3.545 0 12.285 1.58 ;
      RECT 74.39 0 74.56 0.935 ;
      RECT 59.13 0 59.3 0.935 ;
      RECT 43.87 0 44.04 0.935 ;
      RECT 28.61 0 28.78 0.935 ;
      RECT 13.35 0 13.52 0.935 ;
      RECT 78.12 0 78.29 0.93 ;
      RECT 77.13 0 77.3 0.93 ;
      RECT 62.86 0 63.03 0.93 ;
      RECT 61.87 0 62.04 0.93 ;
      RECT 47.6 0 47.77 0.93 ;
      RECT 46.61 0 46.78 0.93 ;
      RECT 32.34 0 32.51 0.93 ;
      RECT 31.35 0 31.52 0.93 ;
      RECT 17.08 0 17.25 0.93 ;
      RECT 16.09 0 16.26 0.93 ;
      RECT 0.295 0.245 0.465 0.335 ;
      RECT 0 0.245 0.805 0.315 ;
      RECT 78.915 0 79.095 0.305 ;
      RECT 63.655 0 76.965 0.305 ;
      RECT 48.395 0 61.705 0.305 ;
      RECT 33.135 0 46.445 0.305 ;
      RECT 17.875 0 31.185 0.305 ;
      RECT 0 0.245 15.925 0.305 ;
      RECT 0.465 0 79.095 0.3 ;
      RECT 0 0 0.295 0.315 ;
      RECT 0 0 79.095 0.075 ;
      RECT 0 8.58 79.095 8.88 ;
      RECT 78.915 8.575 79.095 8.88 ;
      RECT 78.12 7.95 78.29 8.88 ;
      RECT 77.13 7.95 77.3 8.88 ;
      RECT 63.655 8.575 76.965 8.88 ;
      RECT 62.86 7.95 63.03 8.88 ;
      RECT 61.87 7.95 62.04 8.88 ;
      RECT 48.395 8.575 61.705 8.88 ;
      RECT 47.6 7.95 47.77 8.88 ;
      RECT 46.61 7.95 46.78 8.88 ;
      RECT 33.135 8.575 46.445 8.88 ;
      RECT 32.34 7.95 32.51 8.88 ;
      RECT 31.35 7.95 31.52 8.88 ;
      RECT 17.875 8.575 31.185 8.88 ;
      RECT 17.08 7.95 17.25 8.88 ;
      RECT 16.09 7.95 16.26 8.88 ;
      RECT 0 8.575 15.925 8.88 ;
      RECT 74.39 7.945 74.56 8.88 ;
      RECT 68.775 7.945 68.945 8.88 ;
      RECT 59.13 7.945 59.3 8.88 ;
      RECT 53.515 7.945 53.685 8.88 ;
      RECT 43.87 7.945 44.04 8.88 ;
      RECT 38.255 7.945 38.425 8.88 ;
      RECT 28.61 7.945 28.78 8.88 ;
      RECT 22.995 7.945 23.165 8.88 ;
      RECT 13.35 7.945 13.52 8.88 ;
      RECT 7.735 7.945 7.905 8.88 ;
      RECT 0.005 8.565 0.81 8.88 ;
      RECT 0.22 8.545 0.47 8.88 ;
      RECT 0.22 7.945 0.39 8.88 ;
      RECT 78.55 5.02 78.72 6.49 ;
      RECT 78.55 6.315 78.725 6.485 ;
      RECT 78.18 1.74 78.35 2.93 ;
      RECT 78.18 1.74 78.65 1.91 ;
      RECT 78.18 6.97 78.65 7.14 ;
      RECT 78.18 5.95 78.35 7.14 ;
      RECT 77.19 1.74 77.36 2.93 ;
      RECT 77.19 1.74 77.66 1.91 ;
      RECT 77.19 6.97 77.66 7.14 ;
      RECT 77.19 5.95 77.36 7.14 ;
      RECT 75.34 2.635 75.51 3.865 ;
      RECT 75.395 0.855 75.565 2.805 ;
      RECT 75.34 0.575 75.51 1.025 ;
      RECT 75.34 7.855 75.51 8.305 ;
      RECT 75.395 6.075 75.565 8.025 ;
      RECT 75.34 5.015 75.51 6.245 ;
      RECT 74.82 0.575 74.99 3.865 ;
      RECT 74.82 2.075 75.225 2.405 ;
      RECT 74.82 1.235 75.225 1.565 ;
      RECT 74.82 5.015 74.99 8.305 ;
      RECT 74.82 7.315 75.225 7.645 ;
      RECT 74.82 6.475 75.225 6.805 ;
      RECT 72.095 3.61 72.605 3.78 ;
      RECT 72.435 3.22 72.605 3.78 ;
      RECT 72.545 3.14 72.715 3.47 ;
      RECT 72.335 2.53 72.605 2.94 ;
      RECT 72.215 2.53 72.605 2.74 ;
      RECT 70.685 3.14 70.855 3.5 ;
      RECT 70.685 3.22 72.025 3.39 ;
      RECT 71.855 3.05 72.025 3.39 ;
      RECT 70.415 2.57 70.585 2.94 ;
      RECT 69.935 2.57 70.585 2.84 ;
      RECT 69.855 2.57 70.665 2.74 ;
      RECT 69.215 1.81 69.385 2.1 ;
      RECT 69.215 1.81 70.455 1.98 ;
      RECT 69.935 2.15 70.105 2.36 ;
      RECT 69.575 2.15 70.105 2.32 ;
      RECT 69.725 7.855 69.895 8.305 ;
      RECT 69.78 6.075 69.95 8.025 ;
      RECT 69.725 5.015 69.895 6.245 ;
      RECT 69.205 5.015 69.375 8.305 ;
      RECT 69.205 7.315 69.61 7.645 ;
      RECT 69.205 6.475 69.61 6.805 ;
      RECT 68.975 3.22 69.465 3.39 ;
      RECT 68.975 3.05 69.145 3.39 ;
      RECT 68.255 3.22 68.425 3.78 ;
      RECT 68.145 3.22 68.475 3.39 ;
      RECT 68.215 1.83 68.385 2.1 ;
      RECT 68.255 1.75 68.425 2.08 ;
      RECT 68.115 1.83 68.425 2.05 ;
      RECT 66.695 3.22 66.985 3.78 ;
      RECT 66.815 3.14 66.985 3.78 ;
      RECT 66.455 2.57 66.825 2.74 ;
      RECT 66.455 1.93 66.625 2.74 ;
      RECT 66.335 1.93 66.625 2.1 ;
      RECT 63.29 5.02 63.46 6.49 ;
      RECT 63.29 6.315 63.465 6.485 ;
      RECT 62.92 1.74 63.09 2.93 ;
      RECT 62.92 1.74 63.39 1.91 ;
      RECT 62.92 6.97 63.39 7.14 ;
      RECT 62.92 5.95 63.09 7.14 ;
      RECT 61.93 1.74 62.1 2.93 ;
      RECT 61.93 1.74 62.4 1.91 ;
      RECT 61.93 6.97 62.4 7.14 ;
      RECT 61.93 5.95 62.1 7.14 ;
      RECT 60.08 2.635 60.25 3.865 ;
      RECT 60.135 0.855 60.305 2.805 ;
      RECT 60.08 0.575 60.25 1.025 ;
      RECT 60.08 7.855 60.25 8.305 ;
      RECT 60.135 6.075 60.305 8.025 ;
      RECT 60.08 5.015 60.25 6.245 ;
      RECT 59.56 0.575 59.73 3.865 ;
      RECT 59.56 2.075 59.965 2.405 ;
      RECT 59.56 1.235 59.965 1.565 ;
      RECT 59.56 5.015 59.73 8.305 ;
      RECT 59.56 7.315 59.965 7.645 ;
      RECT 59.56 6.475 59.965 6.805 ;
      RECT 56.835 3.61 57.345 3.78 ;
      RECT 57.175 3.22 57.345 3.78 ;
      RECT 57.285 3.14 57.455 3.47 ;
      RECT 57.075 2.53 57.345 2.94 ;
      RECT 56.955 2.53 57.345 2.74 ;
      RECT 55.425 3.14 55.595 3.5 ;
      RECT 55.425 3.22 56.765 3.39 ;
      RECT 56.595 3.05 56.765 3.39 ;
      RECT 55.155 2.57 55.325 2.94 ;
      RECT 54.675 2.57 55.325 2.84 ;
      RECT 54.595 2.57 55.405 2.74 ;
      RECT 53.955 1.81 54.125 2.1 ;
      RECT 53.955 1.81 55.195 1.98 ;
      RECT 54.675 2.15 54.845 2.36 ;
      RECT 54.315 2.15 54.845 2.32 ;
      RECT 54.465 7.855 54.635 8.305 ;
      RECT 54.52 6.075 54.69 8.025 ;
      RECT 54.465 5.015 54.635 6.245 ;
      RECT 53.945 5.015 54.115 8.305 ;
      RECT 53.945 7.315 54.35 7.645 ;
      RECT 53.945 6.475 54.35 6.805 ;
      RECT 53.715 3.22 54.205 3.39 ;
      RECT 53.715 3.05 53.885 3.39 ;
      RECT 52.995 3.22 53.165 3.78 ;
      RECT 52.885 3.22 53.215 3.39 ;
      RECT 52.955 1.83 53.125 2.1 ;
      RECT 52.995 1.75 53.165 2.08 ;
      RECT 52.855 1.83 53.165 2.05 ;
      RECT 51.435 3.22 51.725 3.78 ;
      RECT 51.555 3.14 51.725 3.78 ;
      RECT 51.195 2.57 51.565 2.74 ;
      RECT 51.195 1.93 51.365 2.74 ;
      RECT 51.075 1.93 51.365 2.1 ;
      RECT 48.03 5.02 48.2 6.49 ;
      RECT 48.03 6.315 48.205 6.485 ;
      RECT 47.66 1.74 47.83 2.93 ;
      RECT 47.66 1.74 48.13 1.91 ;
      RECT 47.66 6.97 48.13 7.14 ;
      RECT 47.66 5.95 47.83 7.14 ;
      RECT 46.67 1.74 46.84 2.93 ;
      RECT 46.67 1.74 47.14 1.91 ;
      RECT 46.67 6.97 47.14 7.14 ;
      RECT 46.67 5.95 46.84 7.14 ;
      RECT 44.82 2.635 44.99 3.865 ;
      RECT 44.875 0.855 45.045 2.805 ;
      RECT 44.82 0.575 44.99 1.025 ;
      RECT 44.82 7.855 44.99 8.305 ;
      RECT 44.875 6.075 45.045 8.025 ;
      RECT 44.82 5.015 44.99 6.245 ;
      RECT 44.3 0.575 44.47 3.865 ;
      RECT 44.3 2.075 44.705 2.405 ;
      RECT 44.3 1.235 44.705 1.565 ;
      RECT 44.3 5.015 44.47 8.305 ;
      RECT 44.3 7.315 44.705 7.645 ;
      RECT 44.3 6.475 44.705 6.805 ;
      RECT 41.575 3.61 42.085 3.78 ;
      RECT 41.915 3.22 42.085 3.78 ;
      RECT 42.025 3.14 42.195 3.47 ;
      RECT 41.815 2.53 42.085 2.94 ;
      RECT 41.695 2.53 42.085 2.74 ;
      RECT 40.165 3.14 40.335 3.5 ;
      RECT 40.165 3.22 41.505 3.39 ;
      RECT 41.335 3.05 41.505 3.39 ;
      RECT 39.895 2.57 40.065 2.94 ;
      RECT 39.415 2.57 40.065 2.84 ;
      RECT 39.335 2.57 40.145 2.74 ;
      RECT 38.695 1.81 38.865 2.1 ;
      RECT 38.695 1.81 39.935 1.98 ;
      RECT 39.415 2.15 39.585 2.36 ;
      RECT 39.055 2.15 39.585 2.32 ;
      RECT 39.205 7.855 39.375 8.305 ;
      RECT 39.26 6.075 39.43 8.025 ;
      RECT 39.205 5.015 39.375 6.245 ;
      RECT 38.685 5.015 38.855 8.305 ;
      RECT 38.685 7.315 39.09 7.645 ;
      RECT 38.685 6.475 39.09 6.805 ;
      RECT 38.455 3.22 38.945 3.39 ;
      RECT 38.455 3.05 38.625 3.39 ;
      RECT 37.735 3.22 37.905 3.78 ;
      RECT 37.625 3.22 37.955 3.39 ;
      RECT 37.695 1.83 37.865 2.1 ;
      RECT 37.735 1.75 37.905 2.08 ;
      RECT 37.595 1.83 37.905 2.05 ;
      RECT 36.175 3.22 36.465 3.78 ;
      RECT 36.295 3.14 36.465 3.78 ;
      RECT 35.935 2.57 36.305 2.74 ;
      RECT 35.935 1.93 36.105 2.74 ;
      RECT 35.815 1.93 36.105 2.1 ;
      RECT 32.77 5.02 32.94 6.49 ;
      RECT 32.77 6.315 32.945 6.485 ;
      RECT 32.4 1.74 32.57 2.93 ;
      RECT 32.4 1.74 32.87 1.91 ;
      RECT 32.4 6.97 32.87 7.14 ;
      RECT 32.4 5.95 32.57 7.14 ;
      RECT 31.41 1.74 31.58 2.93 ;
      RECT 31.41 1.74 31.88 1.91 ;
      RECT 31.41 6.97 31.88 7.14 ;
      RECT 31.41 5.95 31.58 7.14 ;
      RECT 29.56 2.635 29.73 3.865 ;
      RECT 29.615 0.855 29.785 2.805 ;
      RECT 29.56 0.575 29.73 1.025 ;
      RECT 29.56 7.855 29.73 8.305 ;
      RECT 29.615 6.075 29.785 8.025 ;
      RECT 29.56 5.015 29.73 6.245 ;
      RECT 29.04 0.575 29.21 3.865 ;
      RECT 29.04 2.075 29.445 2.405 ;
      RECT 29.04 1.235 29.445 1.565 ;
      RECT 29.04 5.015 29.21 8.305 ;
      RECT 29.04 7.315 29.445 7.645 ;
      RECT 29.04 6.475 29.445 6.805 ;
      RECT 26.315 3.61 26.825 3.78 ;
      RECT 26.655 3.22 26.825 3.78 ;
      RECT 26.765 3.14 26.935 3.47 ;
      RECT 26.555 2.53 26.825 2.94 ;
      RECT 26.435 2.53 26.825 2.74 ;
      RECT 24.905 3.14 25.075 3.5 ;
      RECT 24.905 3.22 26.245 3.39 ;
      RECT 26.075 3.05 26.245 3.39 ;
      RECT 24.635 2.57 24.805 2.94 ;
      RECT 24.155 2.57 24.805 2.84 ;
      RECT 24.075 2.57 24.885 2.74 ;
      RECT 23.435 1.81 23.605 2.1 ;
      RECT 23.435 1.81 24.675 1.98 ;
      RECT 24.155 2.15 24.325 2.36 ;
      RECT 23.795 2.15 24.325 2.32 ;
      RECT 23.945 7.855 24.115 8.305 ;
      RECT 24 6.075 24.17 8.025 ;
      RECT 23.945 5.015 24.115 6.245 ;
      RECT 23.425 5.015 23.595 8.305 ;
      RECT 23.425 7.315 23.83 7.645 ;
      RECT 23.425 6.475 23.83 6.805 ;
      RECT 23.195 3.22 23.685 3.39 ;
      RECT 23.195 3.05 23.365 3.39 ;
      RECT 22.475 3.22 22.645 3.78 ;
      RECT 22.365 3.22 22.695 3.39 ;
      RECT 22.435 1.83 22.605 2.1 ;
      RECT 22.475 1.75 22.645 2.08 ;
      RECT 22.335 1.83 22.645 2.05 ;
      RECT 20.915 3.22 21.205 3.78 ;
      RECT 21.035 3.14 21.205 3.78 ;
      RECT 20.675 2.57 21.045 2.74 ;
      RECT 20.675 1.93 20.845 2.74 ;
      RECT 20.555 1.93 20.845 2.1 ;
      RECT 17.51 5.02 17.68 6.49 ;
      RECT 17.51 6.315 17.685 6.485 ;
      RECT 17.14 1.74 17.31 2.93 ;
      RECT 17.14 1.74 17.61 1.91 ;
      RECT 17.14 6.97 17.61 7.14 ;
      RECT 17.14 5.95 17.31 7.14 ;
      RECT 16.15 1.74 16.32 2.93 ;
      RECT 16.15 1.74 16.62 1.91 ;
      RECT 16.15 6.97 16.62 7.14 ;
      RECT 16.15 5.95 16.32 7.14 ;
      RECT 14.3 2.635 14.47 3.865 ;
      RECT 14.355 0.855 14.525 2.805 ;
      RECT 14.3 0.575 14.47 1.025 ;
      RECT 14.3 7.855 14.47 8.305 ;
      RECT 14.355 6.075 14.525 8.025 ;
      RECT 14.3 5.015 14.47 6.245 ;
      RECT 13.78 0.575 13.95 3.865 ;
      RECT 13.78 2.075 14.185 2.405 ;
      RECT 13.78 1.235 14.185 1.565 ;
      RECT 13.78 5.015 13.95 8.305 ;
      RECT 13.78 7.315 14.185 7.645 ;
      RECT 13.78 6.475 14.185 6.805 ;
      RECT 11.055 3.61 11.565 3.78 ;
      RECT 11.395 3.22 11.565 3.78 ;
      RECT 11.505 3.14 11.675 3.47 ;
      RECT 11.295 2.53 11.565 2.94 ;
      RECT 11.175 2.53 11.565 2.74 ;
      RECT 9.645 3.14 9.815 3.5 ;
      RECT 9.645 3.22 10.985 3.39 ;
      RECT 10.815 3.05 10.985 3.39 ;
      RECT 9.375 2.57 9.545 2.94 ;
      RECT 8.895 2.57 9.545 2.84 ;
      RECT 8.815 2.57 9.625 2.74 ;
      RECT 8.175 1.81 8.345 2.1 ;
      RECT 8.175 1.81 9.415 1.98 ;
      RECT 8.895 2.15 9.065 2.36 ;
      RECT 8.535 2.15 9.065 2.32 ;
      RECT 8.685 7.855 8.855 8.305 ;
      RECT 8.74 6.075 8.91 8.025 ;
      RECT 8.685 5.015 8.855 6.245 ;
      RECT 8.165 5.015 8.335 8.305 ;
      RECT 8.165 7.315 8.57 7.645 ;
      RECT 8.165 6.475 8.57 6.805 ;
      RECT 7.935 3.22 8.425 3.39 ;
      RECT 7.935 3.05 8.105 3.39 ;
      RECT 7.215 3.22 7.385 3.78 ;
      RECT 7.105 3.22 7.435 3.39 ;
      RECT 7.175 1.83 7.345 2.1 ;
      RECT 7.215 1.75 7.385 2.08 ;
      RECT 7.075 1.83 7.385 2.05 ;
      RECT 5.655 3.22 5.945 3.78 ;
      RECT 5.775 3.14 5.945 3.78 ;
      RECT 5.415 2.57 5.785 2.74 ;
      RECT 5.415 1.93 5.585 2.74 ;
      RECT 5.295 1.93 5.585 2.1 ;
      RECT 1.17 7.855 1.34 8.305 ;
      RECT 1.225 6.075 1.395 8.025 ;
      RECT 1.17 5.015 1.34 6.245 ;
      RECT 0.65 5.015 0.82 8.305 ;
      RECT 0.65 7.315 1.055 7.645 ;
      RECT 0.65 6.475 1.055 6.805 ;
      RECT 78.55 7.8 78.72 8.31 ;
      RECT 77.56 0.57 77.73 1.08 ;
      RECT 77.56 2.39 77.73 3.86 ;
      RECT 77.56 5.02 77.73 6.49 ;
      RECT 77.56 7.8 77.73 8.31 ;
      RECT 76.2 0.575 76.37 3.865 ;
      RECT 76.2 5.015 76.37 8.305 ;
      RECT 75.77 0.575 75.94 1.085 ;
      RECT 75.77 1.655 75.94 3.865 ;
      RECT 75.77 5.015 75.94 7.225 ;
      RECT 75.77 7.795 75.94 8.305 ;
      RECT 72.095 1.75 72.265 2.1 ;
      RECT 71.855 2.49 72.025 2.82 ;
      RECT 71.375 2.49 71.545 2.94 ;
      RECT 71.135 1.75 71.305 2.1 ;
      RECT 70.895 2.49 71.065 2.82 ;
      RECT 70.585 5.015 70.755 8.305 ;
      RECT 70.155 5.015 70.325 7.225 ;
      RECT 70.155 7.795 70.325 8.305 ;
      RECT 70.145 3.48 70.315 3.81 ;
      RECT 69.455 2.49 69.625 2.94 ;
      RECT 68.975 2.49 69.145 2.82 ;
      RECT 68.495 2.49 68.665 2.82 ;
      RECT 68.015 2.49 68.185 2.94 ;
      RECT 67.775 3.48 67.945 3.81 ;
      RECT 67.535 2.49 67.705 3.22 ;
      RECT 67.055 2.49 67.225 2.82 ;
      RECT 66.815 1.75 66.985 2.1 ;
      RECT 66.335 3.05 66.505 3.47 ;
      RECT 66.095 2.49 66.265 2.82 ;
      RECT 65.855 3.14 66.025 3.5 ;
      RECT 65.615 2.49 65.785 2.94 ;
      RECT 65.135 2.49 65.305 2.94 ;
      RECT 64.925 1.75 65.095 2.1 ;
      RECT 64.925 3.14 65.095 3.5 ;
      RECT 63.29 7.8 63.46 8.31 ;
      RECT 62.3 0.57 62.47 1.08 ;
      RECT 62.3 2.39 62.47 3.86 ;
      RECT 62.3 5.02 62.47 6.49 ;
      RECT 62.3 7.8 62.47 8.31 ;
      RECT 60.94 0.575 61.11 3.865 ;
      RECT 60.94 5.015 61.11 8.305 ;
      RECT 60.51 0.575 60.68 1.085 ;
      RECT 60.51 1.655 60.68 3.865 ;
      RECT 60.51 5.015 60.68 7.225 ;
      RECT 60.51 7.795 60.68 8.305 ;
      RECT 56.835 1.75 57.005 2.1 ;
      RECT 56.595 2.49 56.765 2.82 ;
      RECT 56.115 2.49 56.285 2.94 ;
      RECT 55.875 1.75 56.045 2.1 ;
      RECT 55.635 2.49 55.805 2.82 ;
      RECT 55.325 5.015 55.495 8.305 ;
      RECT 54.895 5.015 55.065 7.225 ;
      RECT 54.895 7.795 55.065 8.305 ;
      RECT 54.885 3.48 55.055 3.81 ;
      RECT 54.195 2.49 54.365 2.94 ;
      RECT 53.715 2.49 53.885 2.82 ;
      RECT 53.235 2.49 53.405 2.82 ;
      RECT 52.755 2.49 52.925 2.94 ;
      RECT 52.515 3.48 52.685 3.81 ;
      RECT 52.275 2.49 52.445 3.22 ;
      RECT 51.795 2.49 51.965 2.82 ;
      RECT 51.555 1.75 51.725 2.1 ;
      RECT 51.075 3.05 51.245 3.47 ;
      RECT 50.835 2.49 51.005 2.82 ;
      RECT 50.595 3.14 50.765 3.5 ;
      RECT 50.355 2.49 50.525 2.94 ;
      RECT 49.875 2.49 50.045 2.94 ;
      RECT 49.665 1.75 49.835 2.1 ;
      RECT 49.665 3.14 49.835 3.5 ;
      RECT 48.03 7.8 48.2 8.31 ;
      RECT 47.04 0.57 47.21 1.08 ;
      RECT 47.04 2.39 47.21 3.86 ;
      RECT 47.04 5.02 47.21 6.49 ;
      RECT 47.04 7.8 47.21 8.31 ;
      RECT 45.68 0.575 45.85 3.865 ;
      RECT 45.68 5.015 45.85 8.305 ;
      RECT 45.25 0.575 45.42 1.085 ;
      RECT 45.25 1.655 45.42 3.865 ;
      RECT 45.25 5.015 45.42 7.225 ;
      RECT 45.25 7.795 45.42 8.305 ;
      RECT 41.575 1.75 41.745 2.1 ;
      RECT 41.335 2.49 41.505 2.82 ;
      RECT 40.855 2.49 41.025 2.94 ;
      RECT 40.615 1.75 40.785 2.1 ;
      RECT 40.375 2.49 40.545 2.82 ;
      RECT 40.065 5.015 40.235 8.305 ;
      RECT 39.635 5.015 39.805 7.225 ;
      RECT 39.635 7.795 39.805 8.305 ;
      RECT 39.625 3.48 39.795 3.81 ;
      RECT 38.935 2.49 39.105 2.94 ;
      RECT 38.455 2.49 38.625 2.82 ;
      RECT 37.975 2.49 38.145 2.82 ;
      RECT 37.495 2.49 37.665 2.94 ;
      RECT 37.255 3.48 37.425 3.81 ;
      RECT 37.015 2.49 37.185 3.22 ;
      RECT 36.535 2.49 36.705 2.82 ;
      RECT 36.295 1.75 36.465 2.1 ;
      RECT 35.815 3.05 35.985 3.47 ;
      RECT 35.575 2.49 35.745 2.82 ;
      RECT 35.335 3.14 35.505 3.5 ;
      RECT 35.095 2.49 35.265 2.94 ;
      RECT 34.615 2.49 34.785 2.94 ;
      RECT 34.405 1.75 34.575 2.1 ;
      RECT 34.405 3.14 34.575 3.5 ;
      RECT 32.77 7.8 32.94 8.31 ;
      RECT 31.78 0.57 31.95 1.08 ;
      RECT 31.78 2.39 31.95 3.86 ;
      RECT 31.78 5.02 31.95 6.49 ;
      RECT 31.78 7.8 31.95 8.31 ;
      RECT 30.42 0.575 30.59 3.865 ;
      RECT 30.42 5.015 30.59 8.305 ;
      RECT 29.99 0.575 30.16 1.085 ;
      RECT 29.99 1.655 30.16 3.865 ;
      RECT 29.99 5.015 30.16 7.225 ;
      RECT 29.99 7.795 30.16 8.305 ;
      RECT 26.315 1.75 26.485 2.1 ;
      RECT 26.075 2.49 26.245 2.82 ;
      RECT 25.595 2.49 25.765 2.94 ;
      RECT 25.355 1.75 25.525 2.1 ;
      RECT 25.115 2.49 25.285 2.82 ;
      RECT 24.805 5.015 24.975 8.305 ;
      RECT 24.375 5.015 24.545 7.225 ;
      RECT 24.375 7.795 24.545 8.305 ;
      RECT 24.365 3.48 24.535 3.81 ;
      RECT 23.675 2.49 23.845 2.94 ;
      RECT 23.195 2.49 23.365 2.82 ;
      RECT 22.715 2.49 22.885 2.82 ;
      RECT 22.235 2.49 22.405 2.94 ;
      RECT 21.995 3.48 22.165 3.81 ;
      RECT 21.755 2.49 21.925 3.22 ;
      RECT 21.275 2.49 21.445 2.82 ;
      RECT 21.035 1.75 21.205 2.1 ;
      RECT 20.555 3.05 20.725 3.47 ;
      RECT 20.315 2.49 20.485 2.82 ;
      RECT 20.075 3.14 20.245 3.5 ;
      RECT 19.835 2.49 20.005 2.94 ;
      RECT 19.355 2.49 19.525 2.94 ;
      RECT 19.145 1.75 19.315 2.1 ;
      RECT 19.145 3.14 19.315 3.5 ;
      RECT 17.51 7.8 17.68 8.31 ;
      RECT 16.52 0.57 16.69 1.08 ;
      RECT 16.52 2.39 16.69 3.86 ;
      RECT 16.52 5.02 16.69 6.49 ;
      RECT 16.52 7.8 16.69 8.31 ;
      RECT 15.16 0.575 15.33 3.865 ;
      RECT 15.16 5.015 15.33 8.305 ;
      RECT 14.73 0.575 14.9 1.085 ;
      RECT 14.73 1.655 14.9 3.865 ;
      RECT 14.73 5.015 14.9 7.225 ;
      RECT 14.73 7.795 14.9 8.305 ;
      RECT 11.055 1.75 11.225 2.1 ;
      RECT 10.815 2.49 10.985 2.82 ;
      RECT 10.335 2.49 10.505 2.94 ;
      RECT 10.095 1.75 10.265 2.1 ;
      RECT 9.855 2.49 10.025 2.82 ;
      RECT 9.545 5.015 9.715 8.305 ;
      RECT 9.115 5.015 9.285 7.225 ;
      RECT 9.115 7.795 9.285 8.305 ;
      RECT 9.105 3.48 9.275 3.81 ;
      RECT 8.415 2.49 8.585 2.94 ;
      RECT 7.935 2.49 8.105 2.82 ;
      RECT 7.455 2.49 7.625 2.82 ;
      RECT 6.975 2.49 7.145 2.94 ;
      RECT 6.735 3.48 6.905 3.81 ;
      RECT 6.495 2.49 6.665 3.22 ;
      RECT 6.015 2.49 6.185 2.82 ;
      RECT 5.775 1.75 5.945 2.1 ;
      RECT 5.295 3.05 5.465 3.47 ;
      RECT 5.055 2.49 5.225 2.82 ;
      RECT 4.815 3.14 4.985 3.5 ;
      RECT 4.575 2.49 4.745 2.94 ;
      RECT 4.095 2.49 4.265 2.94 ;
      RECT 3.885 1.75 4.055 2.1 ;
      RECT 3.885 3.14 4.055 3.5 ;
      RECT 1.6 5.015 1.77 7.225 ;
      RECT 1.6 7.795 1.77 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8_b0r1 ;
  SIZE 79.095 BY 8.89 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 17.515 0.915 17.685 1.085 ;
        RECT 17.51 0.91 17.68 1.08 ;
        RECT 17.51 2.39 17.68 2.56 ;
      LAYER li1 ;
        RECT 17.515 0.915 17.685 1.085 ;
        RECT 17.51 0.57 17.68 1.08 ;
        RECT 17.51 2.39 17.68 3.86 ;
      LAYER met1 ;
        RECT 17.45 2.36 17.74 2.59 ;
        RECT 17.45 0.88 17.74 1.11 ;
        RECT 17.51 0.88 17.68 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 32.775 0.915 32.945 1.085 ;
        RECT 32.77 0.91 32.94 1.08 ;
        RECT 32.77 2.39 32.94 2.56 ;
      LAYER li1 ;
        RECT 32.775 0.915 32.945 1.085 ;
        RECT 32.77 0.57 32.94 1.08 ;
        RECT 32.77 2.39 32.94 3.86 ;
      LAYER met1 ;
        RECT 32.71 2.36 33 2.59 ;
        RECT 32.71 0.88 33 1.11 ;
        RECT 32.77 0.88 32.94 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 48.035 0.915 48.205 1.085 ;
        RECT 48.03 0.91 48.2 1.08 ;
        RECT 48.03 2.39 48.2 2.56 ;
      LAYER li1 ;
        RECT 48.035 0.915 48.205 1.085 ;
        RECT 48.03 0.57 48.2 1.08 ;
        RECT 48.03 2.39 48.2 3.86 ;
      LAYER met1 ;
        RECT 47.97 2.36 48.26 2.59 ;
        RECT 47.97 0.88 48.26 1.11 ;
        RECT 48.03 0.88 48.2 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 63.295 0.915 63.465 1.085 ;
        RECT 63.29 0.91 63.46 1.08 ;
        RECT 63.29 2.39 63.46 2.56 ;
      LAYER li1 ;
        RECT 63.295 0.915 63.465 1.085 ;
        RECT 63.29 0.57 63.46 1.08 ;
        RECT 63.29 2.39 63.46 3.86 ;
      LAYER met1 ;
        RECT 63.23 2.36 63.52 2.59 ;
        RECT 63.23 0.88 63.52 1.11 ;
        RECT 63.29 0.88 63.46 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 78.555 0.915 78.725 1.085 ;
        RECT 78.55 0.91 78.72 1.08 ;
        RECT 78.55 2.39 78.72 2.56 ;
      LAYER li1 ;
        RECT 78.555 0.915 78.725 1.085 ;
        RECT 78.55 0.57 78.72 1.08 ;
        RECT 78.55 2.39 78.72 3.86 ;
      LAYER met1 ;
        RECT 78.49 2.36 78.78 2.59 ;
        RECT 78.49 0.88 78.78 1.11 ;
        RECT 78.55 0.88 78.72 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 13.28 2.705 13.62 3.055 ;
        RECT 13.275 5.86 13.615 6.21 ;
        RECT 13.355 2.705 13.53 6.21 ;
      LAYER li1 ;
        RECT 13.36 1.66 13.53 2.935 ;
        RECT 13.36 5.945 13.53 7.22 ;
        RECT 7.725 5.945 7.895 7.22 ;
      LAYER met1 ;
        RECT 13.28 2.765 13.76 2.935 ;
        RECT 13.28 2.705 13.62 3.055 ;
        RECT 7.665 5.945 13.76 6.115 ;
        RECT 13.275 5.86 13.615 6.21 ;
        RECT 7.665 5.915 7.955 6.145 ;
      LAYER mcon ;
        RECT 7.725 5.945 7.895 6.115 ;
        RECT 13.36 5.945 13.53 6.115 ;
        RECT 13.36 2.765 13.53 2.935 ;
      LAYER via1 ;
        RECT 13.375 5.96 13.525 6.11 ;
        RECT 13.38 2.805 13.53 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 28.54 2.705 28.88 3.055 ;
        RECT 28.535 5.86 28.875 6.21 ;
        RECT 28.615 2.705 28.79 6.21 ;
      LAYER li1 ;
        RECT 28.62 1.66 28.79 2.935 ;
        RECT 28.62 5.945 28.79 7.22 ;
        RECT 22.985 5.945 23.155 7.22 ;
      LAYER met1 ;
        RECT 28.54 2.765 29.02 2.935 ;
        RECT 28.54 2.705 28.88 3.055 ;
        RECT 22.925 5.945 29.02 6.115 ;
        RECT 28.535 5.86 28.875 6.21 ;
        RECT 22.925 5.915 23.215 6.145 ;
      LAYER mcon ;
        RECT 22.985 5.945 23.155 6.115 ;
        RECT 28.62 5.945 28.79 6.115 ;
        RECT 28.62 2.765 28.79 2.935 ;
      LAYER via1 ;
        RECT 28.635 5.96 28.785 6.11 ;
        RECT 28.64 2.805 28.79 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 43.8 2.705 44.14 3.055 ;
        RECT 43.795 5.86 44.135 6.21 ;
        RECT 43.875 2.705 44.05 6.21 ;
      LAYER li1 ;
        RECT 43.88 1.66 44.05 2.935 ;
        RECT 43.88 5.945 44.05 7.22 ;
        RECT 38.245 5.945 38.415 7.22 ;
      LAYER met1 ;
        RECT 43.8 2.765 44.28 2.935 ;
        RECT 43.8 2.705 44.14 3.055 ;
        RECT 38.185 5.945 44.28 6.115 ;
        RECT 43.795 5.86 44.135 6.21 ;
        RECT 38.185 5.915 38.475 6.145 ;
      LAYER mcon ;
        RECT 38.245 5.945 38.415 6.115 ;
        RECT 43.88 5.945 44.05 6.115 ;
        RECT 43.88 2.765 44.05 2.935 ;
      LAYER via1 ;
        RECT 43.895 5.96 44.045 6.11 ;
        RECT 43.9 2.805 44.05 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 59.06 2.705 59.4 3.055 ;
        RECT 59.055 5.86 59.395 6.21 ;
        RECT 59.135 2.705 59.31 6.21 ;
      LAYER li1 ;
        RECT 59.14 1.66 59.31 2.935 ;
        RECT 59.14 5.945 59.31 7.22 ;
        RECT 53.505 5.945 53.675 7.22 ;
      LAYER met1 ;
        RECT 59.06 2.765 59.54 2.935 ;
        RECT 59.06 2.705 59.4 3.055 ;
        RECT 53.445 5.945 59.54 6.115 ;
        RECT 59.055 5.86 59.395 6.21 ;
        RECT 53.445 5.915 53.735 6.145 ;
      LAYER mcon ;
        RECT 53.505 5.945 53.675 6.115 ;
        RECT 59.14 5.945 59.31 6.115 ;
        RECT 59.14 2.765 59.31 2.935 ;
      LAYER via1 ;
        RECT 59.155 5.96 59.305 6.11 ;
        RECT 59.16 2.805 59.31 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 74.32 2.705 74.66 3.055 ;
        RECT 74.315 5.86 74.655 6.21 ;
        RECT 74.395 2.705 74.57 6.21 ;
      LAYER li1 ;
        RECT 74.4 1.66 74.57 2.935 ;
        RECT 74.4 5.945 74.57 7.22 ;
        RECT 68.765 5.945 68.935 7.22 ;
      LAYER met1 ;
        RECT 74.32 2.765 74.8 2.935 ;
        RECT 74.32 2.705 74.66 3.055 ;
        RECT 68.705 5.945 74.8 6.115 ;
        RECT 74.315 5.86 74.655 6.21 ;
        RECT 68.705 5.915 68.995 6.145 ;
      LAYER mcon ;
        RECT 68.765 5.945 68.935 6.115 ;
        RECT 74.4 5.945 74.57 6.115 ;
        RECT 74.4 2.765 74.57 2.935 ;
      LAYER via1 ;
        RECT 74.415 5.96 74.565 6.11 ;
        RECT 74.42 2.805 74.57 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 5.945 0.4 7.22 ;
      LAYER met1 ;
        RECT 0.17 5.945 0.63 6.115 ;
        RECT 0.17 5.915 0.46 6.145 ;
      LAYER mcon ;
        RECT 0.23 5.945 0.4 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.385 4.265 2.19 4.645 ;
      LAYER met2 ;
        RECT 1.575 4.265 1.955 4.645 ;
      LAYER li1 ;
        RECT 0 4.44 79.095 4.745 ;
        RECT 64.585 4.135 79.095 4.745 ;
        RECT 76.96 4.13 78.94 4.75 ;
        RECT 78.12 3.4 78.29 5.48 ;
        RECT 77.13 3.4 77.3 5.48 ;
        RECT 74.39 3.405 74.56 5.475 ;
        RECT 71.615 3.635 71.785 4.745 ;
        RECT 69.695 3.635 69.865 4.745 ;
        RECT 68.755 3.635 68.925 5.475 ;
        RECT 67.295 3.635 67.465 4.745 ;
        RECT 65.375 3.635 65.545 4.745 ;
        RECT 1.85 4.14 79.095 4.745 ;
        RECT 49.325 4.135 63.835 4.745 ;
        RECT 61.7 4.13 63.68 4.75 ;
        RECT 62.86 3.4 63.03 5.48 ;
        RECT 61.87 3.4 62.04 5.48 ;
        RECT 59.13 3.405 59.3 5.475 ;
        RECT 56.355 3.635 56.525 4.745 ;
        RECT 54.435 3.635 54.605 4.745 ;
        RECT 53.495 3.635 53.665 5.475 ;
        RECT 52.035 3.635 52.205 4.745 ;
        RECT 50.115 3.635 50.285 4.745 ;
        RECT 34.065 4.135 48.575 4.745 ;
        RECT 46.44 4.13 48.42 4.75 ;
        RECT 47.6 3.4 47.77 5.48 ;
        RECT 46.61 3.4 46.78 5.48 ;
        RECT 43.87 3.405 44.04 5.475 ;
        RECT 41.095 3.635 41.265 4.745 ;
        RECT 39.175 3.635 39.345 4.745 ;
        RECT 38.235 3.635 38.405 5.475 ;
        RECT 36.775 3.635 36.945 4.745 ;
        RECT 34.855 3.635 35.025 4.745 ;
        RECT 18.805 4.135 33.315 4.745 ;
        RECT 31.18 4.13 33.16 4.75 ;
        RECT 32.34 3.4 32.51 5.48 ;
        RECT 31.35 3.4 31.52 5.48 ;
        RECT 28.61 3.405 28.78 5.475 ;
        RECT 25.835 3.635 26.005 4.745 ;
        RECT 23.915 3.635 24.085 4.745 ;
        RECT 22.975 3.635 23.145 5.475 ;
        RECT 21.515 3.635 21.685 4.745 ;
        RECT 19.595 3.635 19.765 4.745 ;
        RECT 3.545 4.135 18.055 4.745 ;
        RECT 15.92 4.13 17.9 4.75 ;
        RECT 17.08 3.4 17.25 5.48 ;
        RECT 16.09 3.4 16.26 5.48 ;
        RECT 13.35 3.405 13.52 5.475 ;
        RECT 10.575 3.635 10.745 4.745 ;
        RECT 8.655 3.635 8.825 4.745 ;
        RECT 7.715 3.635 7.885 5.475 ;
        RECT 6.255 3.635 6.425 4.745 ;
        RECT 4.335 3.635 4.505 4.745 ;
        RECT 2.03 4.14 2.2 8.305 ;
        RECT 0 4.14 79.095 4.34 ;
        RECT 0 4.14 1.68 4.745 ;
        RECT 0.22 4.14 0.39 5.475 ;
      LAYER met1 ;
        RECT 0 4.14 79.095 4.745 ;
        RECT 64.585 4.135 79.095 4.745 ;
        RECT 76.96 4.13 78.94 4.75 ;
        RECT 64.585 3.98 73.325 4.745 ;
        RECT 49.325 4.135 63.835 4.745 ;
        RECT 61.7 4.13 63.68 4.75 ;
        RECT 49.325 3.98 58.065 4.745 ;
        RECT 34.065 4.135 48.575 4.745 ;
        RECT 46.44 4.13 48.42 4.75 ;
        RECT 34.065 3.98 42.805 4.745 ;
        RECT 18.805 4.135 33.315 4.745 ;
        RECT 31.18 4.13 33.16 4.75 ;
        RECT 18.805 3.98 27.545 4.745 ;
        RECT 3.545 4.135 18.055 4.745 ;
        RECT 15.92 4.13 17.9 4.75 ;
        RECT 3.545 3.98 12.285 4.745 ;
        RECT 1.97 6.655 2.26 6.885 ;
        RECT 1.8 6.685 2.26 6.855 ;
      LAYER via2 ;
        RECT 1.665 4.355 1.865 4.555 ;
      LAYER mcon ;
        RECT 2.03 6.685 2.2 6.855 ;
        RECT 2.34 4.545 2.51 4.715 ;
        RECT 3.69 4.135 3.86 4.305 ;
        RECT 4.15 4.135 4.32 4.305 ;
        RECT 4.61 4.135 4.78 4.305 ;
        RECT 5.07 4.135 5.24 4.305 ;
        RECT 5.53 4.135 5.7 4.305 ;
        RECT 5.99 4.135 6.16 4.305 ;
        RECT 6.45 4.135 6.62 4.305 ;
        RECT 6.91 4.135 7.08 4.305 ;
        RECT 7.37 4.135 7.54 4.305 ;
        RECT 7.83 4.135 8 4.305 ;
        RECT 8.29 4.135 8.46 4.305 ;
        RECT 8.75 4.135 8.92 4.305 ;
        RECT 9.21 4.135 9.38 4.305 ;
        RECT 9.67 4.135 9.84 4.305 ;
        RECT 9.835 4.545 10.005 4.715 ;
        RECT 10.13 4.135 10.3 4.305 ;
        RECT 10.59 4.135 10.76 4.305 ;
        RECT 11.05 4.135 11.22 4.305 ;
        RECT 11.51 4.135 11.68 4.305 ;
        RECT 11.97 4.135 12.14 4.305 ;
        RECT 15.47 4.545 15.64 4.715 ;
        RECT 15.47 4.165 15.64 4.335 ;
        RECT 16.17 4.55 16.34 4.72 ;
        RECT 16.17 4.16 16.34 4.33 ;
        RECT 17.16 4.55 17.33 4.72 ;
        RECT 17.16 4.16 17.33 4.33 ;
        RECT 18.95 4.135 19.12 4.305 ;
        RECT 19.41 4.135 19.58 4.305 ;
        RECT 19.87 4.135 20.04 4.305 ;
        RECT 20.33 4.135 20.5 4.305 ;
        RECT 20.79 4.135 20.96 4.305 ;
        RECT 21.25 4.135 21.42 4.305 ;
        RECT 21.71 4.135 21.88 4.305 ;
        RECT 22.17 4.135 22.34 4.305 ;
        RECT 22.63 4.135 22.8 4.305 ;
        RECT 23.09 4.135 23.26 4.305 ;
        RECT 23.55 4.135 23.72 4.305 ;
        RECT 24.01 4.135 24.18 4.305 ;
        RECT 24.47 4.135 24.64 4.305 ;
        RECT 24.93 4.135 25.1 4.305 ;
        RECT 25.095 4.545 25.265 4.715 ;
        RECT 25.39 4.135 25.56 4.305 ;
        RECT 25.85 4.135 26.02 4.305 ;
        RECT 26.31 4.135 26.48 4.305 ;
        RECT 26.77 4.135 26.94 4.305 ;
        RECT 27.23 4.135 27.4 4.305 ;
        RECT 30.73 4.545 30.9 4.715 ;
        RECT 30.73 4.165 30.9 4.335 ;
        RECT 31.43 4.55 31.6 4.72 ;
        RECT 31.43 4.16 31.6 4.33 ;
        RECT 32.42 4.55 32.59 4.72 ;
        RECT 32.42 4.16 32.59 4.33 ;
        RECT 34.21 4.135 34.38 4.305 ;
        RECT 34.67 4.135 34.84 4.305 ;
        RECT 35.13 4.135 35.3 4.305 ;
        RECT 35.59 4.135 35.76 4.305 ;
        RECT 36.05 4.135 36.22 4.305 ;
        RECT 36.51 4.135 36.68 4.305 ;
        RECT 36.97 4.135 37.14 4.305 ;
        RECT 37.43 4.135 37.6 4.305 ;
        RECT 37.89 4.135 38.06 4.305 ;
        RECT 38.35 4.135 38.52 4.305 ;
        RECT 38.81 4.135 38.98 4.305 ;
        RECT 39.27 4.135 39.44 4.305 ;
        RECT 39.73 4.135 39.9 4.305 ;
        RECT 40.19 4.135 40.36 4.305 ;
        RECT 40.355 4.545 40.525 4.715 ;
        RECT 40.65 4.135 40.82 4.305 ;
        RECT 41.11 4.135 41.28 4.305 ;
        RECT 41.57 4.135 41.74 4.305 ;
        RECT 42.03 4.135 42.2 4.305 ;
        RECT 42.49 4.135 42.66 4.305 ;
        RECT 45.99 4.545 46.16 4.715 ;
        RECT 45.99 4.165 46.16 4.335 ;
        RECT 46.69 4.55 46.86 4.72 ;
        RECT 46.69 4.16 46.86 4.33 ;
        RECT 47.68 4.55 47.85 4.72 ;
        RECT 47.68 4.16 47.85 4.33 ;
        RECT 49.47 4.135 49.64 4.305 ;
        RECT 49.93 4.135 50.1 4.305 ;
        RECT 50.39 4.135 50.56 4.305 ;
        RECT 50.85 4.135 51.02 4.305 ;
        RECT 51.31 4.135 51.48 4.305 ;
        RECT 51.77 4.135 51.94 4.305 ;
        RECT 52.23 4.135 52.4 4.305 ;
        RECT 52.69 4.135 52.86 4.305 ;
        RECT 53.15 4.135 53.32 4.305 ;
        RECT 53.61 4.135 53.78 4.305 ;
        RECT 54.07 4.135 54.24 4.305 ;
        RECT 54.53 4.135 54.7 4.305 ;
        RECT 54.99 4.135 55.16 4.305 ;
        RECT 55.45 4.135 55.62 4.305 ;
        RECT 55.615 4.545 55.785 4.715 ;
        RECT 55.91 4.135 56.08 4.305 ;
        RECT 56.37 4.135 56.54 4.305 ;
        RECT 56.83 4.135 57 4.305 ;
        RECT 57.29 4.135 57.46 4.305 ;
        RECT 57.75 4.135 57.92 4.305 ;
        RECT 61.25 4.545 61.42 4.715 ;
        RECT 61.25 4.165 61.42 4.335 ;
        RECT 61.95 4.55 62.12 4.72 ;
        RECT 61.95 4.16 62.12 4.33 ;
        RECT 62.94 4.55 63.11 4.72 ;
        RECT 62.94 4.16 63.11 4.33 ;
        RECT 64.73 4.135 64.9 4.305 ;
        RECT 65.19 4.135 65.36 4.305 ;
        RECT 65.65 4.135 65.82 4.305 ;
        RECT 66.11 4.135 66.28 4.305 ;
        RECT 66.57 4.135 66.74 4.305 ;
        RECT 67.03 4.135 67.2 4.305 ;
        RECT 67.49 4.135 67.66 4.305 ;
        RECT 67.95 4.135 68.12 4.305 ;
        RECT 68.41 4.135 68.58 4.305 ;
        RECT 68.87 4.135 69.04 4.305 ;
        RECT 69.33 4.135 69.5 4.305 ;
        RECT 69.79 4.135 69.96 4.305 ;
        RECT 70.25 4.135 70.42 4.305 ;
        RECT 70.71 4.135 70.88 4.305 ;
        RECT 70.875 4.545 71.045 4.715 ;
        RECT 71.17 4.135 71.34 4.305 ;
        RECT 71.63 4.135 71.8 4.305 ;
        RECT 72.09 4.135 72.26 4.305 ;
        RECT 72.55 4.135 72.72 4.305 ;
        RECT 73.01 4.135 73.18 4.305 ;
        RECT 76.51 4.545 76.68 4.715 ;
        RECT 76.51 4.165 76.68 4.335 ;
        RECT 77.21 4.55 77.38 4.72 ;
        RECT 77.21 4.16 77.38 4.33 ;
        RECT 78.2 4.55 78.37 4.72 ;
        RECT 78.2 4.16 78.37 4.33 ;
      LAYER via1 ;
        RECT 1.69 4.38 1.84 4.53 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 70.035 7.055 70.405 7.425 ;
      RECT 70.07 4.27 70.37 7.425 ;
      RECT 65.88 4.27 70.37 4.57 ;
      RECT 69.06 1.855 69.36 4.57 ;
      RECT 65.88 2.435 66.18 4.57 ;
      RECT 69.015 2.76 69.36 3.49 ;
      RECT 65.775 2.015 66.105 2.745 ;
      RECT 68.655 1.855 69.385 2.185 ;
      RECT 54.775 7.055 55.145 7.425 ;
      RECT 54.81 4.27 55.11 7.425 ;
      RECT 50.62 4.27 55.11 4.57 ;
      RECT 53.8 1.855 54.1 4.57 ;
      RECT 50.62 2.435 50.92 4.57 ;
      RECT 53.755 2.76 54.1 3.49 ;
      RECT 50.515 2.015 50.845 2.745 ;
      RECT 53.395 1.855 54.125 2.185 ;
      RECT 39.515 7.055 39.885 7.425 ;
      RECT 39.55 4.27 39.85 7.425 ;
      RECT 35.36 4.27 39.85 4.57 ;
      RECT 38.54 1.855 38.84 4.57 ;
      RECT 35.36 2.435 35.66 4.57 ;
      RECT 38.495 2.76 38.84 3.49 ;
      RECT 35.255 2.015 35.585 2.745 ;
      RECT 38.135 1.855 38.865 2.185 ;
      RECT 24.255 7.055 24.625 7.425 ;
      RECT 24.29 4.27 24.59 7.425 ;
      RECT 20.1 4.27 24.59 4.57 ;
      RECT 23.28 1.855 23.58 4.57 ;
      RECT 20.1 2.435 20.4 4.57 ;
      RECT 23.235 2.76 23.58 3.49 ;
      RECT 19.995 2.015 20.325 2.745 ;
      RECT 22.875 1.855 23.605 2.185 ;
      RECT 8.995 7.055 9.365 7.425 ;
      RECT 9.03 4.27 9.33 7.425 ;
      RECT 4.84 4.27 9.33 4.57 ;
      RECT 8.02 1.855 8.32 4.57 ;
      RECT 4.84 2.435 5.14 4.57 ;
      RECT 7.975 2.76 8.32 3.49 ;
      RECT 4.735 2.015 5.065 2.745 ;
      RECT 7.615 1.855 8.345 2.185 ;
      RECT 72.135 2.015 72.465 2.745 ;
      RECT 70.935 2.88 71.265 3.61 ;
      RECT 70.095 1.855 70.825 2.185 ;
      RECT 67.695 1.855 68.025 2.585 ;
      RECT 66.495 2.015 66.825 2.745 ;
      RECT 56.875 2.015 57.205 2.745 ;
      RECT 55.675 2.88 56.005 3.61 ;
      RECT 54.835 1.855 55.565 2.185 ;
      RECT 52.435 1.855 52.765 2.585 ;
      RECT 51.235 2.015 51.565 2.745 ;
      RECT 41.615 2.015 41.945 2.745 ;
      RECT 40.415 2.88 40.745 3.61 ;
      RECT 39.575 1.855 40.305 2.185 ;
      RECT 37.175 1.855 37.505 2.585 ;
      RECT 35.975 2.015 36.305 2.745 ;
      RECT 26.355 2.015 26.685 2.745 ;
      RECT 25.155 2.88 25.485 3.61 ;
      RECT 24.315 1.855 25.045 2.185 ;
      RECT 21.915 1.855 22.245 2.585 ;
      RECT 20.715 2.015 21.045 2.745 ;
      RECT 11.095 2.015 11.425 2.745 ;
      RECT 9.895 2.88 10.225 3.61 ;
      RECT 9.055 1.855 9.785 2.185 ;
      RECT 6.655 1.855 6.985 2.585 ;
      RECT 5.455 2.015 5.785 2.745 ;
      RECT 0.005 8.51 0.81 8.89 ;
    LAYER via2 ;
      RECT 72.2 2.48 72.4 2.68 ;
      RECT 71 3.04 71.2 3.24 ;
      RECT 70.16 1.92 70.36 2.12 ;
      RECT 70.12 7.14 70.32 7.34 ;
      RECT 69.08 2.825 69.28 3.025 ;
      RECT 68.72 1.92 68.92 2.12 ;
      RECT 67.76 1.92 67.96 2.12 ;
      RECT 66.56 2.48 66.76 2.68 ;
      RECT 65.84 2.48 66.04 2.68 ;
      RECT 56.94 2.48 57.14 2.68 ;
      RECT 55.74 3.04 55.94 3.24 ;
      RECT 54.9 1.92 55.1 2.12 ;
      RECT 54.86 7.14 55.06 7.34 ;
      RECT 53.82 2.825 54.02 3.025 ;
      RECT 53.46 1.92 53.66 2.12 ;
      RECT 52.5 1.92 52.7 2.12 ;
      RECT 51.3 2.48 51.5 2.68 ;
      RECT 50.58 2.48 50.78 2.68 ;
      RECT 41.68 2.48 41.88 2.68 ;
      RECT 40.48 3.04 40.68 3.24 ;
      RECT 39.64 1.92 39.84 2.12 ;
      RECT 39.6 7.14 39.8 7.34 ;
      RECT 38.56 2.825 38.76 3.025 ;
      RECT 38.2 1.92 38.4 2.12 ;
      RECT 37.24 1.92 37.44 2.12 ;
      RECT 36.04 2.48 36.24 2.68 ;
      RECT 35.32 2.48 35.52 2.68 ;
      RECT 26.42 2.48 26.62 2.68 ;
      RECT 25.22 3.04 25.42 3.24 ;
      RECT 24.38 1.92 24.58 2.12 ;
      RECT 24.34 7.14 24.54 7.34 ;
      RECT 23.3 2.825 23.5 3.025 ;
      RECT 22.94 1.92 23.14 2.12 ;
      RECT 21.98 1.92 22.18 2.12 ;
      RECT 20.78 2.48 20.98 2.68 ;
      RECT 20.06 2.48 20.26 2.68 ;
      RECT 11.16 2.48 11.36 2.68 ;
      RECT 9.96 3.04 10.16 3.24 ;
      RECT 9.12 1.92 9.32 2.12 ;
      RECT 9.08 7.14 9.28 7.34 ;
      RECT 8.04 2.825 8.24 3.025 ;
      RECT 7.68 1.92 7.88 2.12 ;
      RECT 6.72 1.92 6.92 2.12 ;
      RECT 5.52 2.48 5.72 2.68 ;
      RECT 4.8 2.48 5 2.68 ;
      RECT 0.285 8.6 0.485 8.8 ;
    LAYER met2 ;
      RECT 1.23 8.4 78.725 8.57 ;
      RECT 78.555 7.275 78.725 8.57 ;
      RECT 1.23 6.255 1.4 8.57 ;
      RECT 78.525 7.275 78.875 7.625 ;
      RECT 1.165 6.255 1.455 6.605 ;
      RECT 75.365 6.22 75.685 6.545 ;
      RECT 75.395 5.695 75.565 6.545 ;
      RECT 75.395 5.695 75.57 6.045 ;
      RECT 75.395 5.695 76.37 5.87 ;
      RECT 76.195 1.965 76.37 5.87 ;
      RECT 76.14 1.965 76.49 2.315 ;
      RECT 76.165 6.655 76.49 6.98 ;
      RECT 75.05 6.745 76.49 6.915 ;
      RECT 75.05 2.395 75.21 6.915 ;
      RECT 75.365 2.365 75.685 2.685 ;
      RECT 75.05 2.395 75.685 2.565 ;
      RECT 73.76 2.705 74.1 3.055 ;
      RECT 73.155 2.77 74.1 2.97 ;
      RECT 73.155 2.765 73.37 2.97 ;
      RECT 73.17 2.34 73.37 2.97 ;
      RECT 72.16 2.34 72.44 2.72 ;
      RECT 73.85 2.7 74.02 3.055 ;
      RECT 72.155 2.34 72.44 2.673 ;
      RECT 72.135 2.34 72.44 2.65 ;
      RECT 72.125 2.34 72.44 2.63 ;
      RECT 72.115 2.34 72.44 2.615 ;
      RECT 72.09 2.34 72.44 2.588 ;
      RECT 72.08 2.34 72.44 2.563 ;
      RECT 72.035 2.295 72.315 2.555 ;
      RECT 72.035 2.34 73.37 2.54 ;
      RECT 72.035 2.335 72.36 2.555 ;
      RECT 72.035 2.327 72.355 2.555 ;
      RECT 72.035 2.317 72.35 2.555 ;
      RECT 72.035 2.305 72.345 2.555 ;
      RECT 70.96 3 71.24 3.28 ;
      RECT 70.96 3 71.275 3.26 ;
      RECT 63.24 6.655 63.59 7.005 ;
      RECT 70.705 6.61 71.055 6.96 ;
      RECT 63.24 6.685 71.055 6.885 ;
      RECT 70.995 2.42 71.045 2.68 ;
      RECT 70.785 2.42 70.79 2.68 ;
      RECT 69.98 1.975 70.01 2.235 ;
      RECT 69.75 1.975 69.825 2.235 ;
      RECT 70.97 2.37 70.995 2.68 ;
      RECT 70.965 2.327 70.97 2.68 ;
      RECT 70.96 2.31 70.965 2.68 ;
      RECT 70.955 2.297 70.96 2.68 ;
      RECT 70.88 2.18 70.955 2.68 ;
      RECT 70.835 1.997 70.88 2.68 ;
      RECT 70.83 1.925 70.835 2.68 ;
      RECT 70.815 1.9 70.83 2.68 ;
      RECT 70.79 1.862 70.815 2.68 ;
      RECT 70.78 1.842 70.79 2.402 ;
      RECT 70.765 1.834 70.78 2.357 ;
      RECT 70.76 1.826 70.765 2.328 ;
      RECT 70.755 1.823 70.76 2.308 ;
      RECT 70.75 1.82 70.755 2.288 ;
      RECT 70.745 1.817 70.75 2.268 ;
      RECT 70.715 1.806 70.745 2.205 ;
      RECT 70.695 1.791 70.715 2.12 ;
      RECT 70.69 1.783 70.695 2.083 ;
      RECT 70.68 1.777 70.69 2.05 ;
      RECT 70.665 1.769 70.68 2.01 ;
      RECT 70.66 1.762 70.665 1.97 ;
      RECT 70.655 1.759 70.66 1.948 ;
      RECT 70.65 1.756 70.655 1.935 ;
      RECT 70.645 1.755 70.65 1.925 ;
      RECT 70.63 1.749 70.645 1.915 ;
      RECT 70.605 1.736 70.63 1.9 ;
      RECT 70.555 1.711 70.605 1.871 ;
      RECT 70.54 1.69 70.555 1.846 ;
      RECT 70.53 1.683 70.54 1.835 ;
      RECT 70.475 1.664 70.53 1.808 ;
      RECT 70.45 1.642 70.475 1.781 ;
      RECT 70.445 1.635 70.45 1.776 ;
      RECT 70.43 1.635 70.445 1.774 ;
      RECT 70.405 1.627 70.43 1.77 ;
      RECT 70.39 1.625 70.405 1.766 ;
      RECT 70.36 1.625 70.39 1.763 ;
      RECT 70.35 1.625 70.36 1.758 ;
      RECT 70.305 1.625 70.35 1.756 ;
      RECT 70.276 1.625 70.305 1.757 ;
      RECT 70.19 1.625 70.276 1.759 ;
      RECT 70.176 1.626 70.19 1.761 ;
      RECT 70.09 1.627 70.176 1.763 ;
      RECT 70.075 1.628 70.09 1.773 ;
      RECT 70.07 1.629 70.075 1.782 ;
      RECT 70.05 1.632 70.07 1.792 ;
      RECT 70.035 1.64 70.05 1.807 ;
      RECT 70.015 1.658 70.035 1.822 ;
      RECT 70.005 1.67 70.015 1.845 ;
      RECT 69.995 1.679 70.005 1.875 ;
      RECT 69.98 1.691 69.995 1.92 ;
      RECT 69.925 1.724 69.98 2.235 ;
      RECT 69.92 1.752 69.925 2.235 ;
      RECT 69.9 1.767 69.92 2.235 ;
      RECT 69.865 1.827 69.9 2.235 ;
      RECT 69.863 1.877 69.865 2.235 ;
      RECT 69.86 1.885 69.863 2.235 ;
      RECT 69.85 1.9 69.86 2.235 ;
      RECT 69.845 1.912 69.85 2.235 ;
      RECT 69.835 1.937 69.845 2.235 ;
      RECT 69.825 1.965 69.835 2.235 ;
      RECT 67.73 3.47 67.78 3.73 ;
      RECT 70.64 3.02 70.7 3.28 ;
      RECT 70.625 3.02 70.64 3.29 ;
      RECT 70.606 3.02 70.625 3.323 ;
      RECT 70.52 3.02 70.606 3.448 ;
      RECT 70.44 3.02 70.52 3.63 ;
      RECT 70.435 3.257 70.44 3.715 ;
      RECT 70.41 3.327 70.435 3.743 ;
      RECT 70.405 3.397 70.41 3.77 ;
      RECT 70.385 3.469 70.405 3.792 ;
      RECT 70.38 3.536 70.385 3.815 ;
      RECT 70.37 3.565 70.38 3.83 ;
      RECT 70.36 3.587 70.37 3.847 ;
      RECT 70.355 3.597 70.36 3.858 ;
      RECT 70.35 3.605 70.355 3.866 ;
      RECT 70.34 3.613 70.35 3.878 ;
      RECT 70.335 3.625 70.34 3.888 ;
      RECT 70.33 3.633 70.335 3.893 ;
      RECT 70.31 3.651 70.33 3.903 ;
      RECT 70.305 3.668 70.31 3.91 ;
      RECT 70.3 3.676 70.305 3.911 ;
      RECT 70.295 3.687 70.3 3.913 ;
      RECT 70.255 3.725 70.295 3.923 ;
      RECT 70.25 3.76 70.255 3.934 ;
      RECT 70.245 3.765 70.25 3.937 ;
      RECT 70.22 3.775 70.245 3.944 ;
      RECT 70.21 3.789 70.22 3.953 ;
      RECT 70.19 3.801 70.21 3.956 ;
      RECT 70.14 3.82 70.19 3.96 ;
      RECT 70.095 3.835 70.14 3.965 ;
      RECT 70.03 3.838 70.095 3.971 ;
      RECT 70.015 3.836 70.03 3.978 ;
      RECT 69.985 3.835 70.015 3.978 ;
      RECT 69.946 3.834 69.985 3.974 ;
      RECT 69.86 3.831 69.946 3.97 ;
      RECT 69.843 3.829 69.86 3.967 ;
      RECT 69.757 3.827 69.843 3.964 ;
      RECT 69.671 3.824 69.757 3.958 ;
      RECT 69.585 3.82 69.671 3.953 ;
      RECT 69.507 3.817 69.585 3.949 ;
      RECT 69.421 3.814 69.507 3.947 ;
      RECT 69.335 3.811 69.421 3.944 ;
      RECT 69.277 3.809 69.335 3.941 ;
      RECT 69.191 3.806 69.277 3.939 ;
      RECT 69.105 3.802 69.191 3.937 ;
      RECT 69.019 3.799 69.105 3.934 ;
      RECT 68.933 3.795 69.019 3.932 ;
      RECT 68.847 3.791 68.933 3.929 ;
      RECT 68.761 3.788 68.847 3.927 ;
      RECT 68.675 3.784 68.761 3.924 ;
      RECT 68.589 3.781 68.675 3.922 ;
      RECT 68.503 3.777 68.589 3.919 ;
      RECT 68.417 3.774 68.503 3.917 ;
      RECT 68.331 3.77 68.417 3.914 ;
      RECT 68.245 3.767 68.331 3.912 ;
      RECT 68.235 3.765 68.245 3.908 ;
      RECT 68.23 3.765 68.235 3.906 ;
      RECT 68.19 3.76 68.23 3.9 ;
      RECT 68.176 3.751 68.19 3.893 ;
      RECT 68.09 3.721 68.176 3.878 ;
      RECT 68.07 3.687 68.09 3.863 ;
      RECT 68 3.656 68.07 3.85 ;
      RECT 67.995 3.631 68 3.839 ;
      RECT 67.99 3.625 67.995 3.837 ;
      RECT 67.921 3.47 67.99 3.825 ;
      RECT 67.835 3.47 67.921 3.799 ;
      RECT 67.81 3.47 67.835 3.778 ;
      RECT 67.805 3.47 67.81 3.768 ;
      RECT 67.8 3.47 67.805 3.76 ;
      RECT 67.78 3.47 67.8 3.743 ;
      RECT 70.2 2.04 70.46 2.3 ;
      RECT 70.185 2.04 70.46 2.203 ;
      RECT 70.155 2.04 70.46 2.178 ;
      RECT 70.12 1.88 70.4 2.16 ;
      RECT 70.09 3.37 70.15 3.63 ;
      RECT 69.115 2.06 69.17 2.32 ;
      RECT 70.05 3.327 70.09 3.63 ;
      RECT 70.021 3.248 70.05 3.63 ;
      RECT 69.935 3.12 70.021 3.63 ;
      RECT 69.915 3 69.935 3.63 ;
      RECT 69.89 2.951 69.915 3.63 ;
      RECT 69.885 2.916 69.89 3.48 ;
      RECT 69.855 2.876 69.885 3.418 ;
      RECT 69.83 2.813 69.855 3.333 ;
      RECT 69.82 2.775 69.83 3.27 ;
      RECT 69.805 2.75 69.82 3.231 ;
      RECT 69.762 2.708 69.805 3.137 ;
      RECT 69.76 2.681 69.762 3.064 ;
      RECT 69.755 2.676 69.76 3.055 ;
      RECT 69.75 2.669 69.755 3.03 ;
      RECT 69.745 2.663 69.75 3.015 ;
      RECT 69.74 2.657 69.745 3.003 ;
      RECT 69.73 2.648 69.74 2.985 ;
      RECT 69.725 2.639 69.73 2.963 ;
      RECT 69.7 2.62 69.725 2.913 ;
      RECT 69.695 2.601 69.7 2.863 ;
      RECT 69.68 2.587 69.695 2.823 ;
      RECT 69.675 2.573 69.68 2.79 ;
      RECT 69.67 2.566 69.675 2.783 ;
      RECT 69.655 2.553 69.67 2.775 ;
      RECT 69.61 2.515 69.655 2.748 ;
      RECT 69.58 2.468 69.61 2.713 ;
      RECT 69.56 2.437 69.58 2.69 ;
      RECT 69.48 2.37 69.56 2.643 ;
      RECT 69.45 2.3 69.48 2.59 ;
      RECT 69.445 2.277 69.45 2.573 ;
      RECT 69.415 2.255 69.445 2.558 ;
      RECT 69.385 2.214 69.415 2.53 ;
      RECT 69.38 2.189 69.385 2.515 ;
      RECT 69.375 2.183 69.38 2.508 ;
      RECT 69.365 2.06 69.375 2.5 ;
      RECT 69.355 2.06 69.365 2.493 ;
      RECT 69.35 2.06 69.355 2.485 ;
      RECT 69.33 2.06 69.35 2.473 ;
      RECT 69.28 2.06 69.33 2.443 ;
      RECT 69.225 2.06 69.28 2.393 ;
      RECT 69.195 2.06 69.225 2.353 ;
      RECT 69.17 2.06 69.195 2.33 ;
      RECT 69.04 2.785 69.32 3.065 ;
      RECT 69.005 2.7 69.265 2.96 ;
      RECT 69.005 2.782 69.275 2.96 ;
      RECT 67.205 2.155 67.21 2.64 ;
      RECT 67.095 2.34 67.1 2.64 ;
      RECT 67.005 2.38 67.07 2.64 ;
      RECT 68.68 1.88 68.77 2.51 ;
      RECT 68.645 1.93 68.65 2.51 ;
      RECT 68.59 1.955 68.6 2.51 ;
      RECT 68.545 1.955 68.555 2.51 ;
      RECT 68.915 1.88 68.96 2.16 ;
      RECT 67.765 1.61 67.965 1.75 ;
      RECT 68.881 1.88 68.915 2.172 ;
      RECT 68.795 1.88 68.881 2.212 ;
      RECT 68.78 1.88 68.795 2.253 ;
      RECT 68.775 1.88 68.78 2.273 ;
      RECT 68.77 1.88 68.775 2.293 ;
      RECT 68.65 1.922 68.68 2.51 ;
      RECT 68.6 1.942 68.645 2.51 ;
      RECT 68.585 1.957 68.59 2.51 ;
      RECT 68.555 1.957 68.585 2.51 ;
      RECT 68.51 1.942 68.545 2.51 ;
      RECT 68.505 1.93 68.51 2.29 ;
      RECT 68.5 1.927 68.505 2.27 ;
      RECT 68.485 1.917 68.5 2.223 ;
      RECT 68.48 1.91 68.485 2.186 ;
      RECT 68.475 1.907 68.48 2.169 ;
      RECT 68.46 1.897 68.475 2.125 ;
      RECT 68.455 1.888 68.46 2.085 ;
      RECT 68.45 1.884 68.455 2.07 ;
      RECT 68.44 1.878 68.45 2.053 ;
      RECT 68.4 1.859 68.44 2.028 ;
      RECT 68.395 1.841 68.4 2.008 ;
      RECT 68.385 1.835 68.395 2.003 ;
      RECT 68.355 1.819 68.385 1.99 ;
      RECT 68.34 1.801 68.355 1.973 ;
      RECT 68.325 1.789 68.34 1.96 ;
      RECT 68.32 1.781 68.325 1.953 ;
      RECT 68.29 1.767 68.32 1.94 ;
      RECT 68.285 1.752 68.29 1.928 ;
      RECT 68.275 1.746 68.285 1.92 ;
      RECT 68.255 1.734 68.275 1.908 ;
      RECT 68.245 1.722 68.255 1.895 ;
      RECT 68.215 1.706 68.245 1.88 ;
      RECT 68.195 1.686 68.215 1.863 ;
      RECT 68.19 1.676 68.195 1.853 ;
      RECT 68.165 1.664 68.19 1.84 ;
      RECT 68.16 1.652 68.165 1.828 ;
      RECT 68.155 1.647 68.16 1.824 ;
      RECT 68.14 1.64 68.155 1.816 ;
      RECT 68.13 1.627 68.14 1.806 ;
      RECT 68.125 1.625 68.13 1.8 ;
      RECT 68.1 1.618 68.125 1.789 ;
      RECT 68.095 1.611 68.1 1.778 ;
      RECT 68.07 1.61 68.095 1.765 ;
      RECT 68.051 1.61 68.07 1.755 ;
      RECT 67.965 1.61 68.051 1.752 ;
      RECT 67.735 1.61 67.765 1.755 ;
      RECT 67.695 1.617 67.735 1.768 ;
      RECT 67.67 1.627 67.695 1.781 ;
      RECT 67.655 1.636 67.67 1.791 ;
      RECT 67.625 1.641 67.655 1.81 ;
      RECT 67.62 1.647 67.625 1.828 ;
      RECT 67.6 1.657 67.62 1.843 ;
      RECT 67.59 1.67 67.6 1.863 ;
      RECT 67.575 1.682 67.59 1.88 ;
      RECT 67.57 1.692 67.575 1.89 ;
      RECT 67.565 1.697 67.57 1.895 ;
      RECT 67.555 1.705 67.565 1.908 ;
      RECT 67.505 1.737 67.555 1.945 ;
      RECT 67.49 1.772 67.505 1.986 ;
      RECT 67.485 1.782 67.49 2.001 ;
      RECT 67.48 1.787 67.485 2.008 ;
      RECT 67.455 1.803 67.48 2.028 ;
      RECT 67.44 1.824 67.455 2.053 ;
      RECT 67.415 1.845 67.44 2.078 ;
      RECT 67.405 1.864 67.415 2.101 ;
      RECT 67.38 1.882 67.405 2.124 ;
      RECT 67.365 1.902 67.38 2.148 ;
      RECT 67.36 1.912 67.365 2.16 ;
      RECT 67.345 1.924 67.36 2.18 ;
      RECT 67.335 1.939 67.345 2.22 ;
      RECT 67.33 1.947 67.335 2.248 ;
      RECT 67.32 1.957 67.33 2.268 ;
      RECT 67.315 1.97 67.32 2.293 ;
      RECT 67.31 1.983 67.315 2.313 ;
      RECT 67.305 1.989 67.31 2.335 ;
      RECT 67.295 1.998 67.305 2.355 ;
      RECT 67.29 2.018 67.295 2.378 ;
      RECT 67.285 2.024 67.29 2.398 ;
      RECT 67.28 2.031 67.285 2.42 ;
      RECT 67.275 2.042 67.28 2.433 ;
      RECT 67.265 2.052 67.275 2.458 ;
      RECT 67.245 2.077 67.265 2.64 ;
      RECT 67.215 2.117 67.245 2.64 ;
      RECT 67.21 2.147 67.215 2.64 ;
      RECT 67.185 2.175 67.205 2.64 ;
      RECT 67.155 2.22 67.185 2.64 ;
      RECT 67.15 2.247 67.155 2.64 ;
      RECT 67.13 2.265 67.15 2.64 ;
      RECT 67.12 2.29 67.13 2.64 ;
      RECT 67.115 2.302 67.12 2.64 ;
      RECT 67.1 2.325 67.115 2.64 ;
      RECT 67.08 2.352 67.095 2.64 ;
      RECT 67.07 2.375 67.08 2.64 ;
      RECT 68.86 3.26 68.94 3.52 ;
      RECT 68.095 2.48 68.165 2.74 ;
      RECT 68.826 3.227 68.86 3.52 ;
      RECT 68.74 3.13 68.826 3.52 ;
      RECT 68.72 3.042 68.74 3.52 ;
      RECT 68.71 3.012 68.72 3.52 ;
      RECT 68.7 2.992 68.71 3.52 ;
      RECT 68.68 2.979 68.7 3.52 ;
      RECT 68.665 2.969 68.68 3.348 ;
      RECT 68.66 2.962 68.665 3.303 ;
      RECT 68.65 2.956 68.66 3.293 ;
      RECT 68.64 2.948 68.65 3.275 ;
      RECT 68.635 2.942 68.64 3.263 ;
      RECT 68.625 2.937 68.635 3.25 ;
      RECT 68.605 2.927 68.625 3.223 ;
      RECT 68.565 2.906 68.605 3.175 ;
      RECT 68.55 2.887 68.565 3.133 ;
      RECT 68.525 2.873 68.55 3.103 ;
      RECT 68.515 2.861 68.525 3.07 ;
      RECT 68.51 2.856 68.515 3.06 ;
      RECT 68.48 2.842 68.51 3.04 ;
      RECT 68.47 2.826 68.48 3.013 ;
      RECT 68.465 2.821 68.47 3.003 ;
      RECT 68.44 2.812 68.465 2.983 ;
      RECT 68.43 2.8 68.44 2.963 ;
      RECT 68.36 2.768 68.43 2.938 ;
      RECT 68.355 2.737 68.36 2.915 ;
      RECT 68.306 2.48 68.355 2.898 ;
      RECT 68.22 2.48 68.306 2.857 ;
      RECT 68.165 2.48 68.22 2.785 ;
      RECT 68.255 3.265 68.415 3.525 ;
      RECT 67.78 1.88 67.83 2.565 ;
      RECT 67.57 2.305 67.605 2.565 ;
      RECT 67.885 1.88 67.89 2.34 ;
      RECT 67.975 1.88 68 2.16 ;
      RECT 68.25 3.262 68.255 3.525 ;
      RECT 68.215 3.25 68.25 3.525 ;
      RECT 68.155 3.223 68.215 3.525 ;
      RECT 68.15 3.206 68.155 3.379 ;
      RECT 68.145 3.203 68.15 3.366 ;
      RECT 68.125 3.196 68.145 3.353 ;
      RECT 68.09 3.179 68.125 3.335 ;
      RECT 68.05 3.158 68.09 3.315 ;
      RECT 68.045 3.146 68.05 3.303 ;
      RECT 68.005 3.132 68.045 3.289 ;
      RECT 67.985 3.115 68.005 3.271 ;
      RECT 67.975 3.107 67.985 3.263 ;
      RECT 67.96 1.88 67.975 2.178 ;
      RECT 67.945 3.097 67.975 3.25 ;
      RECT 67.93 1.88 67.96 2.223 ;
      RECT 67.935 3.087 67.945 3.237 ;
      RECT 67.905 3.072 67.935 3.224 ;
      RECT 67.89 1.88 67.93 2.29 ;
      RECT 67.89 3.04 67.905 3.21 ;
      RECT 67.885 3.012 67.89 3.204 ;
      RECT 67.88 1.88 67.885 2.345 ;
      RECT 67.87 2.982 67.885 3.198 ;
      RECT 67.875 1.88 67.88 2.358 ;
      RECT 67.865 1.88 67.875 2.378 ;
      RECT 67.83 2.895 67.87 3.183 ;
      RECT 67.83 1.88 67.865 2.418 ;
      RECT 67.825 2.827 67.83 3.171 ;
      RECT 67.81 2.782 67.825 3.166 ;
      RECT 67.805 2.72 67.81 3.161 ;
      RECT 67.78 2.627 67.805 3.154 ;
      RECT 67.775 1.88 67.78 3.146 ;
      RECT 67.76 1.88 67.775 3.133 ;
      RECT 67.74 1.88 67.76 3.09 ;
      RECT 67.73 1.88 67.74 3.04 ;
      RECT 67.725 1.88 67.73 3.013 ;
      RECT 67.72 1.88 67.725 2.991 ;
      RECT 67.715 2.106 67.72 2.974 ;
      RECT 67.71 2.128 67.715 2.952 ;
      RECT 67.705 2.17 67.71 2.935 ;
      RECT 67.675 2.22 67.705 2.879 ;
      RECT 67.67 2.247 67.675 2.821 ;
      RECT 67.655 2.265 67.67 2.785 ;
      RECT 67.65 2.283 67.655 2.749 ;
      RECT 67.644 2.29 67.65 2.73 ;
      RECT 67.64 2.297 67.644 2.713 ;
      RECT 67.635 2.302 67.64 2.682 ;
      RECT 67.625 2.305 67.635 2.657 ;
      RECT 67.615 2.305 67.625 2.623 ;
      RECT 67.61 2.305 67.615 2.6 ;
      RECT 67.605 2.305 67.61 2.58 ;
      RECT 66.52 2.44 66.8 2.72 ;
      RECT 66.52 2.44 66.82 2.615 ;
      RECT 66.61 2.33 66.87 2.59 ;
      RECT 66.575 2.425 66.87 2.59 ;
      RECT 66.7 0.945 66.865 2.59 ;
      RECT 66.6 0.945 66.97 1.315 ;
      RECT 66.225 3.47 66.485 3.73 ;
      RECT 66.245 3.397 66.425 3.73 ;
      RECT 66.245 3.14 66.42 3.73 ;
      RECT 66.245 2.932 66.41 3.73 ;
      RECT 66.25 2.85 66.41 3.73 ;
      RECT 66.25 2.615 66.4 3.73 ;
      RECT 66.25 2.462 66.395 3.73 ;
      RECT 66.255 2.447 66.395 3.73 ;
      RECT 66.305 2.162 66.395 3.73 ;
      RECT 66.26 2.397 66.395 3.73 ;
      RECT 66.29 2.215 66.395 3.73 ;
      RECT 66.275 2.327 66.395 3.73 ;
      RECT 66.28 2.285 66.395 3.73 ;
      RECT 66.275 2.327 66.41 2.39 ;
      RECT 66.31 1.915 66.415 2.335 ;
      RECT 66.31 1.915 66.43 2.318 ;
      RECT 66.31 1.915 66.465 2.28 ;
      RECT 66.305 2.162 66.515 2.213 ;
      RECT 66.31 1.915 66.57 2.175 ;
      RECT 65.57 2.62 65.83 2.88 ;
      RECT 65.57 2.62 65.84 2.838 ;
      RECT 65.57 2.62 65.926 2.809 ;
      RECT 65.57 2.62 65.995 2.761 ;
      RECT 65.57 2.62 66.03 2.73 ;
      RECT 65.8 2.44 66.08 2.72 ;
      RECT 65.635 2.605 66.08 2.72 ;
      RECT 65.725 2.482 65.83 2.88 ;
      RECT 65.655 2.545 66.08 2.72 ;
      RECT 60.105 6.22 60.425 6.545 ;
      RECT 60.135 5.695 60.305 6.545 ;
      RECT 60.135 5.695 60.31 6.045 ;
      RECT 60.135 5.695 61.11 5.87 ;
      RECT 60.935 1.965 61.11 5.87 ;
      RECT 60.88 1.965 61.23 2.315 ;
      RECT 60.905 6.655 61.23 6.98 ;
      RECT 59.79 6.745 61.23 6.915 ;
      RECT 59.79 2.395 59.95 6.915 ;
      RECT 60.105 2.365 60.425 2.685 ;
      RECT 59.79 2.395 60.425 2.565 ;
      RECT 58.5 2.705 58.84 3.055 ;
      RECT 57.895 2.77 58.84 2.97 ;
      RECT 57.895 2.765 58.11 2.97 ;
      RECT 57.91 2.34 58.11 2.97 ;
      RECT 56.9 2.34 57.18 2.72 ;
      RECT 58.59 2.7 58.76 3.055 ;
      RECT 56.895 2.34 57.18 2.673 ;
      RECT 56.875 2.34 57.18 2.65 ;
      RECT 56.865 2.34 57.18 2.63 ;
      RECT 56.855 2.34 57.18 2.615 ;
      RECT 56.83 2.34 57.18 2.588 ;
      RECT 56.82 2.34 57.18 2.563 ;
      RECT 56.775 2.295 57.055 2.555 ;
      RECT 56.775 2.34 58.11 2.54 ;
      RECT 56.775 2.335 57.1 2.555 ;
      RECT 56.775 2.327 57.095 2.555 ;
      RECT 56.775 2.317 57.09 2.555 ;
      RECT 56.775 2.305 57.085 2.555 ;
      RECT 55.7 3 55.98 3.28 ;
      RECT 55.7 3 56.015 3.26 ;
      RECT 47.98 6.655 48.33 7.005 ;
      RECT 55.445 6.61 55.795 6.96 ;
      RECT 47.98 6.685 55.795 6.885 ;
      RECT 55.735 2.42 55.785 2.68 ;
      RECT 55.525 2.42 55.53 2.68 ;
      RECT 54.72 1.975 54.75 2.235 ;
      RECT 54.49 1.975 54.565 2.235 ;
      RECT 55.71 2.37 55.735 2.68 ;
      RECT 55.705 2.327 55.71 2.68 ;
      RECT 55.7 2.31 55.705 2.68 ;
      RECT 55.695 2.297 55.7 2.68 ;
      RECT 55.62 2.18 55.695 2.68 ;
      RECT 55.575 1.997 55.62 2.68 ;
      RECT 55.57 1.925 55.575 2.68 ;
      RECT 55.555 1.9 55.57 2.68 ;
      RECT 55.53 1.862 55.555 2.68 ;
      RECT 55.52 1.842 55.53 2.402 ;
      RECT 55.505 1.834 55.52 2.357 ;
      RECT 55.5 1.826 55.505 2.328 ;
      RECT 55.495 1.823 55.5 2.308 ;
      RECT 55.49 1.82 55.495 2.288 ;
      RECT 55.485 1.817 55.49 2.268 ;
      RECT 55.455 1.806 55.485 2.205 ;
      RECT 55.435 1.791 55.455 2.12 ;
      RECT 55.43 1.783 55.435 2.083 ;
      RECT 55.42 1.777 55.43 2.05 ;
      RECT 55.405 1.769 55.42 2.01 ;
      RECT 55.4 1.762 55.405 1.97 ;
      RECT 55.395 1.759 55.4 1.948 ;
      RECT 55.39 1.756 55.395 1.935 ;
      RECT 55.385 1.755 55.39 1.925 ;
      RECT 55.37 1.749 55.385 1.915 ;
      RECT 55.345 1.736 55.37 1.9 ;
      RECT 55.295 1.711 55.345 1.871 ;
      RECT 55.28 1.69 55.295 1.846 ;
      RECT 55.27 1.683 55.28 1.835 ;
      RECT 55.215 1.664 55.27 1.808 ;
      RECT 55.19 1.642 55.215 1.781 ;
      RECT 55.185 1.635 55.19 1.776 ;
      RECT 55.17 1.635 55.185 1.774 ;
      RECT 55.145 1.627 55.17 1.77 ;
      RECT 55.13 1.625 55.145 1.766 ;
      RECT 55.1 1.625 55.13 1.763 ;
      RECT 55.09 1.625 55.1 1.758 ;
      RECT 55.045 1.625 55.09 1.756 ;
      RECT 55.016 1.625 55.045 1.757 ;
      RECT 54.93 1.625 55.016 1.759 ;
      RECT 54.916 1.626 54.93 1.761 ;
      RECT 54.83 1.627 54.916 1.763 ;
      RECT 54.815 1.628 54.83 1.773 ;
      RECT 54.81 1.629 54.815 1.782 ;
      RECT 54.79 1.632 54.81 1.792 ;
      RECT 54.775 1.64 54.79 1.807 ;
      RECT 54.755 1.658 54.775 1.822 ;
      RECT 54.745 1.67 54.755 1.845 ;
      RECT 54.735 1.679 54.745 1.875 ;
      RECT 54.72 1.691 54.735 1.92 ;
      RECT 54.665 1.724 54.72 2.235 ;
      RECT 54.66 1.752 54.665 2.235 ;
      RECT 54.64 1.767 54.66 2.235 ;
      RECT 54.605 1.827 54.64 2.235 ;
      RECT 54.603 1.877 54.605 2.235 ;
      RECT 54.6 1.885 54.603 2.235 ;
      RECT 54.59 1.9 54.6 2.235 ;
      RECT 54.585 1.912 54.59 2.235 ;
      RECT 54.575 1.937 54.585 2.235 ;
      RECT 54.565 1.965 54.575 2.235 ;
      RECT 52.47 3.47 52.52 3.73 ;
      RECT 55.38 3.02 55.44 3.28 ;
      RECT 55.365 3.02 55.38 3.29 ;
      RECT 55.346 3.02 55.365 3.323 ;
      RECT 55.26 3.02 55.346 3.448 ;
      RECT 55.18 3.02 55.26 3.63 ;
      RECT 55.175 3.257 55.18 3.715 ;
      RECT 55.15 3.327 55.175 3.743 ;
      RECT 55.145 3.397 55.15 3.77 ;
      RECT 55.125 3.469 55.145 3.792 ;
      RECT 55.12 3.536 55.125 3.815 ;
      RECT 55.11 3.565 55.12 3.83 ;
      RECT 55.1 3.587 55.11 3.847 ;
      RECT 55.095 3.597 55.1 3.858 ;
      RECT 55.09 3.605 55.095 3.866 ;
      RECT 55.08 3.613 55.09 3.878 ;
      RECT 55.075 3.625 55.08 3.888 ;
      RECT 55.07 3.633 55.075 3.893 ;
      RECT 55.05 3.651 55.07 3.903 ;
      RECT 55.045 3.668 55.05 3.91 ;
      RECT 55.04 3.676 55.045 3.911 ;
      RECT 55.035 3.687 55.04 3.913 ;
      RECT 54.995 3.725 55.035 3.923 ;
      RECT 54.99 3.76 54.995 3.934 ;
      RECT 54.985 3.765 54.99 3.937 ;
      RECT 54.96 3.775 54.985 3.944 ;
      RECT 54.95 3.789 54.96 3.953 ;
      RECT 54.93 3.801 54.95 3.956 ;
      RECT 54.88 3.82 54.93 3.96 ;
      RECT 54.835 3.835 54.88 3.965 ;
      RECT 54.77 3.838 54.835 3.971 ;
      RECT 54.755 3.836 54.77 3.978 ;
      RECT 54.725 3.835 54.755 3.978 ;
      RECT 54.686 3.834 54.725 3.974 ;
      RECT 54.6 3.831 54.686 3.97 ;
      RECT 54.583 3.829 54.6 3.967 ;
      RECT 54.497 3.827 54.583 3.964 ;
      RECT 54.411 3.824 54.497 3.958 ;
      RECT 54.325 3.82 54.411 3.953 ;
      RECT 54.247 3.817 54.325 3.949 ;
      RECT 54.161 3.814 54.247 3.947 ;
      RECT 54.075 3.811 54.161 3.944 ;
      RECT 54.017 3.809 54.075 3.941 ;
      RECT 53.931 3.806 54.017 3.939 ;
      RECT 53.845 3.802 53.931 3.937 ;
      RECT 53.759 3.799 53.845 3.934 ;
      RECT 53.673 3.795 53.759 3.932 ;
      RECT 53.587 3.791 53.673 3.929 ;
      RECT 53.501 3.788 53.587 3.927 ;
      RECT 53.415 3.784 53.501 3.924 ;
      RECT 53.329 3.781 53.415 3.922 ;
      RECT 53.243 3.777 53.329 3.919 ;
      RECT 53.157 3.774 53.243 3.917 ;
      RECT 53.071 3.77 53.157 3.914 ;
      RECT 52.985 3.767 53.071 3.912 ;
      RECT 52.975 3.765 52.985 3.908 ;
      RECT 52.97 3.765 52.975 3.906 ;
      RECT 52.93 3.76 52.97 3.9 ;
      RECT 52.916 3.751 52.93 3.893 ;
      RECT 52.83 3.721 52.916 3.878 ;
      RECT 52.81 3.687 52.83 3.863 ;
      RECT 52.74 3.656 52.81 3.85 ;
      RECT 52.735 3.631 52.74 3.839 ;
      RECT 52.73 3.625 52.735 3.837 ;
      RECT 52.661 3.47 52.73 3.825 ;
      RECT 52.575 3.47 52.661 3.799 ;
      RECT 52.55 3.47 52.575 3.778 ;
      RECT 52.545 3.47 52.55 3.768 ;
      RECT 52.54 3.47 52.545 3.76 ;
      RECT 52.52 3.47 52.54 3.743 ;
      RECT 54.94 2.04 55.2 2.3 ;
      RECT 54.925 2.04 55.2 2.203 ;
      RECT 54.895 2.04 55.2 2.178 ;
      RECT 54.86 1.88 55.14 2.16 ;
      RECT 54.83 3.37 54.89 3.63 ;
      RECT 53.855 2.06 53.91 2.32 ;
      RECT 54.79 3.327 54.83 3.63 ;
      RECT 54.761 3.248 54.79 3.63 ;
      RECT 54.675 3.12 54.761 3.63 ;
      RECT 54.655 3 54.675 3.63 ;
      RECT 54.63 2.951 54.655 3.63 ;
      RECT 54.625 2.916 54.63 3.48 ;
      RECT 54.595 2.876 54.625 3.418 ;
      RECT 54.57 2.813 54.595 3.333 ;
      RECT 54.56 2.775 54.57 3.27 ;
      RECT 54.545 2.75 54.56 3.231 ;
      RECT 54.502 2.708 54.545 3.137 ;
      RECT 54.5 2.681 54.502 3.064 ;
      RECT 54.495 2.676 54.5 3.055 ;
      RECT 54.49 2.669 54.495 3.03 ;
      RECT 54.485 2.663 54.49 3.015 ;
      RECT 54.48 2.657 54.485 3.003 ;
      RECT 54.47 2.648 54.48 2.985 ;
      RECT 54.465 2.639 54.47 2.963 ;
      RECT 54.44 2.62 54.465 2.913 ;
      RECT 54.435 2.601 54.44 2.863 ;
      RECT 54.42 2.587 54.435 2.823 ;
      RECT 54.415 2.573 54.42 2.79 ;
      RECT 54.41 2.566 54.415 2.783 ;
      RECT 54.395 2.553 54.41 2.775 ;
      RECT 54.35 2.515 54.395 2.748 ;
      RECT 54.32 2.468 54.35 2.713 ;
      RECT 54.3 2.437 54.32 2.69 ;
      RECT 54.22 2.37 54.3 2.643 ;
      RECT 54.19 2.3 54.22 2.59 ;
      RECT 54.185 2.277 54.19 2.573 ;
      RECT 54.155 2.255 54.185 2.558 ;
      RECT 54.125 2.214 54.155 2.53 ;
      RECT 54.12 2.189 54.125 2.515 ;
      RECT 54.115 2.183 54.12 2.508 ;
      RECT 54.105 2.06 54.115 2.5 ;
      RECT 54.095 2.06 54.105 2.493 ;
      RECT 54.09 2.06 54.095 2.485 ;
      RECT 54.07 2.06 54.09 2.473 ;
      RECT 54.02 2.06 54.07 2.443 ;
      RECT 53.965 2.06 54.02 2.393 ;
      RECT 53.935 2.06 53.965 2.353 ;
      RECT 53.91 2.06 53.935 2.33 ;
      RECT 53.78 2.785 54.06 3.065 ;
      RECT 53.745 2.7 54.005 2.96 ;
      RECT 53.745 2.782 54.015 2.96 ;
      RECT 51.945 2.155 51.95 2.64 ;
      RECT 51.835 2.34 51.84 2.64 ;
      RECT 51.745 2.38 51.81 2.64 ;
      RECT 53.42 1.88 53.51 2.51 ;
      RECT 53.385 1.93 53.39 2.51 ;
      RECT 53.33 1.955 53.34 2.51 ;
      RECT 53.285 1.955 53.295 2.51 ;
      RECT 53.655 1.88 53.7 2.16 ;
      RECT 52.505 1.61 52.705 1.75 ;
      RECT 53.621 1.88 53.655 2.172 ;
      RECT 53.535 1.88 53.621 2.212 ;
      RECT 53.52 1.88 53.535 2.253 ;
      RECT 53.515 1.88 53.52 2.273 ;
      RECT 53.51 1.88 53.515 2.293 ;
      RECT 53.39 1.922 53.42 2.51 ;
      RECT 53.34 1.942 53.385 2.51 ;
      RECT 53.325 1.957 53.33 2.51 ;
      RECT 53.295 1.957 53.325 2.51 ;
      RECT 53.25 1.942 53.285 2.51 ;
      RECT 53.245 1.93 53.25 2.29 ;
      RECT 53.24 1.927 53.245 2.27 ;
      RECT 53.225 1.917 53.24 2.223 ;
      RECT 53.22 1.91 53.225 2.186 ;
      RECT 53.215 1.907 53.22 2.169 ;
      RECT 53.2 1.897 53.215 2.125 ;
      RECT 53.195 1.888 53.2 2.085 ;
      RECT 53.19 1.884 53.195 2.07 ;
      RECT 53.18 1.878 53.19 2.053 ;
      RECT 53.14 1.859 53.18 2.028 ;
      RECT 53.135 1.841 53.14 2.008 ;
      RECT 53.125 1.835 53.135 2.003 ;
      RECT 53.095 1.819 53.125 1.99 ;
      RECT 53.08 1.801 53.095 1.973 ;
      RECT 53.065 1.789 53.08 1.96 ;
      RECT 53.06 1.781 53.065 1.953 ;
      RECT 53.03 1.767 53.06 1.94 ;
      RECT 53.025 1.752 53.03 1.928 ;
      RECT 53.015 1.746 53.025 1.92 ;
      RECT 52.995 1.734 53.015 1.908 ;
      RECT 52.985 1.722 52.995 1.895 ;
      RECT 52.955 1.706 52.985 1.88 ;
      RECT 52.935 1.686 52.955 1.863 ;
      RECT 52.93 1.676 52.935 1.853 ;
      RECT 52.905 1.664 52.93 1.84 ;
      RECT 52.9 1.652 52.905 1.828 ;
      RECT 52.895 1.647 52.9 1.824 ;
      RECT 52.88 1.64 52.895 1.816 ;
      RECT 52.87 1.627 52.88 1.806 ;
      RECT 52.865 1.625 52.87 1.8 ;
      RECT 52.84 1.618 52.865 1.789 ;
      RECT 52.835 1.611 52.84 1.778 ;
      RECT 52.81 1.61 52.835 1.765 ;
      RECT 52.791 1.61 52.81 1.755 ;
      RECT 52.705 1.61 52.791 1.752 ;
      RECT 52.475 1.61 52.505 1.755 ;
      RECT 52.435 1.617 52.475 1.768 ;
      RECT 52.41 1.627 52.435 1.781 ;
      RECT 52.395 1.636 52.41 1.791 ;
      RECT 52.365 1.641 52.395 1.81 ;
      RECT 52.36 1.647 52.365 1.828 ;
      RECT 52.34 1.657 52.36 1.843 ;
      RECT 52.33 1.67 52.34 1.863 ;
      RECT 52.315 1.682 52.33 1.88 ;
      RECT 52.31 1.692 52.315 1.89 ;
      RECT 52.305 1.697 52.31 1.895 ;
      RECT 52.295 1.705 52.305 1.908 ;
      RECT 52.245 1.737 52.295 1.945 ;
      RECT 52.23 1.772 52.245 1.986 ;
      RECT 52.225 1.782 52.23 2.001 ;
      RECT 52.22 1.787 52.225 2.008 ;
      RECT 52.195 1.803 52.22 2.028 ;
      RECT 52.18 1.824 52.195 2.053 ;
      RECT 52.155 1.845 52.18 2.078 ;
      RECT 52.145 1.864 52.155 2.101 ;
      RECT 52.12 1.882 52.145 2.124 ;
      RECT 52.105 1.902 52.12 2.148 ;
      RECT 52.1 1.912 52.105 2.16 ;
      RECT 52.085 1.924 52.1 2.18 ;
      RECT 52.075 1.939 52.085 2.22 ;
      RECT 52.07 1.947 52.075 2.248 ;
      RECT 52.06 1.957 52.07 2.268 ;
      RECT 52.055 1.97 52.06 2.293 ;
      RECT 52.05 1.983 52.055 2.313 ;
      RECT 52.045 1.989 52.05 2.335 ;
      RECT 52.035 1.998 52.045 2.355 ;
      RECT 52.03 2.018 52.035 2.378 ;
      RECT 52.025 2.024 52.03 2.398 ;
      RECT 52.02 2.031 52.025 2.42 ;
      RECT 52.015 2.042 52.02 2.433 ;
      RECT 52.005 2.052 52.015 2.458 ;
      RECT 51.985 2.077 52.005 2.64 ;
      RECT 51.955 2.117 51.985 2.64 ;
      RECT 51.95 2.147 51.955 2.64 ;
      RECT 51.925 2.175 51.945 2.64 ;
      RECT 51.895 2.22 51.925 2.64 ;
      RECT 51.89 2.247 51.895 2.64 ;
      RECT 51.87 2.265 51.89 2.64 ;
      RECT 51.86 2.29 51.87 2.64 ;
      RECT 51.855 2.302 51.86 2.64 ;
      RECT 51.84 2.325 51.855 2.64 ;
      RECT 51.82 2.352 51.835 2.64 ;
      RECT 51.81 2.375 51.82 2.64 ;
      RECT 53.6 3.26 53.68 3.52 ;
      RECT 52.835 2.48 52.905 2.74 ;
      RECT 53.566 3.227 53.6 3.52 ;
      RECT 53.48 3.13 53.566 3.52 ;
      RECT 53.46 3.042 53.48 3.52 ;
      RECT 53.45 3.012 53.46 3.52 ;
      RECT 53.44 2.992 53.45 3.52 ;
      RECT 53.42 2.979 53.44 3.52 ;
      RECT 53.405 2.969 53.42 3.348 ;
      RECT 53.4 2.962 53.405 3.303 ;
      RECT 53.39 2.956 53.4 3.293 ;
      RECT 53.38 2.948 53.39 3.275 ;
      RECT 53.375 2.942 53.38 3.263 ;
      RECT 53.365 2.937 53.375 3.25 ;
      RECT 53.345 2.927 53.365 3.223 ;
      RECT 53.305 2.906 53.345 3.175 ;
      RECT 53.29 2.887 53.305 3.133 ;
      RECT 53.265 2.873 53.29 3.103 ;
      RECT 53.255 2.861 53.265 3.07 ;
      RECT 53.25 2.856 53.255 3.06 ;
      RECT 53.22 2.842 53.25 3.04 ;
      RECT 53.21 2.826 53.22 3.013 ;
      RECT 53.205 2.821 53.21 3.003 ;
      RECT 53.18 2.812 53.205 2.983 ;
      RECT 53.17 2.8 53.18 2.963 ;
      RECT 53.1 2.768 53.17 2.938 ;
      RECT 53.095 2.737 53.1 2.915 ;
      RECT 53.046 2.48 53.095 2.898 ;
      RECT 52.96 2.48 53.046 2.857 ;
      RECT 52.905 2.48 52.96 2.785 ;
      RECT 52.995 3.265 53.155 3.525 ;
      RECT 52.52 1.88 52.57 2.565 ;
      RECT 52.31 2.305 52.345 2.565 ;
      RECT 52.625 1.88 52.63 2.34 ;
      RECT 52.715 1.88 52.74 2.16 ;
      RECT 52.99 3.262 52.995 3.525 ;
      RECT 52.955 3.25 52.99 3.525 ;
      RECT 52.895 3.223 52.955 3.525 ;
      RECT 52.89 3.206 52.895 3.379 ;
      RECT 52.885 3.203 52.89 3.366 ;
      RECT 52.865 3.196 52.885 3.353 ;
      RECT 52.83 3.179 52.865 3.335 ;
      RECT 52.79 3.158 52.83 3.315 ;
      RECT 52.785 3.146 52.79 3.303 ;
      RECT 52.745 3.132 52.785 3.289 ;
      RECT 52.725 3.115 52.745 3.271 ;
      RECT 52.715 3.107 52.725 3.263 ;
      RECT 52.7 1.88 52.715 2.178 ;
      RECT 52.685 3.097 52.715 3.25 ;
      RECT 52.67 1.88 52.7 2.223 ;
      RECT 52.675 3.087 52.685 3.237 ;
      RECT 52.645 3.072 52.675 3.224 ;
      RECT 52.63 1.88 52.67 2.29 ;
      RECT 52.63 3.04 52.645 3.21 ;
      RECT 52.625 3.012 52.63 3.204 ;
      RECT 52.62 1.88 52.625 2.345 ;
      RECT 52.61 2.982 52.625 3.198 ;
      RECT 52.615 1.88 52.62 2.358 ;
      RECT 52.605 1.88 52.615 2.378 ;
      RECT 52.57 2.895 52.61 3.183 ;
      RECT 52.57 1.88 52.605 2.418 ;
      RECT 52.565 2.827 52.57 3.171 ;
      RECT 52.55 2.782 52.565 3.166 ;
      RECT 52.545 2.72 52.55 3.161 ;
      RECT 52.52 2.627 52.545 3.154 ;
      RECT 52.515 1.88 52.52 3.146 ;
      RECT 52.5 1.88 52.515 3.133 ;
      RECT 52.48 1.88 52.5 3.09 ;
      RECT 52.47 1.88 52.48 3.04 ;
      RECT 52.465 1.88 52.47 3.013 ;
      RECT 52.46 1.88 52.465 2.991 ;
      RECT 52.455 2.106 52.46 2.974 ;
      RECT 52.45 2.128 52.455 2.952 ;
      RECT 52.445 2.17 52.45 2.935 ;
      RECT 52.415 2.22 52.445 2.879 ;
      RECT 52.41 2.247 52.415 2.821 ;
      RECT 52.395 2.265 52.41 2.785 ;
      RECT 52.39 2.283 52.395 2.749 ;
      RECT 52.384 2.29 52.39 2.73 ;
      RECT 52.38 2.297 52.384 2.713 ;
      RECT 52.375 2.302 52.38 2.682 ;
      RECT 52.365 2.305 52.375 2.657 ;
      RECT 52.355 2.305 52.365 2.623 ;
      RECT 52.35 2.305 52.355 2.6 ;
      RECT 52.345 2.305 52.35 2.58 ;
      RECT 51.26 2.44 51.54 2.72 ;
      RECT 51.26 2.44 51.56 2.615 ;
      RECT 51.35 2.33 51.61 2.59 ;
      RECT 51.315 2.425 51.61 2.59 ;
      RECT 51.44 0.945 51.605 2.59 ;
      RECT 51.34 0.945 51.71 1.315 ;
      RECT 50.965 3.47 51.225 3.73 ;
      RECT 50.985 3.397 51.165 3.73 ;
      RECT 50.985 3.14 51.16 3.73 ;
      RECT 50.985 2.932 51.15 3.73 ;
      RECT 50.99 2.85 51.15 3.73 ;
      RECT 50.99 2.615 51.14 3.73 ;
      RECT 50.99 2.462 51.135 3.73 ;
      RECT 50.995 2.447 51.135 3.73 ;
      RECT 51.045 2.162 51.135 3.73 ;
      RECT 51 2.397 51.135 3.73 ;
      RECT 51.03 2.215 51.135 3.73 ;
      RECT 51.015 2.327 51.135 3.73 ;
      RECT 51.02 2.285 51.135 3.73 ;
      RECT 51.015 2.327 51.15 2.39 ;
      RECT 51.05 1.915 51.155 2.335 ;
      RECT 51.05 1.915 51.17 2.318 ;
      RECT 51.05 1.915 51.205 2.28 ;
      RECT 51.045 2.162 51.255 2.213 ;
      RECT 51.05 1.915 51.31 2.175 ;
      RECT 50.31 2.62 50.57 2.88 ;
      RECT 50.31 2.62 50.58 2.838 ;
      RECT 50.31 2.62 50.666 2.809 ;
      RECT 50.31 2.62 50.735 2.761 ;
      RECT 50.31 2.62 50.77 2.73 ;
      RECT 50.54 2.44 50.82 2.72 ;
      RECT 50.375 2.605 50.82 2.72 ;
      RECT 50.465 2.482 50.57 2.88 ;
      RECT 50.395 2.545 50.82 2.72 ;
      RECT 44.845 6.22 45.165 6.545 ;
      RECT 44.875 5.695 45.045 6.545 ;
      RECT 44.875 5.695 45.05 6.045 ;
      RECT 44.875 5.695 45.85 5.87 ;
      RECT 45.675 1.965 45.85 5.87 ;
      RECT 45.62 1.965 45.97 2.315 ;
      RECT 45.645 6.655 45.97 6.98 ;
      RECT 44.53 6.745 45.97 6.915 ;
      RECT 44.53 2.395 44.69 6.915 ;
      RECT 44.845 2.365 45.165 2.685 ;
      RECT 44.53 2.395 45.165 2.565 ;
      RECT 43.24 2.705 43.58 3.055 ;
      RECT 42.635 2.77 43.58 2.97 ;
      RECT 42.635 2.765 42.85 2.97 ;
      RECT 42.65 2.34 42.85 2.97 ;
      RECT 41.64 2.34 41.92 2.72 ;
      RECT 43.33 2.7 43.5 3.055 ;
      RECT 41.635 2.34 41.92 2.673 ;
      RECT 41.615 2.34 41.92 2.65 ;
      RECT 41.605 2.34 41.92 2.63 ;
      RECT 41.595 2.34 41.92 2.615 ;
      RECT 41.57 2.34 41.92 2.588 ;
      RECT 41.56 2.34 41.92 2.563 ;
      RECT 41.515 2.295 41.795 2.555 ;
      RECT 41.515 2.34 42.85 2.54 ;
      RECT 41.515 2.335 41.84 2.555 ;
      RECT 41.515 2.327 41.835 2.555 ;
      RECT 41.515 2.317 41.83 2.555 ;
      RECT 41.515 2.305 41.825 2.555 ;
      RECT 40.44 3 40.72 3.28 ;
      RECT 40.44 3 40.755 3.26 ;
      RECT 32.765 6.66 33.115 7.01 ;
      RECT 40.185 6.615 40.535 6.965 ;
      RECT 32.765 6.69 40.535 6.89 ;
      RECT 40.475 2.42 40.525 2.68 ;
      RECT 40.265 2.42 40.27 2.68 ;
      RECT 39.46 1.975 39.49 2.235 ;
      RECT 39.23 1.975 39.305 2.235 ;
      RECT 40.45 2.37 40.475 2.68 ;
      RECT 40.445 2.327 40.45 2.68 ;
      RECT 40.44 2.31 40.445 2.68 ;
      RECT 40.435 2.297 40.44 2.68 ;
      RECT 40.36 2.18 40.435 2.68 ;
      RECT 40.315 1.997 40.36 2.68 ;
      RECT 40.31 1.925 40.315 2.68 ;
      RECT 40.295 1.9 40.31 2.68 ;
      RECT 40.27 1.862 40.295 2.68 ;
      RECT 40.26 1.842 40.27 2.402 ;
      RECT 40.245 1.834 40.26 2.357 ;
      RECT 40.24 1.826 40.245 2.328 ;
      RECT 40.235 1.823 40.24 2.308 ;
      RECT 40.23 1.82 40.235 2.288 ;
      RECT 40.225 1.817 40.23 2.268 ;
      RECT 40.195 1.806 40.225 2.205 ;
      RECT 40.175 1.791 40.195 2.12 ;
      RECT 40.17 1.783 40.175 2.083 ;
      RECT 40.16 1.777 40.17 2.05 ;
      RECT 40.145 1.769 40.16 2.01 ;
      RECT 40.14 1.762 40.145 1.97 ;
      RECT 40.135 1.759 40.14 1.948 ;
      RECT 40.13 1.756 40.135 1.935 ;
      RECT 40.125 1.755 40.13 1.925 ;
      RECT 40.11 1.749 40.125 1.915 ;
      RECT 40.085 1.736 40.11 1.9 ;
      RECT 40.035 1.711 40.085 1.871 ;
      RECT 40.02 1.69 40.035 1.846 ;
      RECT 40.01 1.683 40.02 1.835 ;
      RECT 39.955 1.664 40.01 1.808 ;
      RECT 39.93 1.642 39.955 1.781 ;
      RECT 39.925 1.635 39.93 1.776 ;
      RECT 39.91 1.635 39.925 1.774 ;
      RECT 39.885 1.627 39.91 1.77 ;
      RECT 39.87 1.625 39.885 1.766 ;
      RECT 39.84 1.625 39.87 1.763 ;
      RECT 39.83 1.625 39.84 1.758 ;
      RECT 39.785 1.625 39.83 1.756 ;
      RECT 39.756 1.625 39.785 1.757 ;
      RECT 39.67 1.625 39.756 1.759 ;
      RECT 39.656 1.626 39.67 1.761 ;
      RECT 39.57 1.627 39.656 1.763 ;
      RECT 39.555 1.628 39.57 1.773 ;
      RECT 39.55 1.629 39.555 1.782 ;
      RECT 39.53 1.632 39.55 1.792 ;
      RECT 39.515 1.64 39.53 1.807 ;
      RECT 39.495 1.658 39.515 1.822 ;
      RECT 39.485 1.67 39.495 1.845 ;
      RECT 39.475 1.679 39.485 1.875 ;
      RECT 39.46 1.691 39.475 1.92 ;
      RECT 39.405 1.724 39.46 2.235 ;
      RECT 39.4 1.752 39.405 2.235 ;
      RECT 39.38 1.767 39.4 2.235 ;
      RECT 39.345 1.827 39.38 2.235 ;
      RECT 39.343 1.877 39.345 2.235 ;
      RECT 39.34 1.885 39.343 2.235 ;
      RECT 39.33 1.9 39.34 2.235 ;
      RECT 39.325 1.912 39.33 2.235 ;
      RECT 39.315 1.937 39.325 2.235 ;
      RECT 39.305 1.965 39.315 2.235 ;
      RECT 37.21 3.47 37.26 3.73 ;
      RECT 40.12 3.02 40.18 3.28 ;
      RECT 40.105 3.02 40.12 3.29 ;
      RECT 40.086 3.02 40.105 3.323 ;
      RECT 40 3.02 40.086 3.448 ;
      RECT 39.92 3.02 40 3.63 ;
      RECT 39.915 3.257 39.92 3.715 ;
      RECT 39.89 3.327 39.915 3.743 ;
      RECT 39.885 3.397 39.89 3.77 ;
      RECT 39.865 3.469 39.885 3.792 ;
      RECT 39.86 3.536 39.865 3.815 ;
      RECT 39.85 3.565 39.86 3.83 ;
      RECT 39.84 3.587 39.85 3.847 ;
      RECT 39.835 3.597 39.84 3.858 ;
      RECT 39.83 3.605 39.835 3.866 ;
      RECT 39.82 3.613 39.83 3.878 ;
      RECT 39.815 3.625 39.82 3.888 ;
      RECT 39.81 3.633 39.815 3.893 ;
      RECT 39.79 3.651 39.81 3.903 ;
      RECT 39.785 3.668 39.79 3.91 ;
      RECT 39.78 3.676 39.785 3.911 ;
      RECT 39.775 3.687 39.78 3.913 ;
      RECT 39.735 3.725 39.775 3.923 ;
      RECT 39.73 3.76 39.735 3.934 ;
      RECT 39.725 3.765 39.73 3.937 ;
      RECT 39.7 3.775 39.725 3.944 ;
      RECT 39.69 3.789 39.7 3.953 ;
      RECT 39.67 3.801 39.69 3.956 ;
      RECT 39.62 3.82 39.67 3.96 ;
      RECT 39.575 3.835 39.62 3.965 ;
      RECT 39.51 3.838 39.575 3.971 ;
      RECT 39.495 3.836 39.51 3.978 ;
      RECT 39.465 3.835 39.495 3.978 ;
      RECT 39.426 3.834 39.465 3.974 ;
      RECT 39.34 3.831 39.426 3.97 ;
      RECT 39.323 3.829 39.34 3.967 ;
      RECT 39.237 3.827 39.323 3.964 ;
      RECT 39.151 3.824 39.237 3.958 ;
      RECT 39.065 3.82 39.151 3.953 ;
      RECT 38.987 3.817 39.065 3.949 ;
      RECT 38.901 3.814 38.987 3.947 ;
      RECT 38.815 3.811 38.901 3.944 ;
      RECT 38.757 3.809 38.815 3.941 ;
      RECT 38.671 3.806 38.757 3.939 ;
      RECT 38.585 3.802 38.671 3.937 ;
      RECT 38.499 3.799 38.585 3.934 ;
      RECT 38.413 3.795 38.499 3.932 ;
      RECT 38.327 3.791 38.413 3.929 ;
      RECT 38.241 3.788 38.327 3.927 ;
      RECT 38.155 3.784 38.241 3.924 ;
      RECT 38.069 3.781 38.155 3.922 ;
      RECT 37.983 3.777 38.069 3.919 ;
      RECT 37.897 3.774 37.983 3.917 ;
      RECT 37.811 3.77 37.897 3.914 ;
      RECT 37.725 3.767 37.811 3.912 ;
      RECT 37.715 3.765 37.725 3.908 ;
      RECT 37.71 3.765 37.715 3.906 ;
      RECT 37.67 3.76 37.71 3.9 ;
      RECT 37.656 3.751 37.67 3.893 ;
      RECT 37.57 3.721 37.656 3.878 ;
      RECT 37.55 3.687 37.57 3.863 ;
      RECT 37.48 3.656 37.55 3.85 ;
      RECT 37.475 3.631 37.48 3.839 ;
      RECT 37.47 3.625 37.475 3.837 ;
      RECT 37.401 3.47 37.47 3.825 ;
      RECT 37.315 3.47 37.401 3.799 ;
      RECT 37.29 3.47 37.315 3.778 ;
      RECT 37.285 3.47 37.29 3.768 ;
      RECT 37.28 3.47 37.285 3.76 ;
      RECT 37.26 3.47 37.28 3.743 ;
      RECT 39.68 2.04 39.94 2.3 ;
      RECT 39.665 2.04 39.94 2.203 ;
      RECT 39.635 2.04 39.94 2.178 ;
      RECT 39.6 1.88 39.88 2.16 ;
      RECT 39.57 3.37 39.63 3.63 ;
      RECT 38.595 2.06 38.65 2.32 ;
      RECT 39.53 3.327 39.57 3.63 ;
      RECT 39.501 3.248 39.53 3.63 ;
      RECT 39.415 3.12 39.501 3.63 ;
      RECT 39.395 3 39.415 3.63 ;
      RECT 39.37 2.951 39.395 3.63 ;
      RECT 39.365 2.916 39.37 3.48 ;
      RECT 39.335 2.876 39.365 3.418 ;
      RECT 39.31 2.813 39.335 3.333 ;
      RECT 39.3 2.775 39.31 3.27 ;
      RECT 39.285 2.75 39.3 3.231 ;
      RECT 39.242 2.708 39.285 3.137 ;
      RECT 39.24 2.681 39.242 3.064 ;
      RECT 39.235 2.676 39.24 3.055 ;
      RECT 39.23 2.669 39.235 3.03 ;
      RECT 39.225 2.663 39.23 3.015 ;
      RECT 39.22 2.657 39.225 3.003 ;
      RECT 39.21 2.648 39.22 2.985 ;
      RECT 39.205 2.639 39.21 2.963 ;
      RECT 39.18 2.62 39.205 2.913 ;
      RECT 39.175 2.601 39.18 2.863 ;
      RECT 39.16 2.587 39.175 2.823 ;
      RECT 39.155 2.573 39.16 2.79 ;
      RECT 39.15 2.566 39.155 2.783 ;
      RECT 39.135 2.553 39.15 2.775 ;
      RECT 39.09 2.515 39.135 2.748 ;
      RECT 39.06 2.468 39.09 2.713 ;
      RECT 39.04 2.437 39.06 2.69 ;
      RECT 38.96 2.37 39.04 2.643 ;
      RECT 38.93 2.3 38.96 2.59 ;
      RECT 38.925 2.277 38.93 2.573 ;
      RECT 38.895 2.255 38.925 2.558 ;
      RECT 38.865 2.214 38.895 2.53 ;
      RECT 38.86 2.189 38.865 2.515 ;
      RECT 38.855 2.183 38.86 2.508 ;
      RECT 38.845 2.06 38.855 2.5 ;
      RECT 38.835 2.06 38.845 2.493 ;
      RECT 38.83 2.06 38.835 2.485 ;
      RECT 38.81 2.06 38.83 2.473 ;
      RECT 38.76 2.06 38.81 2.443 ;
      RECT 38.705 2.06 38.76 2.393 ;
      RECT 38.675 2.06 38.705 2.353 ;
      RECT 38.65 2.06 38.675 2.33 ;
      RECT 38.52 2.785 38.8 3.065 ;
      RECT 38.485 2.7 38.745 2.96 ;
      RECT 38.485 2.782 38.755 2.96 ;
      RECT 36.685 2.155 36.69 2.64 ;
      RECT 36.575 2.34 36.58 2.64 ;
      RECT 36.485 2.38 36.55 2.64 ;
      RECT 38.16 1.88 38.25 2.51 ;
      RECT 38.125 1.93 38.13 2.51 ;
      RECT 38.07 1.955 38.08 2.51 ;
      RECT 38.025 1.955 38.035 2.51 ;
      RECT 38.395 1.88 38.44 2.16 ;
      RECT 37.245 1.61 37.445 1.75 ;
      RECT 38.361 1.88 38.395 2.172 ;
      RECT 38.275 1.88 38.361 2.212 ;
      RECT 38.26 1.88 38.275 2.253 ;
      RECT 38.255 1.88 38.26 2.273 ;
      RECT 38.25 1.88 38.255 2.293 ;
      RECT 38.13 1.922 38.16 2.51 ;
      RECT 38.08 1.942 38.125 2.51 ;
      RECT 38.065 1.957 38.07 2.51 ;
      RECT 38.035 1.957 38.065 2.51 ;
      RECT 37.99 1.942 38.025 2.51 ;
      RECT 37.985 1.93 37.99 2.29 ;
      RECT 37.98 1.927 37.985 2.27 ;
      RECT 37.965 1.917 37.98 2.223 ;
      RECT 37.96 1.91 37.965 2.186 ;
      RECT 37.955 1.907 37.96 2.169 ;
      RECT 37.94 1.897 37.955 2.125 ;
      RECT 37.935 1.888 37.94 2.085 ;
      RECT 37.93 1.884 37.935 2.07 ;
      RECT 37.92 1.878 37.93 2.053 ;
      RECT 37.88 1.859 37.92 2.028 ;
      RECT 37.875 1.841 37.88 2.008 ;
      RECT 37.865 1.835 37.875 2.003 ;
      RECT 37.835 1.819 37.865 1.99 ;
      RECT 37.82 1.801 37.835 1.973 ;
      RECT 37.805 1.789 37.82 1.96 ;
      RECT 37.8 1.781 37.805 1.953 ;
      RECT 37.77 1.767 37.8 1.94 ;
      RECT 37.765 1.752 37.77 1.928 ;
      RECT 37.755 1.746 37.765 1.92 ;
      RECT 37.735 1.734 37.755 1.908 ;
      RECT 37.725 1.722 37.735 1.895 ;
      RECT 37.695 1.706 37.725 1.88 ;
      RECT 37.675 1.686 37.695 1.863 ;
      RECT 37.67 1.676 37.675 1.853 ;
      RECT 37.645 1.664 37.67 1.84 ;
      RECT 37.64 1.652 37.645 1.828 ;
      RECT 37.635 1.647 37.64 1.824 ;
      RECT 37.62 1.64 37.635 1.816 ;
      RECT 37.61 1.627 37.62 1.806 ;
      RECT 37.605 1.625 37.61 1.8 ;
      RECT 37.58 1.618 37.605 1.789 ;
      RECT 37.575 1.611 37.58 1.778 ;
      RECT 37.55 1.61 37.575 1.765 ;
      RECT 37.531 1.61 37.55 1.755 ;
      RECT 37.445 1.61 37.531 1.752 ;
      RECT 37.215 1.61 37.245 1.755 ;
      RECT 37.175 1.617 37.215 1.768 ;
      RECT 37.15 1.627 37.175 1.781 ;
      RECT 37.135 1.636 37.15 1.791 ;
      RECT 37.105 1.641 37.135 1.81 ;
      RECT 37.1 1.647 37.105 1.828 ;
      RECT 37.08 1.657 37.1 1.843 ;
      RECT 37.07 1.67 37.08 1.863 ;
      RECT 37.055 1.682 37.07 1.88 ;
      RECT 37.05 1.692 37.055 1.89 ;
      RECT 37.045 1.697 37.05 1.895 ;
      RECT 37.035 1.705 37.045 1.908 ;
      RECT 36.985 1.737 37.035 1.945 ;
      RECT 36.97 1.772 36.985 1.986 ;
      RECT 36.965 1.782 36.97 2.001 ;
      RECT 36.96 1.787 36.965 2.008 ;
      RECT 36.935 1.803 36.96 2.028 ;
      RECT 36.92 1.824 36.935 2.053 ;
      RECT 36.895 1.845 36.92 2.078 ;
      RECT 36.885 1.864 36.895 2.101 ;
      RECT 36.86 1.882 36.885 2.124 ;
      RECT 36.845 1.902 36.86 2.148 ;
      RECT 36.84 1.912 36.845 2.16 ;
      RECT 36.825 1.924 36.84 2.18 ;
      RECT 36.815 1.939 36.825 2.22 ;
      RECT 36.81 1.947 36.815 2.248 ;
      RECT 36.8 1.957 36.81 2.268 ;
      RECT 36.795 1.97 36.8 2.293 ;
      RECT 36.79 1.983 36.795 2.313 ;
      RECT 36.785 1.989 36.79 2.335 ;
      RECT 36.775 1.998 36.785 2.355 ;
      RECT 36.77 2.018 36.775 2.378 ;
      RECT 36.765 2.024 36.77 2.398 ;
      RECT 36.76 2.031 36.765 2.42 ;
      RECT 36.755 2.042 36.76 2.433 ;
      RECT 36.745 2.052 36.755 2.458 ;
      RECT 36.725 2.077 36.745 2.64 ;
      RECT 36.695 2.117 36.725 2.64 ;
      RECT 36.69 2.147 36.695 2.64 ;
      RECT 36.665 2.175 36.685 2.64 ;
      RECT 36.635 2.22 36.665 2.64 ;
      RECT 36.63 2.247 36.635 2.64 ;
      RECT 36.61 2.265 36.63 2.64 ;
      RECT 36.6 2.29 36.61 2.64 ;
      RECT 36.595 2.302 36.6 2.64 ;
      RECT 36.58 2.325 36.595 2.64 ;
      RECT 36.56 2.352 36.575 2.64 ;
      RECT 36.55 2.375 36.56 2.64 ;
      RECT 38.34 3.26 38.42 3.52 ;
      RECT 37.575 2.48 37.645 2.74 ;
      RECT 38.306 3.227 38.34 3.52 ;
      RECT 38.22 3.13 38.306 3.52 ;
      RECT 38.2 3.042 38.22 3.52 ;
      RECT 38.19 3.012 38.2 3.52 ;
      RECT 38.18 2.992 38.19 3.52 ;
      RECT 38.16 2.979 38.18 3.52 ;
      RECT 38.145 2.969 38.16 3.348 ;
      RECT 38.14 2.962 38.145 3.303 ;
      RECT 38.13 2.956 38.14 3.293 ;
      RECT 38.12 2.948 38.13 3.275 ;
      RECT 38.115 2.942 38.12 3.263 ;
      RECT 38.105 2.937 38.115 3.25 ;
      RECT 38.085 2.927 38.105 3.223 ;
      RECT 38.045 2.906 38.085 3.175 ;
      RECT 38.03 2.887 38.045 3.133 ;
      RECT 38.005 2.873 38.03 3.103 ;
      RECT 37.995 2.861 38.005 3.07 ;
      RECT 37.99 2.856 37.995 3.06 ;
      RECT 37.96 2.842 37.99 3.04 ;
      RECT 37.95 2.826 37.96 3.013 ;
      RECT 37.945 2.821 37.95 3.003 ;
      RECT 37.92 2.812 37.945 2.983 ;
      RECT 37.91 2.8 37.92 2.963 ;
      RECT 37.84 2.768 37.91 2.938 ;
      RECT 37.835 2.737 37.84 2.915 ;
      RECT 37.786 2.48 37.835 2.898 ;
      RECT 37.7 2.48 37.786 2.857 ;
      RECT 37.645 2.48 37.7 2.785 ;
      RECT 37.735 3.265 37.895 3.525 ;
      RECT 37.26 1.88 37.31 2.565 ;
      RECT 37.05 2.305 37.085 2.565 ;
      RECT 37.365 1.88 37.37 2.34 ;
      RECT 37.455 1.88 37.48 2.16 ;
      RECT 37.73 3.262 37.735 3.525 ;
      RECT 37.695 3.25 37.73 3.525 ;
      RECT 37.635 3.223 37.695 3.525 ;
      RECT 37.63 3.206 37.635 3.379 ;
      RECT 37.625 3.203 37.63 3.366 ;
      RECT 37.605 3.196 37.625 3.353 ;
      RECT 37.57 3.179 37.605 3.335 ;
      RECT 37.53 3.158 37.57 3.315 ;
      RECT 37.525 3.146 37.53 3.303 ;
      RECT 37.485 3.132 37.525 3.289 ;
      RECT 37.465 3.115 37.485 3.271 ;
      RECT 37.455 3.107 37.465 3.263 ;
      RECT 37.44 1.88 37.455 2.178 ;
      RECT 37.425 3.097 37.455 3.25 ;
      RECT 37.41 1.88 37.44 2.223 ;
      RECT 37.415 3.087 37.425 3.237 ;
      RECT 37.385 3.072 37.415 3.224 ;
      RECT 37.37 1.88 37.41 2.29 ;
      RECT 37.37 3.04 37.385 3.21 ;
      RECT 37.365 3.012 37.37 3.204 ;
      RECT 37.36 1.88 37.365 2.345 ;
      RECT 37.35 2.982 37.365 3.198 ;
      RECT 37.355 1.88 37.36 2.358 ;
      RECT 37.345 1.88 37.355 2.378 ;
      RECT 37.31 2.895 37.35 3.183 ;
      RECT 37.31 1.88 37.345 2.418 ;
      RECT 37.305 2.827 37.31 3.171 ;
      RECT 37.29 2.782 37.305 3.166 ;
      RECT 37.285 2.72 37.29 3.161 ;
      RECT 37.26 2.627 37.285 3.154 ;
      RECT 37.255 1.88 37.26 3.146 ;
      RECT 37.24 1.88 37.255 3.133 ;
      RECT 37.22 1.88 37.24 3.09 ;
      RECT 37.21 1.88 37.22 3.04 ;
      RECT 37.205 1.88 37.21 3.013 ;
      RECT 37.2 1.88 37.205 2.991 ;
      RECT 37.195 2.106 37.2 2.974 ;
      RECT 37.19 2.128 37.195 2.952 ;
      RECT 37.185 2.17 37.19 2.935 ;
      RECT 37.155 2.22 37.185 2.879 ;
      RECT 37.15 2.247 37.155 2.821 ;
      RECT 37.135 2.265 37.15 2.785 ;
      RECT 37.13 2.283 37.135 2.749 ;
      RECT 37.124 2.29 37.13 2.73 ;
      RECT 37.12 2.297 37.124 2.713 ;
      RECT 37.115 2.302 37.12 2.682 ;
      RECT 37.105 2.305 37.115 2.657 ;
      RECT 37.095 2.305 37.105 2.623 ;
      RECT 37.09 2.305 37.095 2.6 ;
      RECT 37.085 2.305 37.09 2.58 ;
      RECT 36 2.44 36.28 2.72 ;
      RECT 36 2.44 36.3 2.615 ;
      RECT 36.09 2.33 36.35 2.59 ;
      RECT 36.055 2.425 36.35 2.59 ;
      RECT 36.18 0.945 36.345 2.59 ;
      RECT 36.08 0.945 36.45 1.315 ;
      RECT 35.705 3.47 35.965 3.73 ;
      RECT 35.725 3.397 35.905 3.73 ;
      RECT 35.725 3.14 35.9 3.73 ;
      RECT 35.725 2.932 35.89 3.73 ;
      RECT 35.73 2.85 35.89 3.73 ;
      RECT 35.73 2.615 35.88 3.73 ;
      RECT 35.73 2.462 35.875 3.73 ;
      RECT 35.735 2.447 35.875 3.73 ;
      RECT 35.785 2.162 35.875 3.73 ;
      RECT 35.74 2.397 35.875 3.73 ;
      RECT 35.77 2.215 35.875 3.73 ;
      RECT 35.755 2.327 35.875 3.73 ;
      RECT 35.76 2.285 35.875 3.73 ;
      RECT 35.755 2.327 35.89 2.39 ;
      RECT 35.79 1.915 35.895 2.335 ;
      RECT 35.79 1.915 35.91 2.318 ;
      RECT 35.79 1.915 35.945 2.28 ;
      RECT 35.785 2.162 35.995 2.213 ;
      RECT 35.79 1.915 36.05 2.175 ;
      RECT 35.05 2.62 35.31 2.88 ;
      RECT 35.05 2.62 35.32 2.838 ;
      RECT 35.05 2.62 35.406 2.809 ;
      RECT 35.05 2.62 35.475 2.761 ;
      RECT 35.05 2.62 35.51 2.73 ;
      RECT 35.28 2.44 35.56 2.72 ;
      RECT 35.115 2.605 35.56 2.72 ;
      RECT 35.205 2.482 35.31 2.88 ;
      RECT 35.135 2.545 35.56 2.72 ;
      RECT 29.585 6.22 29.905 6.545 ;
      RECT 29.615 5.695 29.785 6.545 ;
      RECT 29.615 5.695 29.79 6.045 ;
      RECT 29.615 5.695 30.59 5.87 ;
      RECT 30.415 1.965 30.59 5.87 ;
      RECT 30.36 1.965 30.71 2.315 ;
      RECT 30.385 6.655 30.71 6.98 ;
      RECT 29.27 6.745 30.71 6.915 ;
      RECT 29.27 2.395 29.43 6.915 ;
      RECT 29.585 2.365 29.905 2.685 ;
      RECT 29.27 2.395 29.905 2.565 ;
      RECT 27.98 2.705 28.32 3.055 ;
      RECT 27.375 2.77 28.32 2.97 ;
      RECT 27.375 2.765 27.59 2.97 ;
      RECT 27.39 2.34 27.59 2.97 ;
      RECT 26.38 2.34 26.66 2.72 ;
      RECT 28.07 2.7 28.24 3.055 ;
      RECT 26.375 2.34 26.66 2.673 ;
      RECT 26.355 2.34 26.66 2.65 ;
      RECT 26.345 2.34 26.66 2.63 ;
      RECT 26.335 2.34 26.66 2.615 ;
      RECT 26.31 2.34 26.66 2.588 ;
      RECT 26.3 2.34 26.66 2.563 ;
      RECT 26.255 2.295 26.535 2.555 ;
      RECT 26.255 2.34 27.59 2.54 ;
      RECT 26.255 2.335 26.58 2.555 ;
      RECT 26.255 2.327 26.575 2.555 ;
      RECT 26.255 2.317 26.57 2.555 ;
      RECT 26.255 2.305 26.565 2.555 ;
      RECT 25.18 3 25.46 3.28 ;
      RECT 25.18 3 25.495 3.26 ;
      RECT 17.505 6.655 17.855 7.005 ;
      RECT 24.925 6.61 25.275 6.96 ;
      RECT 17.505 6.685 25.275 6.885 ;
      RECT 25.215 2.42 25.265 2.68 ;
      RECT 25.005 2.42 25.01 2.68 ;
      RECT 24.2 1.975 24.23 2.235 ;
      RECT 23.97 1.975 24.045 2.235 ;
      RECT 25.19 2.37 25.215 2.68 ;
      RECT 25.185 2.327 25.19 2.68 ;
      RECT 25.18 2.31 25.185 2.68 ;
      RECT 25.175 2.297 25.18 2.68 ;
      RECT 25.1 2.18 25.175 2.68 ;
      RECT 25.055 1.997 25.1 2.68 ;
      RECT 25.05 1.925 25.055 2.68 ;
      RECT 25.035 1.9 25.05 2.68 ;
      RECT 25.01 1.862 25.035 2.68 ;
      RECT 25 1.842 25.01 2.402 ;
      RECT 24.985 1.834 25 2.357 ;
      RECT 24.98 1.826 24.985 2.328 ;
      RECT 24.975 1.823 24.98 2.308 ;
      RECT 24.97 1.82 24.975 2.288 ;
      RECT 24.965 1.817 24.97 2.268 ;
      RECT 24.935 1.806 24.965 2.205 ;
      RECT 24.915 1.791 24.935 2.12 ;
      RECT 24.91 1.783 24.915 2.083 ;
      RECT 24.9 1.777 24.91 2.05 ;
      RECT 24.885 1.769 24.9 2.01 ;
      RECT 24.88 1.762 24.885 1.97 ;
      RECT 24.875 1.759 24.88 1.948 ;
      RECT 24.87 1.756 24.875 1.935 ;
      RECT 24.865 1.755 24.87 1.925 ;
      RECT 24.85 1.749 24.865 1.915 ;
      RECT 24.825 1.736 24.85 1.9 ;
      RECT 24.775 1.711 24.825 1.871 ;
      RECT 24.76 1.69 24.775 1.846 ;
      RECT 24.75 1.683 24.76 1.835 ;
      RECT 24.695 1.664 24.75 1.808 ;
      RECT 24.67 1.642 24.695 1.781 ;
      RECT 24.665 1.635 24.67 1.776 ;
      RECT 24.65 1.635 24.665 1.774 ;
      RECT 24.625 1.627 24.65 1.77 ;
      RECT 24.61 1.625 24.625 1.766 ;
      RECT 24.58 1.625 24.61 1.763 ;
      RECT 24.57 1.625 24.58 1.758 ;
      RECT 24.525 1.625 24.57 1.756 ;
      RECT 24.496 1.625 24.525 1.757 ;
      RECT 24.41 1.625 24.496 1.759 ;
      RECT 24.396 1.626 24.41 1.761 ;
      RECT 24.31 1.627 24.396 1.763 ;
      RECT 24.295 1.628 24.31 1.773 ;
      RECT 24.29 1.629 24.295 1.782 ;
      RECT 24.27 1.632 24.29 1.792 ;
      RECT 24.255 1.64 24.27 1.807 ;
      RECT 24.235 1.658 24.255 1.822 ;
      RECT 24.225 1.67 24.235 1.845 ;
      RECT 24.215 1.679 24.225 1.875 ;
      RECT 24.2 1.691 24.215 1.92 ;
      RECT 24.145 1.724 24.2 2.235 ;
      RECT 24.14 1.752 24.145 2.235 ;
      RECT 24.12 1.767 24.14 2.235 ;
      RECT 24.085 1.827 24.12 2.235 ;
      RECT 24.083 1.877 24.085 2.235 ;
      RECT 24.08 1.885 24.083 2.235 ;
      RECT 24.07 1.9 24.08 2.235 ;
      RECT 24.065 1.912 24.07 2.235 ;
      RECT 24.055 1.937 24.065 2.235 ;
      RECT 24.045 1.965 24.055 2.235 ;
      RECT 21.95 3.47 22 3.73 ;
      RECT 24.86 3.02 24.92 3.28 ;
      RECT 24.845 3.02 24.86 3.29 ;
      RECT 24.826 3.02 24.845 3.323 ;
      RECT 24.74 3.02 24.826 3.448 ;
      RECT 24.66 3.02 24.74 3.63 ;
      RECT 24.655 3.257 24.66 3.715 ;
      RECT 24.63 3.327 24.655 3.743 ;
      RECT 24.625 3.397 24.63 3.77 ;
      RECT 24.605 3.469 24.625 3.792 ;
      RECT 24.6 3.536 24.605 3.815 ;
      RECT 24.59 3.565 24.6 3.83 ;
      RECT 24.58 3.587 24.59 3.847 ;
      RECT 24.575 3.597 24.58 3.858 ;
      RECT 24.57 3.605 24.575 3.866 ;
      RECT 24.56 3.613 24.57 3.878 ;
      RECT 24.555 3.625 24.56 3.888 ;
      RECT 24.55 3.633 24.555 3.893 ;
      RECT 24.53 3.651 24.55 3.903 ;
      RECT 24.525 3.668 24.53 3.91 ;
      RECT 24.52 3.676 24.525 3.911 ;
      RECT 24.515 3.687 24.52 3.913 ;
      RECT 24.475 3.725 24.515 3.923 ;
      RECT 24.47 3.76 24.475 3.934 ;
      RECT 24.465 3.765 24.47 3.937 ;
      RECT 24.44 3.775 24.465 3.944 ;
      RECT 24.43 3.789 24.44 3.953 ;
      RECT 24.41 3.801 24.43 3.956 ;
      RECT 24.36 3.82 24.41 3.96 ;
      RECT 24.315 3.835 24.36 3.965 ;
      RECT 24.25 3.838 24.315 3.971 ;
      RECT 24.235 3.836 24.25 3.978 ;
      RECT 24.205 3.835 24.235 3.978 ;
      RECT 24.166 3.834 24.205 3.974 ;
      RECT 24.08 3.831 24.166 3.97 ;
      RECT 24.063 3.829 24.08 3.967 ;
      RECT 23.977 3.827 24.063 3.964 ;
      RECT 23.891 3.824 23.977 3.958 ;
      RECT 23.805 3.82 23.891 3.953 ;
      RECT 23.727 3.817 23.805 3.949 ;
      RECT 23.641 3.814 23.727 3.947 ;
      RECT 23.555 3.811 23.641 3.944 ;
      RECT 23.497 3.809 23.555 3.941 ;
      RECT 23.411 3.806 23.497 3.939 ;
      RECT 23.325 3.802 23.411 3.937 ;
      RECT 23.239 3.799 23.325 3.934 ;
      RECT 23.153 3.795 23.239 3.932 ;
      RECT 23.067 3.791 23.153 3.929 ;
      RECT 22.981 3.788 23.067 3.927 ;
      RECT 22.895 3.784 22.981 3.924 ;
      RECT 22.809 3.781 22.895 3.922 ;
      RECT 22.723 3.777 22.809 3.919 ;
      RECT 22.637 3.774 22.723 3.917 ;
      RECT 22.551 3.77 22.637 3.914 ;
      RECT 22.465 3.767 22.551 3.912 ;
      RECT 22.455 3.765 22.465 3.908 ;
      RECT 22.45 3.765 22.455 3.906 ;
      RECT 22.41 3.76 22.45 3.9 ;
      RECT 22.396 3.751 22.41 3.893 ;
      RECT 22.31 3.721 22.396 3.878 ;
      RECT 22.29 3.687 22.31 3.863 ;
      RECT 22.22 3.656 22.29 3.85 ;
      RECT 22.215 3.631 22.22 3.839 ;
      RECT 22.21 3.625 22.215 3.837 ;
      RECT 22.141 3.47 22.21 3.825 ;
      RECT 22.055 3.47 22.141 3.799 ;
      RECT 22.03 3.47 22.055 3.778 ;
      RECT 22.025 3.47 22.03 3.768 ;
      RECT 22.02 3.47 22.025 3.76 ;
      RECT 22 3.47 22.02 3.743 ;
      RECT 24.42 2.04 24.68 2.3 ;
      RECT 24.405 2.04 24.68 2.203 ;
      RECT 24.375 2.04 24.68 2.178 ;
      RECT 24.34 1.88 24.62 2.16 ;
      RECT 24.31 3.37 24.37 3.63 ;
      RECT 23.335 2.06 23.39 2.32 ;
      RECT 24.27 3.327 24.31 3.63 ;
      RECT 24.241 3.248 24.27 3.63 ;
      RECT 24.155 3.12 24.241 3.63 ;
      RECT 24.135 3 24.155 3.63 ;
      RECT 24.11 2.951 24.135 3.63 ;
      RECT 24.105 2.916 24.11 3.48 ;
      RECT 24.075 2.876 24.105 3.418 ;
      RECT 24.05 2.813 24.075 3.333 ;
      RECT 24.04 2.775 24.05 3.27 ;
      RECT 24.025 2.75 24.04 3.231 ;
      RECT 23.982 2.708 24.025 3.137 ;
      RECT 23.98 2.681 23.982 3.064 ;
      RECT 23.975 2.676 23.98 3.055 ;
      RECT 23.97 2.669 23.975 3.03 ;
      RECT 23.965 2.663 23.97 3.015 ;
      RECT 23.96 2.657 23.965 3.003 ;
      RECT 23.95 2.648 23.96 2.985 ;
      RECT 23.945 2.639 23.95 2.963 ;
      RECT 23.92 2.62 23.945 2.913 ;
      RECT 23.915 2.601 23.92 2.863 ;
      RECT 23.9 2.587 23.915 2.823 ;
      RECT 23.895 2.573 23.9 2.79 ;
      RECT 23.89 2.566 23.895 2.783 ;
      RECT 23.875 2.553 23.89 2.775 ;
      RECT 23.83 2.515 23.875 2.748 ;
      RECT 23.8 2.468 23.83 2.713 ;
      RECT 23.78 2.437 23.8 2.69 ;
      RECT 23.7 2.37 23.78 2.643 ;
      RECT 23.67 2.3 23.7 2.59 ;
      RECT 23.665 2.277 23.67 2.573 ;
      RECT 23.635 2.255 23.665 2.558 ;
      RECT 23.605 2.214 23.635 2.53 ;
      RECT 23.6 2.189 23.605 2.515 ;
      RECT 23.595 2.183 23.6 2.508 ;
      RECT 23.585 2.06 23.595 2.5 ;
      RECT 23.575 2.06 23.585 2.493 ;
      RECT 23.57 2.06 23.575 2.485 ;
      RECT 23.55 2.06 23.57 2.473 ;
      RECT 23.5 2.06 23.55 2.443 ;
      RECT 23.445 2.06 23.5 2.393 ;
      RECT 23.415 2.06 23.445 2.353 ;
      RECT 23.39 2.06 23.415 2.33 ;
      RECT 23.26 2.785 23.54 3.065 ;
      RECT 23.225 2.7 23.485 2.96 ;
      RECT 23.225 2.782 23.495 2.96 ;
      RECT 21.425 2.155 21.43 2.64 ;
      RECT 21.315 2.34 21.32 2.64 ;
      RECT 21.225 2.38 21.29 2.64 ;
      RECT 22.9 1.88 22.99 2.51 ;
      RECT 22.865 1.93 22.87 2.51 ;
      RECT 22.81 1.955 22.82 2.51 ;
      RECT 22.765 1.955 22.775 2.51 ;
      RECT 23.135 1.88 23.18 2.16 ;
      RECT 21.985 1.61 22.185 1.75 ;
      RECT 23.101 1.88 23.135 2.172 ;
      RECT 23.015 1.88 23.101 2.212 ;
      RECT 23 1.88 23.015 2.253 ;
      RECT 22.995 1.88 23 2.273 ;
      RECT 22.99 1.88 22.995 2.293 ;
      RECT 22.87 1.922 22.9 2.51 ;
      RECT 22.82 1.942 22.865 2.51 ;
      RECT 22.805 1.957 22.81 2.51 ;
      RECT 22.775 1.957 22.805 2.51 ;
      RECT 22.73 1.942 22.765 2.51 ;
      RECT 22.725 1.93 22.73 2.29 ;
      RECT 22.72 1.927 22.725 2.27 ;
      RECT 22.705 1.917 22.72 2.223 ;
      RECT 22.7 1.91 22.705 2.186 ;
      RECT 22.695 1.907 22.7 2.169 ;
      RECT 22.68 1.897 22.695 2.125 ;
      RECT 22.675 1.888 22.68 2.085 ;
      RECT 22.67 1.884 22.675 2.07 ;
      RECT 22.66 1.878 22.67 2.053 ;
      RECT 22.62 1.859 22.66 2.028 ;
      RECT 22.615 1.841 22.62 2.008 ;
      RECT 22.605 1.835 22.615 2.003 ;
      RECT 22.575 1.819 22.605 1.99 ;
      RECT 22.56 1.801 22.575 1.973 ;
      RECT 22.545 1.789 22.56 1.96 ;
      RECT 22.54 1.781 22.545 1.953 ;
      RECT 22.51 1.767 22.54 1.94 ;
      RECT 22.505 1.752 22.51 1.928 ;
      RECT 22.495 1.746 22.505 1.92 ;
      RECT 22.475 1.734 22.495 1.908 ;
      RECT 22.465 1.722 22.475 1.895 ;
      RECT 22.435 1.706 22.465 1.88 ;
      RECT 22.415 1.686 22.435 1.863 ;
      RECT 22.41 1.676 22.415 1.853 ;
      RECT 22.385 1.664 22.41 1.84 ;
      RECT 22.38 1.652 22.385 1.828 ;
      RECT 22.375 1.647 22.38 1.824 ;
      RECT 22.36 1.64 22.375 1.816 ;
      RECT 22.35 1.627 22.36 1.806 ;
      RECT 22.345 1.625 22.35 1.8 ;
      RECT 22.32 1.618 22.345 1.789 ;
      RECT 22.315 1.611 22.32 1.778 ;
      RECT 22.29 1.61 22.315 1.765 ;
      RECT 22.271 1.61 22.29 1.755 ;
      RECT 22.185 1.61 22.271 1.752 ;
      RECT 21.955 1.61 21.985 1.755 ;
      RECT 21.915 1.617 21.955 1.768 ;
      RECT 21.89 1.627 21.915 1.781 ;
      RECT 21.875 1.636 21.89 1.791 ;
      RECT 21.845 1.641 21.875 1.81 ;
      RECT 21.84 1.647 21.845 1.828 ;
      RECT 21.82 1.657 21.84 1.843 ;
      RECT 21.81 1.67 21.82 1.863 ;
      RECT 21.795 1.682 21.81 1.88 ;
      RECT 21.79 1.692 21.795 1.89 ;
      RECT 21.785 1.697 21.79 1.895 ;
      RECT 21.775 1.705 21.785 1.908 ;
      RECT 21.725 1.737 21.775 1.945 ;
      RECT 21.71 1.772 21.725 1.986 ;
      RECT 21.705 1.782 21.71 2.001 ;
      RECT 21.7 1.787 21.705 2.008 ;
      RECT 21.675 1.803 21.7 2.028 ;
      RECT 21.66 1.824 21.675 2.053 ;
      RECT 21.635 1.845 21.66 2.078 ;
      RECT 21.625 1.864 21.635 2.101 ;
      RECT 21.6 1.882 21.625 2.124 ;
      RECT 21.585 1.902 21.6 2.148 ;
      RECT 21.58 1.912 21.585 2.16 ;
      RECT 21.565 1.924 21.58 2.18 ;
      RECT 21.555 1.939 21.565 2.22 ;
      RECT 21.55 1.947 21.555 2.248 ;
      RECT 21.54 1.957 21.55 2.268 ;
      RECT 21.535 1.97 21.54 2.293 ;
      RECT 21.53 1.983 21.535 2.313 ;
      RECT 21.525 1.989 21.53 2.335 ;
      RECT 21.515 1.998 21.525 2.355 ;
      RECT 21.51 2.018 21.515 2.378 ;
      RECT 21.505 2.024 21.51 2.398 ;
      RECT 21.5 2.031 21.505 2.42 ;
      RECT 21.495 2.042 21.5 2.433 ;
      RECT 21.485 2.052 21.495 2.458 ;
      RECT 21.465 2.077 21.485 2.64 ;
      RECT 21.435 2.117 21.465 2.64 ;
      RECT 21.43 2.147 21.435 2.64 ;
      RECT 21.405 2.175 21.425 2.64 ;
      RECT 21.375 2.22 21.405 2.64 ;
      RECT 21.37 2.247 21.375 2.64 ;
      RECT 21.35 2.265 21.37 2.64 ;
      RECT 21.34 2.29 21.35 2.64 ;
      RECT 21.335 2.302 21.34 2.64 ;
      RECT 21.32 2.325 21.335 2.64 ;
      RECT 21.3 2.352 21.315 2.64 ;
      RECT 21.29 2.375 21.3 2.64 ;
      RECT 23.08 3.26 23.16 3.52 ;
      RECT 22.315 2.48 22.385 2.74 ;
      RECT 23.046 3.227 23.08 3.52 ;
      RECT 22.96 3.13 23.046 3.52 ;
      RECT 22.94 3.042 22.96 3.52 ;
      RECT 22.93 3.012 22.94 3.52 ;
      RECT 22.92 2.992 22.93 3.52 ;
      RECT 22.9 2.979 22.92 3.52 ;
      RECT 22.885 2.969 22.9 3.348 ;
      RECT 22.88 2.962 22.885 3.303 ;
      RECT 22.87 2.956 22.88 3.293 ;
      RECT 22.86 2.948 22.87 3.275 ;
      RECT 22.855 2.942 22.86 3.263 ;
      RECT 22.845 2.937 22.855 3.25 ;
      RECT 22.825 2.927 22.845 3.223 ;
      RECT 22.785 2.906 22.825 3.175 ;
      RECT 22.77 2.887 22.785 3.133 ;
      RECT 22.745 2.873 22.77 3.103 ;
      RECT 22.735 2.861 22.745 3.07 ;
      RECT 22.73 2.856 22.735 3.06 ;
      RECT 22.7 2.842 22.73 3.04 ;
      RECT 22.69 2.826 22.7 3.013 ;
      RECT 22.685 2.821 22.69 3.003 ;
      RECT 22.66 2.812 22.685 2.983 ;
      RECT 22.65 2.8 22.66 2.963 ;
      RECT 22.58 2.768 22.65 2.938 ;
      RECT 22.575 2.737 22.58 2.915 ;
      RECT 22.526 2.48 22.575 2.898 ;
      RECT 22.44 2.48 22.526 2.857 ;
      RECT 22.385 2.48 22.44 2.785 ;
      RECT 22.475 3.265 22.635 3.525 ;
      RECT 22 1.88 22.05 2.565 ;
      RECT 21.79 2.305 21.825 2.565 ;
      RECT 22.105 1.88 22.11 2.34 ;
      RECT 22.195 1.88 22.22 2.16 ;
      RECT 22.47 3.262 22.475 3.525 ;
      RECT 22.435 3.25 22.47 3.525 ;
      RECT 22.375 3.223 22.435 3.525 ;
      RECT 22.37 3.206 22.375 3.379 ;
      RECT 22.365 3.203 22.37 3.366 ;
      RECT 22.345 3.196 22.365 3.353 ;
      RECT 22.31 3.179 22.345 3.335 ;
      RECT 22.27 3.158 22.31 3.315 ;
      RECT 22.265 3.146 22.27 3.303 ;
      RECT 22.225 3.132 22.265 3.289 ;
      RECT 22.205 3.115 22.225 3.271 ;
      RECT 22.195 3.107 22.205 3.263 ;
      RECT 22.18 1.88 22.195 2.178 ;
      RECT 22.165 3.097 22.195 3.25 ;
      RECT 22.15 1.88 22.18 2.223 ;
      RECT 22.155 3.087 22.165 3.237 ;
      RECT 22.125 3.072 22.155 3.224 ;
      RECT 22.11 1.88 22.15 2.29 ;
      RECT 22.11 3.04 22.125 3.21 ;
      RECT 22.105 3.012 22.11 3.204 ;
      RECT 22.1 1.88 22.105 2.345 ;
      RECT 22.09 2.982 22.105 3.198 ;
      RECT 22.095 1.88 22.1 2.358 ;
      RECT 22.085 1.88 22.095 2.378 ;
      RECT 22.05 2.895 22.09 3.183 ;
      RECT 22.05 1.88 22.085 2.418 ;
      RECT 22.045 2.827 22.05 3.171 ;
      RECT 22.03 2.782 22.045 3.166 ;
      RECT 22.025 2.72 22.03 3.161 ;
      RECT 22 2.627 22.025 3.154 ;
      RECT 21.995 1.88 22 3.146 ;
      RECT 21.98 1.88 21.995 3.133 ;
      RECT 21.96 1.88 21.98 3.09 ;
      RECT 21.95 1.88 21.96 3.04 ;
      RECT 21.945 1.88 21.95 3.013 ;
      RECT 21.94 1.88 21.945 2.991 ;
      RECT 21.935 2.106 21.94 2.974 ;
      RECT 21.93 2.128 21.935 2.952 ;
      RECT 21.925 2.17 21.93 2.935 ;
      RECT 21.895 2.22 21.925 2.879 ;
      RECT 21.89 2.247 21.895 2.821 ;
      RECT 21.875 2.265 21.89 2.785 ;
      RECT 21.87 2.283 21.875 2.749 ;
      RECT 21.864 2.29 21.87 2.73 ;
      RECT 21.86 2.297 21.864 2.713 ;
      RECT 21.855 2.302 21.86 2.682 ;
      RECT 21.845 2.305 21.855 2.657 ;
      RECT 21.835 2.305 21.845 2.623 ;
      RECT 21.83 2.305 21.835 2.6 ;
      RECT 21.825 2.305 21.83 2.58 ;
      RECT 20.74 2.44 21.02 2.72 ;
      RECT 20.74 2.44 21.04 2.615 ;
      RECT 20.83 2.33 21.09 2.59 ;
      RECT 20.795 2.425 21.09 2.59 ;
      RECT 20.92 0.945 21.085 2.59 ;
      RECT 20.82 0.945 21.19 1.315 ;
      RECT 20.445 3.47 20.705 3.73 ;
      RECT 20.465 3.397 20.645 3.73 ;
      RECT 20.465 3.14 20.64 3.73 ;
      RECT 20.465 2.932 20.63 3.73 ;
      RECT 20.47 2.85 20.63 3.73 ;
      RECT 20.47 2.615 20.62 3.73 ;
      RECT 20.47 2.462 20.615 3.73 ;
      RECT 20.475 2.447 20.615 3.73 ;
      RECT 20.525 2.162 20.615 3.73 ;
      RECT 20.48 2.397 20.615 3.73 ;
      RECT 20.51 2.215 20.615 3.73 ;
      RECT 20.495 2.327 20.615 3.73 ;
      RECT 20.5 2.285 20.615 3.73 ;
      RECT 20.495 2.327 20.63 2.39 ;
      RECT 20.53 1.915 20.635 2.335 ;
      RECT 20.53 1.915 20.65 2.318 ;
      RECT 20.53 1.915 20.685 2.28 ;
      RECT 20.525 2.162 20.735 2.213 ;
      RECT 20.53 1.915 20.79 2.175 ;
      RECT 19.79 2.62 20.05 2.88 ;
      RECT 19.79 2.62 20.06 2.838 ;
      RECT 19.79 2.62 20.146 2.809 ;
      RECT 19.79 2.62 20.215 2.761 ;
      RECT 19.79 2.62 20.25 2.73 ;
      RECT 20.02 2.44 20.3 2.72 ;
      RECT 19.855 2.605 20.3 2.72 ;
      RECT 19.945 2.482 20.05 2.88 ;
      RECT 19.875 2.545 20.3 2.72 ;
      RECT 14.325 6.22 14.645 6.545 ;
      RECT 14.355 5.695 14.525 6.545 ;
      RECT 14.355 5.695 14.53 6.045 ;
      RECT 14.355 5.695 15.33 5.87 ;
      RECT 15.155 1.965 15.33 5.87 ;
      RECT 15.1 1.965 15.45 2.315 ;
      RECT 15.125 6.655 15.45 6.98 ;
      RECT 14.01 6.745 15.45 6.915 ;
      RECT 14.01 2.395 14.17 6.915 ;
      RECT 14.325 2.365 14.645 2.685 ;
      RECT 14.01 2.395 14.645 2.565 ;
      RECT 12.72 2.705 13.06 3.055 ;
      RECT 12.115 2.77 13.06 2.97 ;
      RECT 12.115 2.765 12.33 2.97 ;
      RECT 12.13 2.34 12.33 2.97 ;
      RECT 11.12 2.34 11.4 2.72 ;
      RECT 12.81 2.7 12.98 3.055 ;
      RECT 11.115 2.34 11.4 2.673 ;
      RECT 11.095 2.34 11.4 2.65 ;
      RECT 11.085 2.34 11.4 2.63 ;
      RECT 11.075 2.34 11.4 2.615 ;
      RECT 11.05 2.34 11.4 2.588 ;
      RECT 11.04 2.34 11.4 2.563 ;
      RECT 10.995 2.295 11.275 2.555 ;
      RECT 10.995 2.34 12.33 2.54 ;
      RECT 10.995 2.335 11.32 2.555 ;
      RECT 10.995 2.327 11.315 2.555 ;
      RECT 10.995 2.317 11.31 2.555 ;
      RECT 10.995 2.305 11.305 2.555 ;
      RECT 9.92 3 10.2 3.28 ;
      RECT 9.92 3 10.235 3.26 ;
      RECT 1.54 6.995 1.83 7.345 ;
      RECT 1.54 7.055 2.87 7.225 ;
      RECT 2.7 6.685 2.87 7.225 ;
      RECT 9.665 6.605 10.015 6.955 ;
      RECT 2.7 6.685 10.015 6.855 ;
      RECT 9.955 2.42 10.005 2.68 ;
      RECT 9.745 2.42 9.75 2.68 ;
      RECT 8.94 1.975 8.97 2.235 ;
      RECT 8.71 1.975 8.785 2.235 ;
      RECT 9.93 2.37 9.955 2.68 ;
      RECT 9.925 2.327 9.93 2.68 ;
      RECT 9.92 2.31 9.925 2.68 ;
      RECT 9.915 2.297 9.92 2.68 ;
      RECT 9.84 2.18 9.915 2.68 ;
      RECT 9.795 1.997 9.84 2.68 ;
      RECT 9.79 1.925 9.795 2.68 ;
      RECT 9.775 1.9 9.79 2.68 ;
      RECT 9.75 1.862 9.775 2.68 ;
      RECT 9.74 1.842 9.75 2.402 ;
      RECT 9.725 1.834 9.74 2.357 ;
      RECT 9.72 1.826 9.725 2.328 ;
      RECT 9.715 1.823 9.72 2.308 ;
      RECT 9.71 1.82 9.715 2.288 ;
      RECT 9.705 1.817 9.71 2.268 ;
      RECT 9.675 1.806 9.705 2.205 ;
      RECT 9.655 1.791 9.675 2.12 ;
      RECT 9.65 1.783 9.655 2.083 ;
      RECT 9.64 1.777 9.65 2.05 ;
      RECT 9.625 1.769 9.64 2.01 ;
      RECT 9.62 1.762 9.625 1.97 ;
      RECT 9.615 1.759 9.62 1.948 ;
      RECT 9.61 1.756 9.615 1.935 ;
      RECT 9.605 1.755 9.61 1.925 ;
      RECT 9.59 1.749 9.605 1.915 ;
      RECT 9.565 1.736 9.59 1.9 ;
      RECT 9.515 1.711 9.565 1.871 ;
      RECT 9.5 1.69 9.515 1.846 ;
      RECT 9.49 1.683 9.5 1.835 ;
      RECT 9.435 1.664 9.49 1.808 ;
      RECT 9.41 1.642 9.435 1.781 ;
      RECT 9.405 1.635 9.41 1.776 ;
      RECT 9.39 1.635 9.405 1.774 ;
      RECT 9.365 1.627 9.39 1.77 ;
      RECT 9.35 1.625 9.365 1.766 ;
      RECT 9.32 1.625 9.35 1.763 ;
      RECT 9.31 1.625 9.32 1.758 ;
      RECT 9.265 1.625 9.31 1.756 ;
      RECT 9.236 1.625 9.265 1.757 ;
      RECT 9.15 1.625 9.236 1.759 ;
      RECT 9.136 1.626 9.15 1.761 ;
      RECT 9.05 1.627 9.136 1.763 ;
      RECT 9.035 1.628 9.05 1.773 ;
      RECT 9.03 1.629 9.035 1.782 ;
      RECT 9.01 1.632 9.03 1.792 ;
      RECT 8.995 1.64 9.01 1.807 ;
      RECT 8.975 1.658 8.995 1.822 ;
      RECT 8.965 1.67 8.975 1.845 ;
      RECT 8.955 1.679 8.965 1.875 ;
      RECT 8.94 1.691 8.955 1.92 ;
      RECT 8.885 1.724 8.94 2.235 ;
      RECT 8.88 1.752 8.885 2.235 ;
      RECT 8.86 1.767 8.88 2.235 ;
      RECT 8.825 1.827 8.86 2.235 ;
      RECT 8.823 1.877 8.825 2.235 ;
      RECT 8.82 1.885 8.823 2.235 ;
      RECT 8.81 1.9 8.82 2.235 ;
      RECT 8.805 1.912 8.81 2.235 ;
      RECT 8.795 1.937 8.805 2.235 ;
      RECT 8.785 1.965 8.795 2.235 ;
      RECT 6.69 3.47 6.74 3.73 ;
      RECT 9.6 3.02 9.66 3.28 ;
      RECT 9.585 3.02 9.6 3.29 ;
      RECT 9.566 3.02 9.585 3.323 ;
      RECT 9.48 3.02 9.566 3.448 ;
      RECT 9.4 3.02 9.48 3.63 ;
      RECT 9.395 3.257 9.4 3.715 ;
      RECT 9.37 3.327 9.395 3.743 ;
      RECT 9.365 3.397 9.37 3.77 ;
      RECT 9.345 3.469 9.365 3.792 ;
      RECT 9.34 3.536 9.345 3.815 ;
      RECT 9.33 3.565 9.34 3.83 ;
      RECT 9.32 3.587 9.33 3.847 ;
      RECT 9.315 3.597 9.32 3.858 ;
      RECT 9.31 3.605 9.315 3.866 ;
      RECT 9.3 3.613 9.31 3.878 ;
      RECT 9.295 3.625 9.3 3.888 ;
      RECT 9.29 3.633 9.295 3.893 ;
      RECT 9.27 3.651 9.29 3.903 ;
      RECT 9.265 3.668 9.27 3.91 ;
      RECT 9.26 3.676 9.265 3.911 ;
      RECT 9.255 3.687 9.26 3.913 ;
      RECT 9.215 3.725 9.255 3.923 ;
      RECT 9.21 3.76 9.215 3.934 ;
      RECT 9.205 3.765 9.21 3.937 ;
      RECT 9.18 3.775 9.205 3.944 ;
      RECT 9.17 3.789 9.18 3.953 ;
      RECT 9.15 3.801 9.17 3.956 ;
      RECT 9.1 3.82 9.15 3.96 ;
      RECT 9.055 3.835 9.1 3.965 ;
      RECT 8.99 3.838 9.055 3.971 ;
      RECT 8.975 3.836 8.99 3.978 ;
      RECT 8.945 3.835 8.975 3.978 ;
      RECT 8.906 3.834 8.945 3.974 ;
      RECT 8.82 3.831 8.906 3.97 ;
      RECT 8.803 3.829 8.82 3.967 ;
      RECT 8.717 3.827 8.803 3.964 ;
      RECT 8.631 3.824 8.717 3.958 ;
      RECT 8.545 3.82 8.631 3.953 ;
      RECT 8.467 3.817 8.545 3.949 ;
      RECT 8.381 3.814 8.467 3.947 ;
      RECT 8.295 3.811 8.381 3.944 ;
      RECT 8.237 3.809 8.295 3.941 ;
      RECT 8.151 3.806 8.237 3.939 ;
      RECT 8.065 3.802 8.151 3.937 ;
      RECT 7.979 3.799 8.065 3.934 ;
      RECT 7.893 3.795 7.979 3.932 ;
      RECT 7.807 3.791 7.893 3.929 ;
      RECT 7.721 3.788 7.807 3.927 ;
      RECT 7.635 3.784 7.721 3.924 ;
      RECT 7.549 3.781 7.635 3.922 ;
      RECT 7.463 3.777 7.549 3.919 ;
      RECT 7.377 3.774 7.463 3.917 ;
      RECT 7.291 3.77 7.377 3.914 ;
      RECT 7.205 3.767 7.291 3.912 ;
      RECT 7.195 3.765 7.205 3.908 ;
      RECT 7.19 3.765 7.195 3.906 ;
      RECT 7.15 3.76 7.19 3.9 ;
      RECT 7.136 3.751 7.15 3.893 ;
      RECT 7.05 3.721 7.136 3.878 ;
      RECT 7.03 3.687 7.05 3.863 ;
      RECT 6.96 3.656 7.03 3.85 ;
      RECT 6.955 3.631 6.96 3.839 ;
      RECT 6.95 3.625 6.955 3.837 ;
      RECT 6.881 3.47 6.95 3.825 ;
      RECT 6.795 3.47 6.881 3.799 ;
      RECT 6.77 3.47 6.795 3.778 ;
      RECT 6.765 3.47 6.77 3.768 ;
      RECT 6.76 3.47 6.765 3.76 ;
      RECT 6.74 3.47 6.76 3.743 ;
      RECT 9.16 2.04 9.42 2.3 ;
      RECT 9.145 2.04 9.42 2.203 ;
      RECT 9.115 2.04 9.42 2.178 ;
      RECT 9.08 1.88 9.36 2.16 ;
      RECT 9.05 3.37 9.11 3.63 ;
      RECT 8.075 2.06 8.13 2.32 ;
      RECT 9.01 3.327 9.05 3.63 ;
      RECT 8.981 3.248 9.01 3.63 ;
      RECT 8.895 3.12 8.981 3.63 ;
      RECT 8.875 3 8.895 3.63 ;
      RECT 8.85 2.951 8.875 3.63 ;
      RECT 8.845 2.916 8.85 3.48 ;
      RECT 8.815 2.876 8.845 3.418 ;
      RECT 8.79 2.813 8.815 3.333 ;
      RECT 8.78 2.775 8.79 3.27 ;
      RECT 8.765 2.75 8.78 3.231 ;
      RECT 8.722 2.708 8.765 3.137 ;
      RECT 8.72 2.681 8.722 3.064 ;
      RECT 8.715 2.676 8.72 3.055 ;
      RECT 8.71 2.669 8.715 3.03 ;
      RECT 8.705 2.663 8.71 3.015 ;
      RECT 8.7 2.657 8.705 3.003 ;
      RECT 8.69 2.648 8.7 2.985 ;
      RECT 8.685 2.639 8.69 2.963 ;
      RECT 8.66 2.62 8.685 2.913 ;
      RECT 8.655 2.601 8.66 2.863 ;
      RECT 8.64 2.587 8.655 2.823 ;
      RECT 8.635 2.573 8.64 2.79 ;
      RECT 8.63 2.566 8.635 2.783 ;
      RECT 8.615 2.553 8.63 2.775 ;
      RECT 8.57 2.515 8.615 2.748 ;
      RECT 8.54 2.468 8.57 2.713 ;
      RECT 8.52 2.437 8.54 2.69 ;
      RECT 8.44 2.37 8.52 2.643 ;
      RECT 8.41 2.3 8.44 2.59 ;
      RECT 8.405 2.277 8.41 2.573 ;
      RECT 8.375 2.255 8.405 2.558 ;
      RECT 8.345 2.214 8.375 2.53 ;
      RECT 8.34 2.189 8.345 2.515 ;
      RECT 8.335 2.183 8.34 2.508 ;
      RECT 8.325 2.06 8.335 2.5 ;
      RECT 8.315 2.06 8.325 2.493 ;
      RECT 8.31 2.06 8.315 2.485 ;
      RECT 8.29 2.06 8.31 2.473 ;
      RECT 8.24 2.06 8.29 2.443 ;
      RECT 8.185 2.06 8.24 2.393 ;
      RECT 8.155 2.06 8.185 2.353 ;
      RECT 8.13 2.06 8.155 2.33 ;
      RECT 8 2.785 8.28 3.065 ;
      RECT 7.965 2.7 8.225 2.96 ;
      RECT 7.965 2.782 8.235 2.96 ;
      RECT 6.165 2.155 6.17 2.64 ;
      RECT 6.055 2.34 6.06 2.64 ;
      RECT 5.965 2.38 6.03 2.64 ;
      RECT 7.64 1.88 7.73 2.51 ;
      RECT 7.605 1.93 7.61 2.51 ;
      RECT 7.55 1.955 7.56 2.51 ;
      RECT 7.505 1.955 7.515 2.51 ;
      RECT 7.875 1.88 7.92 2.16 ;
      RECT 6.725 1.61 6.925 1.75 ;
      RECT 7.841 1.88 7.875 2.172 ;
      RECT 7.755 1.88 7.841 2.212 ;
      RECT 7.74 1.88 7.755 2.253 ;
      RECT 7.735 1.88 7.74 2.273 ;
      RECT 7.73 1.88 7.735 2.293 ;
      RECT 7.61 1.922 7.64 2.51 ;
      RECT 7.56 1.942 7.605 2.51 ;
      RECT 7.545 1.957 7.55 2.51 ;
      RECT 7.515 1.957 7.545 2.51 ;
      RECT 7.47 1.942 7.505 2.51 ;
      RECT 7.465 1.93 7.47 2.29 ;
      RECT 7.46 1.927 7.465 2.27 ;
      RECT 7.445 1.917 7.46 2.223 ;
      RECT 7.44 1.91 7.445 2.186 ;
      RECT 7.435 1.907 7.44 2.169 ;
      RECT 7.42 1.897 7.435 2.125 ;
      RECT 7.415 1.888 7.42 2.085 ;
      RECT 7.41 1.884 7.415 2.07 ;
      RECT 7.4 1.878 7.41 2.053 ;
      RECT 7.36 1.859 7.4 2.028 ;
      RECT 7.355 1.841 7.36 2.008 ;
      RECT 7.345 1.835 7.355 2.003 ;
      RECT 7.315 1.819 7.345 1.99 ;
      RECT 7.3 1.801 7.315 1.973 ;
      RECT 7.285 1.789 7.3 1.96 ;
      RECT 7.28 1.781 7.285 1.953 ;
      RECT 7.25 1.767 7.28 1.94 ;
      RECT 7.245 1.752 7.25 1.928 ;
      RECT 7.235 1.746 7.245 1.92 ;
      RECT 7.215 1.734 7.235 1.908 ;
      RECT 7.205 1.722 7.215 1.895 ;
      RECT 7.175 1.706 7.205 1.88 ;
      RECT 7.155 1.686 7.175 1.863 ;
      RECT 7.15 1.676 7.155 1.853 ;
      RECT 7.125 1.664 7.15 1.84 ;
      RECT 7.12 1.652 7.125 1.828 ;
      RECT 7.115 1.647 7.12 1.824 ;
      RECT 7.1 1.64 7.115 1.816 ;
      RECT 7.09 1.627 7.1 1.806 ;
      RECT 7.085 1.625 7.09 1.8 ;
      RECT 7.06 1.618 7.085 1.789 ;
      RECT 7.055 1.611 7.06 1.778 ;
      RECT 7.03 1.61 7.055 1.765 ;
      RECT 7.011 1.61 7.03 1.755 ;
      RECT 6.925 1.61 7.011 1.752 ;
      RECT 6.695 1.61 6.725 1.755 ;
      RECT 6.655 1.617 6.695 1.768 ;
      RECT 6.63 1.627 6.655 1.781 ;
      RECT 6.615 1.636 6.63 1.791 ;
      RECT 6.585 1.641 6.615 1.81 ;
      RECT 6.58 1.647 6.585 1.828 ;
      RECT 6.56 1.657 6.58 1.843 ;
      RECT 6.55 1.67 6.56 1.863 ;
      RECT 6.535 1.682 6.55 1.88 ;
      RECT 6.53 1.692 6.535 1.89 ;
      RECT 6.525 1.697 6.53 1.895 ;
      RECT 6.515 1.705 6.525 1.908 ;
      RECT 6.465 1.737 6.515 1.945 ;
      RECT 6.45 1.772 6.465 1.986 ;
      RECT 6.445 1.782 6.45 2.001 ;
      RECT 6.44 1.787 6.445 2.008 ;
      RECT 6.415 1.803 6.44 2.028 ;
      RECT 6.4 1.824 6.415 2.053 ;
      RECT 6.375 1.845 6.4 2.078 ;
      RECT 6.365 1.864 6.375 2.101 ;
      RECT 6.34 1.882 6.365 2.124 ;
      RECT 6.325 1.902 6.34 2.148 ;
      RECT 6.32 1.912 6.325 2.16 ;
      RECT 6.305 1.924 6.32 2.18 ;
      RECT 6.295 1.939 6.305 2.22 ;
      RECT 6.29 1.947 6.295 2.248 ;
      RECT 6.28 1.957 6.29 2.268 ;
      RECT 6.275 1.97 6.28 2.293 ;
      RECT 6.27 1.983 6.275 2.313 ;
      RECT 6.265 1.989 6.27 2.335 ;
      RECT 6.255 1.998 6.265 2.355 ;
      RECT 6.25 2.018 6.255 2.378 ;
      RECT 6.245 2.024 6.25 2.398 ;
      RECT 6.24 2.031 6.245 2.42 ;
      RECT 6.235 2.042 6.24 2.433 ;
      RECT 6.225 2.052 6.235 2.458 ;
      RECT 6.205 2.077 6.225 2.64 ;
      RECT 6.175 2.117 6.205 2.64 ;
      RECT 6.17 2.147 6.175 2.64 ;
      RECT 6.145 2.175 6.165 2.64 ;
      RECT 6.115 2.22 6.145 2.64 ;
      RECT 6.11 2.247 6.115 2.64 ;
      RECT 6.09 2.265 6.11 2.64 ;
      RECT 6.08 2.29 6.09 2.64 ;
      RECT 6.075 2.302 6.08 2.64 ;
      RECT 6.06 2.325 6.075 2.64 ;
      RECT 6.04 2.352 6.055 2.64 ;
      RECT 6.03 2.375 6.04 2.64 ;
      RECT 7.82 3.26 7.9 3.52 ;
      RECT 7.055 2.48 7.125 2.74 ;
      RECT 7.786 3.227 7.82 3.52 ;
      RECT 7.7 3.13 7.786 3.52 ;
      RECT 7.68 3.042 7.7 3.52 ;
      RECT 7.67 3.012 7.68 3.52 ;
      RECT 7.66 2.992 7.67 3.52 ;
      RECT 7.64 2.979 7.66 3.52 ;
      RECT 7.625 2.969 7.64 3.348 ;
      RECT 7.62 2.962 7.625 3.303 ;
      RECT 7.61 2.956 7.62 3.293 ;
      RECT 7.6 2.948 7.61 3.275 ;
      RECT 7.595 2.942 7.6 3.263 ;
      RECT 7.585 2.937 7.595 3.25 ;
      RECT 7.565 2.927 7.585 3.223 ;
      RECT 7.525 2.906 7.565 3.175 ;
      RECT 7.51 2.887 7.525 3.133 ;
      RECT 7.485 2.873 7.51 3.103 ;
      RECT 7.475 2.861 7.485 3.07 ;
      RECT 7.47 2.856 7.475 3.06 ;
      RECT 7.44 2.842 7.47 3.04 ;
      RECT 7.43 2.826 7.44 3.013 ;
      RECT 7.425 2.821 7.43 3.003 ;
      RECT 7.4 2.812 7.425 2.983 ;
      RECT 7.39 2.8 7.4 2.963 ;
      RECT 7.32 2.768 7.39 2.938 ;
      RECT 7.315 2.737 7.32 2.915 ;
      RECT 7.266 2.48 7.315 2.898 ;
      RECT 7.18 2.48 7.266 2.857 ;
      RECT 7.125 2.48 7.18 2.785 ;
      RECT 7.215 3.265 7.375 3.525 ;
      RECT 6.74 1.88 6.79 2.565 ;
      RECT 6.53 2.305 6.565 2.565 ;
      RECT 6.845 1.88 6.85 2.34 ;
      RECT 6.935 1.88 6.96 2.16 ;
      RECT 7.21 3.262 7.215 3.525 ;
      RECT 7.175 3.25 7.21 3.525 ;
      RECT 7.115 3.223 7.175 3.525 ;
      RECT 7.11 3.206 7.115 3.379 ;
      RECT 7.105 3.203 7.11 3.366 ;
      RECT 7.085 3.196 7.105 3.353 ;
      RECT 7.05 3.179 7.085 3.335 ;
      RECT 7.01 3.158 7.05 3.315 ;
      RECT 7.005 3.146 7.01 3.303 ;
      RECT 6.965 3.132 7.005 3.289 ;
      RECT 6.945 3.115 6.965 3.271 ;
      RECT 6.935 3.107 6.945 3.263 ;
      RECT 6.92 1.88 6.935 2.178 ;
      RECT 6.905 3.097 6.935 3.25 ;
      RECT 6.89 1.88 6.92 2.223 ;
      RECT 6.895 3.087 6.905 3.237 ;
      RECT 6.865 3.072 6.895 3.224 ;
      RECT 6.85 1.88 6.89 2.29 ;
      RECT 6.85 3.04 6.865 3.21 ;
      RECT 6.845 3.012 6.85 3.204 ;
      RECT 6.84 1.88 6.845 2.345 ;
      RECT 6.83 2.982 6.845 3.198 ;
      RECT 6.835 1.88 6.84 2.358 ;
      RECT 6.825 1.88 6.835 2.378 ;
      RECT 6.79 2.895 6.83 3.183 ;
      RECT 6.79 1.88 6.825 2.418 ;
      RECT 6.785 2.827 6.79 3.171 ;
      RECT 6.77 2.782 6.785 3.166 ;
      RECT 6.765 2.72 6.77 3.161 ;
      RECT 6.74 2.627 6.765 3.154 ;
      RECT 6.735 1.88 6.74 3.146 ;
      RECT 6.72 1.88 6.735 3.133 ;
      RECT 6.7 1.88 6.72 3.09 ;
      RECT 6.69 1.88 6.7 3.04 ;
      RECT 6.685 1.88 6.69 3.013 ;
      RECT 6.68 1.88 6.685 2.991 ;
      RECT 6.675 2.106 6.68 2.974 ;
      RECT 6.67 2.128 6.675 2.952 ;
      RECT 6.665 2.17 6.67 2.935 ;
      RECT 6.635 2.22 6.665 2.879 ;
      RECT 6.63 2.247 6.635 2.821 ;
      RECT 6.615 2.265 6.63 2.785 ;
      RECT 6.61 2.283 6.615 2.749 ;
      RECT 6.604 2.29 6.61 2.73 ;
      RECT 6.6 2.297 6.604 2.713 ;
      RECT 6.595 2.302 6.6 2.682 ;
      RECT 6.585 2.305 6.595 2.657 ;
      RECT 6.575 2.305 6.585 2.623 ;
      RECT 6.57 2.305 6.575 2.6 ;
      RECT 6.565 2.305 6.57 2.58 ;
      RECT 5.48 2.44 5.76 2.72 ;
      RECT 5.48 2.44 5.78 2.615 ;
      RECT 5.57 2.33 5.83 2.59 ;
      RECT 5.535 2.425 5.83 2.59 ;
      RECT 5.66 0.945 5.825 2.59 ;
      RECT 5.56 0.945 5.93 1.315 ;
      RECT 5.185 3.47 5.445 3.73 ;
      RECT 5.205 3.397 5.385 3.73 ;
      RECT 5.205 3.14 5.38 3.73 ;
      RECT 5.205 2.932 5.37 3.73 ;
      RECT 5.21 2.85 5.37 3.73 ;
      RECT 5.21 2.615 5.36 3.73 ;
      RECT 5.21 2.462 5.355 3.73 ;
      RECT 5.215 2.447 5.355 3.73 ;
      RECT 5.265 2.162 5.355 3.73 ;
      RECT 5.22 2.397 5.355 3.73 ;
      RECT 5.25 2.215 5.355 3.73 ;
      RECT 5.235 2.327 5.355 3.73 ;
      RECT 5.24 2.285 5.355 3.73 ;
      RECT 5.235 2.327 5.37 2.39 ;
      RECT 5.27 1.915 5.375 2.335 ;
      RECT 5.27 1.915 5.39 2.318 ;
      RECT 5.27 1.915 5.425 2.28 ;
      RECT 5.265 2.162 5.475 2.213 ;
      RECT 5.27 1.915 5.53 2.175 ;
      RECT 4.53 2.62 4.79 2.88 ;
      RECT 4.53 2.62 4.8 2.838 ;
      RECT 4.53 2.62 4.886 2.809 ;
      RECT 4.53 2.62 4.955 2.761 ;
      RECT 4.53 2.62 4.99 2.73 ;
      RECT 4.76 2.44 5.04 2.72 ;
      RECT 4.595 2.605 5.04 2.72 ;
      RECT 4.685 2.482 4.79 2.88 ;
      RECT 4.615 2.545 5.04 2.72 ;
      RECT 0.195 8.51 0.575 8.89 ;
      RECT 0.235 8.49 0.405 8.89 ;
      RECT 70.035 7.055 70.405 7.425 ;
      RECT 54.775 7.055 55.145 7.425 ;
      RECT 39.515 7.055 39.885 7.425 ;
      RECT 24.255 7.055 24.625 7.425 ;
      RECT 8.995 7.055 9.365 7.425 ;
    LAYER via1 ;
      RECT 78.625 7.375 78.775 7.525 ;
      RECT 76.255 6.74 76.405 6.89 ;
      RECT 76.24 2.065 76.39 2.215 ;
      RECT 75.45 2.45 75.6 2.6 ;
      RECT 75.45 6.325 75.6 6.475 ;
      RECT 73.86 2.805 74.01 2.955 ;
      RECT 72.09 2.35 72.24 2.5 ;
      RECT 71.07 3.055 71.22 3.205 ;
      RECT 70.84 2.475 70.99 2.625 ;
      RECT 70.805 6.71 70.955 6.86 ;
      RECT 70.495 3.075 70.645 3.225 ;
      RECT 70.255 2.095 70.405 2.245 ;
      RECT 70.145 7.165 70.295 7.315 ;
      RECT 69.945 3.425 70.095 3.575 ;
      RECT 69.805 2.03 69.955 2.18 ;
      RECT 69.17 2.115 69.32 2.265 ;
      RECT 69.06 2.755 69.21 2.905 ;
      RECT 68.735 3.315 68.885 3.465 ;
      RECT 68.565 2.305 68.715 2.455 ;
      RECT 68.21 3.32 68.36 3.47 ;
      RECT 68.15 2.535 68.3 2.685 ;
      RECT 67.785 3.525 67.935 3.675 ;
      RECT 67.625 2.36 67.775 2.51 ;
      RECT 67.06 2.435 67.21 2.585 ;
      RECT 66.71 1.055 66.86 1.205 ;
      RECT 66.665 2.385 66.815 2.535 ;
      RECT 66.365 1.97 66.515 2.12 ;
      RECT 66.28 3.525 66.43 3.675 ;
      RECT 65.625 2.675 65.775 2.825 ;
      RECT 63.34 6.755 63.49 6.905 ;
      RECT 60.995 6.74 61.145 6.89 ;
      RECT 60.98 2.065 61.13 2.215 ;
      RECT 60.19 2.45 60.34 2.6 ;
      RECT 60.19 6.325 60.34 6.475 ;
      RECT 58.6 2.805 58.75 2.955 ;
      RECT 56.83 2.35 56.98 2.5 ;
      RECT 55.81 3.055 55.96 3.205 ;
      RECT 55.58 2.475 55.73 2.625 ;
      RECT 55.545 6.71 55.695 6.86 ;
      RECT 55.235 3.075 55.385 3.225 ;
      RECT 54.995 2.095 55.145 2.245 ;
      RECT 54.885 7.165 55.035 7.315 ;
      RECT 54.685 3.425 54.835 3.575 ;
      RECT 54.545 2.03 54.695 2.18 ;
      RECT 53.91 2.115 54.06 2.265 ;
      RECT 53.8 2.755 53.95 2.905 ;
      RECT 53.475 3.315 53.625 3.465 ;
      RECT 53.305 2.305 53.455 2.455 ;
      RECT 52.95 3.32 53.1 3.47 ;
      RECT 52.89 2.535 53.04 2.685 ;
      RECT 52.525 3.525 52.675 3.675 ;
      RECT 52.365 2.36 52.515 2.51 ;
      RECT 51.8 2.435 51.95 2.585 ;
      RECT 51.45 1.055 51.6 1.205 ;
      RECT 51.405 2.385 51.555 2.535 ;
      RECT 51.105 1.97 51.255 2.12 ;
      RECT 51.02 3.525 51.17 3.675 ;
      RECT 50.365 2.675 50.515 2.825 ;
      RECT 48.08 6.755 48.23 6.905 ;
      RECT 45.735 6.74 45.885 6.89 ;
      RECT 45.72 2.065 45.87 2.215 ;
      RECT 44.93 2.45 45.08 2.6 ;
      RECT 44.93 6.325 45.08 6.475 ;
      RECT 43.34 2.805 43.49 2.955 ;
      RECT 41.57 2.35 41.72 2.5 ;
      RECT 40.55 3.055 40.7 3.205 ;
      RECT 40.32 2.475 40.47 2.625 ;
      RECT 40.285 6.715 40.435 6.865 ;
      RECT 39.975 3.075 40.125 3.225 ;
      RECT 39.735 2.095 39.885 2.245 ;
      RECT 39.625 7.165 39.775 7.315 ;
      RECT 39.425 3.425 39.575 3.575 ;
      RECT 39.285 2.03 39.435 2.18 ;
      RECT 38.65 2.115 38.8 2.265 ;
      RECT 38.54 2.755 38.69 2.905 ;
      RECT 38.215 3.315 38.365 3.465 ;
      RECT 38.045 2.305 38.195 2.455 ;
      RECT 37.69 3.32 37.84 3.47 ;
      RECT 37.63 2.535 37.78 2.685 ;
      RECT 37.265 3.525 37.415 3.675 ;
      RECT 37.105 2.36 37.255 2.51 ;
      RECT 36.54 2.435 36.69 2.585 ;
      RECT 36.19 1.055 36.34 1.205 ;
      RECT 36.145 2.385 36.295 2.535 ;
      RECT 35.845 1.97 35.995 2.12 ;
      RECT 35.76 3.525 35.91 3.675 ;
      RECT 35.105 2.675 35.255 2.825 ;
      RECT 32.865 6.76 33.015 6.91 ;
      RECT 30.475 6.74 30.625 6.89 ;
      RECT 30.46 2.065 30.61 2.215 ;
      RECT 29.67 2.45 29.82 2.6 ;
      RECT 29.67 6.325 29.82 6.475 ;
      RECT 28.08 2.805 28.23 2.955 ;
      RECT 26.31 2.35 26.46 2.5 ;
      RECT 25.29 3.055 25.44 3.205 ;
      RECT 25.06 2.475 25.21 2.625 ;
      RECT 25.025 6.71 25.175 6.86 ;
      RECT 24.715 3.075 24.865 3.225 ;
      RECT 24.475 2.095 24.625 2.245 ;
      RECT 24.365 7.165 24.515 7.315 ;
      RECT 24.165 3.425 24.315 3.575 ;
      RECT 24.025 2.03 24.175 2.18 ;
      RECT 23.39 2.115 23.54 2.265 ;
      RECT 23.28 2.755 23.43 2.905 ;
      RECT 22.955 3.315 23.105 3.465 ;
      RECT 22.785 2.305 22.935 2.455 ;
      RECT 22.43 3.32 22.58 3.47 ;
      RECT 22.37 2.535 22.52 2.685 ;
      RECT 22.005 3.525 22.155 3.675 ;
      RECT 21.845 2.36 21.995 2.51 ;
      RECT 21.28 2.435 21.43 2.585 ;
      RECT 20.93 1.055 21.08 1.205 ;
      RECT 20.885 2.385 21.035 2.535 ;
      RECT 20.585 1.97 20.735 2.12 ;
      RECT 20.5 3.525 20.65 3.675 ;
      RECT 19.845 2.675 19.995 2.825 ;
      RECT 17.605 6.755 17.755 6.905 ;
      RECT 15.215 6.74 15.365 6.89 ;
      RECT 15.2 2.065 15.35 2.215 ;
      RECT 14.41 2.45 14.56 2.6 ;
      RECT 14.41 6.325 14.56 6.475 ;
      RECT 12.82 2.805 12.97 2.955 ;
      RECT 11.05 2.35 11.2 2.5 ;
      RECT 10.03 3.055 10.18 3.205 ;
      RECT 9.8 2.475 9.95 2.625 ;
      RECT 9.765 6.705 9.915 6.855 ;
      RECT 9.455 3.075 9.605 3.225 ;
      RECT 9.215 2.095 9.365 2.245 ;
      RECT 9.105 7.165 9.255 7.315 ;
      RECT 8.905 3.425 9.055 3.575 ;
      RECT 8.765 2.03 8.915 2.18 ;
      RECT 8.13 2.115 8.28 2.265 ;
      RECT 8.02 2.755 8.17 2.905 ;
      RECT 7.695 3.315 7.845 3.465 ;
      RECT 7.525 2.305 7.675 2.455 ;
      RECT 7.17 3.32 7.32 3.47 ;
      RECT 7.11 2.535 7.26 2.685 ;
      RECT 6.745 3.525 6.895 3.675 ;
      RECT 6.585 2.36 6.735 2.51 ;
      RECT 6.02 2.435 6.17 2.585 ;
      RECT 5.67 1.055 5.82 1.205 ;
      RECT 5.625 2.385 5.775 2.535 ;
      RECT 5.325 1.97 5.475 2.12 ;
      RECT 5.24 3.525 5.39 3.675 ;
      RECT 4.585 2.675 4.735 2.825 ;
      RECT 1.61 7.095 1.76 7.245 ;
      RECT 1.235 6.355 1.385 6.505 ;
      RECT 0.31 8.625 0.46 8.775 ;
    LAYER met1 ;
      RECT 64.585 0 73.325 1.74 ;
      RECT 49.325 0 58.065 1.74 ;
      RECT 34.065 0 42.805 1.74 ;
      RECT 18.805 0 27.545 1.74 ;
      RECT 3.545 0 12.285 1.74 ;
      RECT 78.915 0 79.095 0.305 ;
      RECT 63.655 0 76.965 0.305 ;
      RECT 48.395 0 61.705 0.305 ;
      RECT 33.135 0 46.445 0.305 ;
      RECT 17.875 0 31.185 0.305 ;
      RECT 0 0 15.925 0.305 ;
      RECT 0 0 79.095 0.3 ;
      RECT 0.005 8.575 0.81 8.89 ;
      RECT 0 8.58 79.095 8.88 ;
      RECT 78.915 8.575 79.095 8.88 ;
      RECT 63.655 8.575 76.965 8.88 ;
      RECT 48.395 8.575 61.705 8.88 ;
      RECT 33.135 8.575 46.445 8.88 ;
      RECT 17.875 8.575 31.185 8.88 ;
      RECT 0 8.575 15.925 8.88 ;
      RECT 69.53 6.315 69.7 8.88 ;
      RECT 54.27 6.315 54.44 8.88 ;
      RECT 39.01 6.315 39.18 8.88 ;
      RECT 23.75 6.315 23.92 8.88 ;
      RECT 8.49 6.315 8.66 8.88 ;
      RECT 0.21 8.555 0.56 8.89 ;
      RECT 69.7 6.285 69.99 6.515 ;
      RECT 54.44 6.285 54.73 6.515 ;
      RECT 39.18 6.285 39.47 6.515 ;
      RECT 23.92 6.285 24.21 6.515 ;
      RECT 8.66 6.285 8.95 6.515 ;
      RECT 78.49 7.77 78.78 8 ;
      RECT 78.55 6.29 78.72 8 ;
      RECT 78.525 7.275 78.875 7.625 ;
      RECT 78.49 6.29 78.78 6.52 ;
      RECT 78.085 2.395 78.19 2.965 ;
      RECT 78.085 2.73 78.41 2.96 ;
      RECT 78.085 2.76 78.58 2.93 ;
      RECT 78.085 2.395 78.275 2.96 ;
      RECT 77.5 2.36 77.79 2.59 ;
      RECT 77.5 2.395 78.275 2.565 ;
      RECT 77.56 0.88 77.73 2.59 ;
      RECT 77.5 0.88 77.79 1.11 ;
      RECT 77.5 7.77 77.79 8 ;
      RECT 77.56 6.29 77.73 8 ;
      RECT 77.5 6.29 77.79 6.52 ;
      RECT 77.5 6.325 78.355 6.485 ;
      RECT 78.185 5.92 78.355 6.485 ;
      RECT 77.5 6.32 77.895 6.485 ;
      RECT 78.12 5.92 78.41 6.15 ;
      RECT 78.12 5.95 78.58 6.12 ;
      RECT 77.13 2.73 77.42 2.96 ;
      RECT 77.13 2.76 77.59 2.93 ;
      RECT 77.195 1.655 77.36 2.96 ;
      RECT 75.71 1.625 76 1.855 ;
      RECT 75.71 1.655 77.36 1.825 ;
      RECT 75.77 0.885 75.94 1.855 ;
      RECT 75.71 0.885 76 1.115 ;
      RECT 75.71 7.765 76 7.995 ;
      RECT 75.77 7.025 75.94 7.995 ;
      RECT 75.77 7.12 77.36 7.29 ;
      RECT 77.19 5.92 77.36 7.29 ;
      RECT 75.71 7.025 76 7.255 ;
      RECT 77.13 5.92 77.42 6.15 ;
      RECT 77.13 5.95 77.59 6.12 ;
      RECT 73.76 2.705 74.1 3.055 ;
      RECT 73.85 2.025 74.02 3.055 ;
      RECT 76.14 1.965 76.49 2.315 ;
      RECT 73.85 2.025 76.49 2.195 ;
      RECT 76.165 6.655 76.49 6.98 ;
      RECT 70.705 6.61 71.055 6.96 ;
      RECT 76.14 6.655 76.49 6.885 ;
      RECT 70.505 6.655 71.055 6.885 ;
      RECT 70.335 6.685 76.49 6.855 ;
      RECT 75.365 2.365 75.685 2.685 ;
      RECT 75.335 2.365 75.685 2.595 ;
      RECT 75.165 2.395 75.685 2.565 ;
      RECT 75.365 6.255 75.685 6.545 ;
      RECT 75.335 6.285 75.685 6.515 ;
      RECT 75.165 6.315 75.685 6.485 ;
      RECT 71.055 2.985 71.205 3.26 ;
      RECT 71.595 2.065 71.6 2.285 ;
      RECT 72.745 2.265 72.76 2.463 ;
      RECT 72.71 2.257 72.745 2.47 ;
      RECT 72.68 2.25 72.71 2.47 ;
      RECT 72.625 2.215 72.68 2.47 ;
      RECT 72.56 2.152 72.625 2.47 ;
      RECT 72.555 2.117 72.56 2.468 ;
      RECT 72.55 2.112 72.555 2.46 ;
      RECT 72.545 2.107 72.55 2.446 ;
      RECT 72.54 2.104 72.545 2.439 ;
      RECT 72.495 2.094 72.54 2.39 ;
      RECT 72.475 2.081 72.495 2.325 ;
      RECT 72.47 2.076 72.475 2.298 ;
      RECT 72.465 2.075 72.47 2.291 ;
      RECT 72.46 2.074 72.465 2.284 ;
      RECT 72.375 2.059 72.46 2.23 ;
      RECT 72.345 2.04 72.375 2.18 ;
      RECT 72.265 2.023 72.345 2.165 ;
      RECT 72.23 2.01 72.265 2.15 ;
      RECT 72.222 2.01 72.23 2.145 ;
      RECT 72.136 2.011 72.222 2.145 ;
      RECT 72.05 2.013 72.136 2.145 ;
      RECT 72.025 2.014 72.05 2.149 ;
      RECT 71.95 2.02 72.025 2.164 ;
      RECT 71.867 2.032 71.95 2.188 ;
      RECT 71.781 2.045 71.867 2.214 ;
      RECT 71.695 2.058 71.781 2.24 ;
      RECT 71.66 2.067 71.695 2.259 ;
      RECT 71.61 2.067 71.66 2.272 ;
      RECT 71.6 2.065 71.61 2.283 ;
      RECT 71.585 2.062 71.595 2.285 ;
      RECT 71.57 2.054 71.585 2.293 ;
      RECT 71.555 2.046 71.57 2.313 ;
      RECT 71.55 2.041 71.555 2.37 ;
      RECT 71.535 2.036 71.55 2.443 ;
      RECT 71.53 2.031 71.535 2.485 ;
      RECT 71.525 2.029 71.53 2.513 ;
      RECT 71.52 2.027 71.525 2.535 ;
      RECT 71.51 2.023 71.52 2.578 ;
      RECT 71.505 2.02 71.51 2.603 ;
      RECT 71.5 2.018 71.505 2.623 ;
      RECT 71.495 2.016 71.5 2.647 ;
      RECT 71.49 2.012 71.495 2.67 ;
      RECT 71.485 2.008 71.49 2.693 ;
      RECT 71.45 1.998 71.485 2.8 ;
      RECT 71.445 1.988 71.45 2.898 ;
      RECT 71.44 1.986 71.445 2.925 ;
      RECT 71.435 1.985 71.44 2.945 ;
      RECT 71.43 1.977 71.435 2.965 ;
      RECT 71.425 1.972 71.43 3 ;
      RECT 71.42 1.97 71.425 3.018 ;
      RECT 71.415 1.97 71.42 3.043 ;
      RECT 71.41 1.97 71.415 3.065 ;
      RECT 71.375 1.97 71.41 3.108 ;
      RECT 71.35 1.97 71.375 3.137 ;
      RECT 71.34 1.97 71.35 2.323 ;
      RECT 71.343 2.38 71.35 3.147 ;
      RECT 71.34 2.437 71.343 3.15 ;
      RECT 71.335 1.97 71.34 2.295 ;
      RECT 71.335 2.487 71.34 3.153 ;
      RECT 71.325 1.97 71.335 2.285 ;
      RECT 71.33 2.54 71.335 3.156 ;
      RECT 71.325 2.625 71.33 3.16 ;
      RECT 71.315 1.97 71.325 2.273 ;
      RECT 71.32 2.672 71.325 3.164 ;
      RECT 71.315 2.747 71.32 3.168 ;
      RECT 71.28 1.97 71.315 2.248 ;
      RECT 71.305 2.83 71.315 3.173 ;
      RECT 71.295 2.897 71.305 3.18 ;
      RECT 71.29 2.925 71.295 3.185 ;
      RECT 71.28 2.938 71.29 3.191 ;
      RECT 71.235 1.97 71.28 2.205 ;
      RECT 71.275 2.943 71.28 3.198 ;
      RECT 71.235 2.96 71.275 3.26 ;
      RECT 71.23 1.972 71.235 2.178 ;
      RECT 71.205 2.98 71.235 3.26 ;
      RECT 71.225 1.977 71.23 2.15 ;
      RECT 71.015 2.989 71.055 3.26 ;
      RECT 70.99 2.997 71.015 3.23 ;
      RECT 70.945 3.005 70.99 3.23 ;
      RECT 70.93 3.01 70.945 3.225 ;
      RECT 70.92 3.01 70.93 3.219 ;
      RECT 70.91 3.017 70.92 3.216 ;
      RECT 70.905 3.055 70.91 3.205 ;
      RECT 70.9 3.117 70.905 3.183 ;
      RECT 72.17 2.992 72.355 3.215 ;
      RECT 72.17 3.007 72.36 3.211 ;
      RECT 72.16 2.28 72.245 3.21 ;
      RECT 72.16 3.007 72.365 3.204 ;
      RECT 72.155 3.015 72.365 3.203 ;
      RECT 72.36 2.735 72.68 3.055 ;
      RECT 72.155 2.907 72.325 2.998 ;
      RECT 72.15 2.907 72.325 2.98 ;
      RECT 72.14 2.715 72.275 2.955 ;
      RECT 72.135 2.715 72.275 2.9 ;
      RECT 72.095 2.295 72.265 2.8 ;
      RECT 72.08 2.295 72.265 2.67 ;
      RECT 72.075 2.295 72.265 2.623 ;
      RECT 72.07 2.295 72.265 2.603 ;
      RECT 72.065 2.295 72.265 2.578 ;
      RECT 72.035 2.295 72.295 2.555 ;
      RECT 72.045 2.292 72.255 2.555 ;
      RECT 72.17 2.287 72.255 3.215 ;
      RECT 72.055 2.28 72.245 2.555 ;
      RECT 72.05 2.285 72.245 2.555 ;
      RECT 70.88 2.497 71.065 2.71 ;
      RECT 70.88 2.505 71.075 2.703 ;
      RECT 70.86 2.505 71.075 2.7 ;
      RECT 70.855 2.505 71.075 2.685 ;
      RECT 70.785 2.42 71.045 2.68 ;
      RECT 70.785 2.565 71.08 2.593 ;
      RECT 70.44 3.02 70.7 3.28 ;
      RECT 70.465 2.965 70.66 3.28 ;
      RECT 70.46 2.714 70.64 3.008 ;
      RECT 70.46 2.72 70.65 3.008 ;
      RECT 70.44 2.722 70.65 2.953 ;
      RECT 70.435 2.732 70.65 2.82 ;
      RECT 70.465 2.712 70.64 3.28 ;
      RECT 70.551 2.71 70.64 3.28 ;
      RECT 70.41 1.93 70.445 2.3 ;
      RECT 70.2 2.04 70.205 2.3 ;
      RECT 70.445 1.937 70.46 2.3 ;
      RECT 70.335 1.93 70.41 2.378 ;
      RECT 70.325 1.93 70.335 2.463 ;
      RECT 70.3 1.93 70.325 2.498 ;
      RECT 70.26 1.93 70.3 2.566 ;
      RECT 70.25 1.937 70.26 2.618 ;
      RECT 70.22 2.04 70.25 2.659 ;
      RECT 70.215 2.04 70.22 2.698 ;
      RECT 70.205 2.04 70.215 2.718 ;
      RECT 70.2 2.335 70.205 2.755 ;
      RECT 70.195 2.352 70.2 2.775 ;
      RECT 70.18 2.415 70.195 2.815 ;
      RECT 70.175 2.458 70.18 2.85 ;
      RECT 70.17 2.466 70.175 2.863 ;
      RECT 70.16 2.48 70.17 2.885 ;
      RECT 70.135 2.515 70.16 2.95 ;
      RECT 70.125 2.55 70.135 3.013 ;
      RECT 70.105 2.58 70.125 3.074 ;
      RECT 70.09 2.616 70.105 3.141 ;
      RECT 70.08 2.644 70.09 3.18 ;
      RECT 70.07 2.666 70.08 3.2 ;
      RECT 70.065 2.676 70.07 3.211 ;
      RECT 70.06 2.685 70.065 3.214 ;
      RECT 70.05 2.703 70.06 3.218 ;
      RECT 70.04 2.721 70.05 3.219 ;
      RECT 70.015 2.76 70.04 3.216 ;
      RECT 69.995 2.802 70.015 3.213 ;
      RECT 69.98 2.84 69.995 3.212 ;
      RECT 69.945 2.875 69.98 3.209 ;
      RECT 69.94 2.897 69.945 3.207 ;
      RECT 69.875 2.937 69.94 3.204 ;
      RECT 69.87 2.977 69.875 3.2 ;
      RECT 69.855 2.987 69.87 3.191 ;
      RECT 69.845 3.107 69.855 3.176 ;
      RECT 70.325 3.52 70.335 3.78 ;
      RECT 70.325 3.523 70.345 3.779 ;
      RECT 70.315 3.513 70.325 3.778 ;
      RECT 70.305 3.528 70.385 3.774 ;
      RECT 70.29 3.507 70.305 3.772 ;
      RECT 70.265 3.532 70.39 3.768 ;
      RECT 70.25 3.492 70.265 3.763 ;
      RECT 70.25 3.534 70.4 3.762 ;
      RECT 70.25 3.542 70.415 3.755 ;
      RECT 70.19 3.479 70.25 3.745 ;
      RECT 70.18 3.466 70.19 3.727 ;
      RECT 70.155 3.456 70.18 3.717 ;
      RECT 70.15 3.446 70.155 3.709 ;
      RECT 70.085 3.542 70.415 3.691 ;
      RECT 70 3.542 70.415 3.653 ;
      RECT 69.89 3.37 70.15 3.63 ;
      RECT 70.265 3.5 70.29 3.768 ;
      RECT 70.305 3.51 70.315 3.774 ;
      RECT 69.89 3.518 70.33 3.63 ;
      RECT 70.075 7.765 70.365 7.995 ;
      RECT 70.135 7.025 70.305 7.995 ;
      RECT 70.035 7.055 70.405 7.425 ;
      RECT 70.075 7.025 70.365 7.425 ;
      RECT 69.105 3.275 69.135 3.575 ;
      RECT 68.88 3.26 68.885 3.535 ;
      RECT 68.68 3.26 68.835 3.52 ;
      RECT 69.98 1.975 70.01 2.235 ;
      RECT 69.97 1.975 69.98 2.343 ;
      RECT 69.95 1.975 69.97 2.353 ;
      RECT 69.935 1.975 69.95 2.365 ;
      RECT 69.88 1.975 69.935 2.415 ;
      RECT 69.865 1.975 69.88 2.463 ;
      RECT 69.835 1.975 69.865 2.498 ;
      RECT 69.78 1.975 69.835 2.56 ;
      RECT 69.76 1.975 69.78 2.628 ;
      RECT 69.755 1.975 69.76 2.658 ;
      RECT 69.75 1.975 69.755 2.67 ;
      RECT 69.745 2.092 69.75 2.688 ;
      RECT 69.725 2.11 69.745 2.713 ;
      RECT 69.705 2.137 69.725 2.763 ;
      RECT 69.7 2.157 69.705 2.794 ;
      RECT 69.695 2.165 69.7 2.811 ;
      RECT 69.68 2.191 69.695 2.84 ;
      RECT 69.665 2.233 69.68 2.875 ;
      RECT 69.66 2.262 69.665 2.898 ;
      RECT 69.655 2.277 69.66 2.911 ;
      RECT 69.65 2.3 69.655 2.922 ;
      RECT 69.64 2.32 69.65 2.94 ;
      RECT 69.63 2.35 69.64 2.963 ;
      RECT 69.625 2.372 69.63 2.983 ;
      RECT 69.62 2.387 69.625 2.998 ;
      RECT 69.605 2.417 69.62 3.025 ;
      RECT 69.6 2.447 69.605 3.051 ;
      RECT 69.595 2.465 69.6 3.063 ;
      RECT 69.585 2.495 69.595 3.082 ;
      RECT 69.575 2.52 69.585 3.107 ;
      RECT 69.57 2.54 69.575 3.126 ;
      RECT 69.565 2.557 69.57 3.139 ;
      RECT 69.555 2.583 69.565 3.158 ;
      RECT 69.545 2.621 69.555 3.185 ;
      RECT 69.54 2.647 69.545 3.205 ;
      RECT 69.535 2.657 69.54 3.215 ;
      RECT 69.53 2.67 69.535 3.23 ;
      RECT 69.525 2.685 69.53 3.24 ;
      RECT 69.52 2.707 69.525 3.255 ;
      RECT 69.515 2.725 69.52 3.266 ;
      RECT 69.51 2.735 69.515 3.277 ;
      RECT 69.505 2.743 69.51 3.289 ;
      RECT 69.5 2.751 69.505 3.3 ;
      RECT 69.495 2.777 69.5 3.313 ;
      RECT 69.485 2.805 69.495 3.326 ;
      RECT 69.48 2.835 69.485 3.335 ;
      RECT 69.475 2.85 69.48 3.342 ;
      RECT 69.46 2.875 69.475 3.349 ;
      RECT 69.455 2.897 69.46 3.355 ;
      RECT 69.45 2.922 69.455 3.358 ;
      RECT 69.441 2.95 69.45 3.362 ;
      RECT 69.435 2.967 69.441 3.367 ;
      RECT 69.43 2.985 69.435 3.371 ;
      RECT 69.425 2.997 69.43 3.374 ;
      RECT 69.42 3.018 69.425 3.378 ;
      RECT 69.415 3.036 69.42 3.381 ;
      RECT 69.41 3.05 69.415 3.384 ;
      RECT 69.405 3.067 69.41 3.387 ;
      RECT 69.4 3.08 69.405 3.39 ;
      RECT 69.375 3.117 69.4 3.398 ;
      RECT 69.37 3.162 69.375 3.407 ;
      RECT 69.365 3.19 69.37 3.41 ;
      RECT 69.355 3.21 69.365 3.414 ;
      RECT 69.35 3.23 69.355 3.419 ;
      RECT 69.345 3.245 69.35 3.422 ;
      RECT 69.325 3.255 69.345 3.429 ;
      RECT 69.26 3.262 69.325 3.455 ;
      RECT 69.225 3.265 69.26 3.483 ;
      RECT 69.21 3.268 69.225 3.498 ;
      RECT 69.2 3.269 69.21 3.513 ;
      RECT 69.19 3.27 69.2 3.53 ;
      RECT 69.185 3.27 69.19 3.545 ;
      RECT 69.18 3.27 69.185 3.553 ;
      RECT 69.165 3.271 69.18 3.568 ;
      RECT 69.135 3.273 69.165 3.575 ;
      RECT 69.025 3.28 69.105 3.575 ;
      RECT 68.98 3.285 69.025 3.575 ;
      RECT 68.97 3.286 68.98 3.565 ;
      RECT 68.96 3.287 68.97 3.558 ;
      RECT 68.94 3.289 68.96 3.553 ;
      RECT 68.93 3.26 68.94 3.548 ;
      RECT 68.885 3.26 68.93 3.54 ;
      RECT 68.855 3.26 68.88 3.53 ;
      RECT 68.835 3.26 68.855 3.523 ;
      RECT 69.115 2.06 69.375 2.32 ;
      RECT 68.995 2.075 69.005 2.24 ;
      RECT 68.98 2.075 68.985 2.235 ;
      RECT 66.345 1.915 66.53 2.205 ;
      RECT 68.16 2.04 68.175 2.195 ;
      RECT 66.31 1.915 66.335 2.175 ;
      RECT 68.725 1.965 68.73 2.107 ;
      RECT 68.64 1.96 68.665 2.1 ;
      RECT 69.04 2.077 69.115 2.27 ;
      RECT 69.025 2.075 69.04 2.253 ;
      RECT 69.005 2.075 69.025 2.245 ;
      RECT 68.985 2.075 68.995 2.238 ;
      RECT 68.94 2.07 68.98 2.228 ;
      RECT 68.9 2.045 68.94 2.213 ;
      RECT 68.885 2.02 68.9 2.203 ;
      RECT 68.88 2.014 68.885 2.201 ;
      RECT 68.845 2.006 68.88 2.184 ;
      RECT 68.84 1.999 68.845 2.172 ;
      RECT 68.82 1.994 68.84 2.16 ;
      RECT 68.81 1.988 68.82 2.145 ;
      RECT 68.79 1.983 68.81 2.13 ;
      RECT 68.78 1.978 68.79 2.123 ;
      RECT 68.775 1.976 68.78 2.118 ;
      RECT 68.77 1.975 68.775 2.115 ;
      RECT 68.73 1.97 68.77 2.111 ;
      RECT 68.71 1.964 68.725 2.106 ;
      RECT 68.675 1.961 68.71 2.103 ;
      RECT 68.665 1.96 68.675 2.101 ;
      RECT 68.605 1.96 68.64 2.098 ;
      RECT 68.56 1.96 68.605 2.098 ;
      RECT 68.51 1.96 68.56 2.101 ;
      RECT 68.495 1.962 68.51 2.103 ;
      RECT 68.48 1.965 68.495 2.104 ;
      RECT 68.47 1.97 68.48 2.105 ;
      RECT 68.44 1.975 68.47 2.11 ;
      RECT 68.43 1.981 68.44 2.118 ;
      RECT 68.42 1.983 68.43 2.122 ;
      RECT 68.41 1.987 68.42 2.126 ;
      RECT 68.385 1.993 68.41 2.134 ;
      RECT 68.375 1.998 68.385 2.142 ;
      RECT 68.36 2.002 68.375 2.146 ;
      RECT 68.325 2.008 68.36 2.154 ;
      RECT 68.305 2.013 68.325 2.164 ;
      RECT 68.275 2.02 68.305 2.173 ;
      RECT 68.23 2.029 68.275 2.187 ;
      RECT 68.225 2.034 68.23 2.198 ;
      RECT 68.205 2.037 68.225 2.199 ;
      RECT 68.175 2.04 68.205 2.197 ;
      RECT 68.14 2.04 68.16 2.193 ;
      RECT 68.07 2.04 68.14 2.184 ;
      RECT 68.055 2.037 68.07 2.176 ;
      RECT 68.015 2.03 68.055 2.171 ;
      RECT 67.99 2.02 68.015 2.164 ;
      RECT 67.985 2.014 67.99 2.161 ;
      RECT 67.945 2.008 67.985 2.158 ;
      RECT 67.93 2.001 67.945 2.153 ;
      RECT 67.91 1.997 67.93 2.148 ;
      RECT 67.895 1.992 67.91 2.144 ;
      RECT 67.88 1.987 67.895 2.142 ;
      RECT 67.865 1.983 67.88 2.141 ;
      RECT 67.85 1.981 67.865 2.137 ;
      RECT 67.84 1.979 67.85 2.132 ;
      RECT 67.825 1.976 67.84 2.128 ;
      RECT 67.815 1.974 67.825 2.123 ;
      RECT 67.795 1.971 67.815 2.119 ;
      RECT 67.75 1.97 67.795 2.117 ;
      RECT 67.69 1.972 67.75 2.118 ;
      RECT 67.67 1.974 67.69 2.12 ;
      RECT 67.64 1.977 67.67 2.121 ;
      RECT 67.59 1.982 67.64 2.123 ;
      RECT 67.585 1.985 67.59 2.125 ;
      RECT 67.575 1.987 67.585 2.128 ;
      RECT 67.57 1.989 67.575 2.131 ;
      RECT 67.52 1.992 67.57 2.138 ;
      RECT 67.5 1.996 67.52 2.15 ;
      RECT 67.49 1.999 67.5 2.156 ;
      RECT 67.48 2 67.49 2.159 ;
      RECT 67.441 2.003 67.48 2.161 ;
      RECT 67.355 2.01 67.441 2.164 ;
      RECT 67.281 2.02 67.355 2.168 ;
      RECT 67.195 2.031 67.281 2.173 ;
      RECT 67.18 2.038 67.195 2.175 ;
      RECT 67.125 2.042 67.18 2.176 ;
      RECT 67.111 2.045 67.125 2.178 ;
      RECT 67.025 2.045 67.111 2.18 ;
      RECT 66.985 2.042 67.025 2.183 ;
      RECT 66.961 2.038 66.985 2.185 ;
      RECT 66.875 2.028 66.961 2.188 ;
      RECT 66.845 2.017 66.875 2.189 ;
      RECT 66.826 2.013 66.845 2.188 ;
      RECT 66.74 2.006 66.826 2.185 ;
      RECT 66.68 1.995 66.74 2.182 ;
      RECT 66.66 1.987 66.68 2.18 ;
      RECT 66.625 1.982 66.66 2.179 ;
      RECT 66.6 1.977 66.625 2.178 ;
      RECT 66.57 1.972 66.6 2.177 ;
      RECT 66.545 1.915 66.57 2.176 ;
      RECT 66.53 1.915 66.545 2.2 ;
      RECT 66.335 1.915 66.345 2.2 ;
      RECT 68.11 2.935 68.115 3.075 ;
      RECT 67.77 2.935 67.805 3.073 ;
      RECT 67.345 2.92 67.36 3.065 ;
      RECT 69.175 2.7 69.265 2.96 ;
      RECT 69.005 2.565 69.105 2.96 ;
      RECT 66.04 2.54 66.12 2.75 ;
      RECT 69.13 2.677 69.175 2.96 ;
      RECT 69.12 2.647 69.13 2.96 ;
      RECT 69.105 2.57 69.12 2.96 ;
      RECT 68.92 2.565 69.005 2.925 ;
      RECT 68.915 2.567 68.92 2.92 ;
      RECT 68.91 2.572 68.915 2.92 ;
      RECT 68.875 2.672 68.91 2.92 ;
      RECT 68.865 2.7 68.875 2.92 ;
      RECT 68.855 2.715 68.865 2.92 ;
      RECT 68.845 2.727 68.855 2.92 ;
      RECT 68.84 2.737 68.845 2.92 ;
      RECT 68.825 2.747 68.84 2.922 ;
      RECT 68.82 2.762 68.825 2.924 ;
      RECT 68.805 2.775 68.82 2.926 ;
      RECT 68.8 2.79 68.805 2.929 ;
      RECT 68.78 2.8 68.8 2.933 ;
      RECT 68.765 2.81 68.78 2.936 ;
      RECT 68.73 2.817 68.765 2.941 ;
      RECT 68.686 2.824 68.73 2.949 ;
      RECT 68.6 2.836 68.686 2.962 ;
      RECT 68.575 2.847 68.6 2.973 ;
      RECT 68.545 2.852 68.575 2.978 ;
      RECT 68.51 2.857 68.545 2.986 ;
      RECT 68.48 2.862 68.51 2.993 ;
      RECT 68.455 2.867 68.48 2.998 ;
      RECT 68.39 2.874 68.455 3.007 ;
      RECT 68.32 2.887 68.39 3.023 ;
      RECT 68.29 2.897 68.32 3.035 ;
      RECT 68.265 2.902 68.29 3.042 ;
      RECT 68.21 2.909 68.265 3.05 ;
      RECT 68.205 2.916 68.21 3.055 ;
      RECT 68.2 2.918 68.205 3.056 ;
      RECT 68.185 2.92 68.2 3.058 ;
      RECT 68.18 2.92 68.185 3.061 ;
      RECT 68.115 2.927 68.18 3.068 ;
      RECT 68.08 2.937 68.11 3.078 ;
      RECT 68.063 2.94 68.08 3.08 ;
      RECT 67.977 2.939 68.063 3.079 ;
      RECT 67.891 2.937 67.977 3.076 ;
      RECT 67.805 2.936 67.891 3.074 ;
      RECT 67.704 2.934 67.77 3.073 ;
      RECT 67.618 2.931 67.704 3.071 ;
      RECT 67.532 2.927 67.618 3.069 ;
      RECT 67.446 2.924 67.532 3.068 ;
      RECT 67.36 2.921 67.446 3.066 ;
      RECT 67.26 2.92 67.345 3.063 ;
      RECT 67.21 2.918 67.26 3.061 ;
      RECT 67.19 2.915 67.21 3.059 ;
      RECT 67.17 2.913 67.19 3.056 ;
      RECT 67.145 2.909 67.17 3.053 ;
      RECT 67.1 2.903 67.145 3.048 ;
      RECT 67.06 2.897 67.1 3.04 ;
      RECT 67.035 2.892 67.06 3.033 ;
      RECT 66.98 2.885 67.035 3.025 ;
      RECT 66.956 2.878 66.98 3.018 ;
      RECT 66.87 2.869 66.956 3.008 ;
      RECT 66.84 2.861 66.87 2.998 ;
      RECT 66.81 2.857 66.84 2.993 ;
      RECT 66.805 2.854 66.81 2.99 ;
      RECT 66.8 2.853 66.805 2.99 ;
      RECT 66.725 2.846 66.8 2.983 ;
      RECT 66.686 2.837 66.725 2.972 ;
      RECT 66.6 2.827 66.686 2.96 ;
      RECT 66.56 2.817 66.6 2.948 ;
      RECT 66.521 2.812 66.56 2.941 ;
      RECT 66.435 2.802 66.521 2.93 ;
      RECT 66.395 2.79 66.435 2.919 ;
      RECT 66.36 2.775 66.395 2.912 ;
      RECT 66.35 2.765 66.36 2.909 ;
      RECT 66.33 2.75 66.35 2.907 ;
      RECT 66.3 2.72 66.33 2.903 ;
      RECT 66.29 2.7 66.3 2.898 ;
      RECT 66.285 2.692 66.29 2.895 ;
      RECT 66.28 2.685 66.285 2.893 ;
      RECT 66.265 2.672 66.28 2.886 ;
      RECT 66.26 2.662 66.265 2.878 ;
      RECT 66.255 2.655 66.26 2.873 ;
      RECT 66.25 2.65 66.255 2.869 ;
      RECT 66.235 2.637 66.25 2.861 ;
      RECT 66.23 2.547 66.235 2.85 ;
      RECT 66.225 2.542 66.23 2.843 ;
      RECT 66.15 2.54 66.225 2.803 ;
      RECT 66.12 2.54 66.15 2.758 ;
      RECT 66.025 2.545 66.04 2.745 ;
      RECT 68.51 2.25 68.77 2.51 ;
      RECT 68.495 2.238 68.675 2.475 ;
      RECT 68.49 2.239 68.675 2.473 ;
      RECT 68.475 2.243 68.685 2.463 ;
      RECT 68.47 2.248 68.69 2.433 ;
      RECT 68.475 2.245 68.69 2.463 ;
      RECT 68.49 2.24 68.685 2.473 ;
      RECT 68.51 2.237 68.675 2.51 ;
      RECT 68.51 2.236 68.665 2.51 ;
      RECT 68.535 2.235 68.665 2.51 ;
      RECT 68.095 2.48 68.355 2.74 ;
      RECT 67.97 2.525 68.355 2.735 ;
      RECT 67.96 2.53 68.355 2.73 ;
      RECT 67.975 3.47 67.99 3.78 ;
      RECT 66.57 3.24 66.58 3.37 ;
      RECT 66.35 3.235 66.455 3.37 ;
      RECT 66.265 3.24 66.315 3.37 ;
      RECT 64.815 1.975 64.82 3.08 ;
      RECT 68.07 3.562 68.075 3.698 ;
      RECT 68.065 3.557 68.07 3.758 ;
      RECT 68.06 3.555 68.065 3.771 ;
      RECT 68.045 3.552 68.06 3.773 ;
      RECT 68.04 3.547 68.045 3.775 ;
      RECT 68.035 3.543 68.04 3.778 ;
      RECT 68.02 3.538 68.035 3.78 ;
      RECT 67.99 3.53 68.02 3.78 ;
      RECT 67.951 3.47 67.975 3.78 ;
      RECT 67.865 3.47 67.951 3.777 ;
      RECT 67.835 3.47 67.865 3.77 ;
      RECT 67.81 3.47 67.835 3.763 ;
      RECT 67.785 3.47 67.81 3.755 ;
      RECT 67.77 3.47 67.785 3.748 ;
      RECT 67.745 3.47 67.77 3.74 ;
      RECT 67.73 3.47 67.745 3.733 ;
      RECT 67.69 3.48 67.73 3.722 ;
      RECT 67.68 3.475 67.69 3.712 ;
      RECT 67.676 3.474 67.68 3.709 ;
      RECT 67.59 3.466 67.676 3.692 ;
      RECT 67.557 3.455 67.59 3.669 ;
      RECT 67.471 3.444 67.557 3.647 ;
      RECT 67.385 3.428 67.471 3.616 ;
      RECT 67.315 3.413 67.385 3.588 ;
      RECT 67.305 3.406 67.315 3.575 ;
      RECT 67.275 3.403 67.305 3.565 ;
      RECT 67.25 3.399 67.275 3.558 ;
      RECT 67.235 3.396 67.25 3.553 ;
      RECT 67.23 3.395 67.235 3.548 ;
      RECT 67.2 3.39 67.23 3.541 ;
      RECT 67.195 3.385 67.2 3.536 ;
      RECT 67.18 3.382 67.195 3.531 ;
      RECT 67.175 3.377 67.18 3.526 ;
      RECT 67.155 3.372 67.175 3.523 ;
      RECT 67.14 3.367 67.155 3.515 ;
      RECT 67.125 3.361 67.14 3.51 ;
      RECT 67.095 3.352 67.125 3.503 ;
      RECT 67.09 3.345 67.095 3.495 ;
      RECT 67.085 3.343 67.09 3.493 ;
      RECT 67.08 3.342 67.085 3.49 ;
      RECT 67.04 3.335 67.08 3.483 ;
      RECT 67.026 3.325 67.04 3.473 ;
      RECT 66.975 3.314 67.026 3.461 ;
      RECT 66.95 3.3 66.975 3.447 ;
      RECT 66.925 3.289 66.95 3.439 ;
      RECT 66.905 3.278 66.925 3.433 ;
      RECT 66.895 3.272 66.905 3.428 ;
      RECT 66.89 3.27 66.895 3.424 ;
      RECT 66.87 3.265 66.89 3.419 ;
      RECT 66.84 3.255 66.87 3.409 ;
      RECT 66.835 3.247 66.84 3.402 ;
      RECT 66.82 3.245 66.835 3.398 ;
      RECT 66.8 3.245 66.82 3.393 ;
      RECT 66.795 3.244 66.8 3.391 ;
      RECT 66.79 3.244 66.795 3.388 ;
      RECT 66.75 3.243 66.79 3.383 ;
      RECT 66.725 3.242 66.75 3.378 ;
      RECT 66.665 3.241 66.725 3.375 ;
      RECT 66.58 3.24 66.665 3.373 ;
      RECT 66.541 3.239 66.57 3.37 ;
      RECT 66.455 3.237 66.541 3.37 ;
      RECT 66.315 3.237 66.35 3.37 ;
      RECT 66.225 3.241 66.265 3.373 ;
      RECT 66.21 3.244 66.225 3.38 ;
      RECT 66.2 3.245 66.21 3.387 ;
      RECT 66.175 3.248 66.2 3.392 ;
      RECT 66.17 3.25 66.175 3.395 ;
      RECT 66.12 3.252 66.17 3.396 ;
      RECT 66.081 3.256 66.12 3.398 ;
      RECT 65.995 3.258 66.081 3.401 ;
      RECT 65.977 3.26 65.995 3.403 ;
      RECT 65.891 3.263 65.977 3.405 ;
      RECT 65.805 3.267 65.891 3.408 ;
      RECT 65.768 3.271 65.805 3.411 ;
      RECT 65.682 3.274 65.768 3.414 ;
      RECT 65.596 3.278 65.682 3.417 ;
      RECT 65.51 3.283 65.596 3.421 ;
      RECT 65.49 3.285 65.51 3.424 ;
      RECT 65.47 3.284 65.49 3.425 ;
      RECT 65.421 3.281 65.47 3.426 ;
      RECT 65.335 3.276 65.421 3.429 ;
      RECT 65.285 3.271 65.335 3.431 ;
      RECT 65.261 3.269 65.285 3.432 ;
      RECT 65.175 3.264 65.261 3.434 ;
      RECT 65.15 3.26 65.175 3.433 ;
      RECT 65.14 3.257 65.15 3.431 ;
      RECT 65.13 3.25 65.14 3.428 ;
      RECT 65.125 3.23 65.13 3.423 ;
      RECT 65.115 3.2 65.125 3.418 ;
      RECT 65.1 3.07 65.115 3.409 ;
      RECT 65.095 3.062 65.1 3.402 ;
      RECT 65.075 3.055 65.095 3.394 ;
      RECT 65.07 3.037 65.075 3.386 ;
      RECT 65.06 3.017 65.07 3.381 ;
      RECT 65.055 2.99 65.06 3.377 ;
      RECT 65.05 2.967 65.055 3.374 ;
      RECT 65.03 2.925 65.05 3.366 ;
      RECT 64.995 2.84 65.03 3.35 ;
      RECT 64.99 2.772 64.995 3.338 ;
      RECT 64.975 2.742 64.99 3.332 ;
      RECT 64.97 1.987 64.975 2.233 ;
      RECT 64.96 2.712 64.975 3.323 ;
      RECT 64.965 1.982 64.97 2.265 ;
      RECT 64.96 1.977 64.965 2.308 ;
      RECT 64.955 1.975 64.96 2.343 ;
      RECT 64.94 2.675 64.96 3.313 ;
      RECT 64.95 1.975 64.955 2.38 ;
      RECT 64.935 1.975 64.95 2.478 ;
      RECT 64.935 2.648 64.94 3.306 ;
      RECT 64.93 1.975 64.935 2.553 ;
      RECT 64.93 2.636 64.935 3.303 ;
      RECT 64.925 1.975 64.93 2.585 ;
      RECT 64.925 2.615 64.93 3.3 ;
      RECT 64.92 1.975 64.925 3.297 ;
      RECT 64.885 1.975 64.92 3.283 ;
      RECT 64.87 1.975 64.885 3.265 ;
      RECT 64.85 1.975 64.87 3.255 ;
      RECT 64.825 1.975 64.85 3.238 ;
      RECT 64.82 1.975 64.825 3.188 ;
      RECT 64.81 1.975 64.815 3.018 ;
      RECT 64.805 1.975 64.81 2.925 ;
      RECT 64.8 1.975 64.805 2.838 ;
      RECT 64.795 1.975 64.8 2.77 ;
      RECT 64.79 1.975 64.795 2.713 ;
      RECT 64.78 1.975 64.79 2.608 ;
      RECT 64.775 1.975 64.78 2.48 ;
      RECT 64.77 1.975 64.775 2.398 ;
      RECT 64.765 1.977 64.77 2.315 ;
      RECT 64.76 1.982 64.765 2.248 ;
      RECT 64.755 1.987 64.76 2.175 ;
      RECT 67.57 2.305 67.83 2.565 ;
      RECT 67.59 2.272 67.8 2.565 ;
      RECT 67.59 2.27 67.79 2.565 ;
      RECT 67.6 2.257 67.79 2.565 ;
      RECT 67.6 2.255 67.715 2.565 ;
      RECT 67.075 2.38 67.25 2.66 ;
      RECT 67.07 2.38 67.25 2.658 ;
      RECT 67.07 2.38 67.265 2.655 ;
      RECT 67.06 2.38 67.265 2.653 ;
      RECT 67.005 2.38 67.265 2.64 ;
      RECT 67.005 2.455 67.27 2.618 ;
      RECT 66.55 2.392 66.57 2.635 ;
      RECT 66.55 2.392 66.61 2.634 ;
      RECT 66.545 2.394 66.61 2.633 ;
      RECT 66.545 2.394 66.696 2.632 ;
      RECT 66.545 2.394 66.765 2.631 ;
      RECT 66.545 2.394 66.785 2.623 ;
      RECT 66.525 2.397 66.785 2.621 ;
      RECT 66.51 2.407 66.785 2.606 ;
      RECT 66.51 2.407 66.8 2.605 ;
      RECT 66.505 2.416 66.8 2.597 ;
      RECT 66.505 2.416 66.805 2.593 ;
      RECT 66.61 2.33 66.87 2.59 ;
      RECT 66.5 2.418 66.87 2.475 ;
      RECT 66.57 2.385 66.87 2.59 ;
      RECT 66.535 3.578 66.54 3.785 ;
      RECT 66.485 3.572 66.535 3.784 ;
      RECT 66.452 3.586 66.545 3.783 ;
      RECT 66.366 3.586 66.545 3.782 ;
      RECT 66.28 3.586 66.545 3.781 ;
      RECT 66.28 3.685 66.55 3.778 ;
      RECT 66.275 3.685 66.55 3.773 ;
      RECT 66.27 3.685 66.55 3.755 ;
      RECT 66.265 3.685 66.55 3.738 ;
      RECT 66.225 3.47 66.485 3.73 ;
      RECT 65.685 2.62 65.771 3.034 ;
      RECT 65.685 2.62 65.81 3.031 ;
      RECT 65.685 2.62 65.83 3.021 ;
      RECT 65.64 2.62 65.83 3.018 ;
      RECT 65.64 2.772 65.84 3.008 ;
      RECT 65.64 2.793 65.845 3.002 ;
      RECT 65.64 2.811 65.85 2.998 ;
      RECT 65.64 2.831 65.86 2.993 ;
      RECT 65.615 2.831 65.86 2.99 ;
      RECT 65.605 2.831 65.86 2.968 ;
      RECT 65.605 2.847 65.865 2.938 ;
      RECT 65.57 2.62 65.83 2.925 ;
      RECT 65.57 2.859 65.87 2.88 ;
      RECT 63.23 7.77 63.52 8 ;
      RECT 63.29 6.29 63.46 8 ;
      RECT 63.24 6.655 63.59 7.005 ;
      RECT 63.23 6.29 63.52 6.52 ;
      RECT 62.825 2.395 62.93 2.965 ;
      RECT 62.825 2.73 63.15 2.96 ;
      RECT 62.825 2.76 63.32 2.93 ;
      RECT 62.825 2.395 63.015 2.96 ;
      RECT 62.24 2.36 62.53 2.59 ;
      RECT 62.24 2.395 63.015 2.565 ;
      RECT 62.3 0.88 62.47 2.59 ;
      RECT 62.24 0.88 62.53 1.11 ;
      RECT 62.24 7.77 62.53 8 ;
      RECT 62.3 6.29 62.47 8 ;
      RECT 62.24 6.29 62.53 6.52 ;
      RECT 62.24 6.325 63.095 6.485 ;
      RECT 62.925 5.92 63.095 6.485 ;
      RECT 62.24 6.32 62.635 6.485 ;
      RECT 62.86 5.92 63.15 6.15 ;
      RECT 62.86 5.95 63.32 6.12 ;
      RECT 61.87 2.73 62.16 2.96 ;
      RECT 61.87 2.76 62.33 2.93 ;
      RECT 61.935 1.655 62.1 2.96 ;
      RECT 60.45 1.625 60.74 1.855 ;
      RECT 60.45 1.655 62.1 1.825 ;
      RECT 60.51 0.885 60.68 1.855 ;
      RECT 60.45 0.885 60.74 1.115 ;
      RECT 60.45 7.765 60.74 7.995 ;
      RECT 60.51 7.025 60.68 7.995 ;
      RECT 60.51 7.12 62.1 7.29 ;
      RECT 61.93 5.92 62.1 7.29 ;
      RECT 60.45 7.025 60.74 7.255 ;
      RECT 61.87 5.92 62.16 6.15 ;
      RECT 61.87 5.95 62.33 6.12 ;
      RECT 58.5 2.705 58.84 3.055 ;
      RECT 58.59 2.025 58.76 3.055 ;
      RECT 60.88 1.965 61.23 2.315 ;
      RECT 58.59 2.025 61.23 2.195 ;
      RECT 60.905 6.655 61.23 6.98 ;
      RECT 55.445 6.61 55.795 6.96 ;
      RECT 60.88 6.655 61.23 6.885 ;
      RECT 55.245 6.655 55.795 6.885 ;
      RECT 55.075 6.685 61.23 6.855 ;
      RECT 60.105 2.365 60.425 2.685 ;
      RECT 60.075 2.365 60.425 2.595 ;
      RECT 59.905 2.395 60.425 2.565 ;
      RECT 60.105 6.255 60.425 6.545 ;
      RECT 60.075 6.285 60.425 6.515 ;
      RECT 59.905 6.315 60.425 6.485 ;
      RECT 55.795 2.985 55.945 3.26 ;
      RECT 56.335 2.065 56.34 2.285 ;
      RECT 57.485 2.265 57.5 2.463 ;
      RECT 57.45 2.257 57.485 2.47 ;
      RECT 57.42 2.25 57.45 2.47 ;
      RECT 57.365 2.215 57.42 2.47 ;
      RECT 57.3 2.152 57.365 2.47 ;
      RECT 57.295 2.117 57.3 2.468 ;
      RECT 57.29 2.112 57.295 2.46 ;
      RECT 57.285 2.107 57.29 2.446 ;
      RECT 57.28 2.104 57.285 2.439 ;
      RECT 57.235 2.094 57.28 2.39 ;
      RECT 57.215 2.081 57.235 2.325 ;
      RECT 57.21 2.076 57.215 2.298 ;
      RECT 57.205 2.075 57.21 2.291 ;
      RECT 57.2 2.074 57.205 2.284 ;
      RECT 57.115 2.059 57.2 2.23 ;
      RECT 57.085 2.04 57.115 2.18 ;
      RECT 57.005 2.023 57.085 2.165 ;
      RECT 56.97 2.01 57.005 2.15 ;
      RECT 56.962 2.01 56.97 2.145 ;
      RECT 56.876 2.011 56.962 2.145 ;
      RECT 56.79 2.013 56.876 2.145 ;
      RECT 56.765 2.014 56.79 2.149 ;
      RECT 56.69 2.02 56.765 2.164 ;
      RECT 56.607 2.032 56.69 2.188 ;
      RECT 56.521 2.045 56.607 2.214 ;
      RECT 56.435 2.058 56.521 2.24 ;
      RECT 56.4 2.067 56.435 2.259 ;
      RECT 56.35 2.067 56.4 2.272 ;
      RECT 56.34 2.065 56.35 2.283 ;
      RECT 56.325 2.062 56.335 2.285 ;
      RECT 56.31 2.054 56.325 2.293 ;
      RECT 56.295 2.046 56.31 2.313 ;
      RECT 56.29 2.041 56.295 2.37 ;
      RECT 56.275 2.036 56.29 2.443 ;
      RECT 56.27 2.031 56.275 2.485 ;
      RECT 56.265 2.029 56.27 2.513 ;
      RECT 56.26 2.027 56.265 2.535 ;
      RECT 56.25 2.023 56.26 2.578 ;
      RECT 56.245 2.02 56.25 2.603 ;
      RECT 56.24 2.018 56.245 2.623 ;
      RECT 56.235 2.016 56.24 2.647 ;
      RECT 56.23 2.012 56.235 2.67 ;
      RECT 56.225 2.008 56.23 2.693 ;
      RECT 56.19 1.998 56.225 2.8 ;
      RECT 56.185 1.988 56.19 2.898 ;
      RECT 56.18 1.986 56.185 2.925 ;
      RECT 56.175 1.985 56.18 2.945 ;
      RECT 56.17 1.977 56.175 2.965 ;
      RECT 56.165 1.972 56.17 3 ;
      RECT 56.16 1.97 56.165 3.018 ;
      RECT 56.155 1.97 56.16 3.043 ;
      RECT 56.15 1.97 56.155 3.065 ;
      RECT 56.115 1.97 56.15 3.108 ;
      RECT 56.09 1.97 56.115 3.137 ;
      RECT 56.08 1.97 56.09 2.323 ;
      RECT 56.083 2.38 56.09 3.147 ;
      RECT 56.08 2.437 56.083 3.15 ;
      RECT 56.075 1.97 56.08 2.295 ;
      RECT 56.075 2.487 56.08 3.153 ;
      RECT 56.065 1.97 56.075 2.285 ;
      RECT 56.07 2.54 56.075 3.156 ;
      RECT 56.065 2.625 56.07 3.16 ;
      RECT 56.055 1.97 56.065 2.273 ;
      RECT 56.06 2.672 56.065 3.164 ;
      RECT 56.055 2.747 56.06 3.168 ;
      RECT 56.02 1.97 56.055 2.248 ;
      RECT 56.045 2.83 56.055 3.173 ;
      RECT 56.035 2.897 56.045 3.18 ;
      RECT 56.03 2.925 56.035 3.185 ;
      RECT 56.02 2.938 56.03 3.191 ;
      RECT 55.975 1.97 56.02 2.205 ;
      RECT 56.015 2.943 56.02 3.198 ;
      RECT 55.975 2.96 56.015 3.26 ;
      RECT 55.97 1.972 55.975 2.178 ;
      RECT 55.945 2.98 55.975 3.26 ;
      RECT 55.965 1.977 55.97 2.15 ;
      RECT 55.755 2.989 55.795 3.26 ;
      RECT 55.73 2.997 55.755 3.23 ;
      RECT 55.685 3.005 55.73 3.23 ;
      RECT 55.67 3.01 55.685 3.225 ;
      RECT 55.66 3.01 55.67 3.219 ;
      RECT 55.65 3.017 55.66 3.216 ;
      RECT 55.645 3.055 55.65 3.205 ;
      RECT 55.64 3.117 55.645 3.183 ;
      RECT 56.91 2.992 57.095 3.215 ;
      RECT 56.91 3.007 57.1 3.211 ;
      RECT 56.9 2.28 56.985 3.21 ;
      RECT 56.9 3.007 57.105 3.204 ;
      RECT 56.895 3.015 57.105 3.203 ;
      RECT 57.1 2.735 57.42 3.055 ;
      RECT 56.895 2.907 57.065 2.998 ;
      RECT 56.89 2.907 57.065 2.98 ;
      RECT 56.88 2.715 57.015 2.955 ;
      RECT 56.875 2.715 57.015 2.9 ;
      RECT 56.835 2.295 57.005 2.8 ;
      RECT 56.82 2.295 57.005 2.67 ;
      RECT 56.815 2.295 57.005 2.623 ;
      RECT 56.81 2.295 57.005 2.603 ;
      RECT 56.805 2.295 57.005 2.578 ;
      RECT 56.775 2.295 57.035 2.555 ;
      RECT 56.785 2.292 56.995 2.555 ;
      RECT 56.91 2.287 56.995 3.215 ;
      RECT 56.795 2.28 56.985 2.555 ;
      RECT 56.79 2.285 56.985 2.555 ;
      RECT 55.62 2.497 55.805 2.71 ;
      RECT 55.62 2.505 55.815 2.703 ;
      RECT 55.6 2.505 55.815 2.7 ;
      RECT 55.595 2.505 55.815 2.685 ;
      RECT 55.525 2.42 55.785 2.68 ;
      RECT 55.525 2.565 55.82 2.593 ;
      RECT 55.18 3.02 55.44 3.28 ;
      RECT 55.205 2.965 55.4 3.28 ;
      RECT 55.2 2.714 55.38 3.008 ;
      RECT 55.2 2.72 55.39 3.008 ;
      RECT 55.18 2.722 55.39 2.953 ;
      RECT 55.175 2.732 55.39 2.82 ;
      RECT 55.205 2.712 55.38 3.28 ;
      RECT 55.291 2.71 55.38 3.28 ;
      RECT 55.15 1.93 55.185 2.3 ;
      RECT 54.94 2.04 54.945 2.3 ;
      RECT 55.185 1.937 55.2 2.3 ;
      RECT 55.075 1.93 55.15 2.378 ;
      RECT 55.065 1.93 55.075 2.463 ;
      RECT 55.04 1.93 55.065 2.498 ;
      RECT 55 1.93 55.04 2.566 ;
      RECT 54.99 1.937 55 2.618 ;
      RECT 54.96 2.04 54.99 2.659 ;
      RECT 54.955 2.04 54.96 2.698 ;
      RECT 54.945 2.04 54.955 2.718 ;
      RECT 54.94 2.335 54.945 2.755 ;
      RECT 54.935 2.352 54.94 2.775 ;
      RECT 54.92 2.415 54.935 2.815 ;
      RECT 54.915 2.458 54.92 2.85 ;
      RECT 54.91 2.466 54.915 2.863 ;
      RECT 54.9 2.48 54.91 2.885 ;
      RECT 54.875 2.515 54.9 2.95 ;
      RECT 54.865 2.55 54.875 3.013 ;
      RECT 54.845 2.58 54.865 3.074 ;
      RECT 54.83 2.616 54.845 3.141 ;
      RECT 54.82 2.644 54.83 3.18 ;
      RECT 54.81 2.666 54.82 3.2 ;
      RECT 54.805 2.676 54.81 3.211 ;
      RECT 54.8 2.685 54.805 3.214 ;
      RECT 54.79 2.703 54.8 3.218 ;
      RECT 54.78 2.721 54.79 3.219 ;
      RECT 54.755 2.76 54.78 3.216 ;
      RECT 54.735 2.802 54.755 3.213 ;
      RECT 54.72 2.84 54.735 3.212 ;
      RECT 54.685 2.875 54.72 3.209 ;
      RECT 54.68 2.897 54.685 3.207 ;
      RECT 54.615 2.937 54.68 3.204 ;
      RECT 54.61 2.977 54.615 3.2 ;
      RECT 54.595 2.987 54.61 3.191 ;
      RECT 54.585 3.107 54.595 3.176 ;
      RECT 55.065 3.52 55.075 3.78 ;
      RECT 55.065 3.523 55.085 3.779 ;
      RECT 55.055 3.513 55.065 3.778 ;
      RECT 55.045 3.528 55.125 3.774 ;
      RECT 55.03 3.507 55.045 3.772 ;
      RECT 55.005 3.532 55.13 3.768 ;
      RECT 54.99 3.492 55.005 3.763 ;
      RECT 54.99 3.534 55.14 3.762 ;
      RECT 54.99 3.542 55.155 3.755 ;
      RECT 54.93 3.479 54.99 3.745 ;
      RECT 54.92 3.466 54.93 3.727 ;
      RECT 54.895 3.456 54.92 3.717 ;
      RECT 54.89 3.446 54.895 3.709 ;
      RECT 54.825 3.542 55.155 3.691 ;
      RECT 54.74 3.542 55.155 3.653 ;
      RECT 54.63 3.37 54.89 3.63 ;
      RECT 55.005 3.5 55.03 3.768 ;
      RECT 55.045 3.51 55.055 3.774 ;
      RECT 54.63 3.518 55.07 3.63 ;
      RECT 54.815 7.765 55.105 7.995 ;
      RECT 54.875 7.025 55.045 7.995 ;
      RECT 54.775 7.055 55.145 7.425 ;
      RECT 54.815 7.025 55.105 7.425 ;
      RECT 53.845 3.275 53.875 3.575 ;
      RECT 53.62 3.26 53.625 3.535 ;
      RECT 53.42 3.26 53.575 3.52 ;
      RECT 54.72 1.975 54.75 2.235 ;
      RECT 54.71 1.975 54.72 2.343 ;
      RECT 54.69 1.975 54.71 2.353 ;
      RECT 54.675 1.975 54.69 2.365 ;
      RECT 54.62 1.975 54.675 2.415 ;
      RECT 54.605 1.975 54.62 2.463 ;
      RECT 54.575 1.975 54.605 2.498 ;
      RECT 54.52 1.975 54.575 2.56 ;
      RECT 54.5 1.975 54.52 2.628 ;
      RECT 54.495 1.975 54.5 2.658 ;
      RECT 54.49 1.975 54.495 2.67 ;
      RECT 54.485 2.092 54.49 2.688 ;
      RECT 54.465 2.11 54.485 2.713 ;
      RECT 54.445 2.137 54.465 2.763 ;
      RECT 54.44 2.157 54.445 2.794 ;
      RECT 54.435 2.165 54.44 2.811 ;
      RECT 54.42 2.191 54.435 2.84 ;
      RECT 54.405 2.233 54.42 2.875 ;
      RECT 54.4 2.262 54.405 2.898 ;
      RECT 54.395 2.277 54.4 2.911 ;
      RECT 54.39 2.3 54.395 2.922 ;
      RECT 54.38 2.32 54.39 2.94 ;
      RECT 54.37 2.35 54.38 2.963 ;
      RECT 54.365 2.372 54.37 2.983 ;
      RECT 54.36 2.387 54.365 2.998 ;
      RECT 54.345 2.417 54.36 3.025 ;
      RECT 54.34 2.447 54.345 3.051 ;
      RECT 54.335 2.465 54.34 3.063 ;
      RECT 54.325 2.495 54.335 3.082 ;
      RECT 54.315 2.52 54.325 3.107 ;
      RECT 54.31 2.54 54.315 3.126 ;
      RECT 54.305 2.557 54.31 3.139 ;
      RECT 54.295 2.583 54.305 3.158 ;
      RECT 54.285 2.621 54.295 3.185 ;
      RECT 54.28 2.647 54.285 3.205 ;
      RECT 54.275 2.657 54.28 3.215 ;
      RECT 54.27 2.67 54.275 3.23 ;
      RECT 54.265 2.685 54.27 3.24 ;
      RECT 54.26 2.707 54.265 3.255 ;
      RECT 54.255 2.725 54.26 3.266 ;
      RECT 54.25 2.735 54.255 3.277 ;
      RECT 54.245 2.743 54.25 3.289 ;
      RECT 54.24 2.751 54.245 3.3 ;
      RECT 54.235 2.777 54.24 3.313 ;
      RECT 54.225 2.805 54.235 3.326 ;
      RECT 54.22 2.835 54.225 3.335 ;
      RECT 54.215 2.85 54.22 3.342 ;
      RECT 54.2 2.875 54.215 3.349 ;
      RECT 54.195 2.897 54.2 3.355 ;
      RECT 54.19 2.922 54.195 3.358 ;
      RECT 54.181 2.95 54.19 3.362 ;
      RECT 54.175 2.967 54.181 3.367 ;
      RECT 54.17 2.985 54.175 3.371 ;
      RECT 54.165 2.997 54.17 3.374 ;
      RECT 54.16 3.018 54.165 3.378 ;
      RECT 54.155 3.036 54.16 3.381 ;
      RECT 54.15 3.05 54.155 3.384 ;
      RECT 54.145 3.067 54.15 3.387 ;
      RECT 54.14 3.08 54.145 3.39 ;
      RECT 54.115 3.117 54.14 3.398 ;
      RECT 54.11 3.162 54.115 3.407 ;
      RECT 54.105 3.19 54.11 3.41 ;
      RECT 54.095 3.21 54.105 3.414 ;
      RECT 54.09 3.23 54.095 3.419 ;
      RECT 54.085 3.245 54.09 3.422 ;
      RECT 54.065 3.255 54.085 3.429 ;
      RECT 54 3.262 54.065 3.455 ;
      RECT 53.965 3.265 54 3.483 ;
      RECT 53.95 3.268 53.965 3.498 ;
      RECT 53.94 3.269 53.95 3.513 ;
      RECT 53.93 3.27 53.94 3.53 ;
      RECT 53.925 3.27 53.93 3.545 ;
      RECT 53.92 3.27 53.925 3.553 ;
      RECT 53.905 3.271 53.92 3.568 ;
      RECT 53.875 3.273 53.905 3.575 ;
      RECT 53.765 3.28 53.845 3.575 ;
      RECT 53.72 3.285 53.765 3.575 ;
      RECT 53.71 3.286 53.72 3.565 ;
      RECT 53.7 3.287 53.71 3.558 ;
      RECT 53.68 3.289 53.7 3.553 ;
      RECT 53.67 3.26 53.68 3.548 ;
      RECT 53.625 3.26 53.67 3.54 ;
      RECT 53.595 3.26 53.62 3.53 ;
      RECT 53.575 3.26 53.595 3.523 ;
      RECT 53.855 2.06 54.115 2.32 ;
      RECT 53.735 2.075 53.745 2.24 ;
      RECT 53.72 2.075 53.725 2.235 ;
      RECT 51.085 1.915 51.27 2.205 ;
      RECT 52.9 2.04 52.915 2.195 ;
      RECT 51.05 1.915 51.075 2.175 ;
      RECT 53.465 1.965 53.47 2.107 ;
      RECT 53.38 1.96 53.405 2.1 ;
      RECT 53.78 2.077 53.855 2.27 ;
      RECT 53.765 2.075 53.78 2.253 ;
      RECT 53.745 2.075 53.765 2.245 ;
      RECT 53.725 2.075 53.735 2.238 ;
      RECT 53.68 2.07 53.72 2.228 ;
      RECT 53.64 2.045 53.68 2.213 ;
      RECT 53.625 2.02 53.64 2.203 ;
      RECT 53.62 2.014 53.625 2.201 ;
      RECT 53.585 2.006 53.62 2.184 ;
      RECT 53.58 1.999 53.585 2.172 ;
      RECT 53.56 1.994 53.58 2.16 ;
      RECT 53.55 1.988 53.56 2.145 ;
      RECT 53.53 1.983 53.55 2.13 ;
      RECT 53.52 1.978 53.53 2.123 ;
      RECT 53.515 1.976 53.52 2.118 ;
      RECT 53.51 1.975 53.515 2.115 ;
      RECT 53.47 1.97 53.51 2.111 ;
      RECT 53.45 1.964 53.465 2.106 ;
      RECT 53.415 1.961 53.45 2.103 ;
      RECT 53.405 1.96 53.415 2.101 ;
      RECT 53.345 1.96 53.38 2.098 ;
      RECT 53.3 1.96 53.345 2.098 ;
      RECT 53.25 1.96 53.3 2.101 ;
      RECT 53.235 1.962 53.25 2.103 ;
      RECT 53.22 1.965 53.235 2.104 ;
      RECT 53.21 1.97 53.22 2.105 ;
      RECT 53.18 1.975 53.21 2.11 ;
      RECT 53.17 1.981 53.18 2.118 ;
      RECT 53.16 1.983 53.17 2.122 ;
      RECT 53.15 1.987 53.16 2.126 ;
      RECT 53.125 1.993 53.15 2.134 ;
      RECT 53.115 1.998 53.125 2.142 ;
      RECT 53.1 2.002 53.115 2.146 ;
      RECT 53.065 2.008 53.1 2.154 ;
      RECT 53.045 2.013 53.065 2.164 ;
      RECT 53.015 2.02 53.045 2.173 ;
      RECT 52.97 2.029 53.015 2.187 ;
      RECT 52.965 2.034 52.97 2.198 ;
      RECT 52.945 2.037 52.965 2.199 ;
      RECT 52.915 2.04 52.945 2.197 ;
      RECT 52.88 2.04 52.9 2.193 ;
      RECT 52.81 2.04 52.88 2.184 ;
      RECT 52.795 2.037 52.81 2.176 ;
      RECT 52.755 2.03 52.795 2.171 ;
      RECT 52.73 2.02 52.755 2.164 ;
      RECT 52.725 2.014 52.73 2.161 ;
      RECT 52.685 2.008 52.725 2.158 ;
      RECT 52.67 2.001 52.685 2.153 ;
      RECT 52.65 1.997 52.67 2.148 ;
      RECT 52.635 1.992 52.65 2.144 ;
      RECT 52.62 1.987 52.635 2.142 ;
      RECT 52.605 1.983 52.62 2.141 ;
      RECT 52.59 1.981 52.605 2.137 ;
      RECT 52.58 1.979 52.59 2.132 ;
      RECT 52.565 1.976 52.58 2.128 ;
      RECT 52.555 1.974 52.565 2.123 ;
      RECT 52.535 1.971 52.555 2.119 ;
      RECT 52.49 1.97 52.535 2.117 ;
      RECT 52.43 1.972 52.49 2.118 ;
      RECT 52.41 1.974 52.43 2.12 ;
      RECT 52.38 1.977 52.41 2.121 ;
      RECT 52.33 1.982 52.38 2.123 ;
      RECT 52.325 1.985 52.33 2.125 ;
      RECT 52.315 1.987 52.325 2.128 ;
      RECT 52.31 1.989 52.315 2.131 ;
      RECT 52.26 1.992 52.31 2.138 ;
      RECT 52.24 1.996 52.26 2.15 ;
      RECT 52.23 1.999 52.24 2.156 ;
      RECT 52.22 2 52.23 2.159 ;
      RECT 52.181 2.003 52.22 2.161 ;
      RECT 52.095 2.01 52.181 2.164 ;
      RECT 52.021 2.02 52.095 2.168 ;
      RECT 51.935 2.031 52.021 2.173 ;
      RECT 51.92 2.038 51.935 2.175 ;
      RECT 51.865 2.042 51.92 2.176 ;
      RECT 51.851 2.045 51.865 2.178 ;
      RECT 51.765 2.045 51.851 2.18 ;
      RECT 51.725 2.042 51.765 2.183 ;
      RECT 51.701 2.038 51.725 2.185 ;
      RECT 51.615 2.028 51.701 2.188 ;
      RECT 51.585 2.017 51.615 2.189 ;
      RECT 51.566 2.013 51.585 2.188 ;
      RECT 51.48 2.006 51.566 2.185 ;
      RECT 51.42 1.995 51.48 2.182 ;
      RECT 51.4 1.987 51.42 2.18 ;
      RECT 51.365 1.982 51.4 2.179 ;
      RECT 51.34 1.977 51.365 2.178 ;
      RECT 51.31 1.972 51.34 2.177 ;
      RECT 51.285 1.915 51.31 2.176 ;
      RECT 51.27 1.915 51.285 2.2 ;
      RECT 51.075 1.915 51.085 2.2 ;
      RECT 52.85 2.935 52.855 3.075 ;
      RECT 52.51 2.935 52.545 3.073 ;
      RECT 52.085 2.92 52.1 3.065 ;
      RECT 53.915 2.7 54.005 2.96 ;
      RECT 53.745 2.565 53.845 2.96 ;
      RECT 50.78 2.54 50.86 2.75 ;
      RECT 53.87 2.677 53.915 2.96 ;
      RECT 53.86 2.647 53.87 2.96 ;
      RECT 53.845 2.57 53.86 2.96 ;
      RECT 53.66 2.565 53.745 2.925 ;
      RECT 53.655 2.567 53.66 2.92 ;
      RECT 53.65 2.572 53.655 2.92 ;
      RECT 53.615 2.672 53.65 2.92 ;
      RECT 53.605 2.7 53.615 2.92 ;
      RECT 53.595 2.715 53.605 2.92 ;
      RECT 53.585 2.727 53.595 2.92 ;
      RECT 53.58 2.737 53.585 2.92 ;
      RECT 53.565 2.747 53.58 2.922 ;
      RECT 53.56 2.762 53.565 2.924 ;
      RECT 53.545 2.775 53.56 2.926 ;
      RECT 53.54 2.79 53.545 2.929 ;
      RECT 53.52 2.8 53.54 2.933 ;
      RECT 53.505 2.81 53.52 2.936 ;
      RECT 53.47 2.817 53.505 2.941 ;
      RECT 53.426 2.824 53.47 2.949 ;
      RECT 53.34 2.836 53.426 2.962 ;
      RECT 53.315 2.847 53.34 2.973 ;
      RECT 53.285 2.852 53.315 2.978 ;
      RECT 53.25 2.857 53.285 2.986 ;
      RECT 53.22 2.862 53.25 2.993 ;
      RECT 53.195 2.867 53.22 2.998 ;
      RECT 53.13 2.874 53.195 3.007 ;
      RECT 53.06 2.887 53.13 3.023 ;
      RECT 53.03 2.897 53.06 3.035 ;
      RECT 53.005 2.902 53.03 3.042 ;
      RECT 52.95 2.909 53.005 3.05 ;
      RECT 52.945 2.916 52.95 3.055 ;
      RECT 52.94 2.918 52.945 3.056 ;
      RECT 52.925 2.92 52.94 3.058 ;
      RECT 52.92 2.92 52.925 3.061 ;
      RECT 52.855 2.927 52.92 3.068 ;
      RECT 52.82 2.937 52.85 3.078 ;
      RECT 52.803 2.94 52.82 3.08 ;
      RECT 52.717 2.939 52.803 3.079 ;
      RECT 52.631 2.937 52.717 3.076 ;
      RECT 52.545 2.936 52.631 3.074 ;
      RECT 52.444 2.934 52.51 3.073 ;
      RECT 52.358 2.931 52.444 3.071 ;
      RECT 52.272 2.927 52.358 3.069 ;
      RECT 52.186 2.924 52.272 3.068 ;
      RECT 52.1 2.921 52.186 3.066 ;
      RECT 52 2.92 52.085 3.063 ;
      RECT 51.95 2.918 52 3.061 ;
      RECT 51.93 2.915 51.95 3.059 ;
      RECT 51.91 2.913 51.93 3.056 ;
      RECT 51.885 2.909 51.91 3.053 ;
      RECT 51.84 2.903 51.885 3.048 ;
      RECT 51.8 2.897 51.84 3.04 ;
      RECT 51.775 2.892 51.8 3.033 ;
      RECT 51.72 2.885 51.775 3.025 ;
      RECT 51.696 2.878 51.72 3.018 ;
      RECT 51.61 2.869 51.696 3.008 ;
      RECT 51.58 2.861 51.61 2.998 ;
      RECT 51.55 2.857 51.58 2.993 ;
      RECT 51.545 2.854 51.55 2.99 ;
      RECT 51.54 2.853 51.545 2.99 ;
      RECT 51.465 2.846 51.54 2.983 ;
      RECT 51.426 2.837 51.465 2.972 ;
      RECT 51.34 2.827 51.426 2.96 ;
      RECT 51.3 2.817 51.34 2.948 ;
      RECT 51.261 2.812 51.3 2.941 ;
      RECT 51.175 2.802 51.261 2.93 ;
      RECT 51.135 2.79 51.175 2.919 ;
      RECT 51.1 2.775 51.135 2.912 ;
      RECT 51.09 2.765 51.1 2.909 ;
      RECT 51.07 2.75 51.09 2.907 ;
      RECT 51.04 2.72 51.07 2.903 ;
      RECT 51.03 2.7 51.04 2.898 ;
      RECT 51.025 2.692 51.03 2.895 ;
      RECT 51.02 2.685 51.025 2.893 ;
      RECT 51.005 2.672 51.02 2.886 ;
      RECT 51 2.662 51.005 2.878 ;
      RECT 50.995 2.655 51 2.873 ;
      RECT 50.99 2.65 50.995 2.869 ;
      RECT 50.975 2.637 50.99 2.861 ;
      RECT 50.97 2.547 50.975 2.85 ;
      RECT 50.965 2.542 50.97 2.843 ;
      RECT 50.89 2.54 50.965 2.803 ;
      RECT 50.86 2.54 50.89 2.758 ;
      RECT 50.765 2.545 50.78 2.745 ;
      RECT 53.25 2.25 53.51 2.51 ;
      RECT 53.235 2.238 53.415 2.475 ;
      RECT 53.23 2.239 53.415 2.473 ;
      RECT 53.215 2.243 53.425 2.463 ;
      RECT 53.21 2.248 53.43 2.433 ;
      RECT 53.215 2.245 53.43 2.463 ;
      RECT 53.23 2.24 53.425 2.473 ;
      RECT 53.25 2.237 53.415 2.51 ;
      RECT 53.25 2.236 53.405 2.51 ;
      RECT 53.275 2.235 53.405 2.51 ;
      RECT 52.835 2.48 53.095 2.74 ;
      RECT 52.71 2.525 53.095 2.735 ;
      RECT 52.7 2.53 53.095 2.73 ;
      RECT 52.715 3.47 52.73 3.78 ;
      RECT 51.31 3.24 51.32 3.37 ;
      RECT 51.09 3.235 51.195 3.37 ;
      RECT 51.005 3.24 51.055 3.37 ;
      RECT 49.555 1.975 49.56 3.08 ;
      RECT 52.81 3.562 52.815 3.698 ;
      RECT 52.805 3.557 52.81 3.758 ;
      RECT 52.8 3.555 52.805 3.771 ;
      RECT 52.785 3.552 52.8 3.773 ;
      RECT 52.78 3.547 52.785 3.775 ;
      RECT 52.775 3.543 52.78 3.778 ;
      RECT 52.76 3.538 52.775 3.78 ;
      RECT 52.73 3.53 52.76 3.78 ;
      RECT 52.691 3.47 52.715 3.78 ;
      RECT 52.605 3.47 52.691 3.777 ;
      RECT 52.575 3.47 52.605 3.77 ;
      RECT 52.55 3.47 52.575 3.763 ;
      RECT 52.525 3.47 52.55 3.755 ;
      RECT 52.51 3.47 52.525 3.748 ;
      RECT 52.485 3.47 52.51 3.74 ;
      RECT 52.47 3.47 52.485 3.733 ;
      RECT 52.43 3.48 52.47 3.722 ;
      RECT 52.42 3.475 52.43 3.712 ;
      RECT 52.416 3.474 52.42 3.709 ;
      RECT 52.33 3.466 52.416 3.692 ;
      RECT 52.297 3.455 52.33 3.669 ;
      RECT 52.211 3.444 52.297 3.647 ;
      RECT 52.125 3.428 52.211 3.616 ;
      RECT 52.055 3.413 52.125 3.588 ;
      RECT 52.045 3.406 52.055 3.575 ;
      RECT 52.015 3.403 52.045 3.565 ;
      RECT 51.99 3.399 52.015 3.558 ;
      RECT 51.975 3.396 51.99 3.553 ;
      RECT 51.97 3.395 51.975 3.548 ;
      RECT 51.94 3.39 51.97 3.541 ;
      RECT 51.935 3.385 51.94 3.536 ;
      RECT 51.92 3.382 51.935 3.531 ;
      RECT 51.915 3.377 51.92 3.526 ;
      RECT 51.895 3.372 51.915 3.523 ;
      RECT 51.88 3.367 51.895 3.515 ;
      RECT 51.865 3.361 51.88 3.51 ;
      RECT 51.835 3.352 51.865 3.503 ;
      RECT 51.83 3.345 51.835 3.495 ;
      RECT 51.825 3.343 51.83 3.493 ;
      RECT 51.82 3.342 51.825 3.49 ;
      RECT 51.78 3.335 51.82 3.483 ;
      RECT 51.766 3.325 51.78 3.473 ;
      RECT 51.715 3.314 51.766 3.461 ;
      RECT 51.69 3.3 51.715 3.447 ;
      RECT 51.665 3.289 51.69 3.439 ;
      RECT 51.645 3.278 51.665 3.433 ;
      RECT 51.635 3.272 51.645 3.428 ;
      RECT 51.63 3.27 51.635 3.424 ;
      RECT 51.61 3.265 51.63 3.419 ;
      RECT 51.58 3.255 51.61 3.409 ;
      RECT 51.575 3.247 51.58 3.402 ;
      RECT 51.56 3.245 51.575 3.398 ;
      RECT 51.54 3.245 51.56 3.393 ;
      RECT 51.535 3.244 51.54 3.391 ;
      RECT 51.53 3.244 51.535 3.388 ;
      RECT 51.49 3.243 51.53 3.383 ;
      RECT 51.465 3.242 51.49 3.378 ;
      RECT 51.405 3.241 51.465 3.375 ;
      RECT 51.32 3.24 51.405 3.373 ;
      RECT 51.281 3.239 51.31 3.37 ;
      RECT 51.195 3.237 51.281 3.37 ;
      RECT 51.055 3.237 51.09 3.37 ;
      RECT 50.965 3.241 51.005 3.373 ;
      RECT 50.95 3.244 50.965 3.38 ;
      RECT 50.94 3.245 50.95 3.387 ;
      RECT 50.915 3.248 50.94 3.392 ;
      RECT 50.91 3.25 50.915 3.395 ;
      RECT 50.86 3.252 50.91 3.396 ;
      RECT 50.821 3.256 50.86 3.398 ;
      RECT 50.735 3.258 50.821 3.401 ;
      RECT 50.717 3.26 50.735 3.403 ;
      RECT 50.631 3.263 50.717 3.405 ;
      RECT 50.545 3.267 50.631 3.408 ;
      RECT 50.508 3.271 50.545 3.411 ;
      RECT 50.422 3.274 50.508 3.414 ;
      RECT 50.336 3.278 50.422 3.417 ;
      RECT 50.25 3.283 50.336 3.421 ;
      RECT 50.23 3.285 50.25 3.424 ;
      RECT 50.21 3.284 50.23 3.425 ;
      RECT 50.161 3.281 50.21 3.426 ;
      RECT 50.075 3.276 50.161 3.429 ;
      RECT 50.025 3.271 50.075 3.431 ;
      RECT 50.001 3.269 50.025 3.432 ;
      RECT 49.915 3.264 50.001 3.434 ;
      RECT 49.89 3.26 49.915 3.433 ;
      RECT 49.88 3.257 49.89 3.431 ;
      RECT 49.87 3.25 49.88 3.428 ;
      RECT 49.865 3.23 49.87 3.423 ;
      RECT 49.855 3.2 49.865 3.418 ;
      RECT 49.84 3.07 49.855 3.409 ;
      RECT 49.835 3.062 49.84 3.402 ;
      RECT 49.815 3.055 49.835 3.394 ;
      RECT 49.81 3.037 49.815 3.386 ;
      RECT 49.8 3.017 49.81 3.381 ;
      RECT 49.795 2.99 49.8 3.377 ;
      RECT 49.79 2.967 49.795 3.374 ;
      RECT 49.77 2.925 49.79 3.366 ;
      RECT 49.735 2.84 49.77 3.35 ;
      RECT 49.73 2.772 49.735 3.338 ;
      RECT 49.715 2.742 49.73 3.332 ;
      RECT 49.71 1.987 49.715 2.233 ;
      RECT 49.7 2.712 49.715 3.323 ;
      RECT 49.705 1.982 49.71 2.265 ;
      RECT 49.7 1.977 49.705 2.308 ;
      RECT 49.695 1.975 49.7 2.343 ;
      RECT 49.68 2.675 49.7 3.313 ;
      RECT 49.69 1.975 49.695 2.38 ;
      RECT 49.675 1.975 49.69 2.478 ;
      RECT 49.675 2.648 49.68 3.306 ;
      RECT 49.67 1.975 49.675 2.553 ;
      RECT 49.67 2.636 49.675 3.303 ;
      RECT 49.665 1.975 49.67 2.585 ;
      RECT 49.665 2.615 49.67 3.3 ;
      RECT 49.66 1.975 49.665 3.297 ;
      RECT 49.625 1.975 49.66 3.283 ;
      RECT 49.61 1.975 49.625 3.265 ;
      RECT 49.59 1.975 49.61 3.255 ;
      RECT 49.565 1.975 49.59 3.238 ;
      RECT 49.56 1.975 49.565 3.188 ;
      RECT 49.55 1.975 49.555 3.018 ;
      RECT 49.545 1.975 49.55 2.925 ;
      RECT 49.54 1.975 49.545 2.838 ;
      RECT 49.535 1.975 49.54 2.77 ;
      RECT 49.53 1.975 49.535 2.713 ;
      RECT 49.52 1.975 49.53 2.608 ;
      RECT 49.515 1.975 49.52 2.48 ;
      RECT 49.51 1.975 49.515 2.398 ;
      RECT 49.505 1.977 49.51 2.315 ;
      RECT 49.5 1.982 49.505 2.248 ;
      RECT 49.495 1.987 49.5 2.175 ;
      RECT 52.31 2.305 52.57 2.565 ;
      RECT 52.33 2.272 52.54 2.565 ;
      RECT 52.33 2.27 52.53 2.565 ;
      RECT 52.34 2.257 52.53 2.565 ;
      RECT 52.34 2.255 52.455 2.565 ;
      RECT 51.815 2.38 51.99 2.66 ;
      RECT 51.81 2.38 51.99 2.658 ;
      RECT 51.81 2.38 52.005 2.655 ;
      RECT 51.8 2.38 52.005 2.653 ;
      RECT 51.745 2.38 52.005 2.64 ;
      RECT 51.745 2.455 52.01 2.618 ;
      RECT 51.29 2.392 51.31 2.635 ;
      RECT 51.29 2.392 51.35 2.634 ;
      RECT 51.285 2.394 51.35 2.633 ;
      RECT 51.285 2.394 51.436 2.632 ;
      RECT 51.285 2.394 51.505 2.631 ;
      RECT 51.285 2.394 51.525 2.623 ;
      RECT 51.265 2.397 51.525 2.621 ;
      RECT 51.25 2.407 51.525 2.606 ;
      RECT 51.25 2.407 51.54 2.605 ;
      RECT 51.245 2.416 51.54 2.597 ;
      RECT 51.245 2.416 51.545 2.593 ;
      RECT 51.35 2.33 51.61 2.59 ;
      RECT 51.24 2.418 51.61 2.475 ;
      RECT 51.31 2.385 51.61 2.59 ;
      RECT 51.275 3.578 51.28 3.785 ;
      RECT 51.225 3.572 51.275 3.784 ;
      RECT 51.192 3.586 51.285 3.783 ;
      RECT 51.106 3.586 51.285 3.782 ;
      RECT 51.02 3.586 51.285 3.781 ;
      RECT 51.02 3.685 51.29 3.778 ;
      RECT 51.015 3.685 51.29 3.773 ;
      RECT 51.01 3.685 51.29 3.755 ;
      RECT 51.005 3.685 51.29 3.738 ;
      RECT 50.965 3.47 51.225 3.73 ;
      RECT 50.425 2.62 50.511 3.034 ;
      RECT 50.425 2.62 50.55 3.031 ;
      RECT 50.425 2.62 50.57 3.021 ;
      RECT 50.38 2.62 50.57 3.018 ;
      RECT 50.38 2.772 50.58 3.008 ;
      RECT 50.38 2.793 50.585 3.002 ;
      RECT 50.38 2.811 50.59 2.998 ;
      RECT 50.38 2.831 50.6 2.993 ;
      RECT 50.355 2.831 50.6 2.99 ;
      RECT 50.345 2.831 50.6 2.968 ;
      RECT 50.345 2.847 50.605 2.938 ;
      RECT 50.31 2.62 50.57 2.925 ;
      RECT 50.31 2.859 50.61 2.88 ;
      RECT 47.97 7.77 48.26 8 ;
      RECT 48.03 6.29 48.2 8 ;
      RECT 47.98 6.655 48.33 7.005 ;
      RECT 47.97 6.29 48.26 6.52 ;
      RECT 47.565 2.395 47.67 2.965 ;
      RECT 47.565 2.73 47.89 2.96 ;
      RECT 47.565 2.76 48.06 2.93 ;
      RECT 47.565 2.395 47.755 2.96 ;
      RECT 46.98 2.36 47.27 2.59 ;
      RECT 46.98 2.395 47.755 2.565 ;
      RECT 47.04 0.88 47.21 2.59 ;
      RECT 46.98 0.88 47.27 1.11 ;
      RECT 46.98 7.77 47.27 8 ;
      RECT 47.04 6.29 47.21 8 ;
      RECT 46.98 6.29 47.27 6.52 ;
      RECT 46.98 6.325 47.835 6.485 ;
      RECT 47.665 5.92 47.835 6.485 ;
      RECT 46.98 6.32 47.375 6.485 ;
      RECT 47.6 5.92 47.89 6.15 ;
      RECT 47.6 5.95 48.06 6.12 ;
      RECT 46.61 2.73 46.9 2.96 ;
      RECT 46.61 2.76 47.07 2.93 ;
      RECT 46.675 1.655 46.84 2.96 ;
      RECT 45.19 1.625 45.48 1.855 ;
      RECT 45.19 1.655 46.84 1.825 ;
      RECT 45.25 0.885 45.42 1.855 ;
      RECT 45.19 0.885 45.48 1.115 ;
      RECT 45.19 7.765 45.48 7.995 ;
      RECT 45.25 7.025 45.42 7.995 ;
      RECT 45.25 7.12 46.84 7.29 ;
      RECT 46.67 5.92 46.84 7.29 ;
      RECT 45.19 7.025 45.48 7.255 ;
      RECT 46.61 5.92 46.9 6.15 ;
      RECT 46.61 5.95 47.07 6.12 ;
      RECT 43.24 2.705 43.58 3.055 ;
      RECT 43.33 2.025 43.5 3.055 ;
      RECT 45.62 1.965 45.97 2.315 ;
      RECT 43.33 2.025 45.97 2.195 ;
      RECT 45.645 6.655 45.97 6.98 ;
      RECT 40.185 6.615 40.535 6.965 ;
      RECT 45.62 6.655 45.97 6.885 ;
      RECT 39.985 6.655 40.535 6.885 ;
      RECT 39.815 6.685 45.97 6.855 ;
      RECT 44.845 2.365 45.165 2.685 ;
      RECT 44.815 2.365 45.165 2.595 ;
      RECT 44.645 2.395 45.165 2.565 ;
      RECT 44.845 6.255 45.165 6.545 ;
      RECT 44.815 6.285 45.165 6.515 ;
      RECT 44.645 6.315 45.165 6.485 ;
      RECT 40.535 2.985 40.685 3.26 ;
      RECT 41.075 2.065 41.08 2.285 ;
      RECT 42.225 2.265 42.24 2.463 ;
      RECT 42.19 2.257 42.225 2.47 ;
      RECT 42.16 2.25 42.19 2.47 ;
      RECT 42.105 2.215 42.16 2.47 ;
      RECT 42.04 2.152 42.105 2.47 ;
      RECT 42.035 2.117 42.04 2.468 ;
      RECT 42.03 2.112 42.035 2.46 ;
      RECT 42.025 2.107 42.03 2.446 ;
      RECT 42.02 2.104 42.025 2.439 ;
      RECT 41.975 2.094 42.02 2.39 ;
      RECT 41.955 2.081 41.975 2.325 ;
      RECT 41.95 2.076 41.955 2.298 ;
      RECT 41.945 2.075 41.95 2.291 ;
      RECT 41.94 2.074 41.945 2.284 ;
      RECT 41.855 2.059 41.94 2.23 ;
      RECT 41.825 2.04 41.855 2.18 ;
      RECT 41.745 2.023 41.825 2.165 ;
      RECT 41.71 2.01 41.745 2.15 ;
      RECT 41.702 2.01 41.71 2.145 ;
      RECT 41.616 2.011 41.702 2.145 ;
      RECT 41.53 2.013 41.616 2.145 ;
      RECT 41.505 2.014 41.53 2.149 ;
      RECT 41.43 2.02 41.505 2.164 ;
      RECT 41.347 2.032 41.43 2.188 ;
      RECT 41.261 2.045 41.347 2.214 ;
      RECT 41.175 2.058 41.261 2.24 ;
      RECT 41.14 2.067 41.175 2.259 ;
      RECT 41.09 2.067 41.14 2.272 ;
      RECT 41.08 2.065 41.09 2.283 ;
      RECT 41.065 2.062 41.075 2.285 ;
      RECT 41.05 2.054 41.065 2.293 ;
      RECT 41.035 2.046 41.05 2.313 ;
      RECT 41.03 2.041 41.035 2.37 ;
      RECT 41.015 2.036 41.03 2.443 ;
      RECT 41.01 2.031 41.015 2.485 ;
      RECT 41.005 2.029 41.01 2.513 ;
      RECT 41 2.027 41.005 2.535 ;
      RECT 40.99 2.023 41 2.578 ;
      RECT 40.985 2.02 40.99 2.603 ;
      RECT 40.98 2.018 40.985 2.623 ;
      RECT 40.975 2.016 40.98 2.647 ;
      RECT 40.97 2.012 40.975 2.67 ;
      RECT 40.965 2.008 40.97 2.693 ;
      RECT 40.93 1.998 40.965 2.8 ;
      RECT 40.925 1.988 40.93 2.898 ;
      RECT 40.92 1.986 40.925 2.925 ;
      RECT 40.915 1.985 40.92 2.945 ;
      RECT 40.91 1.977 40.915 2.965 ;
      RECT 40.905 1.972 40.91 3 ;
      RECT 40.9 1.97 40.905 3.018 ;
      RECT 40.895 1.97 40.9 3.043 ;
      RECT 40.89 1.97 40.895 3.065 ;
      RECT 40.855 1.97 40.89 3.108 ;
      RECT 40.83 1.97 40.855 3.137 ;
      RECT 40.82 1.97 40.83 2.323 ;
      RECT 40.823 2.38 40.83 3.147 ;
      RECT 40.82 2.437 40.823 3.15 ;
      RECT 40.815 1.97 40.82 2.295 ;
      RECT 40.815 2.487 40.82 3.153 ;
      RECT 40.805 1.97 40.815 2.285 ;
      RECT 40.81 2.54 40.815 3.156 ;
      RECT 40.805 2.625 40.81 3.16 ;
      RECT 40.795 1.97 40.805 2.273 ;
      RECT 40.8 2.672 40.805 3.164 ;
      RECT 40.795 2.747 40.8 3.168 ;
      RECT 40.76 1.97 40.795 2.248 ;
      RECT 40.785 2.83 40.795 3.173 ;
      RECT 40.775 2.897 40.785 3.18 ;
      RECT 40.77 2.925 40.775 3.185 ;
      RECT 40.76 2.938 40.77 3.191 ;
      RECT 40.715 1.97 40.76 2.205 ;
      RECT 40.755 2.943 40.76 3.198 ;
      RECT 40.715 2.96 40.755 3.26 ;
      RECT 40.71 1.972 40.715 2.178 ;
      RECT 40.685 2.98 40.715 3.26 ;
      RECT 40.705 1.977 40.71 2.15 ;
      RECT 40.495 2.989 40.535 3.26 ;
      RECT 40.47 2.997 40.495 3.23 ;
      RECT 40.425 3.005 40.47 3.23 ;
      RECT 40.41 3.01 40.425 3.225 ;
      RECT 40.4 3.01 40.41 3.219 ;
      RECT 40.39 3.017 40.4 3.216 ;
      RECT 40.385 3.055 40.39 3.205 ;
      RECT 40.38 3.117 40.385 3.183 ;
      RECT 41.65 2.992 41.835 3.215 ;
      RECT 41.65 3.007 41.84 3.211 ;
      RECT 41.64 2.28 41.725 3.21 ;
      RECT 41.64 3.007 41.845 3.204 ;
      RECT 41.635 3.015 41.845 3.203 ;
      RECT 41.84 2.735 42.16 3.055 ;
      RECT 41.635 2.907 41.805 2.998 ;
      RECT 41.63 2.907 41.805 2.98 ;
      RECT 41.62 2.715 41.755 2.955 ;
      RECT 41.615 2.715 41.755 2.9 ;
      RECT 41.575 2.295 41.745 2.8 ;
      RECT 41.56 2.295 41.745 2.67 ;
      RECT 41.555 2.295 41.745 2.623 ;
      RECT 41.55 2.295 41.745 2.603 ;
      RECT 41.545 2.295 41.745 2.578 ;
      RECT 41.515 2.295 41.775 2.555 ;
      RECT 41.525 2.292 41.735 2.555 ;
      RECT 41.65 2.287 41.735 3.215 ;
      RECT 41.535 2.28 41.725 2.555 ;
      RECT 41.53 2.285 41.725 2.555 ;
      RECT 40.36 2.497 40.545 2.71 ;
      RECT 40.36 2.505 40.555 2.703 ;
      RECT 40.34 2.505 40.555 2.7 ;
      RECT 40.335 2.505 40.555 2.685 ;
      RECT 40.265 2.42 40.525 2.68 ;
      RECT 40.265 2.565 40.56 2.593 ;
      RECT 39.92 3.02 40.18 3.28 ;
      RECT 39.945 2.965 40.14 3.28 ;
      RECT 39.94 2.714 40.12 3.008 ;
      RECT 39.94 2.72 40.13 3.008 ;
      RECT 39.92 2.722 40.13 2.953 ;
      RECT 39.915 2.732 40.13 2.82 ;
      RECT 39.945 2.712 40.12 3.28 ;
      RECT 40.031 2.71 40.12 3.28 ;
      RECT 39.89 1.93 39.925 2.3 ;
      RECT 39.68 2.04 39.685 2.3 ;
      RECT 39.925 1.937 39.94 2.3 ;
      RECT 39.815 1.93 39.89 2.378 ;
      RECT 39.805 1.93 39.815 2.463 ;
      RECT 39.78 1.93 39.805 2.498 ;
      RECT 39.74 1.93 39.78 2.566 ;
      RECT 39.73 1.937 39.74 2.618 ;
      RECT 39.7 2.04 39.73 2.659 ;
      RECT 39.695 2.04 39.7 2.698 ;
      RECT 39.685 2.04 39.695 2.718 ;
      RECT 39.68 2.335 39.685 2.755 ;
      RECT 39.675 2.352 39.68 2.775 ;
      RECT 39.66 2.415 39.675 2.815 ;
      RECT 39.655 2.458 39.66 2.85 ;
      RECT 39.65 2.466 39.655 2.863 ;
      RECT 39.64 2.48 39.65 2.885 ;
      RECT 39.615 2.515 39.64 2.95 ;
      RECT 39.605 2.55 39.615 3.013 ;
      RECT 39.585 2.58 39.605 3.074 ;
      RECT 39.57 2.616 39.585 3.141 ;
      RECT 39.56 2.644 39.57 3.18 ;
      RECT 39.55 2.666 39.56 3.2 ;
      RECT 39.545 2.676 39.55 3.211 ;
      RECT 39.54 2.685 39.545 3.214 ;
      RECT 39.53 2.703 39.54 3.218 ;
      RECT 39.52 2.721 39.53 3.219 ;
      RECT 39.495 2.76 39.52 3.216 ;
      RECT 39.475 2.802 39.495 3.213 ;
      RECT 39.46 2.84 39.475 3.212 ;
      RECT 39.425 2.875 39.46 3.209 ;
      RECT 39.42 2.897 39.425 3.207 ;
      RECT 39.355 2.937 39.42 3.204 ;
      RECT 39.35 2.977 39.355 3.2 ;
      RECT 39.335 2.987 39.35 3.191 ;
      RECT 39.325 3.107 39.335 3.176 ;
      RECT 39.805 3.52 39.815 3.78 ;
      RECT 39.805 3.523 39.825 3.779 ;
      RECT 39.795 3.513 39.805 3.778 ;
      RECT 39.785 3.528 39.865 3.774 ;
      RECT 39.77 3.507 39.785 3.772 ;
      RECT 39.745 3.532 39.87 3.768 ;
      RECT 39.73 3.492 39.745 3.763 ;
      RECT 39.73 3.534 39.88 3.762 ;
      RECT 39.73 3.542 39.895 3.755 ;
      RECT 39.67 3.479 39.73 3.745 ;
      RECT 39.66 3.466 39.67 3.727 ;
      RECT 39.635 3.456 39.66 3.717 ;
      RECT 39.63 3.446 39.635 3.709 ;
      RECT 39.565 3.542 39.895 3.691 ;
      RECT 39.48 3.542 39.895 3.653 ;
      RECT 39.37 3.37 39.63 3.63 ;
      RECT 39.745 3.5 39.77 3.768 ;
      RECT 39.785 3.51 39.795 3.774 ;
      RECT 39.37 3.518 39.81 3.63 ;
      RECT 39.555 7.765 39.845 7.995 ;
      RECT 39.615 7.025 39.785 7.995 ;
      RECT 39.515 7.055 39.885 7.425 ;
      RECT 39.555 7.025 39.845 7.425 ;
      RECT 38.585 3.275 38.615 3.575 ;
      RECT 38.36 3.26 38.365 3.535 ;
      RECT 38.16 3.26 38.315 3.52 ;
      RECT 39.46 1.975 39.49 2.235 ;
      RECT 39.45 1.975 39.46 2.343 ;
      RECT 39.43 1.975 39.45 2.353 ;
      RECT 39.415 1.975 39.43 2.365 ;
      RECT 39.36 1.975 39.415 2.415 ;
      RECT 39.345 1.975 39.36 2.463 ;
      RECT 39.315 1.975 39.345 2.498 ;
      RECT 39.26 1.975 39.315 2.56 ;
      RECT 39.24 1.975 39.26 2.628 ;
      RECT 39.235 1.975 39.24 2.658 ;
      RECT 39.23 1.975 39.235 2.67 ;
      RECT 39.225 2.092 39.23 2.688 ;
      RECT 39.205 2.11 39.225 2.713 ;
      RECT 39.185 2.137 39.205 2.763 ;
      RECT 39.18 2.157 39.185 2.794 ;
      RECT 39.175 2.165 39.18 2.811 ;
      RECT 39.16 2.191 39.175 2.84 ;
      RECT 39.145 2.233 39.16 2.875 ;
      RECT 39.14 2.262 39.145 2.898 ;
      RECT 39.135 2.277 39.14 2.911 ;
      RECT 39.13 2.3 39.135 2.922 ;
      RECT 39.12 2.32 39.13 2.94 ;
      RECT 39.11 2.35 39.12 2.963 ;
      RECT 39.105 2.372 39.11 2.983 ;
      RECT 39.1 2.387 39.105 2.998 ;
      RECT 39.085 2.417 39.1 3.025 ;
      RECT 39.08 2.447 39.085 3.051 ;
      RECT 39.075 2.465 39.08 3.063 ;
      RECT 39.065 2.495 39.075 3.082 ;
      RECT 39.055 2.52 39.065 3.107 ;
      RECT 39.05 2.54 39.055 3.126 ;
      RECT 39.045 2.557 39.05 3.139 ;
      RECT 39.035 2.583 39.045 3.158 ;
      RECT 39.025 2.621 39.035 3.185 ;
      RECT 39.02 2.647 39.025 3.205 ;
      RECT 39.015 2.657 39.02 3.215 ;
      RECT 39.01 2.67 39.015 3.23 ;
      RECT 39.005 2.685 39.01 3.24 ;
      RECT 39 2.707 39.005 3.255 ;
      RECT 38.995 2.725 39 3.266 ;
      RECT 38.99 2.735 38.995 3.277 ;
      RECT 38.985 2.743 38.99 3.289 ;
      RECT 38.98 2.751 38.985 3.3 ;
      RECT 38.975 2.777 38.98 3.313 ;
      RECT 38.965 2.805 38.975 3.326 ;
      RECT 38.96 2.835 38.965 3.335 ;
      RECT 38.955 2.85 38.96 3.342 ;
      RECT 38.94 2.875 38.955 3.349 ;
      RECT 38.935 2.897 38.94 3.355 ;
      RECT 38.93 2.922 38.935 3.358 ;
      RECT 38.921 2.95 38.93 3.362 ;
      RECT 38.915 2.967 38.921 3.367 ;
      RECT 38.91 2.985 38.915 3.371 ;
      RECT 38.905 2.997 38.91 3.374 ;
      RECT 38.9 3.018 38.905 3.378 ;
      RECT 38.895 3.036 38.9 3.381 ;
      RECT 38.89 3.05 38.895 3.384 ;
      RECT 38.885 3.067 38.89 3.387 ;
      RECT 38.88 3.08 38.885 3.39 ;
      RECT 38.855 3.117 38.88 3.398 ;
      RECT 38.85 3.162 38.855 3.407 ;
      RECT 38.845 3.19 38.85 3.41 ;
      RECT 38.835 3.21 38.845 3.414 ;
      RECT 38.83 3.23 38.835 3.419 ;
      RECT 38.825 3.245 38.83 3.422 ;
      RECT 38.805 3.255 38.825 3.429 ;
      RECT 38.74 3.262 38.805 3.455 ;
      RECT 38.705 3.265 38.74 3.483 ;
      RECT 38.69 3.268 38.705 3.498 ;
      RECT 38.68 3.269 38.69 3.513 ;
      RECT 38.67 3.27 38.68 3.53 ;
      RECT 38.665 3.27 38.67 3.545 ;
      RECT 38.66 3.27 38.665 3.553 ;
      RECT 38.645 3.271 38.66 3.568 ;
      RECT 38.615 3.273 38.645 3.575 ;
      RECT 38.505 3.28 38.585 3.575 ;
      RECT 38.46 3.285 38.505 3.575 ;
      RECT 38.45 3.286 38.46 3.565 ;
      RECT 38.44 3.287 38.45 3.558 ;
      RECT 38.42 3.289 38.44 3.553 ;
      RECT 38.41 3.26 38.42 3.548 ;
      RECT 38.365 3.26 38.41 3.54 ;
      RECT 38.335 3.26 38.36 3.53 ;
      RECT 38.315 3.26 38.335 3.523 ;
      RECT 38.595 2.06 38.855 2.32 ;
      RECT 38.475 2.075 38.485 2.24 ;
      RECT 38.46 2.075 38.465 2.235 ;
      RECT 35.825 1.915 36.01 2.205 ;
      RECT 37.64 2.04 37.655 2.195 ;
      RECT 35.79 1.915 35.815 2.175 ;
      RECT 38.205 1.965 38.21 2.107 ;
      RECT 38.12 1.96 38.145 2.1 ;
      RECT 38.52 2.077 38.595 2.27 ;
      RECT 38.505 2.075 38.52 2.253 ;
      RECT 38.485 2.075 38.505 2.245 ;
      RECT 38.465 2.075 38.475 2.238 ;
      RECT 38.42 2.07 38.46 2.228 ;
      RECT 38.38 2.045 38.42 2.213 ;
      RECT 38.365 2.02 38.38 2.203 ;
      RECT 38.36 2.014 38.365 2.201 ;
      RECT 38.325 2.006 38.36 2.184 ;
      RECT 38.32 1.999 38.325 2.172 ;
      RECT 38.3 1.994 38.32 2.16 ;
      RECT 38.29 1.988 38.3 2.145 ;
      RECT 38.27 1.983 38.29 2.13 ;
      RECT 38.26 1.978 38.27 2.123 ;
      RECT 38.255 1.976 38.26 2.118 ;
      RECT 38.25 1.975 38.255 2.115 ;
      RECT 38.21 1.97 38.25 2.111 ;
      RECT 38.19 1.964 38.205 2.106 ;
      RECT 38.155 1.961 38.19 2.103 ;
      RECT 38.145 1.96 38.155 2.101 ;
      RECT 38.085 1.96 38.12 2.098 ;
      RECT 38.04 1.96 38.085 2.098 ;
      RECT 37.99 1.96 38.04 2.101 ;
      RECT 37.975 1.962 37.99 2.103 ;
      RECT 37.96 1.965 37.975 2.104 ;
      RECT 37.95 1.97 37.96 2.105 ;
      RECT 37.92 1.975 37.95 2.11 ;
      RECT 37.91 1.981 37.92 2.118 ;
      RECT 37.9 1.983 37.91 2.122 ;
      RECT 37.89 1.987 37.9 2.126 ;
      RECT 37.865 1.993 37.89 2.134 ;
      RECT 37.855 1.998 37.865 2.142 ;
      RECT 37.84 2.002 37.855 2.146 ;
      RECT 37.805 2.008 37.84 2.154 ;
      RECT 37.785 2.013 37.805 2.164 ;
      RECT 37.755 2.02 37.785 2.173 ;
      RECT 37.71 2.029 37.755 2.187 ;
      RECT 37.705 2.034 37.71 2.198 ;
      RECT 37.685 2.037 37.705 2.199 ;
      RECT 37.655 2.04 37.685 2.197 ;
      RECT 37.62 2.04 37.64 2.193 ;
      RECT 37.55 2.04 37.62 2.184 ;
      RECT 37.535 2.037 37.55 2.176 ;
      RECT 37.495 2.03 37.535 2.171 ;
      RECT 37.47 2.02 37.495 2.164 ;
      RECT 37.465 2.014 37.47 2.161 ;
      RECT 37.425 2.008 37.465 2.158 ;
      RECT 37.41 2.001 37.425 2.153 ;
      RECT 37.39 1.997 37.41 2.148 ;
      RECT 37.375 1.992 37.39 2.144 ;
      RECT 37.36 1.987 37.375 2.142 ;
      RECT 37.345 1.983 37.36 2.141 ;
      RECT 37.33 1.981 37.345 2.137 ;
      RECT 37.32 1.979 37.33 2.132 ;
      RECT 37.305 1.976 37.32 2.128 ;
      RECT 37.295 1.974 37.305 2.123 ;
      RECT 37.275 1.971 37.295 2.119 ;
      RECT 37.23 1.97 37.275 2.117 ;
      RECT 37.17 1.972 37.23 2.118 ;
      RECT 37.15 1.974 37.17 2.12 ;
      RECT 37.12 1.977 37.15 2.121 ;
      RECT 37.07 1.982 37.12 2.123 ;
      RECT 37.065 1.985 37.07 2.125 ;
      RECT 37.055 1.987 37.065 2.128 ;
      RECT 37.05 1.989 37.055 2.131 ;
      RECT 37 1.992 37.05 2.138 ;
      RECT 36.98 1.996 37 2.15 ;
      RECT 36.97 1.999 36.98 2.156 ;
      RECT 36.96 2 36.97 2.159 ;
      RECT 36.921 2.003 36.96 2.161 ;
      RECT 36.835 2.01 36.921 2.164 ;
      RECT 36.761 2.02 36.835 2.168 ;
      RECT 36.675 2.031 36.761 2.173 ;
      RECT 36.66 2.038 36.675 2.175 ;
      RECT 36.605 2.042 36.66 2.176 ;
      RECT 36.591 2.045 36.605 2.178 ;
      RECT 36.505 2.045 36.591 2.18 ;
      RECT 36.465 2.042 36.505 2.183 ;
      RECT 36.441 2.038 36.465 2.185 ;
      RECT 36.355 2.028 36.441 2.188 ;
      RECT 36.325 2.017 36.355 2.189 ;
      RECT 36.306 2.013 36.325 2.188 ;
      RECT 36.22 2.006 36.306 2.185 ;
      RECT 36.16 1.995 36.22 2.182 ;
      RECT 36.14 1.987 36.16 2.18 ;
      RECT 36.105 1.982 36.14 2.179 ;
      RECT 36.08 1.977 36.105 2.178 ;
      RECT 36.05 1.972 36.08 2.177 ;
      RECT 36.025 1.915 36.05 2.176 ;
      RECT 36.01 1.915 36.025 2.2 ;
      RECT 35.815 1.915 35.825 2.2 ;
      RECT 37.59 2.935 37.595 3.075 ;
      RECT 37.25 2.935 37.285 3.073 ;
      RECT 36.825 2.92 36.84 3.065 ;
      RECT 38.655 2.7 38.745 2.96 ;
      RECT 38.485 2.565 38.585 2.96 ;
      RECT 35.52 2.54 35.6 2.75 ;
      RECT 38.61 2.677 38.655 2.96 ;
      RECT 38.6 2.647 38.61 2.96 ;
      RECT 38.585 2.57 38.6 2.96 ;
      RECT 38.4 2.565 38.485 2.925 ;
      RECT 38.395 2.567 38.4 2.92 ;
      RECT 38.39 2.572 38.395 2.92 ;
      RECT 38.355 2.672 38.39 2.92 ;
      RECT 38.345 2.7 38.355 2.92 ;
      RECT 38.335 2.715 38.345 2.92 ;
      RECT 38.325 2.727 38.335 2.92 ;
      RECT 38.32 2.737 38.325 2.92 ;
      RECT 38.305 2.747 38.32 2.922 ;
      RECT 38.3 2.762 38.305 2.924 ;
      RECT 38.285 2.775 38.3 2.926 ;
      RECT 38.28 2.79 38.285 2.929 ;
      RECT 38.26 2.8 38.28 2.933 ;
      RECT 38.245 2.81 38.26 2.936 ;
      RECT 38.21 2.817 38.245 2.941 ;
      RECT 38.166 2.824 38.21 2.949 ;
      RECT 38.08 2.836 38.166 2.962 ;
      RECT 38.055 2.847 38.08 2.973 ;
      RECT 38.025 2.852 38.055 2.978 ;
      RECT 37.99 2.857 38.025 2.986 ;
      RECT 37.96 2.862 37.99 2.993 ;
      RECT 37.935 2.867 37.96 2.998 ;
      RECT 37.87 2.874 37.935 3.007 ;
      RECT 37.8 2.887 37.87 3.023 ;
      RECT 37.77 2.897 37.8 3.035 ;
      RECT 37.745 2.902 37.77 3.042 ;
      RECT 37.69 2.909 37.745 3.05 ;
      RECT 37.685 2.916 37.69 3.055 ;
      RECT 37.68 2.918 37.685 3.056 ;
      RECT 37.665 2.92 37.68 3.058 ;
      RECT 37.66 2.92 37.665 3.061 ;
      RECT 37.595 2.927 37.66 3.068 ;
      RECT 37.56 2.937 37.59 3.078 ;
      RECT 37.543 2.94 37.56 3.08 ;
      RECT 37.457 2.939 37.543 3.079 ;
      RECT 37.371 2.937 37.457 3.076 ;
      RECT 37.285 2.936 37.371 3.074 ;
      RECT 37.184 2.934 37.25 3.073 ;
      RECT 37.098 2.931 37.184 3.071 ;
      RECT 37.012 2.927 37.098 3.069 ;
      RECT 36.926 2.924 37.012 3.068 ;
      RECT 36.84 2.921 36.926 3.066 ;
      RECT 36.74 2.92 36.825 3.063 ;
      RECT 36.69 2.918 36.74 3.061 ;
      RECT 36.67 2.915 36.69 3.059 ;
      RECT 36.65 2.913 36.67 3.056 ;
      RECT 36.625 2.909 36.65 3.053 ;
      RECT 36.58 2.903 36.625 3.048 ;
      RECT 36.54 2.897 36.58 3.04 ;
      RECT 36.515 2.892 36.54 3.033 ;
      RECT 36.46 2.885 36.515 3.025 ;
      RECT 36.436 2.878 36.46 3.018 ;
      RECT 36.35 2.869 36.436 3.008 ;
      RECT 36.32 2.861 36.35 2.998 ;
      RECT 36.29 2.857 36.32 2.993 ;
      RECT 36.285 2.854 36.29 2.99 ;
      RECT 36.28 2.853 36.285 2.99 ;
      RECT 36.205 2.846 36.28 2.983 ;
      RECT 36.166 2.837 36.205 2.972 ;
      RECT 36.08 2.827 36.166 2.96 ;
      RECT 36.04 2.817 36.08 2.948 ;
      RECT 36.001 2.812 36.04 2.941 ;
      RECT 35.915 2.802 36.001 2.93 ;
      RECT 35.875 2.79 35.915 2.919 ;
      RECT 35.84 2.775 35.875 2.912 ;
      RECT 35.83 2.765 35.84 2.909 ;
      RECT 35.81 2.75 35.83 2.907 ;
      RECT 35.78 2.72 35.81 2.903 ;
      RECT 35.77 2.7 35.78 2.898 ;
      RECT 35.765 2.692 35.77 2.895 ;
      RECT 35.76 2.685 35.765 2.893 ;
      RECT 35.745 2.672 35.76 2.886 ;
      RECT 35.74 2.662 35.745 2.878 ;
      RECT 35.735 2.655 35.74 2.873 ;
      RECT 35.73 2.65 35.735 2.869 ;
      RECT 35.715 2.637 35.73 2.861 ;
      RECT 35.71 2.547 35.715 2.85 ;
      RECT 35.705 2.542 35.71 2.843 ;
      RECT 35.63 2.54 35.705 2.803 ;
      RECT 35.6 2.54 35.63 2.758 ;
      RECT 35.505 2.545 35.52 2.745 ;
      RECT 37.99 2.25 38.25 2.51 ;
      RECT 37.975 2.238 38.155 2.475 ;
      RECT 37.97 2.239 38.155 2.473 ;
      RECT 37.955 2.243 38.165 2.463 ;
      RECT 37.95 2.248 38.17 2.433 ;
      RECT 37.955 2.245 38.17 2.463 ;
      RECT 37.97 2.24 38.165 2.473 ;
      RECT 37.99 2.237 38.155 2.51 ;
      RECT 37.99 2.236 38.145 2.51 ;
      RECT 38.015 2.235 38.145 2.51 ;
      RECT 37.575 2.48 37.835 2.74 ;
      RECT 37.45 2.525 37.835 2.735 ;
      RECT 37.44 2.53 37.835 2.73 ;
      RECT 37.455 3.47 37.47 3.78 ;
      RECT 36.05 3.24 36.06 3.37 ;
      RECT 35.83 3.235 35.935 3.37 ;
      RECT 35.745 3.24 35.795 3.37 ;
      RECT 34.295 1.975 34.3 3.08 ;
      RECT 37.55 3.562 37.555 3.698 ;
      RECT 37.545 3.557 37.55 3.758 ;
      RECT 37.54 3.555 37.545 3.771 ;
      RECT 37.525 3.552 37.54 3.773 ;
      RECT 37.52 3.547 37.525 3.775 ;
      RECT 37.515 3.543 37.52 3.778 ;
      RECT 37.5 3.538 37.515 3.78 ;
      RECT 37.47 3.53 37.5 3.78 ;
      RECT 37.431 3.47 37.455 3.78 ;
      RECT 37.345 3.47 37.431 3.777 ;
      RECT 37.315 3.47 37.345 3.77 ;
      RECT 37.29 3.47 37.315 3.763 ;
      RECT 37.265 3.47 37.29 3.755 ;
      RECT 37.25 3.47 37.265 3.748 ;
      RECT 37.225 3.47 37.25 3.74 ;
      RECT 37.21 3.47 37.225 3.733 ;
      RECT 37.17 3.48 37.21 3.722 ;
      RECT 37.16 3.475 37.17 3.712 ;
      RECT 37.156 3.474 37.16 3.709 ;
      RECT 37.07 3.466 37.156 3.692 ;
      RECT 37.037 3.455 37.07 3.669 ;
      RECT 36.951 3.444 37.037 3.647 ;
      RECT 36.865 3.428 36.951 3.616 ;
      RECT 36.795 3.413 36.865 3.588 ;
      RECT 36.785 3.406 36.795 3.575 ;
      RECT 36.755 3.403 36.785 3.565 ;
      RECT 36.73 3.399 36.755 3.558 ;
      RECT 36.715 3.396 36.73 3.553 ;
      RECT 36.71 3.395 36.715 3.548 ;
      RECT 36.68 3.39 36.71 3.541 ;
      RECT 36.675 3.385 36.68 3.536 ;
      RECT 36.66 3.382 36.675 3.531 ;
      RECT 36.655 3.377 36.66 3.526 ;
      RECT 36.635 3.372 36.655 3.523 ;
      RECT 36.62 3.367 36.635 3.515 ;
      RECT 36.605 3.361 36.62 3.51 ;
      RECT 36.575 3.352 36.605 3.503 ;
      RECT 36.57 3.345 36.575 3.495 ;
      RECT 36.565 3.343 36.57 3.493 ;
      RECT 36.56 3.342 36.565 3.49 ;
      RECT 36.52 3.335 36.56 3.483 ;
      RECT 36.506 3.325 36.52 3.473 ;
      RECT 36.455 3.314 36.506 3.461 ;
      RECT 36.43 3.3 36.455 3.447 ;
      RECT 36.405 3.289 36.43 3.439 ;
      RECT 36.385 3.278 36.405 3.433 ;
      RECT 36.375 3.272 36.385 3.428 ;
      RECT 36.37 3.27 36.375 3.424 ;
      RECT 36.35 3.265 36.37 3.419 ;
      RECT 36.32 3.255 36.35 3.409 ;
      RECT 36.315 3.247 36.32 3.402 ;
      RECT 36.3 3.245 36.315 3.398 ;
      RECT 36.28 3.245 36.3 3.393 ;
      RECT 36.275 3.244 36.28 3.391 ;
      RECT 36.27 3.244 36.275 3.388 ;
      RECT 36.23 3.243 36.27 3.383 ;
      RECT 36.205 3.242 36.23 3.378 ;
      RECT 36.145 3.241 36.205 3.375 ;
      RECT 36.06 3.24 36.145 3.373 ;
      RECT 36.021 3.239 36.05 3.37 ;
      RECT 35.935 3.237 36.021 3.37 ;
      RECT 35.795 3.237 35.83 3.37 ;
      RECT 35.705 3.241 35.745 3.373 ;
      RECT 35.69 3.244 35.705 3.38 ;
      RECT 35.68 3.245 35.69 3.387 ;
      RECT 35.655 3.248 35.68 3.392 ;
      RECT 35.65 3.25 35.655 3.395 ;
      RECT 35.6 3.252 35.65 3.396 ;
      RECT 35.561 3.256 35.6 3.398 ;
      RECT 35.475 3.258 35.561 3.401 ;
      RECT 35.457 3.26 35.475 3.403 ;
      RECT 35.371 3.263 35.457 3.405 ;
      RECT 35.285 3.267 35.371 3.408 ;
      RECT 35.248 3.271 35.285 3.411 ;
      RECT 35.162 3.274 35.248 3.414 ;
      RECT 35.076 3.278 35.162 3.417 ;
      RECT 34.99 3.283 35.076 3.421 ;
      RECT 34.97 3.285 34.99 3.424 ;
      RECT 34.95 3.284 34.97 3.425 ;
      RECT 34.901 3.281 34.95 3.426 ;
      RECT 34.815 3.276 34.901 3.429 ;
      RECT 34.765 3.271 34.815 3.431 ;
      RECT 34.741 3.269 34.765 3.432 ;
      RECT 34.655 3.264 34.741 3.434 ;
      RECT 34.63 3.26 34.655 3.433 ;
      RECT 34.62 3.257 34.63 3.431 ;
      RECT 34.61 3.25 34.62 3.428 ;
      RECT 34.605 3.23 34.61 3.423 ;
      RECT 34.595 3.2 34.605 3.418 ;
      RECT 34.58 3.07 34.595 3.409 ;
      RECT 34.575 3.062 34.58 3.402 ;
      RECT 34.555 3.055 34.575 3.394 ;
      RECT 34.55 3.037 34.555 3.386 ;
      RECT 34.54 3.017 34.55 3.381 ;
      RECT 34.535 2.99 34.54 3.377 ;
      RECT 34.53 2.967 34.535 3.374 ;
      RECT 34.51 2.925 34.53 3.366 ;
      RECT 34.475 2.84 34.51 3.35 ;
      RECT 34.47 2.772 34.475 3.338 ;
      RECT 34.455 2.742 34.47 3.332 ;
      RECT 34.45 1.987 34.455 2.233 ;
      RECT 34.44 2.712 34.455 3.323 ;
      RECT 34.445 1.982 34.45 2.265 ;
      RECT 34.44 1.977 34.445 2.308 ;
      RECT 34.435 1.975 34.44 2.343 ;
      RECT 34.42 2.675 34.44 3.313 ;
      RECT 34.43 1.975 34.435 2.38 ;
      RECT 34.415 1.975 34.43 2.478 ;
      RECT 34.415 2.648 34.42 3.306 ;
      RECT 34.41 1.975 34.415 2.553 ;
      RECT 34.41 2.636 34.415 3.303 ;
      RECT 34.405 1.975 34.41 2.585 ;
      RECT 34.405 2.615 34.41 3.3 ;
      RECT 34.4 1.975 34.405 3.297 ;
      RECT 34.365 1.975 34.4 3.283 ;
      RECT 34.35 1.975 34.365 3.265 ;
      RECT 34.33 1.975 34.35 3.255 ;
      RECT 34.305 1.975 34.33 3.238 ;
      RECT 34.3 1.975 34.305 3.188 ;
      RECT 34.29 1.975 34.295 3.018 ;
      RECT 34.285 1.975 34.29 2.925 ;
      RECT 34.28 1.975 34.285 2.838 ;
      RECT 34.275 1.975 34.28 2.77 ;
      RECT 34.27 1.975 34.275 2.713 ;
      RECT 34.26 1.975 34.27 2.608 ;
      RECT 34.255 1.975 34.26 2.48 ;
      RECT 34.25 1.975 34.255 2.398 ;
      RECT 34.245 1.977 34.25 2.315 ;
      RECT 34.24 1.982 34.245 2.248 ;
      RECT 34.235 1.987 34.24 2.175 ;
      RECT 37.05 2.305 37.31 2.565 ;
      RECT 37.07 2.272 37.28 2.565 ;
      RECT 37.07 2.27 37.27 2.565 ;
      RECT 37.08 2.257 37.27 2.565 ;
      RECT 37.08 2.255 37.195 2.565 ;
      RECT 36.555 2.38 36.73 2.66 ;
      RECT 36.55 2.38 36.73 2.658 ;
      RECT 36.55 2.38 36.745 2.655 ;
      RECT 36.54 2.38 36.745 2.653 ;
      RECT 36.485 2.38 36.745 2.64 ;
      RECT 36.485 2.455 36.75 2.618 ;
      RECT 36.03 2.392 36.05 2.635 ;
      RECT 36.03 2.392 36.09 2.634 ;
      RECT 36.025 2.394 36.09 2.633 ;
      RECT 36.025 2.394 36.176 2.632 ;
      RECT 36.025 2.394 36.245 2.631 ;
      RECT 36.025 2.394 36.265 2.623 ;
      RECT 36.005 2.397 36.265 2.621 ;
      RECT 35.99 2.407 36.265 2.606 ;
      RECT 35.99 2.407 36.28 2.605 ;
      RECT 35.985 2.416 36.28 2.597 ;
      RECT 35.985 2.416 36.285 2.593 ;
      RECT 36.09 2.33 36.35 2.59 ;
      RECT 35.98 2.418 36.35 2.475 ;
      RECT 36.05 2.385 36.35 2.59 ;
      RECT 36.015 3.578 36.02 3.785 ;
      RECT 35.965 3.572 36.015 3.784 ;
      RECT 35.932 3.586 36.025 3.783 ;
      RECT 35.846 3.586 36.025 3.782 ;
      RECT 35.76 3.586 36.025 3.781 ;
      RECT 35.76 3.685 36.03 3.778 ;
      RECT 35.755 3.685 36.03 3.773 ;
      RECT 35.75 3.685 36.03 3.755 ;
      RECT 35.745 3.685 36.03 3.738 ;
      RECT 35.705 3.47 35.965 3.73 ;
      RECT 35.165 2.62 35.251 3.034 ;
      RECT 35.165 2.62 35.29 3.031 ;
      RECT 35.165 2.62 35.31 3.021 ;
      RECT 35.12 2.62 35.31 3.018 ;
      RECT 35.12 2.772 35.32 3.008 ;
      RECT 35.12 2.793 35.325 3.002 ;
      RECT 35.12 2.811 35.33 2.998 ;
      RECT 35.12 2.831 35.34 2.993 ;
      RECT 35.095 2.831 35.34 2.99 ;
      RECT 35.085 2.831 35.34 2.968 ;
      RECT 35.085 2.847 35.345 2.938 ;
      RECT 35.05 2.62 35.31 2.925 ;
      RECT 35.05 2.859 35.35 2.88 ;
      RECT 32.71 7.77 33 8 ;
      RECT 32.77 6.29 32.94 8 ;
      RECT 32.76 6.66 33.115 7.015 ;
      RECT 32.71 6.29 33 6.52 ;
      RECT 32.305 2.395 32.41 2.965 ;
      RECT 32.305 2.73 32.63 2.96 ;
      RECT 32.305 2.76 32.8 2.93 ;
      RECT 32.305 2.395 32.495 2.96 ;
      RECT 31.72 2.36 32.01 2.59 ;
      RECT 31.72 2.395 32.495 2.565 ;
      RECT 31.78 0.88 31.95 2.59 ;
      RECT 31.72 0.88 32.01 1.11 ;
      RECT 31.72 7.77 32.01 8 ;
      RECT 31.78 6.29 31.95 8 ;
      RECT 31.72 6.29 32.01 6.52 ;
      RECT 31.72 6.325 32.575 6.485 ;
      RECT 32.405 5.92 32.575 6.485 ;
      RECT 31.72 6.32 32.115 6.485 ;
      RECT 32.34 5.92 32.63 6.15 ;
      RECT 32.34 5.95 32.8 6.12 ;
      RECT 31.35 2.73 31.64 2.96 ;
      RECT 31.35 2.76 31.81 2.93 ;
      RECT 31.415 1.655 31.58 2.96 ;
      RECT 29.93 1.625 30.22 1.855 ;
      RECT 29.93 1.655 31.58 1.825 ;
      RECT 29.99 0.885 30.16 1.855 ;
      RECT 29.93 0.885 30.22 1.115 ;
      RECT 29.93 7.765 30.22 7.995 ;
      RECT 29.99 7.025 30.16 7.995 ;
      RECT 29.99 7.12 31.58 7.29 ;
      RECT 31.41 5.92 31.58 7.29 ;
      RECT 29.93 7.025 30.22 7.255 ;
      RECT 31.35 5.92 31.64 6.15 ;
      RECT 31.35 5.95 31.81 6.12 ;
      RECT 27.98 2.705 28.32 3.055 ;
      RECT 28.07 2.025 28.24 3.055 ;
      RECT 30.36 1.965 30.71 2.315 ;
      RECT 28.07 2.025 30.71 2.195 ;
      RECT 30.385 6.655 30.71 6.98 ;
      RECT 24.925 6.61 25.275 6.96 ;
      RECT 30.36 6.655 30.71 6.885 ;
      RECT 24.725 6.655 25.275 6.885 ;
      RECT 24.555 6.685 30.71 6.855 ;
      RECT 29.585 2.365 29.905 2.685 ;
      RECT 29.555 2.365 29.905 2.595 ;
      RECT 29.385 2.395 29.905 2.565 ;
      RECT 29.585 6.255 29.905 6.545 ;
      RECT 29.555 6.285 29.905 6.515 ;
      RECT 29.385 6.315 29.905 6.485 ;
      RECT 25.275 2.985 25.425 3.26 ;
      RECT 25.815 2.065 25.82 2.285 ;
      RECT 26.965 2.265 26.98 2.463 ;
      RECT 26.93 2.257 26.965 2.47 ;
      RECT 26.9 2.25 26.93 2.47 ;
      RECT 26.845 2.215 26.9 2.47 ;
      RECT 26.78 2.152 26.845 2.47 ;
      RECT 26.775 2.117 26.78 2.468 ;
      RECT 26.77 2.112 26.775 2.46 ;
      RECT 26.765 2.107 26.77 2.446 ;
      RECT 26.76 2.104 26.765 2.439 ;
      RECT 26.715 2.094 26.76 2.39 ;
      RECT 26.695 2.081 26.715 2.325 ;
      RECT 26.69 2.076 26.695 2.298 ;
      RECT 26.685 2.075 26.69 2.291 ;
      RECT 26.68 2.074 26.685 2.284 ;
      RECT 26.595 2.059 26.68 2.23 ;
      RECT 26.565 2.04 26.595 2.18 ;
      RECT 26.485 2.023 26.565 2.165 ;
      RECT 26.45 2.01 26.485 2.15 ;
      RECT 26.442 2.01 26.45 2.145 ;
      RECT 26.356 2.011 26.442 2.145 ;
      RECT 26.27 2.013 26.356 2.145 ;
      RECT 26.245 2.014 26.27 2.149 ;
      RECT 26.17 2.02 26.245 2.164 ;
      RECT 26.087 2.032 26.17 2.188 ;
      RECT 26.001 2.045 26.087 2.214 ;
      RECT 25.915 2.058 26.001 2.24 ;
      RECT 25.88 2.067 25.915 2.259 ;
      RECT 25.83 2.067 25.88 2.272 ;
      RECT 25.82 2.065 25.83 2.283 ;
      RECT 25.805 2.062 25.815 2.285 ;
      RECT 25.79 2.054 25.805 2.293 ;
      RECT 25.775 2.046 25.79 2.313 ;
      RECT 25.77 2.041 25.775 2.37 ;
      RECT 25.755 2.036 25.77 2.443 ;
      RECT 25.75 2.031 25.755 2.485 ;
      RECT 25.745 2.029 25.75 2.513 ;
      RECT 25.74 2.027 25.745 2.535 ;
      RECT 25.73 2.023 25.74 2.578 ;
      RECT 25.725 2.02 25.73 2.603 ;
      RECT 25.72 2.018 25.725 2.623 ;
      RECT 25.715 2.016 25.72 2.647 ;
      RECT 25.71 2.012 25.715 2.67 ;
      RECT 25.705 2.008 25.71 2.693 ;
      RECT 25.67 1.998 25.705 2.8 ;
      RECT 25.665 1.988 25.67 2.898 ;
      RECT 25.66 1.986 25.665 2.925 ;
      RECT 25.655 1.985 25.66 2.945 ;
      RECT 25.65 1.977 25.655 2.965 ;
      RECT 25.645 1.972 25.65 3 ;
      RECT 25.64 1.97 25.645 3.018 ;
      RECT 25.635 1.97 25.64 3.043 ;
      RECT 25.63 1.97 25.635 3.065 ;
      RECT 25.595 1.97 25.63 3.108 ;
      RECT 25.57 1.97 25.595 3.137 ;
      RECT 25.56 1.97 25.57 2.323 ;
      RECT 25.563 2.38 25.57 3.147 ;
      RECT 25.56 2.437 25.563 3.15 ;
      RECT 25.555 1.97 25.56 2.295 ;
      RECT 25.555 2.487 25.56 3.153 ;
      RECT 25.545 1.97 25.555 2.285 ;
      RECT 25.55 2.54 25.555 3.156 ;
      RECT 25.545 2.625 25.55 3.16 ;
      RECT 25.535 1.97 25.545 2.273 ;
      RECT 25.54 2.672 25.545 3.164 ;
      RECT 25.535 2.747 25.54 3.168 ;
      RECT 25.5 1.97 25.535 2.248 ;
      RECT 25.525 2.83 25.535 3.173 ;
      RECT 25.515 2.897 25.525 3.18 ;
      RECT 25.51 2.925 25.515 3.185 ;
      RECT 25.5 2.938 25.51 3.191 ;
      RECT 25.455 1.97 25.5 2.205 ;
      RECT 25.495 2.943 25.5 3.198 ;
      RECT 25.455 2.96 25.495 3.26 ;
      RECT 25.45 1.972 25.455 2.178 ;
      RECT 25.425 2.98 25.455 3.26 ;
      RECT 25.445 1.977 25.45 2.15 ;
      RECT 25.235 2.989 25.275 3.26 ;
      RECT 25.21 2.997 25.235 3.23 ;
      RECT 25.165 3.005 25.21 3.23 ;
      RECT 25.15 3.01 25.165 3.225 ;
      RECT 25.14 3.01 25.15 3.219 ;
      RECT 25.13 3.017 25.14 3.216 ;
      RECT 25.125 3.055 25.13 3.205 ;
      RECT 25.12 3.117 25.125 3.183 ;
      RECT 26.39 2.992 26.575 3.215 ;
      RECT 26.39 3.007 26.58 3.211 ;
      RECT 26.38 2.28 26.465 3.21 ;
      RECT 26.38 3.007 26.585 3.204 ;
      RECT 26.375 3.015 26.585 3.203 ;
      RECT 26.58 2.735 26.9 3.055 ;
      RECT 26.375 2.907 26.545 2.998 ;
      RECT 26.37 2.907 26.545 2.98 ;
      RECT 26.36 2.715 26.495 2.955 ;
      RECT 26.355 2.715 26.495 2.9 ;
      RECT 26.315 2.295 26.485 2.8 ;
      RECT 26.3 2.295 26.485 2.67 ;
      RECT 26.295 2.295 26.485 2.623 ;
      RECT 26.29 2.295 26.485 2.603 ;
      RECT 26.285 2.295 26.485 2.578 ;
      RECT 26.255 2.295 26.515 2.555 ;
      RECT 26.265 2.292 26.475 2.555 ;
      RECT 26.39 2.287 26.475 3.215 ;
      RECT 26.275 2.28 26.465 2.555 ;
      RECT 26.27 2.285 26.465 2.555 ;
      RECT 25.1 2.497 25.285 2.71 ;
      RECT 25.1 2.505 25.295 2.703 ;
      RECT 25.08 2.505 25.295 2.7 ;
      RECT 25.075 2.505 25.295 2.685 ;
      RECT 25.005 2.42 25.265 2.68 ;
      RECT 25.005 2.565 25.3 2.593 ;
      RECT 24.66 3.02 24.92 3.28 ;
      RECT 24.685 2.965 24.88 3.28 ;
      RECT 24.68 2.714 24.86 3.008 ;
      RECT 24.68 2.72 24.87 3.008 ;
      RECT 24.66 2.722 24.87 2.953 ;
      RECT 24.655 2.732 24.87 2.82 ;
      RECT 24.685 2.712 24.86 3.28 ;
      RECT 24.771 2.71 24.86 3.28 ;
      RECT 24.63 1.93 24.665 2.3 ;
      RECT 24.42 2.04 24.425 2.3 ;
      RECT 24.665 1.937 24.68 2.3 ;
      RECT 24.555 1.93 24.63 2.378 ;
      RECT 24.545 1.93 24.555 2.463 ;
      RECT 24.52 1.93 24.545 2.498 ;
      RECT 24.48 1.93 24.52 2.566 ;
      RECT 24.47 1.937 24.48 2.618 ;
      RECT 24.44 2.04 24.47 2.659 ;
      RECT 24.435 2.04 24.44 2.698 ;
      RECT 24.425 2.04 24.435 2.718 ;
      RECT 24.42 2.335 24.425 2.755 ;
      RECT 24.415 2.352 24.42 2.775 ;
      RECT 24.4 2.415 24.415 2.815 ;
      RECT 24.395 2.458 24.4 2.85 ;
      RECT 24.39 2.466 24.395 2.863 ;
      RECT 24.38 2.48 24.39 2.885 ;
      RECT 24.355 2.515 24.38 2.95 ;
      RECT 24.345 2.55 24.355 3.013 ;
      RECT 24.325 2.58 24.345 3.074 ;
      RECT 24.31 2.616 24.325 3.141 ;
      RECT 24.3 2.644 24.31 3.18 ;
      RECT 24.29 2.666 24.3 3.2 ;
      RECT 24.285 2.676 24.29 3.211 ;
      RECT 24.28 2.685 24.285 3.214 ;
      RECT 24.27 2.703 24.28 3.218 ;
      RECT 24.26 2.721 24.27 3.219 ;
      RECT 24.235 2.76 24.26 3.216 ;
      RECT 24.215 2.802 24.235 3.213 ;
      RECT 24.2 2.84 24.215 3.212 ;
      RECT 24.165 2.875 24.2 3.209 ;
      RECT 24.16 2.897 24.165 3.207 ;
      RECT 24.095 2.937 24.16 3.204 ;
      RECT 24.09 2.977 24.095 3.2 ;
      RECT 24.075 2.987 24.09 3.191 ;
      RECT 24.065 3.107 24.075 3.176 ;
      RECT 24.545 3.52 24.555 3.78 ;
      RECT 24.545 3.523 24.565 3.779 ;
      RECT 24.535 3.513 24.545 3.778 ;
      RECT 24.525 3.528 24.605 3.774 ;
      RECT 24.51 3.507 24.525 3.772 ;
      RECT 24.485 3.532 24.61 3.768 ;
      RECT 24.47 3.492 24.485 3.763 ;
      RECT 24.47 3.534 24.62 3.762 ;
      RECT 24.47 3.542 24.635 3.755 ;
      RECT 24.41 3.479 24.47 3.745 ;
      RECT 24.4 3.466 24.41 3.727 ;
      RECT 24.375 3.456 24.4 3.717 ;
      RECT 24.37 3.446 24.375 3.709 ;
      RECT 24.305 3.542 24.635 3.691 ;
      RECT 24.22 3.542 24.635 3.653 ;
      RECT 24.11 3.37 24.37 3.63 ;
      RECT 24.485 3.5 24.51 3.768 ;
      RECT 24.525 3.51 24.535 3.774 ;
      RECT 24.11 3.518 24.55 3.63 ;
      RECT 24.295 7.765 24.585 7.995 ;
      RECT 24.355 7.025 24.525 7.995 ;
      RECT 24.255 7.055 24.625 7.425 ;
      RECT 24.295 7.025 24.585 7.425 ;
      RECT 23.325 3.275 23.355 3.575 ;
      RECT 23.1 3.26 23.105 3.535 ;
      RECT 22.9 3.26 23.055 3.52 ;
      RECT 24.2 1.975 24.23 2.235 ;
      RECT 24.19 1.975 24.2 2.343 ;
      RECT 24.17 1.975 24.19 2.353 ;
      RECT 24.155 1.975 24.17 2.365 ;
      RECT 24.1 1.975 24.155 2.415 ;
      RECT 24.085 1.975 24.1 2.463 ;
      RECT 24.055 1.975 24.085 2.498 ;
      RECT 24 1.975 24.055 2.56 ;
      RECT 23.98 1.975 24 2.628 ;
      RECT 23.975 1.975 23.98 2.658 ;
      RECT 23.97 1.975 23.975 2.67 ;
      RECT 23.965 2.092 23.97 2.688 ;
      RECT 23.945 2.11 23.965 2.713 ;
      RECT 23.925 2.137 23.945 2.763 ;
      RECT 23.92 2.157 23.925 2.794 ;
      RECT 23.915 2.165 23.92 2.811 ;
      RECT 23.9 2.191 23.915 2.84 ;
      RECT 23.885 2.233 23.9 2.875 ;
      RECT 23.88 2.262 23.885 2.898 ;
      RECT 23.875 2.277 23.88 2.911 ;
      RECT 23.87 2.3 23.875 2.922 ;
      RECT 23.86 2.32 23.87 2.94 ;
      RECT 23.85 2.35 23.86 2.963 ;
      RECT 23.845 2.372 23.85 2.983 ;
      RECT 23.84 2.387 23.845 2.998 ;
      RECT 23.825 2.417 23.84 3.025 ;
      RECT 23.82 2.447 23.825 3.051 ;
      RECT 23.815 2.465 23.82 3.063 ;
      RECT 23.805 2.495 23.815 3.082 ;
      RECT 23.795 2.52 23.805 3.107 ;
      RECT 23.79 2.54 23.795 3.126 ;
      RECT 23.785 2.557 23.79 3.139 ;
      RECT 23.775 2.583 23.785 3.158 ;
      RECT 23.765 2.621 23.775 3.185 ;
      RECT 23.76 2.647 23.765 3.205 ;
      RECT 23.755 2.657 23.76 3.215 ;
      RECT 23.75 2.67 23.755 3.23 ;
      RECT 23.745 2.685 23.75 3.24 ;
      RECT 23.74 2.707 23.745 3.255 ;
      RECT 23.735 2.725 23.74 3.266 ;
      RECT 23.73 2.735 23.735 3.277 ;
      RECT 23.725 2.743 23.73 3.289 ;
      RECT 23.72 2.751 23.725 3.3 ;
      RECT 23.715 2.777 23.72 3.313 ;
      RECT 23.705 2.805 23.715 3.326 ;
      RECT 23.7 2.835 23.705 3.335 ;
      RECT 23.695 2.85 23.7 3.342 ;
      RECT 23.68 2.875 23.695 3.349 ;
      RECT 23.675 2.897 23.68 3.355 ;
      RECT 23.67 2.922 23.675 3.358 ;
      RECT 23.661 2.95 23.67 3.362 ;
      RECT 23.655 2.967 23.661 3.367 ;
      RECT 23.65 2.985 23.655 3.371 ;
      RECT 23.645 2.997 23.65 3.374 ;
      RECT 23.64 3.018 23.645 3.378 ;
      RECT 23.635 3.036 23.64 3.381 ;
      RECT 23.63 3.05 23.635 3.384 ;
      RECT 23.625 3.067 23.63 3.387 ;
      RECT 23.62 3.08 23.625 3.39 ;
      RECT 23.595 3.117 23.62 3.398 ;
      RECT 23.59 3.162 23.595 3.407 ;
      RECT 23.585 3.19 23.59 3.41 ;
      RECT 23.575 3.21 23.585 3.414 ;
      RECT 23.57 3.23 23.575 3.419 ;
      RECT 23.565 3.245 23.57 3.422 ;
      RECT 23.545 3.255 23.565 3.429 ;
      RECT 23.48 3.262 23.545 3.455 ;
      RECT 23.445 3.265 23.48 3.483 ;
      RECT 23.43 3.268 23.445 3.498 ;
      RECT 23.42 3.269 23.43 3.513 ;
      RECT 23.41 3.27 23.42 3.53 ;
      RECT 23.405 3.27 23.41 3.545 ;
      RECT 23.4 3.27 23.405 3.553 ;
      RECT 23.385 3.271 23.4 3.568 ;
      RECT 23.355 3.273 23.385 3.575 ;
      RECT 23.245 3.28 23.325 3.575 ;
      RECT 23.2 3.285 23.245 3.575 ;
      RECT 23.19 3.286 23.2 3.565 ;
      RECT 23.18 3.287 23.19 3.558 ;
      RECT 23.16 3.289 23.18 3.553 ;
      RECT 23.15 3.26 23.16 3.548 ;
      RECT 23.105 3.26 23.15 3.54 ;
      RECT 23.075 3.26 23.1 3.53 ;
      RECT 23.055 3.26 23.075 3.523 ;
      RECT 23.335 2.06 23.595 2.32 ;
      RECT 23.215 2.075 23.225 2.24 ;
      RECT 23.2 2.075 23.205 2.235 ;
      RECT 20.565 1.915 20.75 2.205 ;
      RECT 22.38 2.04 22.395 2.195 ;
      RECT 20.53 1.915 20.555 2.175 ;
      RECT 22.945 1.965 22.95 2.107 ;
      RECT 22.86 1.96 22.885 2.1 ;
      RECT 23.26 2.077 23.335 2.27 ;
      RECT 23.245 2.075 23.26 2.253 ;
      RECT 23.225 2.075 23.245 2.245 ;
      RECT 23.205 2.075 23.215 2.238 ;
      RECT 23.16 2.07 23.2 2.228 ;
      RECT 23.12 2.045 23.16 2.213 ;
      RECT 23.105 2.02 23.12 2.203 ;
      RECT 23.1 2.014 23.105 2.201 ;
      RECT 23.065 2.006 23.1 2.184 ;
      RECT 23.06 1.999 23.065 2.172 ;
      RECT 23.04 1.994 23.06 2.16 ;
      RECT 23.03 1.988 23.04 2.145 ;
      RECT 23.01 1.983 23.03 2.13 ;
      RECT 23 1.978 23.01 2.123 ;
      RECT 22.995 1.976 23 2.118 ;
      RECT 22.99 1.975 22.995 2.115 ;
      RECT 22.95 1.97 22.99 2.111 ;
      RECT 22.93 1.964 22.945 2.106 ;
      RECT 22.895 1.961 22.93 2.103 ;
      RECT 22.885 1.96 22.895 2.101 ;
      RECT 22.825 1.96 22.86 2.098 ;
      RECT 22.78 1.96 22.825 2.098 ;
      RECT 22.73 1.96 22.78 2.101 ;
      RECT 22.715 1.962 22.73 2.103 ;
      RECT 22.7 1.965 22.715 2.104 ;
      RECT 22.69 1.97 22.7 2.105 ;
      RECT 22.66 1.975 22.69 2.11 ;
      RECT 22.65 1.981 22.66 2.118 ;
      RECT 22.64 1.983 22.65 2.122 ;
      RECT 22.63 1.987 22.64 2.126 ;
      RECT 22.605 1.993 22.63 2.134 ;
      RECT 22.595 1.998 22.605 2.142 ;
      RECT 22.58 2.002 22.595 2.146 ;
      RECT 22.545 2.008 22.58 2.154 ;
      RECT 22.525 2.013 22.545 2.164 ;
      RECT 22.495 2.02 22.525 2.173 ;
      RECT 22.45 2.029 22.495 2.187 ;
      RECT 22.445 2.034 22.45 2.198 ;
      RECT 22.425 2.037 22.445 2.199 ;
      RECT 22.395 2.04 22.425 2.197 ;
      RECT 22.36 2.04 22.38 2.193 ;
      RECT 22.29 2.04 22.36 2.184 ;
      RECT 22.275 2.037 22.29 2.176 ;
      RECT 22.235 2.03 22.275 2.171 ;
      RECT 22.21 2.02 22.235 2.164 ;
      RECT 22.205 2.014 22.21 2.161 ;
      RECT 22.165 2.008 22.205 2.158 ;
      RECT 22.15 2.001 22.165 2.153 ;
      RECT 22.13 1.997 22.15 2.148 ;
      RECT 22.115 1.992 22.13 2.144 ;
      RECT 22.1 1.987 22.115 2.142 ;
      RECT 22.085 1.983 22.1 2.141 ;
      RECT 22.07 1.981 22.085 2.137 ;
      RECT 22.06 1.979 22.07 2.132 ;
      RECT 22.045 1.976 22.06 2.128 ;
      RECT 22.035 1.974 22.045 2.123 ;
      RECT 22.015 1.971 22.035 2.119 ;
      RECT 21.97 1.97 22.015 2.117 ;
      RECT 21.91 1.972 21.97 2.118 ;
      RECT 21.89 1.974 21.91 2.12 ;
      RECT 21.86 1.977 21.89 2.121 ;
      RECT 21.81 1.982 21.86 2.123 ;
      RECT 21.805 1.985 21.81 2.125 ;
      RECT 21.795 1.987 21.805 2.128 ;
      RECT 21.79 1.989 21.795 2.131 ;
      RECT 21.74 1.992 21.79 2.138 ;
      RECT 21.72 1.996 21.74 2.15 ;
      RECT 21.71 1.999 21.72 2.156 ;
      RECT 21.7 2 21.71 2.159 ;
      RECT 21.661 2.003 21.7 2.161 ;
      RECT 21.575 2.01 21.661 2.164 ;
      RECT 21.501 2.02 21.575 2.168 ;
      RECT 21.415 2.031 21.501 2.173 ;
      RECT 21.4 2.038 21.415 2.175 ;
      RECT 21.345 2.042 21.4 2.176 ;
      RECT 21.331 2.045 21.345 2.178 ;
      RECT 21.245 2.045 21.331 2.18 ;
      RECT 21.205 2.042 21.245 2.183 ;
      RECT 21.181 2.038 21.205 2.185 ;
      RECT 21.095 2.028 21.181 2.188 ;
      RECT 21.065 2.017 21.095 2.189 ;
      RECT 21.046 2.013 21.065 2.188 ;
      RECT 20.96 2.006 21.046 2.185 ;
      RECT 20.9 1.995 20.96 2.182 ;
      RECT 20.88 1.987 20.9 2.18 ;
      RECT 20.845 1.982 20.88 2.179 ;
      RECT 20.82 1.977 20.845 2.178 ;
      RECT 20.79 1.972 20.82 2.177 ;
      RECT 20.765 1.915 20.79 2.176 ;
      RECT 20.75 1.915 20.765 2.2 ;
      RECT 20.555 1.915 20.565 2.2 ;
      RECT 22.33 2.935 22.335 3.075 ;
      RECT 21.99 2.935 22.025 3.073 ;
      RECT 21.565 2.92 21.58 3.065 ;
      RECT 23.395 2.7 23.485 2.96 ;
      RECT 23.225 2.565 23.325 2.96 ;
      RECT 20.26 2.54 20.34 2.75 ;
      RECT 23.35 2.677 23.395 2.96 ;
      RECT 23.34 2.647 23.35 2.96 ;
      RECT 23.325 2.57 23.34 2.96 ;
      RECT 23.14 2.565 23.225 2.925 ;
      RECT 23.135 2.567 23.14 2.92 ;
      RECT 23.13 2.572 23.135 2.92 ;
      RECT 23.095 2.672 23.13 2.92 ;
      RECT 23.085 2.7 23.095 2.92 ;
      RECT 23.075 2.715 23.085 2.92 ;
      RECT 23.065 2.727 23.075 2.92 ;
      RECT 23.06 2.737 23.065 2.92 ;
      RECT 23.045 2.747 23.06 2.922 ;
      RECT 23.04 2.762 23.045 2.924 ;
      RECT 23.025 2.775 23.04 2.926 ;
      RECT 23.02 2.79 23.025 2.929 ;
      RECT 23 2.8 23.02 2.933 ;
      RECT 22.985 2.81 23 2.936 ;
      RECT 22.95 2.817 22.985 2.941 ;
      RECT 22.906 2.824 22.95 2.949 ;
      RECT 22.82 2.836 22.906 2.962 ;
      RECT 22.795 2.847 22.82 2.973 ;
      RECT 22.765 2.852 22.795 2.978 ;
      RECT 22.73 2.857 22.765 2.986 ;
      RECT 22.7 2.862 22.73 2.993 ;
      RECT 22.675 2.867 22.7 2.998 ;
      RECT 22.61 2.874 22.675 3.007 ;
      RECT 22.54 2.887 22.61 3.023 ;
      RECT 22.51 2.897 22.54 3.035 ;
      RECT 22.485 2.902 22.51 3.042 ;
      RECT 22.43 2.909 22.485 3.05 ;
      RECT 22.425 2.916 22.43 3.055 ;
      RECT 22.42 2.918 22.425 3.056 ;
      RECT 22.405 2.92 22.42 3.058 ;
      RECT 22.4 2.92 22.405 3.061 ;
      RECT 22.335 2.927 22.4 3.068 ;
      RECT 22.3 2.937 22.33 3.078 ;
      RECT 22.283 2.94 22.3 3.08 ;
      RECT 22.197 2.939 22.283 3.079 ;
      RECT 22.111 2.937 22.197 3.076 ;
      RECT 22.025 2.936 22.111 3.074 ;
      RECT 21.924 2.934 21.99 3.073 ;
      RECT 21.838 2.931 21.924 3.071 ;
      RECT 21.752 2.927 21.838 3.069 ;
      RECT 21.666 2.924 21.752 3.068 ;
      RECT 21.58 2.921 21.666 3.066 ;
      RECT 21.48 2.92 21.565 3.063 ;
      RECT 21.43 2.918 21.48 3.061 ;
      RECT 21.41 2.915 21.43 3.059 ;
      RECT 21.39 2.913 21.41 3.056 ;
      RECT 21.365 2.909 21.39 3.053 ;
      RECT 21.32 2.903 21.365 3.048 ;
      RECT 21.28 2.897 21.32 3.04 ;
      RECT 21.255 2.892 21.28 3.033 ;
      RECT 21.2 2.885 21.255 3.025 ;
      RECT 21.176 2.878 21.2 3.018 ;
      RECT 21.09 2.869 21.176 3.008 ;
      RECT 21.06 2.861 21.09 2.998 ;
      RECT 21.03 2.857 21.06 2.993 ;
      RECT 21.025 2.854 21.03 2.99 ;
      RECT 21.02 2.853 21.025 2.99 ;
      RECT 20.945 2.846 21.02 2.983 ;
      RECT 20.906 2.837 20.945 2.972 ;
      RECT 20.82 2.827 20.906 2.96 ;
      RECT 20.78 2.817 20.82 2.948 ;
      RECT 20.741 2.812 20.78 2.941 ;
      RECT 20.655 2.802 20.741 2.93 ;
      RECT 20.615 2.79 20.655 2.919 ;
      RECT 20.58 2.775 20.615 2.912 ;
      RECT 20.57 2.765 20.58 2.909 ;
      RECT 20.55 2.75 20.57 2.907 ;
      RECT 20.52 2.72 20.55 2.903 ;
      RECT 20.51 2.7 20.52 2.898 ;
      RECT 20.505 2.692 20.51 2.895 ;
      RECT 20.5 2.685 20.505 2.893 ;
      RECT 20.485 2.672 20.5 2.886 ;
      RECT 20.48 2.662 20.485 2.878 ;
      RECT 20.475 2.655 20.48 2.873 ;
      RECT 20.47 2.65 20.475 2.869 ;
      RECT 20.455 2.637 20.47 2.861 ;
      RECT 20.45 2.547 20.455 2.85 ;
      RECT 20.445 2.542 20.45 2.843 ;
      RECT 20.37 2.54 20.445 2.803 ;
      RECT 20.34 2.54 20.37 2.758 ;
      RECT 20.245 2.545 20.26 2.745 ;
      RECT 22.73 2.25 22.99 2.51 ;
      RECT 22.715 2.238 22.895 2.475 ;
      RECT 22.71 2.239 22.895 2.473 ;
      RECT 22.695 2.243 22.905 2.463 ;
      RECT 22.69 2.248 22.91 2.433 ;
      RECT 22.695 2.245 22.91 2.463 ;
      RECT 22.71 2.24 22.905 2.473 ;
      RECT 22.73 2.237 22.895 2.51 ;
      RECT 22.73 2.236 22.885 2.51 ;
      RECT 22.755 2.235 22.885 2.51 ;
      RECT 22.315 2.48 22.575 2.74 ;
      RECT 22.19 2.525 22.575 2.735 ;
      RECT 22.18 2.53 22.575 2.73 ;
      RECT 22.195 3.47 22.21 3.78 ;
      RECT 20.79 3.24 20.8 3.37 ;
      RECT 20.57 3.235 20.675 3.37 ;
      RECT 20.485 3.24 20.535 3.37 ;
      RECT 19.035 1.975 19.04 3.08 ;
      RECT 22.29 3.562 22.295 3.698 ;
      RECT 22.285 3.557 22.29 3.758 ;
      RECT 22.28 3.555 22.285 3.771 ;
      RECT 22.265 3.552 22.28 3.773 ;
      RECT 22.26 3.547 22.265 3.775 ;
      RECT 22.255 3.543 22.26 3.778 ;
      RECT 22.24 3.538 22.255 3.78 ;
      RECT 22.21 3.53 22.24 3.78 ;
      RECT 22.171 3.47 22.195 3.78 ;
      RECT 22.085 3.47 22.171 3.777 ;
      RECT 22.055 3.47 22.085 3.77 ;
      RECT 22.03 3.47 22.055 3.763 ;
      RECT 22.005 3.47 22.03 3.755 ;
      RECT 21.99 3.47 22.005 3.748 ;
      RECT 21.965 3.47 21.99 3.74 ;
      RECT 21.95 3.47 21.965 3.733 ;
      RECT 21.91 3.48 21.95 3.722 ;
      RECT 21.9 3.475 21.91 3.712 ;
      RECT 21.896 3.474 21.9 3.709 ;
      RECT 21.81 3.466 21.896 3.692 ;
      RECT 21.777 3.455 21.81 3.669 ;
      RECT 21.691 3.444 21.777 3.647 ;
      RECT 21.605 3.428 21.691 3.616 ;
      RECT 21.535 3.413 21.605 3.588 ;
      RECT 21.525 3.406 21.535 3.575 ;
      RECT 21.495 3.403 21.525 3.565 ;
      RECT 21.47 3.399 21.495 3.558 ;
      RECT 21.455 3.396 21.47 3.553 ;
      RECT 21.45 3.395 21.455 3.548 ;
      RECT 21.42 3.39 21.45 3.541 ;
      RECT 21.415 3.385 21.42 3.536 ;
      RECT 21.4 3.382 21.415 3.531 ;
      RECT 21.395 3.377 21.4 3.526 ;
      RECT 21.375 3.372 21.395 3.523 ;
      RECT 21.36 3.367 21.375 3.515 ;
      RECT 21.345 3.361 21.36 3.51 ;
      RECT 21.315 3.352 21.345 3.503 ;
      RECT 21.31 3.345 21.315 3.495 ;
      RECT 21.305 3.343 21.31 3.493 ;
      RECT 21.3 3.342 21.305 3.49 ;
      RECT 21.26 3.335 21.3 3.483 ;
      RECT 21.246 3.325 21.26 3.473 ;
      RECT 21.195 3.314 21.246 3.461 ;
      RECT 21.17 3.3 21.195 3.447 ;
      RECT 21.145 3.289 21.17 3.439 ;
      RECT 21.125 3.278 21.145 3.433 ;
      RECT 21.115 3.272 21.125 3.428 ;
      RECT 21.11 3.27 21.115 3.424 ;
      RECT 21.09 3.265 21.11 3.419 ;
      RECT 21.06 3.255 21.09 3.409 ;
      RECT 21.055 3.247 21.06 3.402 ;
      RECT 21.04 3.245 21.055 3.398 ;
      RECT 21.02 3.245 21.04 3.393 ;
      RECT 21.015 3.244 21.02 3.391 ;
      RECT 21.01 3.244 21.015 3.388 ;
      RECT 20.97 3.243 21.01 3.383 ;
      RECT 20.945 3.242 20.97 3.378 ;
      RECT 20.885 3.241 20.945 3.375 ;
      RECT 20.8 3.24 20.885 3.373 ;
      RECT 20.761 3.239 20.79 3.37 ;
      RECT 20.675 3.237 20.761 3.37 ;
      RECT 20.535 3.237 20.57 3.37 ;
      RECT 20.445 3.241 20.485 3.373 ;
      RECT 20.43 3.244 20.445 3.38 ;
      RECT 20.42 3.245 20.43 3.387 ;
      RECT 20.395 3.248 20.42 3.392 ;
      RECT 20.39 3.25 20.395 3.395 ;
      RECT 20.34 3.252 20.39 3.396 ;
      RECT 20.301 3.256 20.34 3.398 ;
      RECT 20.215 3.258 20.301 3.401 ;
      RECT 20.197 3.26 20.215 3.403 ;
      RECT 20.111 3.263 20.197 3.405 ;
      RECT 20.025 3.267 20.111 3.408 ;
      RECT 19.988 3.271 20.025 3.411 ;
      RECT 19.902 3.274 19.988 3.414 ;
      RECT 19.816 3.278 19.902 3.417 ;
      RECT 19.73 3.283 19.816 3.421 ;
      RECT 19.71 3.285 19.73 3.424 ;
      RECT 19.69 3.284 19.71 3.425 ;
      RECT 19.641 3.281 19.69 3.426 ;
      RECT 19.555 3.276 19.641 3.429 ;
      RECT 19.505 3.271 19.555 3.431 ;
      RECT 19.481 3.269 19.505 3.432 ;
      RECT 19.395 3.264 19.481 3.434 ;
      RECT 19.37 3.26 19.395 3.433 ;
      RECT 19.36 3.257 19.37 3.431 ;
      RECT 19.35 3.25 19.36 3.428 ;
      RECT 19.345 3.23 19.35 3.423 ;
      RECT 19.335 3.2 19.345 3.418 ;
      RECT 19.32 3.07 19.335 3.409 ;
      RECT 19.315 3.062 19.32 3.402 ;
      RECT 19.295 3.055 19.315 3.394 ;
      RECT 19.29 3.037 19.295 3.386 ;
      RECT 19.28 3.017 19.29 3.381 ;
      RECT 19.275 2.99 19.28 3.377 ;
      RECT 19.27 2.967 19.275 3.374 ;
      RECT 19.25 2.925 19.27 3.366 ;
      RECT 19.215 2.84 19.25 3.35 ;
      RECT 19.21 2.772 19.215 3.338 ;
      RECT 19.195 2.742 19.21 3.332 ;
      RECT 19.19 1.987 19.195 2.233 ;
      RECT 19.18 2.712 19.195 3.323 ;
      RECT 19.185 1.982 19.19 2.265 ;
      RECT 19.18 1.977 19.185 2.308 ;
      RECT 19.175 1.975 19.18 2.343 ;
      RECT 19.16 2.675 19.18 3.313 ;
      RECT 19.17 1.975 19.175 2.38 ;
      RECT 19.155 1.975 19.17 2.478 ;
      RECT 19.155 2.648 19.16 3.306 ;
      RECT 19.15 1.975 19.155 2.553 ;
      RECT 19.15 2.636 19.155 3.303 ;
      RECT 19.145 1.975 19.15 2.585 ;
      RECT 19.145 2.615 19.15 3.3 ;
      RECT 19.14 1.975 19.145 3.297 ;
      RECT 19.105 1.975 19.14 3.283 ;
      RECT 19.09 1.975 19.105 3.265 ;
      RECT 19.07 1.975 19.09 3.255 ;
      RECT 19.045 1.975 19.07 3.238 ;
      RECT 19.04 1.975 19.045 3.188 ;
      RECT 19.03 1.975 19.035 3.018 ;
      RECT 19.025 1.975 19.03 2.925 ;
      RECT 19.02 1.975 19.025 2.838 ;
      RECT 19.015 1.975 19.02 2.77 ;
      RECT 19.01 1.975 19.015 2.713 ;
      RECT 19 1.975 19.01 2.608 ;
      RECT 18.995 1.975 19 2.48 ;
      RECT 18.99 1.975 18.995 2.398 ;
      RECT 18.985 1.977 18.99 2.315 ;
      RECT 18.98 1.982 18.985 2.248 ;
      RECT 18.975 1.987 18.98 2.175 ;
      RECT 21.79 2.305 22.05 2.565 ;
      RECT 21.81 2.272 22.02 2.565 ;
      RECT 21.81 2.27 22.01 2.565 ;
      RECT 21.82 2.257 22.01 2.565 ;
      RECT 21.82 2.255 21.935 2.565 ;
      RECT 21.295 2.38 21.47 2.66 ;
      RECT 21.29 2.38 21.47 2.658 ;
      RECT 21.29 2.38 21.485 2.655 ;
      RECT 21.28 2.38 21.485 2.653 ;
      RECT 21.225 2.38 21.485 2.64 ;
      RECT 21.225 2.455 21.49 2.618 ;
      RECT 20.77 2.392 20.79 2.635 ;
      RECT 20.77 2.392 20.83 2.634 ;
      RECT 20.765 2.394 20.83 2.633 ;
      RECT 20.765 2.394 20.916 2.632 ;
      RECT 20.765 2.394 20.985 2.631 ;
      RECT 20.765 2.394 21.005 2.623 ;
      RECT 20.745 2.397 21.005 2.621 ;
      RECT 20.73 2.407 21.005 2.606 ;
      RECT 20.73 2.407 21.02 2.605 ;
      RECT 20.725 2.416 21.02 2.597 ;
      RECT 20.725 2.416 21.025 2.593 ;
      RECT 20.83 2.33 21.09 2.59 ;
      RECT 20.72 2.418 21.09 2.475 ;
      RECT 20.79 2.385 21.09 2.59 ;
      RECT 20.755 3.578 20.76 3.785 ;
      RECT 20.705 3.572 20.755 3.784 ;
      RECT 20.672 3.586 20.765 3.783 ;
      RECT 20.586 3.586 20.765 3.782 ;
      RECT 20.5 3.586 20.765 3.781 ;
      RECT 20.5 3.685 20.77 3.778 ;
      RECT 20.495 3.685 20.77 3.773 ;
      RECT 20.49 3.685 20.77 3.755 ;
      RECT 20.485 3.685 20.77 3.738 ;
      RECT 20.445 3.47 20.705 3.73 ;
      RECT 19.905 2.62 19.991 3.034 ;
      RECT 19.905 2.62 20.03 3.031 ;
      RECT 19.905 2.62 20.05 3.021 ;
      RECT 19.86 2.62 20.05 3.018 ;
      RECT 19.86 2.772 20.06 3.008 ;
      RECT 19.86 2.793 20.065 3.002 ;
      RECT 19.86 2.811 20.07 2.998 ;
      RECT 19.86 2.831 20.08 2.993 ;
      RECT 19.835 2.831 20.08 2.99 ;
      RECT 19.825 2.831 20.08 2.968 ;
      RECT 19.825 2.847 20.085 2.938 ;
      RECT 19.79 2.62 20.05 2.925 ;
      RECT 19.79 2.859 20.09 2.88 ;
      RECT 17.45 7.77 17.74 8 ;
      RECT 17.51 6.29 17.68 8 ;
      RECT 17.505 6.655 17.855 7.005 ;
      RECT 17.45 6.29 17.74 6.52 ;
      RECT 17.045 2.395 17.15 2.965 ;
      RECT 17.045 2.73 17.37 2.96 ;
      RECT 17.045 2.76 17.54 2.93 ;
      RECT 17.045 2.395 17.235 2.96 ;
      RECT 16.46 2.36 16.75 2.59 ;
      RECT 16.46 2.395 17.235 2.565 ;
      RECT 16.52 0.88 16.69 2.59 ;
      RECT 16.46 0.88 16.75 1.11 ;
      RECT 16.46 7.77 16.75 8 ;
      RECT 16.52 6.29 16.69 8 ;
      RECT 16.46 6.29 16.75 6.52 ;
      RECT 16.46 6.325 17.315 6.485 ;
      RECT 17.145 5.92 17.315 6.485 ;
      RECT 16.46 6.32 16.855 6.485 ;
      RECT 17.08 5.92 17.37 6.15 ;
      RECT 17.08 5.95 17.54 6.12 ;
      RECT 16.09 2.73 16.38 2.96 ;
      RECT 16.09 2.76 16.55 2.93 ;
      RECT 16.155 1.655 16.32 2.96 ;
      RECT 14.67 1.625 14.96 1.855 ;
      RECT 14.67 1.655 16.32 1.825 ;
      RECT 14.73 0.885 14.9 1.855 ;
      RECT 14.67 0.885 14.96 1.115 ;
      RECT 14.67 7.765 14.96 7.995 ;
      RECT 14.73 7.025 14.9 7.995 ;
      RECT 14.73 7.12 16.32 7.29 ;
      RECT 16.15 5.92 16.32 7.29 ;
      RECT 14.67 7.025 14.96 7.255 ;
      RECT 16.09 5.92 16.38 6.15 ;
      RECT 16.09 5.95 16.55 6.12 ;
      RECT 12.72 2.705 13.06 3.055 ;
      RECT 12.81 2.025 12.98 3.055 ;
      RECT 15.1 1.965 15.45 2.315 ;
      RECT 12.81 2.025 15.45 2.195 ;
      RECT 15.125 6.655 15.45 6.98 ;
      RECT 9.665 6.605 10.015 6.955 ;
      RECT 15.1 6.655 15.45 6.885 ;
      RECT 9.465 6.655 10.015 6.885 ;
      RECT 9.295 6.685 15.45 6.855 ;
      RECT 14.325 2.365 14.645 2.685 ;
      RECT 14.295 2.365 14.645 2.595 ;
      RECT 14.125 2.395 14.645 2.565 ;
      RECT 14.325 6.255 14.645 6.545 ;
      RECT 14.295 6.285 14.645 6.515 ;
      RECT 14.125 6.315 14.645 6.485 ;
      RECT 10.015 2.985 10.165 3.26 ;
      RECT 10.555 2.065 10.56 2.285 ;
      RECT 11.705 2.265 11.72 2.463 ;
      RECT 11.67 2.257 11.705 2.47 ;
      RECT 11.64 2.25 11.67 2.47 ;
      RECT 11.585 2.215 11.64 2.47 ;
      RECT 11.52 2.152 11.585 2.47 ;
      RECT 11.515 2.117 11.52 2.468 ;
      RECT 11.51 2.112 11.515 2.46 ;
      RECT 11.505 2.107 11.51 2.446 ;
      RECT 11.5 2.104 11.505 2.439 ;
      RECT 11.455 2.094 11.5 2.39 ;
      RECT 11.435 2.081 11.455 2.325 ;
      RECT 11.43 2.076 11.435 2.298 ;
      RECT 11.425 2.075 11.43 2.291 ;
      RECT 11.42 2.074 11.425 2.284 ;
      RECT 11.335 2.059 11.42 2.23 ;
      RECT 11.305 2.04 11.335 2.18 ;
      RECT 11.225 2.023 11.305 2.165 ;
      RECT 11.19 2.01 11.225 2.15 ;
      RECT 11.182 2.01 11.19 2.145 ;
      RECT 11.096 2.011 11.182 2.145 ;
      RECT 11.01 2.013 11.096 2.145 ;
      RECT 10.985 2.014 11.01 2.149 ;
      RECT 10.91 2.02 10.985 2.164 ;
      RECT 10.827 2.032 10.91 2.188 ;
      RECT 10.741 2.045 10.827 2.214 ;
      RECT 10.655 2.058 10.741 2.24 ;
      RECT 10.62 2.067 10.655 2.259 ;
      RECT 10.57 2.067 10.62 2.272 ;
      RECT 10.56 2.065 10.57 2.283 ;
      RECT 10.545 2.062 10.555 2.285 ;
      RECT 10.53 2.054 10.545 2.293 ;
      RECT 10.515 2.046 10.53 2.313 ;
      RECT 10.51 2.041 10.515 2.37 ;
      RECT 10.495 2.036 10.51 2.443 ;
      RECT 10.49 2.031 10.495 2.485 ;
      RECT 10.485 2.029 10.49 2.513 ;
      RECT 10.48 2.027 10.485 2.535 ;
      RECT 10.47 2.023 10.48 2.578 ;
      RECT 10.465 2.02 10.47 2.603 ;
      RECT 10.46 2.018 10.465 2.623 ;
      RECT 10.455 2.016 10.46 2.647 ;
      RECT 10.45 2.012 10.455 2.67 ;
      RECT 10.445 2.008 10.45 2.693 ;
      RECT 10.41 1.998 10.445 2.8 ;
      RECT 10.405 1.988 10.41 2.898 ;
      RECT 10.4 1.986 10.405 2.925 ;
      RECT 10.395 1.985 10.4 2.945 ;
      RECT 10.39 1.977 10.395 2.965 ;
      RECT 10.385 1.972 10.39 3 ;
      RECT 10.38 1.97 10.385 3.018 ;
      RECT 10.375 1.97 10.38 3.043 ;
      RECT 10.37 1.97 10.375 3.065 ;
      RECT 10.335 1.97 10.37 3.108 ;
      RECT 10.31 1.97 10.335 3.137 ;
      RECT 10.3 1.97 10.31 2.323 ;
      RECT 10.303 2.38 10.31 3.147 ;
      RECT 10.3 2.437 10.303 3.15 ;
      RECT 10.295 1.97 10.3 2.295 ;
      RECT 10.295 2.487 10.3 3.153 ;
      RECT 10.285 1.97 10.295 2.285 ;
      RECT 10.29 2.54 10.295 3.156 ;
      RECT 10.285 2.625 10.29 3.16 ;
      RECT 10.275 1.97 10.285 2.273 ;
      RECT 10.28 2.672 10.285 3.164 ;
      RECT 10.275 2.747 10.28 3.168 ;
      RECT 10.24 1.97 10.275 2.248 ;
      RECT 10.265 2.83 10.275 3.173 ;
      RECT 10.255 2.897 10.265 3.18 ;
      RECT 10.25 2.925 10.255 3.185 ;
      RECT 10.24 2.938 10.25 3.191 ;
      RECT 10.195 1.97 10.24 2.205 ;
      RECT 10.235 2.943 10.24 3.198 ;
      RECT 10.195 2.96 10.235 3.26 ;
      RECT 10.19 1.972 10.195 2.178 ;
      RECT 10.165 2.98 10.195 3.26 ;
      RECT 10.185 1.977 10.19 2.15 ;
      RECT 9.975 2.989 10.015 3.26 ;
      RECT 9.95 2.997 9.975 3.23 ;
      RECT 9.905 3.005 9.95 3.23 ;
      RECT 9.89 3.01 9.905 3.225 ;
      RECT 9.88 3.01 9.89 3.219 ;
      RECT 9.87 3.017 9.88 3.216 ;
      RECT 9.865 3.055 9.87 3.205 ;
      RECT 9.86 3.117 9.865 3.183 ;
      RECT 11.13 2.992 11.315 3.215 ;
      RECT 11.13 3.007 11.32 3.211 ;
      RECT 11.12 2.28 11.205 3.21 ;
      RECT 11.12 3.007 11.325 3.204 ;
      RECT 11.115 3.015 11.325 3.203 ;
      RECT 11.32 2.735 11.64 3.055 ;
      RECT 11.115 2.907 11.285 2.998 ;
      RECT 11.11 2.907 11.285 2.98 ;
      RECT 11.1 2.715 11.235 2.955 ;
      RECT 11.095 2.715 11.235 2.9 ;
      RECT 11.055 2.295 11.225 2.8 ;
      RECT 11.04 2.295 11.225 2.67 ;
      RECT 11.035 2.295 11.225 2.623 ;
      RECT 11.03 2.295 11.225 2.603 ;
      RECT 11.025 2.295 11.225 2.578 ;
      RECT 10.995 2.295 11.255 2.555 ;
      RECT 11.005 2.292 11.215 2.555 ;
      RECT 11.13 2.287 11.215 3.215 ;
      RECT 11.015 2.28 11.205 2.555 ;
      RECT 11.01 2.285 11.205 2.555 ;
      RECT 9.84 2.497 10.025 2.71 ;
      RECT 9.84 2.505 10.035 2.703 ;
      RECT 9.82 2.505 10.035 2.7 ;
      RECT 9.815 2.505 10.035 2.685 ;
      RECT 9.745 2.42 10.005 2.68 ;
      RECT 9.745 2.565 10.04 2.593 ;
      RECT 9.4 3.02 9.66 3.28 ;
      RECT 9.425 2.965 9.62 3.28 ;
      RECT 9.42 2.714 9.6 3.008 ;
      RECT 9.42 2.72 9.61 3.008 ;
      RECT 9.4 2.722 9.61 2.953 ;
      RECT 9.395 2.732 9.61 2.82 ;
      RECT 9.425 2.712 9.6 3.28 ;
      RECT 9.511 2.71 9.6 3.28 ;
      RECT 9.37 1.93 9.405 2.3 ;
      RECT 9.16 2.04 9.165 2.3 ;
      RECT 9.405 1.937 9.42 2.3 ;
      RECT 9.295 1.93 9.37 2.378 ;
      RECT 9.285 1.93 9.295 2.463 ;
      RECT 9.26 1.93 9.285 2.498 ;
      RECT 9.22 1.93 9.26 2.566 ;
      RECT 9.21 1.937 9.22 2.618 ;
      RECT 9.18 2.04 9.21 2.659 ;
      RECT 9.175 2.04 9.18 2.698 ;
      RECT 9.165 2.04 9.175 2.718 ;
      RECT 9.16 2.335 9.165 2.755 ;
      RECT 9.155 2.352 9.16 2.775 ;
      RECT 9.14 2.415 9.155 2.815 ;
      RECT 9.135 2.458 9.14 2.85 ;
      RECT 9.13 2.466 9.135 2.863 ;
      RECT 9.12 2.48 9.13 2.885 ;
      RECT 9.095 2.515 9.12 2.95 ;
      RECT 9.085 2.55 9.095 3.013 ;
      RECT 9.065 2.58 9.085 3.074 ;
      RECT 9.05 2.616 9.065 3.141 ;
      RECT 9.04 2.644 9.05 3.18 ;
      RECT 9.03 2.666 9.04 3.2 ;
      RECT 9.025 2.676 9.03 3.211 ;
      RECT 9.02 2.685 9.025 3.214 ;
      RECT 9.01 2.703 9.02 3.218 ;
      RECT 9 2.721 9.01 3.219 ;
      RECT 8.975 2.76 9 3.216 ;
      RECT 8.955 2.802 8.975 3.213 ;
      RECT 8.94 2.84 8.955 3.212 ;
      RECT 8.905 2.875 8.94 3.209 ;
      RECT 8.9 2.897 8.905 3.207 ;
      RECT 8.835 2.937 8.9 3.204 ;
      RECT 8.83 2.977 8.835 3.2 ;
      RECT 8.815 2.987 8.83 3.191 ;
      RECT 8.805 3.107 8.815 3.176 ;
      RECT 9.285 3.52 9.295 3.78 ;
      RECT 9.285 3.523 9.305 3.779 ;
      RECT 9.275 3.513 9.285 3.778 ;
      RECT 9.265 3.528 9.345 3.774 ;
      RECT 9.25 3.507 9.265 3.772 ;
      RECT 9.225 3.532 9.35 3.768 ;
      RECT 9.21 3.492 9.225 3.763 ;
      RECT 9.21 3.534 9.36 3.762 ;
      RECT 9.21 3.542 9.375 3.755 ;
      RECT 9.15 3.479 9.21 3.745 ;
      RECT 9.14 3.466 9.15 3.727 ;
      RECT 9.115 3.456 9.14 3.717 ;
      RECT 9.11 3.446 9.115 3.709 ;
      RECT 9.045 3.542 9.375 3.691 ;
      RECT 8.96 3.542 9.375 3.653 ;
      RECT 8.85 3.37 9.11 3.63 ;
      RECT 9.225 3.5 9.25 3.768 ;
      RECT 9.265 3.51 9.275 3.774 ;
      RECT 8.85 3.518 9.29 3.63 ;
      RECT 9.035 7.765 9.325 7.995 ;
      RECT 9.095 7.025 9.265 7.995 ;
      RECT 8.995 7.055 9.365 7.425 ;
      RECT 9.035 7.025 9.325 7.425 ;
      RECT 8.065 3.275 8.095 3.575 ;
      RECT 7.84 3.26 7.845 3.535 ;
      RECT 7.64 3.26 7.795 3.52 ;
      RECT 8.94 1.975 8.97 2.235 ;
      RECT 8.93 1.975 8.94 2.343 ;
      RECT 8.91 1.975 8.93 2.353 ;
      RECT 8.895 1.975 8.91 2.365 ;
      RECT 8.84 1.975 8.895 2.415 ;
      RECT 8.825 1.975 8.84 2.463 ;
      RECT 8.795 1.975 8.825 2.498 ;
      RECT 8.74 1.975 8.795 2.56 ;
      RECT 8.72 1.975 8.74 2.628 ;
      RECT 8.715 1.975 8.72 2.658 ;
      RECT 8.71 1.975 8.715 2.67 ;
      RECT 8.705 2.092 8.71 2.688 ;
      RECT 8.685 2.11 8.705 2.713 ;
      RECT 8.665 2.137 8.685 2.763 ;
      RECT 8.66 2.157 8.665 2.794 ;
      RECT 8.655 2.165 8.66 2.811 ;
      RECT 8.64 2.191 8.655 2.84 ;
      RECT 8.625 2.233 8.64 2.875 ;
      RECT 8.62 2.262 8.625 2.898 ;
      RECT 8.615 2.277 8.62 2.911 ;
      RECT 8.61 2.3 8.615 2.922 ;
      RECT 8.6 2.32 8.61 2.94 ;
      RECT 8.59 2.35 8.6 2.963 ;
      RECT 8.585 2.372 8.59 2.983 ;
      RECT 8.58 2.387 8.585 2.998 ;
      RECT 8.565 2.417 8.58 3.025 ;
      RECT 8.56 2.447 8.565 3.051 ;
      RECT 8.555 2.465 8.56 3.063 ;
      RECT 8.545 2.495 8.555 3.082 ;
      RECT 8.535 2.52 8.545 3.107 ;
      RECT 8.53 2.54 8.535 3.126 ;
      RECT 8.525 2.557 8.53 3.139 ;
      RECT 8.515 2.583 8.525 3.158 ;
      RECT 8.505 2.621 8.515 3.185 ;
      RECT 8.5 2.647 8.505 3.205 ;
      RECT 8.495 2.657 8.5 3.215 ;
      RECT 8.49 2.67 8.495 3.23 ;
      RECT 8.485 2.685 8.49 3.24 ;
      RECT 8.48 2.707 8.485 3.255 ;
      RECT 8.475 2.725 8.48 3.266 ;
      RECT 8.47 2.735 8.475 3.277 ;
      RECT 8.465 2.743 8.47 3.289 ;
      RECT 8.46 2.751 8.465 3.3 ;
      RECT 8.455 2.777 8.46 3.313 ;
      RECT 8.445 2.805 8.455 3.326 ;
      RECT 8.44 2.835 8.445 3.335 ;
      RECT 8.435 2.85 8.44 3.342 ;
      RECT 8.42 2.875 8.435 3.349 ;
      RECT 8.415 2.897 8.42 3.355 ;
      RECT 8.41 2.922 8.415 3.358 ;
      RECT 8.401 2.95 8.41 3.362 ;
      RECT 8.395 2.967 8.401 3.367 ;
      RECT 8.39 2.985 8.395 3.371 ;
      RECT 8.385 2.997 8.39 3.374 ;
      RECT 8.38 3.018 8.385 3.378 ;
      RECT 8.375 3.036 8.38 3.381 ;
      RECT 8.37 3.05 8.375 3.384 ;
      RECT 8.365 3.067 8.37 3.387 ;
      RECT 8.36 3.08 8.365 3.39 ;
      RECT 8.335 3.117 8.36 3.398 ;
      RECT 8.33 3.162 8.335 3.407 ;
      RECT 8.325 3.19 8.33 3.41 ;
      RECT 8.315 3.21 8.325 3.414 ;
      RECT 8.31 3.23 8.315 3.419 ;
      RECT 8.305 3.245 8.31 3.422 ;
      RECT 8.285 3.255 8.305 3.429 ;
      RECT 8.22 3.262 8.285 3.455 ;
      RECT 8.185 3.265 8.22 3.483 ;
      RECT 8.17 3.268 8.185 3.498 ;
      RECT 8.16 3.269 8.17 3.513 ;
      RECT 8.15 3.27 8.16 3.53 ;
      RECT 8.145 3.27 8.15 3.545 ;
      RECT 8.14 3.27 8.145 3.553 ;
      RECT 8.125 3.271 8.14 3.568 ;
      RECT 8.095 3.273 8.125 3.575 ;
      RECT 7.985 3.28 8.065 3.575 ;
      RECT 7.94 3.285 7.985 3.575 ;
      RECT 7.93 3.286 7.94 3.565 ;
      RECT 7.92 3.287 7.93 3.558 ;
      RECT 7.9 3.289 7.92 3.553 ;
      RECT 7.89 3.26 7.9 3.548 ;
      RECT 7.845 3.26 7.89 3.54 ;
      RECT 7.815 3.26 7.84 3.53 ;
      RECT 7.795 3.26 7.815 3.523 ;
      RECT 8.075 2.06 8.335 2.32 ;
      RECT 7.955 2.075 7.965 2.24 ;
      RECT 7.94 2.075 7.945 2.235 ;
      RECT 5.305 1.915 5.49 2.205 ;
      RECT 7.12 2.04 7.135 2.195 ;
      RECT 5.27 1.915 5.295 2.175 ;
      RECT 7.685 1.965 7.69 2.107 ;
      RECT 7.6 1.96 7.625 2.1 ;
      RECT 8 2.077 8.075 2.27 ;
      RECT 7.985 2.075 8 2.253 ;
      RECT 7.965 2.075 7.985 2.245 ;
      RECT 7.945 2.075 7.955 2.238 ;
      RECT 7.9 2.07 7.94 2.228 ;
      RECT 7.86 2.045 7.9 2.213 ;
      RECT 7.845 2.02 7.86 2.203 ;
      RECT 7.84 2.014 7.845 2.201 ;
      RECT 7.805 2.006 7.84 2.184 ;
      RECT 7.8 1.999 7.805 2.172 ;
      RECT 7.78 1.994 7.8 2.16 ;
      RECT 7.77 1.988 7.78 2.145 ;
      RECT 7.75 1.983 7.77 2.13 ;
      RECT 7.74 1.978 7.75 2.123 ;
      RECT 7.735 1.976 7.74 2.118 ;
      RECT 7.73 1.975 7.735 2.115 ;
      RECT 7.69 1.97 7.73 2.111 ;
      RECT 7.67 1.964 7.685 2.106 ;
      RECT 7.635 1.961 7.67 2.103 ;
      RECT 7.625 1.96 7.635 2.101 ;
      RECT 7.565 1.96 7.6 2.098 ;
      RECT 7.52 1.96 7.565 2.098 ;
      RECT 7.47 1.96 7.52 2.101 ;
      RECT 7.455 1.962 7.47 2.103 ;
      RECT 7.44 1.965 7.455 2.104 ;
      RECT 7.43 1.97 7.44 2.105 ;
      RECT 7.4 1.975 7.43 2.11 ;
      RECT 7.39 1.981 7.4 2.118 ;
      RECT 7.38 1.983 7.39 2.122 ;
      RECT 7.37 1.987 7.38 2.126 ;
      RECT 7.345 1.993 7.37 2.134 ;
      RECT 7.335 1.998 7.345 2.142 ;
      RECT 7.32 2.002 7.335 2.146 ;
      RECT 7.285 2.008 7.32 2.154 ;
      RECT 7.265 2.013 7.285 2.164 ;
      RECT 7.235 2.02 7.265 2.173 ;
      RECT 7.19 2.029 7.235 2.187 ;
      RECT 7.185 2.034 7.19 2.198 ;
      RECT 7.165 2.037 7.185 2.199 ;
      RECT 7.135 2.04 7.165 2.197 ;
      RECT 7.1 2.04 7.12 2.193 ;
      RECT 7.03 2.04 7.1 2.184 ;
      RECT 7.015 2.037 7.03 2.176 ;
      RECT 6.975 2.03 7.015 2.171 ;
      RECT 6.95 2.02 6.975 2.164 ;
      RECT 6.945 2.014 6.95 2.161 ;
      RECT 6.905 2.008 6.945 2.158 ;
      RECT 6.89 2.001 6.905 2.153 ;
      RECT 6.87 1.997 6.89 2.148 ;
      RECT 6.855 1.992 6.87 2.144 ;
      RECT 6.84 1.987 6.855 2.142 ;
      RECT 6.825 1.983 6.84 2.141 ;
      RECT 6.81 1.981 6.825 2.137 ;
      RECT 6.8 1.979 6.81 2.132 ;
      RECT 6.785 1.976 6.8 2.128 ;
      RECT 6.775 1.974 6.785 2.123 ;
      RECT 6.755 1.971 6.775 2.119 ;
      RECT 6.71 1.97 6.755 2.117 ;
      RECT 6.65 1.972 6.71 2.118 ;
      RECT 6.63 1.974 6.65 2.12 ;
      RECT 6.6 1.977 6.63 2.121 ;
      RECT 6.55 1.982 6.6 2.123 ;
      RECT 6.545 1.985 6.55 2.125 ;
      RECT 6.535 1.987 6.545 2.128 ;
      RECT 6.53 1.989 6.535 2.131 ;
      RECT 6.48 1.992 6.53 2.138 ;
      RECT 6.46 1.996 6.48 2.15 ;
      RECT 6.45 1.999 6.46 2.156 ;
      RECT 6.44 2 6.45 2.159 ;
      RECT 6.401 2.003 6.44 2.161 ;
      RECT 6.315 2.01 6.401 2.164 ;
      RECT 6.241 2.02 6.315 2.168 ;
      RECT 6.155 2.031 6.241 2.173 ;
      RECT 6.14 2.038 6.155 2.175 ;
      RECT 6.085 2.042 6.14 2.176 ;
      RECT 6.071 2.045 6.085 2.178 ;
      RECT 5.985 2.045 6.071 2.18 ;
      RECT 5.945 2.042 5.985 2.183 ;
      RECT 5.921 2.038 5.945 2.185 ;
      RECT 5.835 2.028 5.921 2.188 ;
      RECT 5.805 2.017 5.835 2.189 ;
      RECT 5.786 2.013 5.805 2.188 ;
      RECT 5.7 2.006 5.786 2.185 ;
      RECT 5.64 1.995 5.7 2.182 ;
      RECT 5.62 1.987 5.64 2.18 ;
      RECT 5.585 1.982 5.62 2.179 ;
      RECT 5.56 1.977 5.585 2.178 ;
      RECT 5.53 1.972 5.56 2.177 ;
      RECT 5.505 1.915 5.53 2.176 ;
      RECT 5.49 1.915 5.505 2.2 ;
      RECT 5.295 1.915 5.305 2.2 ;
      RECT 7.07 2.935 7.075 3.075 ;
      RECT 6.73 2.935 6.765 3.073 ;
      RECT 6.305 2.92 6.32 3.065 ;
      RECT 8.135 2.7 8.225 2.96 ;
      RECT 7.965 2.565 8.065 2.96 ;
      RECT 5 2.54 5.08 2.75 ;
      RECT 8.09 2.677 8.135 2.96 ;
      RECT 8.08 2.647 8.09 2.96 ;
      RECT 8.065 2.57 8.08 2.96 ;
      RECT 7.88 2.565 7.965 2.925 ;
      RECT 7.875 2.567 7.88 2.92 ;
      RECT 7.87 2.572 7.875 2.92 ;
      RECT 7.835 2.672 7.87 2.92 ;
      RECT 7.825 2.7 7.835 2.92 ;
      RECT 7.815 2.715 7.825 2.92 ;
      RECT 7.805 2.727 7.815 2.92 ;
      RECT 7.8 2.737 7.805 2.92 ;
      RECT 7.785 2.747 7.8 2.922 ;
      RECT 7.78 2.762 7.785 2.924 ;
      RECT 7.765 2.775 7.78 2.926 ;
      RECT 7.76 2.79 7.765 2.929 ;
      RECT 7.74 2.8 7.76 2.933 ;
      RECT 7.725 2.81 7.74 2.936 ;
      RECT 7.69 2.817 7.725 2.941 ;
      RECT 7.646 2.824 7.69 2.949 ;
      RECT 7.56 2.836 7.646 2.962 ;
      RECT 7.535 2.847 7.56 2.973 ;
      RECT 7.505 2.852 7.535 2.978 ;
      RECT 7.47 2.857 7.505 2.986 ;
      RECT 7.44 2.862 7.47 2.993 ;
      RECT 7.415 2.867 7.44 2.998 ;
      RECT 7.35 2.874 7.415 3.007 ;
      RECT 7.28 2.887 7.35 3.023 ;
      RECT 7.25 2.897 7.28 3.035 ;
      RECT 7.225 2.902 7.25 3.042 ;
      RECT 7.17 2.909 7.225 3.05 ;
      RECT 7.165 2.916 7.17 3.055 ;
      RECT 7.16 2.918 7.165 3.056 ;
      RECT 7.145 2.92 7.16 3.058 ;
      RECT 7.14 2.92 7.145 3.061 ;
      RECT 7.075 2.927 7.14 3.068 ;
      RECT 7.04 2.937 7.07 3.078 ;
      RECT 7.023 2.94 7.04 3.08 ;
      RECT 6.937 2.939 7.023 3.079 ;
      RECT 6.851 2.937 6.937 3.076 ;
      RECT 6.765 2.936 6.851 3.074 ;
      RECT 6.664 2.934 6.73 3.073 ;
      RECT 6.578 2.931 6.664 3.071 ;
      RECT 6.492 2.927 6.578 3.069 ;
      RECT 6.406 2.924 6.492 3.068 ;
      RECT 6.32 2.921 6.406 3.066 ;
      RECT 6.22 2.92 6.305 3.063 ;
      RECT 6.17 2.918 6.22 3.061 ;
      RECT 6.15 2.915 6.17 3.059 ;
      RECT 6.13 2.913 6.15 3.056 ;
      RECT 6.105 2.909 6.13 3.053 ;
      RECT 6.06 2.903 6.105 3.048 ;
      RECT 6.02 2.897 6.06 3.04 ;
      RECT 5.995 2.892 6.02 3.033 ;
      RECT 5.94 2.885 5.995 3.025 ;
      RECT 5.916 2.878 5.94 3.018 ;
      RECT 5.83 2.869 5.916 3.008 ;
      RECT 5.8 2.861 5.83 2.998 ;
      RECT 5.77 2.857 5.8 2.993 ;
      RECT 5.765 2.854 5.77 2.99 ;
      RECT 5.76 2.853 5.765 2.99 ;
      RECT 5.685 2.846 5.76 2.983 ;
      RECT 5.646 2.837 5.685 2.972 ;
      RECT 5.56 2.827 5.646 2.96 ;
      RECT 5.52 2.817 5.56 2.948 ;
      RECT 5.481 2.812 5.52 2.941 ;
      RECT 5.395 2.802 5.481 2.93 ;
      RECT 5.355 2.79 5.395 2.919 ;
      RECT 5.32 2.775 5.355 2.912 ;
      RECT 5.31 2.765 5.32 2.909 ;
      RECT 5.29 2.75 5.31 2.907 ;
      RECT 5.26 2.72 5.29 2.903 ;
      RECT 5.25 2.7 5.26 2.898 ;
      RECT 5.245 2.692 5.25 2.895 ;
      RECT 5.24 2.685 5.245 2.893 ;
      RECT 5.225 2.672 5.24 2.886 ;
      RECT 5.22 2.662 5.225 2.878 ;
      RECT 5.215 2.655 5.22 2.873 ;
      RECT 5.21 2.65 5.215 2.869 ;
      RECT 5.195 2.637 5.21 2.861 ;
      RECT 5.19 2.547 5.195 2.85 ;
      RECT 5.185 2.542 5.19 2.843 ;
      RECT 5.11 2.54 5.185 2.803 ;
      RECT 5.08 2.54 5.11 2.758 ;
      RECT 4.985 2.545 5 2.745 ;
      RECT 7.47 2.25 7.73 2.51 ;
      RECT 7.455 2.238 7.635 2.475 ;
      RECT 7.45 2.239 7.635 2.473 ;
      RECT 7.435 2.243 7.645 2.463 ;
      RECT 7.43 2.248 7.65 2.433 ;
      RECT 7.435 2.245 7.65 2.463 ;
      RECT 7.45 2.24 7.645 2.473 ;
      RECT 7.47 2.237 7.635 2.51 ;
      RECT 7.47 2.236 7.625 2.51 ;
      RECT 7.495 2.235 7.625 2.51 ;
      RECT 7.055 2.48 7.315 2.74 ;
      RECT 6.93 2.525 7.315 2.735 ;
      RECT 6.92 2.53 7.315 2.73 ;
      RECT 6.935 3.47 6.95 3.78 ;
      RECT 5.53 3.24 5.54 3.37 ;
      RECT 5.31 3.235 5.415 3.37 ;
      RECT 5.225 3.24 5.275 3.37 ;
      RECT 3.775 1.975 3.78 3.08 ;
      RECT 7.03 3.562 7.035 3.698 ;
      RECT 7.025 3.557 7.03 3.758 ;
      RECT 7.02 3.555 7.025 3.771 ;
      RECT 7.005 3.552 7.02 3.773 ;
      RECT 7 3.547 7.005 3.775 ;
      RECT 6.995 3.543 7 3.778 ;
      RECT 6.98 3.538 6.995 3.78 ;
      RECT 6.95 3.53 6.98 3.78 ;
      RECT 6.911 3.47 6.935 3.78 ;
      RECT 6.825 3.47 6.911 3.777 ;
      RECT 6.795 3.47 6.825 3.77 ;
      RECT 6.77 3.47 6.795 3.763 ;
      RECT 6.745 3.47 6.77 3.755 ;
      RECT 6.73 3.47 6.745 3.748 ;
      RECT 6.705 3.47 6.73 3.74 ;
      RECT 6.69 3.47 6.705 3.733 ;
      RECT 6.65 3.48 6.69 3.722 ;
      RECT 6.64 3.475 6.65 3.712 ;
      RECT 6.636 3.474 6.64 3.709 ;
      RECT 6.55 3.466 6.636 3.692 ;
      RECT 6.517 3.455 6.55 3.669 ;
      RECT 6.431 3.444 6.517 3.647 ;
      RECT 6.345 3.428 6.431 3.616 ;
      RECT 6.275 3.413 6.345 3.588 ;
      RECT 6.265 3.406 6.275 3.575 ;
      RECT 6.235 3.403 6.265 3.565 ;
      RECT 6.21 3.399 6.235 3.558 ;
      RECT 6.195 3.396 6.21 3.553 ;
      RECT 6.19 3.395 6.195 3.548 ;
      RECT 6.16 3.39 6.19 3.541 ;
      RECT 6.155 3.385 6.16 3.536 ;
      RECT 6.14 3.382 6.155 3.531 ;
      RECT 6.135 3.377 6.14 3.526 ;
      RECT 6.115 3.372 6.135 3.523 ;
      RECT 6.1 3.367 6.115 3.515 ;
      RECT 6.085 3.361 6.1 3.51 ;
      RECT 6.055 3.352 6.085 3.503 ;
      RECT 6.05 3.345 6.055 3.495 ;
      RECT 6.045 3.343 6.05 3.493 ;
      RECT 6.04 3.342 6.045 3.49 ;
      RECT 6 3.335 6.04 3.483 ;
      RECT 5.986 3.325 6 3.473 ;
      RECT 5.935 3.314 5.986 3.461 ;
      RECT 5.91 3.3 5.935 3.447 ;
      RECT 5.885 3.289 5.91 3.439 ;
      RECT 5.865 3.278 5.885 3.433 ;
      RECT 5.855 3.272 5.865 3.428 ;
      RECT 5.85 3.27 5.855 3.424 ;
      RECT 5.83 3.265 5.85 3.419 ;
      RECT 5.8 3.255 5.83 3.409 ;
      RECT 5.795 3.247 5.8 3.402 ;
      RECT 5.78 3.245 5.795 3.398 ;
      RECT 5.76 3.245 5.78 3.393 ;
      RECT 5.755 3.244 5.76 3.391 ;
      RECT 5.75 3.244 5.755 3.388 ;
      RECT 5.71 3.243 5.75 3.383 ;
      RECT 5.685 3.242 5.71 3.378 ;
      RECT 5.625 3.241 5.685 3.375 ;
      RECT 5.54 3.24 5.625 3.373 ;
      RECT 5.501 3.239 5.53 3.37 ;
      RECT 5.415 3.237 5.501 3.37 ;
      RECT 5.275 3.237 5.31 3.37 ;
      RECT 5.185 3.241 5.225 3.373 ;
      RECT 5.17 3.244 5.185 3.38 ;
      RECT 5.16 3.245 5.17 3.387 ;
      RECT 5.135 3.248 5.16 3.392 ;
      RECT 5.13 3.25 5.135 3.395 ;
      RECT 5.08 3.252 5.13 3.396 ;
      RECT 5.041 3.256 5.08 3.398 ;
      RECT 4.955 3.258 5.041 3.401 ;
      RECT 4.937 3.26 4.955 3.403 ;
      RECT 4.851 3.263 4.937 3.405 ;
      RECT 4.765 3.267 4.851 3.408 ;
      RECT 4.728 3.271 4.765 3.411 ;
      RECT 4.642 3.274 4.728 3.414 ;
      RECT 4.556 3.278 4.642 3.417 ;
      RECT 4.47 3.283 4.556 3.421 ;
      RECT 4.45 3.285 4.47 3.424 ;
      RECT 4.43 3.284 4.45 3.425 ;
      RECT 4.381 3.281 4.43 3.426 ;
      RECT 4.295 3.276 4.381 3.429 ;
      RECT 4.245 3.271 4.295 3.431 ;
      RECT 4.221 3.269 4.245 3.432 ;
      RECT 4.135 3.264 4.221 3.434 ;
      RECT 4.11 3.26 4.135 3.433 ;
      RECT 4.1 3.257 4.11 3.431 ;
      RECT 4.09 3.25 4.1 3.428 ;
      RECT 4.085 3.23 4.09 3.423 ;
      RECT 4.075 3.2 4.085 3.418 ;
      RECT 4.06 3.07 4.075 3.409 ;
      RECT 4.055 3.062 4.06 3.402 ;
      RECT 4.035 3.055 4.055 3.394 ;
      RECT 4.03 3.037 4.035 3.386 ;
      RECT 4.02 3.017 4.03 3.381 ;
      RECT 4.015 2.99 4.02 3.377 ;
      RECT 4.01 2.967 4.015 3.374 ;
      RECT 3.99 2.925 4.01 3.366 ;
      RECT 3.955 2.84 3.99 3.35 ;
      RECT 3.95 2.772 3.955 3.338 ;
      RECT 3.935 2.742 3.95 3.332 ;
      RECT 3.93 1.987 3.935 2.233 ;
      RECT 3.92 2.712 3.935 3.323 ;
      RECT 3.925 1.982 3.93 2.265 ;
      RECT 3.92 1.977 3.925 2.308 ;
      RECT 3.915 1.975 3.92 2.343 ;
      RECT 3.9 2.675 3.92 3.313 ;
      RECT 3.91 1.975 3.915 2.38 ;
      RECT 3.895 1.975 3.91 2.478 ;
      RECT 3.895 2.648 3.9 3.306 ;
      RECT 3.89 1.975 3.895 2.553 ;
      RECT 3.89 2.636 3.895 3.303 ;
      RECT 3.885 1.975 3.89 2.585 ;
      RECT 3.885 2.615 3.89 3.3 ;
      RECT 3.88 1.975 3.885 3.297 ;
      RECT 3.845 1.975 3.88 3.283 ;
      RECT 3.83 1.975 3.845 3.265 ;
      RECT 3.81 1.975 3.83 3.255 ;
      RECT 3.785 1.975 3.81 3.238 ;
      RECT 3.78 1.975 3.785 3.188 ;
      RECT 3.77 1.975 3.775 3.018 ;
      RECT 3.765 1.975 3.77 2.925 ;
      RECT 3.76 1.975 3.765 2.838 ;
      RECT 3.755 1.975 3.76 2.77 ;
      RECT 3.75 1.975 3.755 2.713 ;
      RECT 3.74 1.975 3.75 2.608 ;
      RECT 3.735 1.975 3.74 2.48 ;
      RECT 3.73 1.975 3.735 2.398 ;
      RECT 3.725 1.977 3.73 2.315 ;
      RECT 3.72 1.982 3.725 2.248 ;
      RECT 3.715 1.987 3.72 2.175 ;
      RECT 6.53 2.305 6.79 2.565 ;
      RECT 6.55 2.272 6.76 2.565 ;
      RECT 6.55 2.27 6.75 2.565 ;
      RECT 6.56 2.257 6.75 2.565 ;
      RECT 6.56 2.255 6.675 2.565 ;
      RECT 6.035 2.38 6.21 2.66 ;
      RECT 6.03 2.38 6.21 2.658 ;
      RECT 6.03 2.38 6.225 2.655 ;
      RECT 6.02 2.38 6.225 2.653 ;
      RECT 5.965 2.38 6.225 2.64 ;
      RECT 5.965 2.455 6.23 2.618 ;
      RECT 5.51 2.392 5.53 2.635 ;
      RECT 5.51 2.392 5.57 2.634 ;
      RECT 5.505 2.394 5.57 2.633 ;
      RECT 5.505 2.394 5.656 2.632 ;
      RECT 5.505 2.394 5.725 2.631 ;
      RECT 5.505 2.394 5.745 2.623 ;
      RECT 5.485 2.397 5.745 2.621 ;
      RECT 5.47 2.407 5.745 2.606 ;
      RECT 5.47 2.407 5.76 2.605 ;
      RECT 5.465 2.416 5.76 2.597 ;
      RECT 5.465 2.416 5.765 2.593 ;
      RECT 5.57 2.33 5.83 2.59 ;
      RECT 5.46 2.418 5.83 2.475 ;
      RECT 5.53 2.385 5.83 2.59 ;
      RECT 5.495 3.578 5.5 3.785 ;
      RECT 5.445 3.572 5.495 3.784 ;
      RECT 5.412 3.586 5.505 3.783 ;
      RECT 5.326 3.586 5.505 3.782 ;
      RECT 5.24 3.586 5.505 3.781 ;
      RECT 5.24 3.685 5.51 3.778 ;
      RECT 5.235 3.685 5.51 3.773 ;
      RECT 5.23 3.685 5.51 3.755 ;
      RECT 5.225 3.685 5.51 3.738 ;
      RECT 5.185 3.47 5.445 3.73 ;
      RECT 4.645 2.62 4.731 3.034 ;
      RECT 4.645 2.62 4.77 3.031 ;
      RECT 4.645 2.62 4.79 3.021 ;
      RECT 4.6 2.62 4.79 3.018 ;
      RECT 4.6 2.772 4.8 3.008 ;
      RECT 4.6 2.793 4.805 3.002 ;
      RECT 4.6 2.811 4.81 2.998 ;
      RECT 4.6 2.831 4.82 2.993 ;
      RECT 4.575 2.831 4.82 2.99 ;
      RECT 4.565 2.831 4.82 2.968 ;
      RECT 4.565 2.847 4.825 2.938 ;
      RECT 4.53 2.62 4.79 2.925 ;
      RECT 4.53 2.859 4.83 2.88 ;
      RECT 1.54 7.765 1.83 7.995 ;
      RECT 1.6 7.025 1.77 7.995 ;
      RECT 1.51 7.025 1.86 7.315 ;
      RECT 1.135 6.285 1.485 6.575 ;
      RECT 0.995 6.315 1.485 6.485 ;
      RECT 68.155 3.265 68.415 3.525 ;
      RECT 52.895 3.265 53.155 3.525 ;
      RECT 37.635 3.265 37.895 3.525 ;
      RECT 22.375 3.265 22.635 3.525 ;
      RECT 7.115 3.265 7.375 3.525 ;
    LAYER mcon ;
      RECT 78.55 6.32 78.72 6.49 ;
      RECT 78.555 6.315 78.725 6.485 ;
      RECT 63.29 6.32 63.46 6.49 ;
      RECT 63.295 6.315 63.465 6.485 ;
      RECT 48.03 6.32 48.2 6.49 ;
      RECT 48.035 6.315 48.205 6.485 ;
      RECT 32.77 6.32 32.94 6.49 ;
      RECT 32.775 6.315 32.945 6.485 ;
      RECT 17.51 6.32 17.68 6.49 ;
      RECT 17.515 6.315 17.685 6.485 ;
      RECT 78.55 7.8 78.72 7.97 ;
      RECT 78.2 0.1 78.37 0.27 ;
      RECT 78.2 8.61 78.37 8.78 ;
      RECT 78.18 2.76 78.35 2.93 ;
      RECT 78.18 5.95 78.35 6.12 ;
      RECT 77.56 0.91 77.73 1.08 ;
      RECT 77.56 2.39 77.73 2.56 ;
      RECT 77.56 6.32 77.73 6.49 ;
      RECT 77.56 7.8 77.73 7.97 ;
      RECT 77.21 0.1 77.38 0.27 ;
      RECT 77.21 8.61 77.38 8.78 ;
      RECT 77.19 2.76 77.36 2.93 ;
      RECT 77.19 5.95 77.36 6.12 ;
      RECT 76.51 0.105 76.68 0.275 ;
      RECT 76.51 8.605 76.68 8.775 ;
      RECT 76.2 2.025 76.37 2.195 ;
      RECT 76.2 6.685 76.37 6.855 ;
      RECT 75.83 0.105 76 0.275 ;
      RECT 75.83 8.605 76 8.775 ;
      RECT 75.77 0.915 75.94 1.085 ;
      RECT 75.77 1.655 75.94 1.825 ;
      RECT 75.77 7.055 75.94 7.225 ;
      RECT 75.77 7.795 75.94 7.965 ;
      RECT 75.395 2.395 75.565 2.565 ;
      RECT 75.395 6.315 75.565 6.485 ;
      RECT 75.15 0.105 75.32 0.275 ;
      RECT 75.15 8.605 75.32 8.775 ;
      RECT 74.47 0.105 74.64 0.275 ;
      RECT 74.47 8.605 74.64 8.775 ;
      RECT 73.01 1.415 73.18 1.585 ;
      RECT 72.57 2.28 72.74 2.45 ;
      RECT 72.55 1.415 72.72 1.585 ;
      RECT 72.175 3.025 72.345 3.195 ;
      RECT 72.09 1.415 72.26 1.585 ;
      RECT 72.065 2.3 72.235 2.47 ;
      RECT 71.63 1.415 71.8 1.585 ;
      RECT 71.245 1.99 71.415 2.16 ;
      RECT 71.17 1.415 71.34 1.585 ;
      RECT 70.93 3.03 71.1 3.2 ;
      RECT 70.885 2.52 71.055 2.69 ;
      RECT 70.875 8.605 71.045 8.775 ;
      RECT 70.71 1.415 70.88 1.585 ;
      RECT 70.565 6.685 70.735 6.855 ;
      RECT 70.46 2.73 70.63 2.9 ;
      RECT 70.27 1.95 70.44 2.12 ;
      RECT 70.25 1.415 70.42 1.585 ;
      RECT 70.22 3.56 70.39 3.73 ;
      RECT 70.195 8.605 70.365 8.775 ;
      RECT 70.135 7.055 70.305 7.225 ;
      RECT 70.135 7.795 70.305 7.965 ;
      RECT 69.885 3 70.055 3.17 ;
      RECT 69.79 1.415 69.96 1.585 ;
      RECT 69.79 2.16 69.96 2.33 ;
      RECT 69.76 6.315 69.93 6.485 ;
      RECT 69.515 8.605 69.685 8.775 ;
      RECT 69.33 1.415 69.5 1.585 ;
      RECT 68.99 3.385 69.16 3.555 ;
      RECT 68.93 2.585 69.1 2.755 ;
      RECT 68.87 1.415 69.04 1.585 ;
      RECT 68.835 8.605 69.005 8.775 ;
      RECT 68.49 2.255 68.66 2.425 ;
      RECT 68.41 1.415 68.58 1.585 ;
      RECT 68.225 3.305 68.395 3.475 ;
      RECT 67.98 2.545 68.15 2.715 ;
      RECT 67.95 1.415 68.12 1.585 ;
      RECT 67.885 3.575 68.055 3.745 ;
      RECT 67.61 2.27 67.78 2.44 ;
      RECT 67.49 1.415 67.66 1.585 ;
      RECT 67.08 2.47 67.25 2.64 ;
      RECT 67.03 1.415 67.2 1.585 ;
      RECT 66.57 1.415 66.74 1.585 ;
      RECT 66.56 2.415 66.73 2.585 ;
      RECT 66.355 2.015 66.525 2.185 ;
      RECT 66.355 3.595 66.525 3.765 ;
      RECT 66.11 1.415 66.28 1.585 ;
      RECT 66.045 2.56 66.215 2.73 ;
      RECT 65.65 1.415 65.82 1.585 ;
      RECT 65.635 2.785 65.805 2.955 ;
      RECT 65.19 1.415 65.36 1.585 ;
      RECT 64.925 3.085 65.095 3.255 ;
      RECT 64.78 1.995 64.95 2.165 ;
      RECT 64.73 1.415 64.9 1.585 ;
      RECT 63.29 7.8 63.46 7.97 ;
      RECT 62.94 0.1 63.11 0.27 ;
      RECT 62.94 8.61 63.11 8.78 ;
      RECT 62.92 2.76 63.09 2.93 ;
      RECT 62.92 5.95 63.09 6.12 ;
      RECT 62.3 0.91 62.47 1.08 ;
      RECT 62.3 2.39 62.47 2.56 ;
      RECT 62.3 6.32 62.47 6.49 ;
      RECT 62.3 7.8 62.47 7.97 ;
      RECT 61.95 0.1 62.12 0.27 ;
      RECT 61.95 8.61 62.12 8.78 ;
      RECT 61.93 2.76 62.1 2.93 ;
      RECT 61.93 5.95 62.1 6.12 ;
      RECT 61.25 0.105 61.42 0.275 ;
      RECT 61.25 8.605 61.42 8.775 ;
      RECT 60.94 2.025 61.11 2.195 ;
      RECT 60.94 6.685 61.11 6.855 ;
      RECT 60.57 0.105 60.74 0.275 ;
      RECT 60.57 8.605 60.74 8.775 ;
      RECT 60.51 0.915 60.68 1.085 ;
      RECT 60.51 1.655 60.68 1.825 ;
      RECT 60.51 7.055 60.68 7.225 ;
      RECT 60.51 7.795 60.68 7.965 ;
      RECT 60.135 2.395 60.305 2.565 ;
      RECT 60.135 6.315 60.305 6.485 ;
      RECT 59.89 0.105 60.06 0.275 ;
      RECT 59.89 8.605 60.06 8.775 ;
      RECT 59.21 0.105 59.38 0.275 ;
      RECT 59.21 8.605 59.38 8.775 ;
      RECT 57.75 1.415 57.92 1.585 ;
      RECT 57.31 2.28 57.48 2.45 ;
      RECT 57.29 1.415 57.46 1.585 ;
      RECT 56.915 3.025 57.085 3.195 ;
      RECT 56.83 1.415 57 1.585 ;
      RECT 56.805 2.3 56.975 2.47 ;
      RECT 56.37 1.415 56.54 1.585 ;
      RECT 55.985 1.99 56.155 2.16 ;
      RECT 55.91 1.415 56.08 1.585 ;
      RECT 55.67 3.03 55.84 3.2 ;
      RECT 55.625 2.52 55.795 2.69 ;
      RECT 55.615 8.605 55.785 8.775 ;
      RECT 55.45 1.415 55.62 1.585 ;
      RECT 55.305 6.685 55.475 6.855 ;
      RECT 55.2 2.73 55.37 2.9 ;
      RECT 55.01 1.95 55.18 2.12 ;
      RECT 54.99 1.415 55.16 1.585 ;
      RECT 54.96 3.56 55.13 3.73 ;
      RECT 54.935 8.605 55.105 8.775 ;
      RECT 54.875 7.055 55.045 7.225 ;
      RECT 54.875 7.795 55.045 7.965 ;
      RECT 54.625 3 54.795 3.17 ;
      RECT 54.53 1.415 54.7 1.585 ;
      RECT 54.53 2.16 54.7 2.33 ;
      RECT 54.5 6.315 54.67 6.485 ;
      RECT 54.255 8.605 54.425 8.775 ;
      RECT 54.07 1.415 54.24 1.585 ;
      RECT 53.73 3.385 53.9 3.555 ;
      RECT 53.67 2.585 53.84 2.755 ;
      RECT 53.61 1.415 53.78 1.585 ;
      RECT 53.575 8.605 53.745 8.775 ;
      RECT 53.23 2.255 53.4 2.425 ;
      RECT 53.15 1.415 53.32 1.585 ;
      RECT 52.965 3.305 53.135 3.475 ;
      RECT 52.72 2.545 52.89 2.715 ;
      RECT 52.69 1.415 52.86 1.585 ;
      RECT 52.625 3.575 52.795 3.745 ;
      RECT 52.35 2.27 52.52 2.44 ;
      RECT 52.23 1.415 52.4 1.585 ;
      RECT 51.82 2.47 51.99 2.64 ;
      RECT 51.77 1.415 51.94 1.585 ;
      RECT 51.31 1.415 51.48 1.585 ;
      RECT 51.3 2.415 51.47 2.585 ;
      RECT 51.095 2.015 51.265 2.185 ;
      RECT 51.095 3.595 51.265 3.765 ;
      RECT 50.85 1.415 51.02 1.585 ;
      RECT 50.785 2.56 50.955 2.73 ;
      RECT 50.39 1.415 50.56 1.585 ;
      RECT 50.375 2.785 50.545 2.955 ;
      RECT 49.93 1.415 50.1 1.585 ;
      RECT 49.665 3.085 49.835 3.255 ;
      RECT 49.52 1.995 49.69 2.165 ;
      RECT 49.47 1.415 49.64 1.585 ;
      RECT 48.03 7.8 48.2 7.97 ;
      RECT 47.68 0.1 47.85 0.27 ;
      RECT 47.68 8.61 47.85 8.78 ;
      RECT 47.66 2.76 47.83 2.93 ;
      RECT 47.66 5.95 47.83 6.12 ;
      RECT 47.04 0.91 47.21 1.08 ;
      RECT 47.04 2.39 47.21 2.56 ;
      RECT 47.04 6.32 47.21 6.49 ;
      RECT 47.04 7.8 47.21 7.97 ;
      RECT 46.69 0.1 46.86 0.27 ;
      RECT 46.69 8.61 46.86 8.78 ;
      RECT 46.67 2.76 46.84 2.93 ;
      RECT 46.67 5.95 46.84 6.12 ;
      RECT 45.99 0.105 46.16 0.275 ;
      RECT 45.99 8.605 46.16 8.775 ;
      RECT 45.68 2.025 45.85 2.195 ;
      RECT 45.68 6.685 45.85 6.855 ;
      RECT 45.31 0.105 45.48 0.275 ;
      RECT 45.31 8.605 45.48 8.775 ;
      RECT 45.25 0.915 45.42 1.085 ;
      RECT 45.25 1.655 45.42 1.825 ;
      RECT 45.25 7.055 45.42 7.225 ;
      RECT 45.25 7.795 45.42 7.965 ;
      RECT 44.875 2.395 45.045 2.565 ;
      RECT 44.875 6.315 45.045 6.485 ;
      RECT 44.63 0.105 44.8 0.275 ;
      RECT 44.63 8.605 44.8 8.775 ;
      RECT 43.95 0.105 44.12 0.275 ;
      RECT 43.95 8.605 44.12 8.775 ;
      RECT 42.49 1.415 42.66 1.585 ;
      RECT 42.05 2.28 42.22 2.45 ;
      RECT 42.03 1.415 42.2 1.585 ;
      RECT 41.655 3.025 41.825 3.195 ;
      RECT 41.57 1.415 41.74 1.585 ;
      RECT 41.545 2.3 41.715 2.47 ;
      RECT 41.11 1.415 41.28 1.585 ;
      RECT 40.725 1.99 40.895 2.16 ;
      RECT 40.65 1.415 40.82 1.585 ;
      RECT 40.41 3.03 40.58 3.2 ;
      RECT 40.365 2.52 40.535 2.69 ;
      RECT 40.355 8.605 40.525 8.775 ;
      RECT 40.19 1.415 40.36 1.585 ;
      RECT 40.045 6.685 40.215 6.855 ;
      RECT 39.94 2.73 40.11 2.9 ;
      RECT 39.75 1.95 39.92 2.12 ;
      RECT 39.73 1.415 39.9 1.585 ;
      RECT 39.7 3.56 39.87 3.73 ;
      RECT 39.675 8.605 39.845 8.775 ;
      RECT 39.615 7.055 39.785 7.225 ;
      RECT 39.615 7.795 39.785 7.965 ;
      RECT 39.365 3 39.535 3.17 ;
      RECT 39.27 1.415 39.44 1.585 ;
      RECT 39.27 2.16 39.44 2.33 ;
      RECT 39.24 6.315 39.41 6.485 ;
      RECT 38.995 8.605 39.165 8.775 ;
      RECT 38.81 1.415 38.98 1.585 ;
      RECT 38.47 3.385 38.64 3.555 ;
      RECT 38.41 2.585 38.58 2.755 ;
      RECT 38.35 1.415 38.52 1.585 ;
      RECT 38.315 8.605 38.485 8.775 ;
      RECT 37.97 2.255 38.14 2.425 ;
      RECT 37.89 1.415 38.06 1.585 ;
      RECT 37.705 3.305 37.875 3.475 ;
      RECT 37.46 2.545 37.63 2.715 ;
      RECT 37.43 1.415 37.6 1.585 ;
      RECT 37.365 3.575 37.535 3.745 ;
      RECT 37.09 2.27 37.26 2.44 ;
      RECT 36.97 1.415 37.14 1.585 ;
      RECT 36.56 2.47 36.73 2.64 ;
      RECT 36.51 1.415 36.68 1.585 ;
      RECT 36.05 1.415 36.22 1.585 ;
      RECT 36.04 2.415 36.21 2.585 ;
      RECT 35.835 2.015 36.005 2.185 ;
      RECT 35.835 3.595 36.005 3.765 ;
      RECT 35.59 1.415 35.76 1.585 ;
      RECT 35.525 2.56 35.695 2.73 ;
      RECT 35.13 1.415 35.3 1.585 ;
      RECT 35.115 2.785 35.285 2.955 ;
      RECT 34.67 1.415 34.84 1.585 ;
      RECT 34.405 3.085 34.575 3.255 ;
      RECT 34.26 1.995 34.43 2.165 ;
      RECT 34.21 1.415 34.38 1.585 ;
      RECT 32.77 7.8 32.94 7.97 ;
      RECT 32.42 0.1 32.59 0.27 ;
      RECT 32.42 8.61 32.59 8.78 ;
      RECT 32.4 2.76 32.57 2.93 ;
      RECT 32.4 5.95 32.57 6.12 ;
      RECT 31.78 0.91 31.95 1.08 ;
      RECT 31.78 2.39 31.95 2.56 ;
      RECT 31.78 6.32 31.95 6.49 ;
      RECT 31.78 7.8 31.95 7.97 ;
      RECT 31.43 0.1 31.6 0.27 ;
      RECT 31.43 8.61 31.6 8.78 ;
      RECT 31.41 2.76 31.58 2.93 ;
      RECT 31.41 5.95 31.58 6.12 ;
      RECT 30.73 0.105 30.9 0.275 ;
      RECT 30.73 8.605 30.9 8.775 ;
      RECT 30.42 2.025 30.59 2.195 ;
      RECT 30.42 6.685 30.59 6.855 ;
      RECT 30.05 0.105 30.22 0.275 ;
      RECT 30.05 8.605 30.22 8.775 ;
      RECT 29.99 0.915 30.16 1.085 ;
      RECT 29.99 1.655 30.16 1.825 ;
      RECT 29.99 7.055 30.16 7.225 ;
      RECT 29.99 7.795 30.16 7.965 ;
      RECT 29.615 2.395 29.785 2.565 ;
      RECT 29.615 6.315 29.785 6.485 ;
      RECT 29.37 0.105 29.54 0.275 ;
      RECT 29.37 8.605 29.54 8.775 ;
      RECT 28.69 0.105 28.86 0.275 ;
      RECT 28.69 8.605 28.86 8.775 ;
      RECT 27.23 1.415 27.4 1.585 ;
      RECT 26.79 2.28 26.96 2.45 ;
      RECT 26.77 1.415 26.94 1.585 ;
      RECT 26.395 3.025 26.565 3.195 ;
      RECT 26.31 1.415 26.48 1.585 ;
      RECT 26.285 2.3 26.455 2.47 ;
      RECT 25.85 1.415 26.02 1.585 ;
      RECT 25.465 1.99 25.635 2.16 ;
      RECT 25.39 1.415 25.56 1.585 ;
      RECT 25.15 3.03 25.32 3.2 ;
      RECT 25.105 2.52 25.275 2.69 ;
      RECT 25.095 8.605 25.265 8.775 ;
      RECT 24.93 1.415 25.1 1.585 ;
      RECT 24.785 6.685 24.955 6.855 ;
      RECT 24.68 2.73 24.85 2.9 ;
      RECT 24.49 1.95 24.66 2.12 ;
      RECT 24.47 1.415 24.64 1.585 ;
      RECT 24.44 3.56 24.61 3.73 ;
      RECT 24.415 8.605 24.585 8.775 ;
      RECT 24.355 7.055 24.525 7.225 ;
      RECT 24.355 7.795 24.525 7.965 ;
      RECT 24.105 3 24.275 3.17 ;
      RECT 24.01 1.415 24.18 1.585 ;
      RECT 24.01 2.16 24.18 2.33 ;
      RECT 23.98 6.315 24.15 6.485 ;
      RECT 23.735 8.605 23.905 8.775 ;
      RECT 23.55 1.415 23.72 1.585 ;
      RECT 23.21 3.385 23.38 3.555 ;
      RECT 23.15 2.585 23.32 2.755 ;
      RECT 23.09 1.415 23.26 1.585 ;
      RECT 23.055 8.605 23.225 8.775 ;
      RECT 22.71 2.255 22.88 2.425 ;
      RECT 22.63 1.415 22.8 1.585 ;
      RECT 22.445 3.305 22.615 3.475 ;
      RECT 22.2 2.545 22.37 2.715 ;
      RECT 22.17 1.415 22.34 1.585 ;
      RECT 22.105 3.575 22.275 3.745 ;
      RECT 21.83 2.27 22 2.44 ;
      RECT 21.71 1.415 21.88 1.585 ;
      RECT 21.3 2.47 21.47 2.64 ;
      RECT 21.25 1.415 21.42 1.585 ;
      RECT 20.79 1.415 20.96 1.585 ;
      RECT 20.78 2.415 20.95 2.585 ;
      RECT 20.575 2.015 20.745 2.185 ;
      RECT 20.575 3.595 20.745 3.765 ;
      RECT 20.33 1.415 20.5 1.585 ;
      RECT 20.265 2.56 20.435 2.73 ;
      RECT 19.87 1.415 20.04 1.585 ;
      RECT 19.855 2.785 20.025 2.955 ;
      RECT 19.41 1.415 19.58 1.585 ;
      RECT 19.145 3.085 19.315 3.255 ;
      RECT 19 1.995 19.17 2.165 ;
      RECT 18.95 1.415 19.12 1.585 ;
      RECT 17.51 7.8 17.68 7.97 ;
      RECT 17.16 0.1 17.33 0.27 ;
      RECT 17.16 8.61 17.33 8.78 ;
      RECT 17.14 2.76 17.31 2.93 ;
      RECT 17.14 5.95 17.31 6.12 ;
      RECT 16.52 0.91 16.69 1.08 ;
      RECT 16.52 2.39 16.69 2.56 ;
      RECT 16.52 6.32 16.69 6.49 ;
      RECT 16.52 7.8 16.69 7.97 ;
      RECT 16.17 0.1 16.34 0.27 ;
      RECT 16.17 8.61 16.34 8.78 ;
      RECT 16.15 2.76 16.32 2.93 ;
      RECT 16.15 5.95 16.32 6.12 ;
      RECT 15.47 0.105 15.64 0.275 ;
      RECT 15.47 8.605 15.64 8.775 ;
      RECT 15.16 2.025 15.33 2.195 ;
      RECT 15.16 6.685 15.33 6.855 ;
      RECT 14.79 0.105 14.96 0.275 ;
      RECT 14.79 8.605 14.96 8.775 ;
      RECT 14.73 0.915 14.9 1.085 ;
      RECT 14.73 1.655 14.9 1.825 ;
      RECT 14.73 7.055 14.9 7.225 ;
      RECT 14.73 7.795 14.9 7.965 ;
      RECT 14.355 2.395 14.525 2.565 ;
      RECT 14.355 6.315 14.525 6.485 ;
      RECT 14.11 0.105 14.28 0.275 ;
      RECT 14.11 8.605 14.28 8.775 ;
      RECT 13.43 0.105 13.6 0.275 ;
      RECT 13.43 8.605 13.6 8.775 ;
      RECT 11.97 1.415 12.14 1.585 ;
      RECT 11.53 2.28 11.7 2.45 ;
      RECT 11.51 1.415 11.68 1.585 ;
      RECT 11.135 3.025 11.305 3.195 ;
      RECT 11.05 1.415 11.22 1.585 ;
      RECT 11.025 2.3 11.195 2.47 ;
      RECT 10.59 1.415 10.76 1.585 ;
      RECT 10.205 1.99 10.375 2.16 ;
      RECT 10.13 1.415 10.3 1.585 ;
      RECT 9.89 3.03 10.06 3.2 ;
      RECT 9.845 2.52 10.015 2.69 ;
      RECT 9.835 8.605 10.005 8.775 ;
      RECT 9.67 1.415 9.84 1.585 ;
      RECT 9.525 6.685 9.695 6.855 ;
      RECT 9.42 2.73 9.59 2.9 ;
      RECT 9.23 1.95 9.4 2.12 ;
      RECT 9.21 1.415 9.38 1.585 ;
      RECT 9.18 3.56 9.35 3.73 ;
      RECT 9.155 8.605 9.325 8.775 ;
      RECT 9.095 7.055 9.265 7.225 ;
      RECT 9.095 7.795 9.265 7.965 ;
      RECT 8.845 3 9.015 3.17 ;
      RECT 8.75 1.415 8.92 1.585 ;
      RECT 8.75 2.16 8.92 2.33 ;
      RECT 8.72 6.315 8.89 6.485 ;
      RECT 8.475 8.605 8.645 8.775 ;
      RECT 8.29 1.415 8.46 1.585 ;
      RECT 7.95 3.385 8.12 3.555 ;
      RECT 7.89 2.585 8.06 2.755 ;
      RECT 7.83 1.415 8 1.585 ;
      RECT 7.795 8.605 7.965 8.775 ;
      RECT 7.45 2.255 7.62 2.425 ;
      RECT 7.37 1.415 7.54 1.585 ;
      RECT 7.185 3.305 7.355 3.475 ;
      RECT 6.94 2.545 7.11 2.715 ;
      RECT 6.91 1.415 7.08 1.585 ;
      RECT 6.845 3.575 7.015 3.745 ;
      RECT 6.57 2.27 6.74 2.44 ;
      RECT 6.45 1.415 6.62 1.585 ;
      RECT 6.04 2.47 6.21 2.64 ;
      RECT 5.99 1.415 6.16 1.585 ;
      RECT 5.53 1.415 5.7 1.585 ;
      RECT 5.52 2.415 5.69 2.585 ;
      RECT 5.315 2.015 5.485 2.185 ;
      RECT 5.315 3.595 5.485 3.765 ;
      RECT 5.07 1.415 5.24 1.585 ;
      RECT 5.005 2.56 5.175 2.73 ;
      RECT 4.61 1.415 4.78 1.585 ;
      RECT 4.595 2.785 4.765 2.955 ;
      RECT 4.15 1.415 4.32 1.585 ;
      RECT 3.885 3.085 4.055 3.255 ;
      RECT 3.74 1.995 3.91 2.165 ;
      RECT 3.69 1.415 3.86 1.585 ;
      RECT 2.34 8.605 2.51 8.775 ;
      RECT 1.66 8.605 1.83 8.775 ;
      RECT 1.6 7.055 1.77 7.225 ;
      RECT 1.6 7.795 1.77 7.965 ;
      RECT 1.225 6.315 1.395 6.485 ;
      RECT 0.98 8.605 1.15 8.775 ;
      RECT 0.3 8.605 0.47 8.775 ;
    LAYER li1 ;
      RECT 72.555 0 72.725 2.085 ;
      RECT 71.615 0 71.785 2.085 ;
      RECT 70.655 0 70.825 2.085 ;
      RECT 68.735 0 68.905 2.085 ;
      RECT 67.775 0 67.945 2.085 ;
      RECT 65.855 0 66.025 2.085 ;
      RECT 57.295 0 57.465 2.085 ;
      RECT 56.355 0 56.525 2.085 ;
      RECT 55.395 0 55.565 2.085 ;
      RECT 53.475 0 53.645 2.085 ;
      RECT 52.515 0 52.685 2.085 ;
      RECT 50.595 0 50.765 2.085 ;
      RECT 42.035 0 42.205 2.085 ;
      RECT 41.095 0 41.265 2.085 ;
      RECT 40.135 0 40.305 2.085 ;
      RECT 38.215 0 38.385 2.085 ;
      RECT 37.255 0 37.425 2.085 ;
      RECT 35.335 0 35.505 2.085 ;
      RECT 26.775 0 26.945 2.085 ;
      RECT 25.835 0 26.005 2.085 ;
      RECT 24.875 0 25.045 2.085 ;
      RECT 22.955 0 23.125 2.085 ;
      RECT 21.995 0 22.165 2.085 ;
      RECT 20.075 0 20.245 2.085 ;
      RECT 11.515 0 11.685 2.085 ;
      RECT 10.575 0 10.745 2.085 ;
      RECT 9.615 0 9.785 2.085 ;
      RECT 7.695 0 7.865 2.085 ;
      RECT 6.735 0 6.905 2.085 ;
      RECT 4.815 0 4.985 2.085 ;
      RECT 69.61 0 69.805 1.595 ;
      RECT 65.855 0 66.13 1.595 ;
      RECT 54.35 0 54.545 1.595 ;
      RECT 50.595 0 50.87 1.595 ;
      RECT 39.09 0 39.285 1.595 ;
      RECT 35.335 0 35.61 1.595 ;
      RECT 23.83 0 24.025 1.595 ;
      RECT 20.075 0 20.35 1.595 ;
      RECT 8.57 0 8.765 1.595 ;
      RECT 4.815 0 5.09 1.595 ;
      RECT 64.585 0 73.325 1.585 ;
      RECT 49.325 0 58.065 1.585 ;
      RECT 34.065 0 42.805 1.585 ;
      RECT 18.805 0 27.545 1.585 ;
      RECT 3.545 0 12.285 1.585 ;
      RECT 74.39 0 74.56 0.935 ;
      RECT 59.13 0 59.3 0.935 ;
      RECT 43.87 0 44.04 0.935 ;
      RECT 28.61 0 28.78 0.935 ;
      RECT 13.35 0 13.52 0.935 ;
      RECT 78.12 0 78.29 0.93 ;
      RECT 77.13 0 77.3 0.93 ;
      RECT 62.86 0 63.03 0.93 ;
      RECT 61.87 0 62.04 0.93 ;
      RECT 47.6 0 47.77 0.93 ;
      RECT 46.61 0 46.78 0.93 ;
      RECT 32.34 0 32.51 0.93 ;
      RECT 31.35 0 31.52 0.93 ;
      RECT 17.08 0 17.25 0.93 ;
      RECT 16.09 0 16.26 0.93 ;
      RECT 78.915 0 79.095 0.305 ;
      RECT 63.655 0 76.965 0.305 ;
      RECT 48.395 0 61.705 0.305 ;
      RECT 33.135 0 46.445 0.305 ;
      RECT 17.875 0 31.185 0.305 ;
      RECT 0 0 15.925 0.305 ;
      RECT 0 0 79.095 0.3 ;
      RECT 0.005 8.575 0.81 8.89 ;
      RECT 0 8.58 79.095 8.88 ;
      RECT 78.915 8.575 79.095 8.88 ;
      RECT 78.12 7.95 78.29 8.88 ;
      RECT 77.13 7.95 77.3 8.88 ;
      RECT 63.655 8.575 76.965 8.88 ;
      RECT 62.86 7.95 63.03 8.88 ;
      RECT 61.87 7.95 62.04 8.88 ;
      RECT 48.395 8.575 61.705 8.88 ;
      RECT 47.6 7.95 47.77 8.88 ;
      RECT 46.61 7.95 46.78 8.88 ;
      RECT 33.135 8.575 46.445 8.88 ;
      RECT 32.34 7.95 32.51 8.88 ;
      RECT 31.35 7.95 31.52 8.88 ;
      RECT 17.875 8.575 31.185 8.88 ;
      RECT 17.08 7.95 17.25 8.88 ;
      RECT 16.09 7.95 16.26 8.88 ;
      RECT 0 8.575 15.925 8.88 ;
      RECT 74.39 7.945 74.56 8.88 ;
      RECT 68.755 7.945 68.925 8.88 ;
      RECT 59.13 7.945 59.3 8.88 ;
      RECT 53.495 7.945 53.665 8.88 ;
      RECT 43.87 7.945 44.04 8.88 ;
      RECT 38.235 7.945 38.405 8.88 ;
      RECT 28.61 7.945 28.78 8.88 ;
      RECT 22.975 7.945 23.145 8.88 ;
      RECT 13.35 7.945 13.52 8.88 ;
      RECT 7.715 7.945 7.885 8.88 ;
      RECT 0.22 8.555 0.47 8.89 ;
      RECT 0.22 7.945 0.39 8.89 ;
      RECT 78.55 5.02 78.72 6.49 ;
      RECT 78.55 6.315 78.725 6.485 ;
      RECT 78.18 1.74 78.35 2.93 ;
      RECT 78.18 1.74 78.65 1.91 ;
      RECT 78.18 6.97 78.65 7.14 ;
      RECT 78.18 5.95 78.35 7.14 ;
      RECT 77.19 1.74 77.36 2.93 ;
      RECT 77.19 1.74 77.66 1.91 ;
      RECT 77.19 6.97 77.66 7.14 ;
      RECT 77.19 5.95 77.36 7.14 ;
      RECT 75.34 2.635 75.51 3.865 ;
      RECT 75.395 0.855 75.565 2.805 ;
      RECT 75.34 0.575 75.51 1.025 ;
      RECT 75.34 7.855 75.51 8.305 ;
      RECT 75.395 6.075 75.565 8.025 ;
      RECT 75.34 5.015 75.51 6.245 ;
      RECT 74.82 0.575 74.99 3.865 ;
      RECT 74.82 2.075 75.225 2.405 ;
      RECT 74.82 1.235 75.225 1.565 ;
      RECT 74.82 5.015 74.99 8.305 ;
      RECT 74.82 7.315 75.225 7.645 ;
      RECT 74.82 6.475 75.225 6.805 ;
      RECT 72.745 3.126 72.75 3.298 ;
      RECT 72.74 3.119 72.745 3.388 ;
      RECT 72.735 3.113 72.74 3.407 ;
      RECT 72.715 3.107 72.735 3.417 ;
      RECT 72.7 3.102 72.715 3.425 ;
      RECT 72.663 3.096 72.7 3.423 ;
      RECT 72.577 3.082 72.663 3.419 ;
      RECT 72.491 3.064 72.577 3.414 ;
      RECT 72.405 3.045 72.491 3.408 ;
      RECT 72.375 3.033 72.405 3.404 ;
      RECT 72.355 3.027 72.375 3.403 ;
      RECT 72.29 3.025 72.355 3.401 ;
      RECT 72.275 3.025 72.29 3.393 ;
      RECT 72.26 3.025 72.275 3.38 ;
      RECT 72.255 3.025 72.26 3.37 ;
      RECT 72.24 3.025 72.255 3.348 ;
      RECT 72.225 3.025 72.24 3.315 ;
      RECT 72.22 3.025 72.225 3.293 ;
      RECT 72.21 3.025 72.22 3.275 ;
      RECT 72.195 3.025 72.21 3.253 ;
      RECT 72.175 3.025 72.195 3.215 ;
      RECT 72.525 2.31 72.56 2.749 ;
      RECT 72.525 2.31 72.565 2.748 ;
      RECT 72.47 2.37 72.565 2.747 ;
      RECT 72.335 2.542 72.565 2.746 ;
      RECT 72.445 2.42 72.565 2.746 ;
      RECT 72.335 2.542 72.59 2.736 ;
      RECT 72.39 2.487 72.67 2.653 ;
      RECT 72.565 2.281 72.57 2.744 ;
      RECT 72.42 2.457 72.71 2.53 ;
      RECT 72.435 2.44 72.565 2.746 ;
      RECT 72.57 2.28 72.74 2.468 ;
      RECT 72.56 2.283 72.74 2.468 ;
      RECT 72.065 2.16 72.235 2.47 ;
      RECT 72.065 2.16 72.24 2.443 ;
      RECT 72.065 2.16 72.245 2.42 ;
      RECT 72.065 2.16 72.255 2.37 ;
      RECT 72.06 2.265 72.255 2.34 ;
      RECT 72.095 1.835 72.265 2.313 ;
      RECT 72.095 1.835 72.28 2.234 ;
      RECT 72.085 2.045 72.28 2.234 ;
      RECT 72.095 1.845 72.29 2.149 ;
      RECT 72.025 2.587 72.03 2.79 ;
      RECT 72.015 2.575 72.025 2.9 ;
      RECT 71.99 2.575 72.015 2.94 ;
      RECT 71.91 2.575 71.99 3.025 ;
      RECT 71.9 2.575 71.91 3.095 ;
      RECT 71.875 2.575 71.9 3.118 ;
      RECT 71.855 2.575 71.875 3.153 ;
      RECT 71.81 2.585 71.855 3.196 ;
      RECT 71.8 2.597 71.81 3.233 ;
      RECT 71.78 2.611 71.8 3.253 ;
      RECT 71.77 2.629 71.78 3.269 ;
      RECT 71.755 2.655 71.77 3.279 ;
      RECT 71.74 2.696 71.755 3.293 ;
      RECT 71.73 2.731 71.74 3.303 ;
      RECT 71.725 2.747 71.73 3.308 ;
      RECT 71.715 2.762 71.725 3.313 ;
      RECT 71.695 2.805 71.715 3.323 ;
      RECT 71.675 2.842 71.695 3.336 ;
      RECT 71.64 2.865 71.675 3.354 ;
      RECT 71.63 2.879 71.64 3.37 ;
      RECT 71.61 2.889 71.63 3.38 ;
      RECT 71.605 2.898 71.61 3.388 ;
      RECT 71.595 2.905 71.605 3.395 ;
      RECT 71.585 2.912 71.595 3.403 ;
      RECT 71.57 2.922 71.585 3.411 ;
      RECT 71.56 2.936 71.57 3.421 ;
      RECT 71.55 2.948 71.56 3.433 ;
      RECT 71.535 2.97 71.55 3.446 ;
      RECT 71.525 2.992 71.535 3.457 ;
      RECT 71.515 3.012 71.525 3.466 ;
      RECT 71.51 3.027 71.515 3.473 ;
      RECT 71.48 3.06 71.51 3.487 ;
      RECT 71.47 3.095 71.48 3.502 ;
      RECT 71.465 3.102 71.47 3.508 ;
      RECT 71.445 3.117 71.465 3.515 ;
      RECT 71.44 3.132 71.445 3.523 ;
      RECT 71.435 3.141 71.44 3.528 ;
      RECT 71.42 3.147 71.435 3.535 ;
      RECT 71.415 3.153 71.42 3.543 ;
      RECT 71.41 3.157 71.415 3.55 ;
      RECT 71.405 3.161 71.41 3.56 ;
      RECT 71.395 3.166 71.405 3.57 ;
      RECT 71.375 3.177 71.395 3.598 ;
      RECT 71.36 3.189 71.375 3.625 ;
      RECT 71.34 3.202 71.36 3.65 ;
      RECT 71.32 3.217 71.34 3.674 ;
      RECT 71.305 3.232 71.32 3.689 ;
      RECT 71.3 3.243 71.305 3.698 ;
      RECT 71.235 3.288 71.3 3.708 ;
      RECT 71.2 3.347 71.235 3.721 ;
      RECT 71.195 3.37 71.2 3.727 ;
      RECT 71.19 3.377 71.195 3.729 ;
      RECT 71.175 3.387 71.19 3.732 ;
      RECT 71.145 3.412 71.175 3.736 ;
      RECT 71.14 3.43 71.145 3.74 ;
      RECT 71.135 3.437 71.14 3.741 ;
      RECT 71.115 3.445 71.135 3.745 ;
      RECT 71.105 3.452 71.115 3.749 ;
      RECT 71.061 3.463 71.105 3.756 ;
      RECT 70.975 3.491 71.061 3.772 ;
      RECT 70.915 3.515 70.975 3.79 ;
      RECT 70.87 3.525 70.915 3.804 ;
      RECT 70.811 3.533 70.87 3.818 ;
      RECT 70.725 3.54 70.811 3.837 ;
      RECT 70.7 3.545 70.725 3.852 ;
      RECT 70.62 3.548 70.7 3.855 ;
      RECT 70.54 3.552 70.62 3.842 ;
      RECT 70.531 3.555 70.54 3.827 ;
      RECT 70.445 3.555 70.531 3.812 ;
      RECT 70.385 3.557 70.445 3.789 ;
      RECT 70.381 3.56 70.385 3.779 ;
      RECT 70.295 3.56 70.381 3.764 ;
      RECT 70.22 3.56 70.295 3.74 ;
      RECT 71.535 2.569 71.545 2.745 ;
      RECT 71.49 2.536 71.535 2.745 ;
      RECT 71.445 2.487 71.49 2.745 ;
      RECT 71.415 2.457 71.445 2.746 ;
      RECT 71.41 2.44 71.415 2.747 ;
      RECT 71.385 2.42 71.41 2.748 ;
      RECT 71.37 2.395 71.385 2.749 ;
      RECT 71.365 2.382 71.37 2.75 ;
      RECT 71.36 2.376 71.365 2.748 ;
      RECT 71.355 2.368 71.36 2.742 ;
      RECT 71.33 2.36 71.355 2.722 ;
      RECT 71.31 2.349 71.33 2.693 ;
      RECT 71.28 2.334 71.31 2.664 ;
      RECT 71.26 2.32 71.28 2.636 ;
      RECT 71.25 2.314 71.26 2.615 ;
      RECT 71.245 2.311 71.25 2.598 ;
      RECT 71.24 2.308 71.245 2.583 ;
      RECT 71.225 2.303 71.24 2.548 ;
      RECT 71.22 2.299 71.225 2.515 ;
      RECT 71.2 2.294 71.22 2.491 ;
      RECT 71.17 2.286 71.2 2.456 ;
      RECT 71.155 2.28 71.17 2.433 ;
      RECT 71.115 2.273 71.155 2.418 ;
      RECT 71.09 2.265 71.115 2.398 ;
      RECT 71.07 2.26 71.09 2.388 ;
      RECT 71.035 2.254 71.07 2.383 ;
      RECT 70.99 2.245 71.035 2.382 ;
      RECT 70.96 2.241 70.99 2.384 ;
      RECT 70.875 2.249 70.96 2.388 ;
      RECT 70.805 2.26 70.875 2.41 ;
      RECT 70.792 2.266 70.805 2.433 ;
      RECT 70.706 2.273 70.792 2.455 ;
      RECT 70.62 2.285 70.706 2.492 ;
      RECT 70.62 2.662 70.63 2.9 ;
      RECT 70.615 2.291 70.62 2.515 ;
      RECT 70.61 2.547 70.62 2.9 ;
      RECT 70.61 2.292 70.615 2.52 ;
      RECT 70.605 2.293 70.61 2.9 ;
      RECT 70.581 2.295 70.605 2.901 ;
      RECT 70.495 2.303 70.581 2.903 ;
      RECT 70.475 2.317 70.495 2.906 ;
      RECT 70.47 2.345 70.475 2.907 ;
      RECT 70.465 2.357 70.47 2.908 ;
      RECT 70.46 2.372 70.465 2.909 ;
      RECT 70.45 2.402 70.46 2.91 ;
      RECT 70.445 2.44 70.45 2.908 ;
      RECT 70.44 2.46 70.445 2.903 ;
      RECT 70.425 2.495 70.44 2.888 ;
      RECT 70.415 2.547 70.425 2.868 ;
      RECT 70.41 2.577 70.415 2.856 ;
      RECT 70.395 2.59 70.41 2.839 ;
      RECT 70.37 2.594 70.395 2.806 ;
      RECT 70.355 2.592 70.37 2.783 ;
      RECT 70.34 2.591 70.355 2.78 ;
      RECT 70.28 2.589 70.34 2.778 ;
      RECT 70.27 2.587 70.28 2.773 ;
      RECT 70.23 2.586 70.27 2.77 ;
      RECT 70.16 2.583 70.23 2.768 ;
      RECT 70.105 2.581 70.16 2.763 ;
      RECT 70.035 2.575 70.105 2.758 ;
      RECT 70.026 2.575 70.035 2.755 ;
      RECT 69.94 2.575 70.026 2.75 ;
      RECT 69.935 2.575 69.94 2.745 ;
      RECT 71.24 1.81 71.415 2.16 ;
      RECT 71.24 1.825 71.425 2.158 ;
      RECT 71.215 1.775 71.36 2.155 ;
      RECT 71.195 1.776 71.36 2.148 ;
      RECT 71.185 1.777 71.37 2.143 ;
      RECT 71.155 1.778 71.37 2.13 ;
      RECT 71.105 1.779 71.37 2.106 ;
      RECT 71.1 1.781 71.37 2.091 ;
      RECT 71.1 1.847 71.43 2.085 ;
      RECT 71.08 1.788 71.385 2.065 ;
      RECT 71.07 1.797 71.395 1.92 ;
      RECT 71.08 1.792 71.395 2.065 ;
      RECT 71.1 1.782 71.385 2.091 ;
      RECT 70.685 3.107 70.855 3.395 ;
      RECT 70.68 3.125 70.865 3.39 ;
      RECT 70.645 3.133 70.93 3.31 ;
      RECT 70.645 3.133 71.016 3.3 ;
      RECT 70.645 3.133 71.07 3.246 ;
      RECT 70.93 3.03 71.1 3.214 ;
      RECT 70.645 3.185 71.105 3.202 ;
      RECT 70.63 3.155 71.1 3.198 ;
      RECT 70.89 3.037 70.93 3.349 ;
      RECT 70.77 3.074 71.1 3.214 ;
      RECT 70.865 3.049 70.89 3.375 ;
      RECT 70.855 3.056 71.1 3.214 ;
      RECT 70.986 2.52 71.055 2.779 ;
      RECT 70.986 2.575 71.06 2.778 ;
      RECT 70.9 2.575 71.06 2.777 ;
      RECT 70.895 2.575 71.065 2.77 ;
      RECT 70.885 2.52 71.055 2.765 ;
      RECT 70.265 1.819 70.44 2.12 ;
      RECT 70.25 1.807 70.265 2.105 ;
      RECT 70.22 1.806 70.25 2.058 ;
      RECT 70.22 1.824 70.445 2.053 ;
      RECT 70.205 1.808 70.265 2.018 ;
      RECT 70.2 1.83 70.455 1.918 ;
      RECT 70.2 1.813 70.351 1.918 ;
      RECT 70.2 1.815 70.355 1.918 ;
      RECT 70.205 1.811 70.351 2.018 ;
      RECT 70.31 3.047 70.315 3.395 ;
      RECT 70.3 3.037 70.31 3.401 ;
      RECT 70.265 3.027 70.3 3.403 ;
      RECT 70.227 3.022 70.265 3.407 ;
      RECT 70.141 3.015 70.227 3.414 ;
      RECT 70.055 3.005 70.141 3.424 ;
      RECT 70.01 3 70.055 3.432 ;
      RECT 70.006 3 70.01 3.436 ;
      RECT 69.92 3 70.006 3.443 ;
      RECT 69.905 3 69.92 3.443 ;
      RECT 69.895 2.998 69.905 3.415 ;
      RECT 69.885 2.994 69.895 3.358 ;
      RECT 69.865 2.988 69.885 3.29 ;
      RECT 69.86 2.984 69.865 3.238 ;
      RECT 69.85 2.983 69.86 3.205 ;
      RECT 69.8 2.981 69.85 3.19 ;
      RECT 69.775 2.979 69.8 3.185 ;
      RECT 69.732 2.977 69.775 3.181 ;
      RECT 69.646 2.973 69.732 3.169 ;
      RECT 69.56 2.968 69.646 3.153 ;
      RECT 69.53 2.965 69.56 3.14 ;
      RECT 69.505 2.964 69.53 3.128 ;
      RECT 69.5 2.964 69.505 3.118 ;
      RECT 69.46 2.963 69.5 3.11 ;
      RECT 69.445 2.962 69.46 3.103 ;
      RECT 69.395 2.961 69.445 3.095 ;
      RECT 69.393 2.96 69.395 3.09 ;
      RECT 69.307 2.958 69.393 3.09 ;
      RECT 69.221 2.953 69.307 3.09 ;
      RECT 69.135 2.949 69.221 3.09 ;
      RECT 69.086 2.945 69.135 3.088 ;
      RECT 69 2.942 69.086 3.083 ;
      RECT 68.977 2.939 69 3.079 ;
      RECT 68.891 2.936 68.977 3.074 ;
      RECT 68.805 2.932 68.891 3.065 ;
      RECT 68.78 2.925 68.805 3.06 ;
      RECT 68.72 2.89 68.78 3.057 ;
      RECT 68.7 2.815 68.72 3.054 ;
      RECT 68.695 2.757 68.7 3.053 ;
      RECT 68.67 2.697 68.695 3.052 ;
      RECT 68.595 2.575 68.67 3.048 ;
      RECT 68.585 2.575 68.595 3.04 ;
      RECT 68.57 2.575 68.585 3.03 ;
      RECT 68.555 2.575 68.57 3 ;
      RECT 68.54 2.575 68.555 2.945 ;
      RECT 68.525 2.575 68.54 2.883 ;
      RECT 68.5 2.575 68.525 2.808 ;
      RECT 68.495 2.575 68.5 2.758 ;
      RECT 69.84 2.12 69.86 2.429 ;
      RECT 69.826 2.122 69.875 2.426 ;
      RECT 69.826 2.127 69.895 2.417 ;
      RECT 69.74 2.125 69.875 2.411 ;
      RECT 69.74 2.133 69.93 2.394 ;
      RECT 69.705 2.135 69.93 2.393 ;
      RECT 69.675 2.143 69.93 2.384 ;
      RECT 69.665 2.148 69.95 2.37 ;
      RECT 69.705 2.138 69.95 2.37 ;
      RECT 69.705 2.141 69.96 2.358 ;
      RECT 69.675 2.143 69.97 2.345 ;
      RECT 69.675 2.147 69.98 2.288 ;
      RECT 69.665 2.152 69.985 2.203 ;
      RECT 69.826 2.12 69.86 2.426 ;
      RECT 69.705 7.855 69.875 8.305 ;
      RECT 69.76 6.075 69.93 8.025 ;
      RECT 69.705 5.015 69.875 6.245 ;
      RECT 69.265 2.223 69.27 2.435 ;
      RECT 69.14 2.22 69.155 2.435 ;
      RECT 68.605 2.25 68.675 2.435 ;
      RECT 68.49 2.25 68.525 2.43 ;
      RECT 69.611 2.552 69.63 2.746 ;
      RECT 69.525 2.507 69.611 2.747 ;
      RECT 69.515 2.46 69.525 2.749 ;
      RECT 69.51 2.44 69.515 2.75 ;
      RECT 69.49 2.405 69.51 2.751 ;
      RECT 69.475 2.355 69.49 2.752 ;
      RECT 69.455 2.292 69.475 2.753 ;
      RECT 69.445 2.255 69.455 2.754 ;
      RECT 69.43 2.244 69.445 2.755 ;
      RECT 69.425 2.236 69.43 2.753 ;
      RECT 69.415 2.235 69.425 2.745 ;
      RECT 69.385 2.232 69.415 2.724 ;
      RECT 69.31 2.227 69.385 2.669 ;
      RECT 69.295 2.223 69.31 2.615 ;
      RECT 69.285 2.223 69.295 2.51 ;
      RECT 69.27 2.223 69.285 2.443 ;
      RECT 69.255 2.223 69.265 2.433 ;
      RECT 69.2 2.222 69.255 2.43 ;
      RECT 69.155 2.22 69.2 2.433 ;
      RECT 69.127 2.22 69.14 2.436 ;
      RECT 69.041 2.224 69.127 2.438 ;
      RECT 68.955 2.23 69.041 2.443 ;
      RECT 68.935 2.234 68.955 2.445 ;
      RECT 68.933 2.235 68.935 2.444 ;
      RECT 68.847 2.237 68.933 2.443 ;
      RECT 68.761 2.242 68.847 2.44 ;
      RECT 68.675 2.247 68.761 2.437 ;
      RECT 68.525 2.25 68.605 2.433 ;
      RECT 69.185 5.015 69.355 8.305 ;
      RECT 69.185 7.315 69.59 7.645 ;
      RECT 69.185 6.475 69.59 6.805 ;
      RECT 69.301 3.225 69.35 3.559 ;
      RECT 69.301 3.225 69.355 3.558 ;
      RECT 69.215 3.225 69.355 3.557 ;
      RECT 68.99 3.333 69.36 3.555 ;
      RECT 69.215 3.225 69.385 3.548 ;
      RECT 69.185 3.237 69.39 3.539 ;
      RECT 69.17 3.255 69.395 3.536 ;
      RECT 68.985 3.339 69.395 3.463 ;
      RECT 68.98 3.346 69.395 3.423 ;
      RECT 68.995 3.312 69.395 3.536 ;
      RECT 69.156 3.258 69.36 3.555 ;
      RECT 69.07 3.278 69.395 3.536 ;
      RECT 69.17 3.252 69.39 3.539 ;
      RECT 68.94 2.576 69.13 2.77 ;
      RECT 68.935 2.578 69.13 2.769 ;
      RECT 68.93 2.582 69.145 2.766 ;
      RECT 68.945 2.575 69.145 2.766 ;
      RECT 68.93 2.685 69.15 2.761 ;
      RECT 68.225 3.185 68.316 3.483 ;
      RECT 68.22 3.187 68.395 3.478 ;
      RECT 68.225 3.185 68.395 3.478 ;
      RECT 68.22 3.191 68.415 3.476 ;
      RECT 68.22 3.246 68.455 3.475 ;
      RECT 68.22 3.281 68.47 3.469 ;
      RECT 68.22 3.315 68.48 3.459 ;
      RECT 68.21 3.195 68.415 3.31 ;
      RECT 68.21 3.215 68.43 3.31 ;
      RECT 68.21 3.198 68.42 3.31 ;
      RECT 68.435 1.966 68.44 2.028 ;
      RECT 68.43 1.888 68.435 2.051 ;
      RECT 68.425 1.845 68.43 2.062 ;
      RECT 68.42 1.835 68.425 2.074 ;
      RECT 68.415 1.835 68.42 2.083 ;
      RECT 68.39 1.835 68.415 2.115 ;
      RECT 68.385 1.835 68.39 2.148 ;
      RECT 68.37 1.835 68.385 2.173 ;
      RECT 68.36 1.835 68.37 2.2 ;
      RECT 68.355 1.835 68.36 2.213 ;
      RECT 68.35 1.835 68.355 2.228 ;
      RECT 68.34 1.835 68.35 2.243 ;
      RECT 68.335 1.835 68.34 2.263 ;
      RECT 68.31 1.835 68.335 2.298 ;
      RECT 68.265 1.835 68.31 2.343 ;
      RECT 68.255 1.835 68.265 2.356 ;
      RECT 68.17 1.92 68.255 2.363 ;
      RECT 68.135 2.042 68.17 2.372 ;
      RECT 68.13 2.082 68.135 2.376 ;
      RECT 68.11 2.105 68.13 2.378 ;
      RECT 68.105 2.135 68.11 2.381 ;
      RECT 68.095 2.147 68.105 2.382 ;
      RECT 68.05 2.17 68.095 2.387 ;
      RECT 68.01 2.2 68.05 2.395 ;
      RECT 67.975 2.212 68.01 2.401 ;
      RECT 67.97 2.217 67.975 2.405 ;
      RECT 67.9 2.227 67.97 2.412 ;
      RECT 67.86 2.237 67.9 2.422 ;
      RECT 67.84 2.242 67.86 2.428 ;
      RECT 67.83 2.246 67.84 2.433 ;
      RECT 67.825 2.249 67.83 2.436 ;
      RECT 67.815 2.25 67.825 2.437 ;
      RECT 67.79 2.252 67.815 2.441 ;
      RECT 67.78 2.257 67.79 2.444 ;
      RECT 67.735 2.265 67.78 2.445 ;
      RECT 67.61 2.27 67.735 2.445 ;
      RECT 68.165 2.567 68.185 2.749 ;
      RECT 68.116 2.552 68.165 2.748 ;
      RECT 68.03 2.567 68.185 2.746 ;
      RECT 68.015 2.567 68.185 2.745 ;
      RECT 67.98 2.545 68.15 2.73 ;
      RECT 68.05 3.565 68.065 3.774 ;
      RECT 68.05 3.573 68.07 3.773 ;
      RECT 67.995 3.573 68.07 3.772 ;
      RECT 67.975 3.577 68.075 3.77 ;
      RECT 67.955 3.527 67.995 3.769 ;
      RECT 67.9 3.585 68.08 3.767 ;
      RECT 67.865 3.542 67.995 3.765 ;
      RECT 67.861 3.545 68.05 3.764 ;
      RECT 67.775 3.553 68.05 3.762 ;
      RECT 67.775 3.597 68.085 3.755 ;
      RECT 67.765 3.69 68.085 3.753 ;
      RECT 67.775 3.609 68.09 3.738 ;
      RECT 67.775 3.63 68.105 3.708 ;
      RECT 67.775 3.657 68.11 3.678 ;
      RECT 67.9 3.535 67.995 3.767 ;
      RECT 67.53 2.58 67.535 3.118 ;
      RECT 67.335 2.91 67.34 3.105 ;
      RECT 65.635 2.575 65.65 2.955 ;
      RECT 67.7 2.575 67.705 2.745 ;
      RECT 67.695 2.575 67.7 2.755 ;
      RECT 67.69 2.575 67.695 2.768 ;
      RECT 67.665 2.575 67.69 2.81 ;
      RECT 67.64 2.575 67.665 2.883 ;
      RECT 67.625 2.575 67.64 2.935 ;
      RECT 67.62 2.575 67.625 2.965 ;
      RECT 67.595 2.575 67.62 3.005 ;
      RECT 67.58 2.575 67.595 3.06 ;
      RECT 67.575 2.575 67.58 3.093 ;
      RECT 67.55 2.575 67.575 3.113 ;
      RECT 67.535 2.575 67.55 3.119 ;
      RECT 67.465 2.61 67.53 3.115 ;
      RECT 67.415 2.665 67.465 3.11 ;
      RECT 67.405 2.697 67.415 3.108 ;
      RECT 67.4 2.722 67.405 3.108 ;
      RECT 67.38 2.795 67.4 3.108 ;
      RECT 67.37 2.875 67.38 3.107 ;
      RECT 67.355 2.905 67.37 3.107 ;
      RECT 67.34 2.91 67.355 3.106 ;
      RECT 67.28 2.912 67.335 3.103 ;
      RECT 67.25 2.917 67.28 3.099 ;
      RECT 67.248 2.92 67.25 3.098 ;
      RECT 67.162 2.922 67.248 3.095 ;
      RECT 67.076 2.928 67.162 3.089 ;
      RECT 66.99 2.933 67.076 3.083 ;
      RECT 66.917 2.938 66.99 3.084 ;
      RECT 66.831 2.944 66.917 3.092 ;
      RECT 66.745 2.95 66.831 3.101 ;
      RECT 66.725 2.954 66.745 3.106 ;
      RECT 66.678 2.956 66.725 3.109 ;
      RECT 66.592 2.961 66.678 3.115 ;
      RECT 66.506 2.966 66.592 3.124 ;
      RECT 66.42 2.972 66.506 3.132 ;
      RECT 66.335 2.97 66.42 3.141 ;
      RECT 66.331 2.965 66.335 3.145 ;
      RECT 66.245 2.96 66.331 3.137 ;
      RECT 66.181 2.951 66.245 3.125 ;
      RECT 66.095 2.942 66.181 3.112 ;
      RECT 66.071 2.935 66.095 3.103 ;
      RECT 65.985 2.929 66.071 3.09 ;
      RECT 65.945 2.922 65.985 3.076 ;
      RECT 65.94 2.912 65.945 3.072 ;
      RECT 65.93 2.9 65.94 3.071 ;
      RECT 65.91 2.87 65.93 3.068 ;
      RECT 65.855 2.79 65.91 3.062 ;
      RECT 65.835 2.709 65.855 3.057 ;
      RECT 65.815 2.667 65.835 3.053 ;
      RECT 65.79 2.62 65.815 3.047 ;
      RECT 65.785 2.595 65.79 3.044 ;
      RECT 65.75 2.575 65.785 3.039 ;
      RECT 65.741 2.575 65.75 3.032 ;
      RECT 65.655 2.575 65.741 3.002 ;
      RECT 65.65 2.575 65.655 2.965 ;
      RECT 65.615 2.575 65.635 2.887 ;
      RECT 65.61 2.617 65.615 2.852 ;
      RECT 65.605 2.692 65.61 2.808 ;
      RECT 67.055 2.497 67.23 2.745 ;
      RECT 67.055 2.497 67.235 2.743 ;
      RECT 67.05 2.529 67.235 2.703 ;
      RECT 67.08 2.47 67.25 2.69 ;
      RECT 67.045 2.547 67.25 2.623 ;
      RECT 66.355 2.01 66.525 2.185 ;
      RECT 66.355 2.01 66.697 2.177 ;
      RECT 66.355 2.01 66.78 2.171 ;
      RECT 66.355 2.01 66.815 2.167 ;
      RECT 66.355 2.01 66.835 2.166 ;
      RECT 66.355 2.01 66.921 2.162 ;
      RECT 66.815 1.835 66.985 2.157 ;
      RECT 66.39 1.942 67.015 2.155 ;
      RECT 66.38 1.997 67.02 2.153 ;
      RECT 66.355 2.033 67.03 2.148 ;
      RECT 66.355 2.06 67.035 2.078 ;
      RECT 66.42 1.885 66.995 2.155 ;
      RECT 66.611 1.87 66.995 2.155 ;
      RECT 66.445 1.873 66.995 2.155 ;
      RECT 66.525 1.871 66.611 2.182 ;
      RECT 66.611 1.868 66.99 2.155 ;
      RECT 66.795 1.845 66.99 2.155 ;
      RECT 66.697 1.866 66.99 2.155 ;
      RECT 66.78 1.86 66.795 2.168 ;
      RECT 66.93 3.225 66.935 3.425 ;
      RECT 66.395 3.29 66.44 3.425 ;
      RECT 66.965 3.225 66.985 3.398 ;
      RECT 66.935 3.225 66.965 3.413 ;
      RECT 66.87 3.225 66.93 3.45 ;
      RECT 66.855 3.225 66.87 3.48 ;
      RECT 66.84 3.225 66.855 3.493 ;
      RECT 66.82 3.225 66.84 3.508 ;
      RECT 66.815 3.225 66.82 3.517 ;
      RECT 66.805 3.229 66.815 3.522 ;
      RECT 66.79 3.239 66.805 3.533 ;
      RECT 66.765 3.255 66.79 3.543 ;
      RECT 66.755 3.269 66.765 3.545 ;
      RECT 66.735 3.281 66.755 3.542 ;
      RECT 66.705 3.302 66.735 3.536 ;
      RECT 66.695 3.314 66.705 3.531 ;
      RECT 66.685 3.312 66.695 3.528 ;
      RECT 66.67 3.311 66.685 3.523 ;
      RECT 66.665 3.31 66.67 3.518 ;
      RECT 66.63 3.308 66.665 3.508 ;
      RECT 66.61 3.305 66.63 3.49 ;
      RECT 66.6 3.303 66.61 3.485 ;
      RECT 66.59 3.302 66.6 3.48 ;
      RECT 66.555 3.3 66.59 3.468 ;
      RECT 66.5 3.296 66.555 3.448 ;
      RECT 66.49 3.294 66.5 3.433 ;
      RECT 66.485 3.294 66.49 3.428 ;
      RECT 66.44 3.292 66.485 3.425 ;
      RECT 66.345 3.29 66.395 3.429 ;
      RECT 66.335 3.291 66.345 3.434 ;
      RECT 66.275 3.298 66.335 3.448 ;
      RECT 66.25 3.306 66.275 3.468 ;
      RECT 66.24 3.31 66.25 3.48 ;
      RECT 66.235 3.311 66.24 3.485 ;
      RECT 66.22 3.313 66.235 3.488 ;
      RECT 66.205 3.315 66.22 3.493 ;
      RECT 66.2 3.315 66.205 3.496 ;
      RECT 66.155 3.32 66.2 3.507 ;
      RECT 66.15 3.324 66.155 3.519 ;
      RECT 66.125 3.32 66.15 3.523 ;
      RECT 66.115 3.316 66.125 3.527 ;
      RECT 66.105 3.315 66.115 3.531 ;
      RECT 66.09 3.305 66.105 3.537 ;
      RECT 66.085 3.293 66.09 3.541 ;
      RECT 66.08 3.29 66.085 3.542 ;
      RECT 66.075 3.287 66.08 3.544 ;
      RECT 66.06 3.275 66.075 3.543 ;
      RECT 66.045 3.257 66.06 3.54 ;
      RECT 66.025 3.236 66.045 3.533 ;
      RECT 65.96 3.225 66.025 3.505 ;
      RECT 65.956 3.225 65.96 3.484 ;
      RECT 65.87 3.225 65.956 3.454 ;
      RECT 65.855 3.225 65.87 3.41 ;
      RECT 66.43 2.325 66.435 2.56 ;
      RECT 65.56 2.241 65.565 2.445 ;
      RECT 66.14 2.27 66.145 2.425 ;
      RECT 66.06 2.25 66.065 2.425 ;
      RECT 66.73 2.392 66.745 2.745 ;
      RECT 66.656 2.377 66.73 2.745 ;
      RECT 66.57 2.36 66.656 2.745 ;
      RECT 66.56 2.35 66.57 2.743 ;
      RECT 66.555 2.348 66.56 2.738 ;
      RECT 66.54 2.346 66.555 2.724 ;
      RECT 66.47 2.338 66.54 2.664 ;
      RECT 66.45 2.329 66.47 2.598 ;
      RECT 66.445 2.326 66.45 2.578 ;
      RECT 66.435 2.325 66.445 2.568 ;
      RECT 66.425 2.325 66.43 2.552 ;
      RECT 66.415 2.324 66.425 2.542 ;
      RECT 66.405 2.322 66.415 2.53 ;
      RECT 66.39 2.319 66.405 2.51 ;
      RECT 66.38 2.317 66.39 2.495 ;
      RECT 66.36 2.314 66.38 2.483 ;
      RECT 66.355 2.312 66.36 2.473 ;
      RECT 66.33 2.31 66.355 2.46 ;
      RECT 66.3 2.305 66.33 2.445 ;
      RECT 66.22 2.296 66.3 2.436 ;
      RECT 66.175 2.285 66.22 2.429 ;
      RECT 66.155 2.276 66.175 2.426 ;
      RECT 66.145 2.271 66.155 2.425 ;
      RECT 66.1 2.265 66.14 2.425 ;
      RECT 66.085 2.257 66.1 2.425 ;
      RECT 66.065 2.252 66.085 2.425 ;
      RECT 66.045 2.249 66.06 2.425 ;
      RECT 65.962 2.248 66.045 2.424 ;
      RECT 65.876 2.247 65.962 2.42 ;
      RECT 65.79 2.245 65.876 2.417 ;
      RECT 65.737 2.244 65.79 2.419 ;
      RECT 65.651 2.243 65.737 2.428 ;
      RECT 65.565 2.242 65.651 2.44 ;
      RECT 65.545 2.241 65.56 2.448 ;
      RECT 65.465 2.24 65.545 2.46 ;
      RECT 65.44 2.24 65.465 2.473 ;
      RECT 65.415 2.24 65.44 2.488 ;
      RECT 65.41 2.24 65.415 2.51 ;
      RECT 65.405 2.24 65.41 2.528 ;
      RECT 65.4 2.24 65.405 2.545 ;
      RECT 65.395 2.24 65.4 2.558 ;
      RECT 65.39 2.24 65.395 2.568 ;
      RECT 65.35 2.24 65.39 2.653 ;
      RECT 65.335 2.24 65.35 2.738 ;
      RECT 65.325 2.241 65.335 2.75 ;
      RECT 65.29 2.246 65.325 2.755 ;
      RECT 65.25 2.255 65.29 2.755 ;
      RECT 65.235 2.265 65.25 2.755 ;
      RECT 65.23 2.275 65.235 2.755 ;
      RECT 65.21 2.302 65.23 2.755 ;
      RECT 65.16 2.385 65.21 2.755 ;
      RECT 65.155 2.447 65.16 2.755 ;
      RECT 65.145 2.46 65.155 2.755 ;
      RECT 65.135 2.482 65.145 2.755 ;
      RECT 65.125 2.507 65.135 2.75 ;
      RECT 65.12 2.545 65.125 2.743 ;
      RECT 65.11 2.655 65.12 2.738 ;
      RECT 66.505 3.576 66.52 3.835 ;
      RECT 66.505 3.591 66.525 3.834 ;
      RECT 66.421 3.591 66.525 3.832 ;
      RECT 66.421 3.605 66.53 3.831 ;
      RECT 66.335 3.647 66.535 3.828 ;
      RECT 66.33 3.59 66.52 3.823 ;
      RECT 66.33 3.661 66.54 3.82 ;
      RECT 66.325 3.692 66.54 3.818 ;
      RECT 66.33 3.689 66.555 3.808 ;
      RECT 66.325 3.735 66.57 3.793 ;
      RECT 66.325 3.763 66.575 3.778 ;
      RECT 66.335 3.565 66.505 3.828 ;
      RECT 66.095 2.575 66.265 2.745 ;
      RECT 66.06 2.575 66.265 2.74 ;
      RECT 66.05 2.575 66.265 2.733 ;
      RECT 66.045 2.56 66.215 2.73 ;
      RECT 64.875 3.097 65.14 3.54 ;
      RECT 64.87 3.068 65.085 3.538 ;
      RECT 64.865 3.222 65.145 3.533 ;
      RECT 64.87 3.117 65.145 3.533 ;
      RECT 64.87 3.128 65.155 3.52 ;
      RECT 64.87 3.075 65.115 3.538 ;
      RECT 64.875 3.062 65.085 3.54 ;
      RECT 64.875 3.06 65.035 3.54 ;
      RECT 64.976 3.052 65.035 3.54 ;
      RECT 64.89 3.053 65.035 3.54 ;
      RECT 64.976 3.051 65.025 3.54 ;
      RECT 64.78 1.866 64.955 2.165 ;
      RECT 64.83 1.828 64.955 2.165 ;
      RECT 64.815 1.83 65.041 2.157 ;
      RECT 64.815 1.833 65.08 2.144 ;
      RECT 64.815 1.834 65.09 2.13 ;
      RECT 64.77 1.885 65.09 2.12 ;
      RECT 64.815 1.835 65.095 2.115 ;
      RECT 64.77 2.045 65.1 2.105 ;
      RECT 64.755 1.905 65.095 2.045 ;
      RECT 64.75 1.921 65.095 1.985 ;
      RECT 64.795 1.845 65.095 2.115 ;
      RECT 64.83 1.826 64.916 2.165 ;
      RECT 63.29 5.02 63.46 6.49 ;
      RECT 63.29 6.315 63.465 6.485 ;
      RECT 62.92 1.74 63.09 2.93 ;
      RECT 62.92 1.74 63.39 1.91 ;
      RECT 62.92 6.97 63.39 7.14 ;
      RECT 62.92 5.95 63.09 7.14 ;
      RECT 61.93 1.74 62.1 2.93 ;
      RECT 61.93 1.74 62.4 1.91 ;
      RECT 61.93 6.97 62.4 7.14 ;
      RECT 61.93 5.95 62.1 7.14 ;
      RECT 60.08 2.635 60.25 3.865 ;
      RECT 60.135 0.855 60.305 2.805 ;
      RECT 60.08 0.575 60.25 1.025 ;
      RECT 60.08 7.855 60.25 8.305 ;
      RECT 60.135 6.075 60.305 8.025 ;
      RECT 60.08 5.015 60.25 6.245 ;
      RECT 59.56 0.575 59.73 3.865 ;
      RECT 59.56 2.075 59.965 2.405 ;
      RECT 59.56 1.235 59.965 1.565 ;
      RECT 59.56 5.015 59.73 8.305 ;
      RECT 59.56 7.315 59.965 7.645 ;
      RECT 59.56 6.475 59.965 6.805 ;
      RECT 57.485 3.126 57.49 3.298 ;
      RECT 57.48 3.119 57.485 3.388 ;
      RECT 57.475 3.113 57.48 3.407 ;
      RECT 57.455 3.107 57.475 3.417 ;
      RECT 57.44 3.102 57.455 3.425 ;
      RECT 57.403 3.096 57.44 3.423 ;
      RECT 57.317 3.082 57.403 3.419 ;
      RECT 57.231 3.064 57.317 3.414 ;
      RECT 57.145 3.045 57.231 3.408 ;
      RECT 57.115 3.033 57.145 3.404 ;
      RECT 57.095 3.027 57.115 3.403 ;
      RECT 57.03 3.025 57.095 3.401 ;
      RECT 57.015 3.025 57.03 3.393 ;
      RECT 57 3.025 57.015 3.38 ;
      RECT 56.995 3.025 57 3.37 ;
      RECT 56.98 3.025 56.995 3.348 ;
      RECT 56.965 3.025 56.98 3.315 ;
      RECT 56.96 3.025 56.965 3.293 ;
      RECT 56.95 3.025 56.96 3.275 ;
      RECT 56.935 3.025 56.95 3.253 ;
      RECT 56.915 3.025 56.935 3.215 ;
      RECT 57.265 2.31 57.3 2.749 ;
      RECT 57.265 2.31 57.305 2.748 ;
      RECT 57.21 2.37 57.305 2.747 ;
      RECT 57.075 2.542 57.305 2.746 ;
      RECT 57.185 2.42 57.305 2.746 ;
      RECT 57.075 2.542 57.33 2.736 ;
      RECT 57.13 2.487 57.41 2.653 ;
      RECT 57.305 2.281 57.31 2.744 ;
      RECT 57.16 2.457 57.45 2.53 ;
      RECT 57.175 2.44 57.305 2.746 ;
      RECT 57.31 2.28 57.48 2.468 ;
      RECT 57.3 2.283 57.48 2.468 ;
      RECT 56.805 2.16 56.975 2.47 ;
      RECT 56.805 2.16 56.98 2.443 ;
      RECT 56.805 2.16 56.985 2.42 ;
      RECT 56.805 2.16 56.995 2.37 ;
      RECT 56.8 2.265 56.995 2.34 ;
      RECT 56.835 1.835 57.005 2.313 ;
      RECT 56.835 1.835 57.02 2.234 ;
      RECT 56.825 2.045 57.02 2.234 ;
      RECT 56.835 1.845 57.03 2.149 ;
      RECT 56.765 2.587 56.77 2.79 ;
      RECT 56.755 2.575 56.765 2.9 ;
      RECT 56.73 2.575 56.755 2.94 ;
      RECT 56.65 2.575 56.73 3.025 ;
      RECT 56.64 2.575 56.65 3.095 ;
      RECT 56.615 2.575 56.64 3.118 ;
      RECT 56.595 2.575 56.615 3.153 ;
      RECT 56.55 2.585 56.595 3.196 ;
      RECT 56.54 2.597 56.55 3.233 ;
      RECT 56.52 2.611 56.54 3.253 ;
      RECT 56.51 2.629 56.52 3.269 ;
      RECT 56.495 2.655 56.51 3.279 ;
      RECT 56.48 2.696 56.495 3.293 ;
      RECT 56.47 2.731 56.48 3.303 ;
      RECT 56.465 2.747 56.47 3.308 ;
      RECT 56.455 2.762 56.465 3.313 ;
      RECT 56.435 2.805 56.455 3.323 ;
      RECT 56.415 2.842 56.435 3.336 ;
      RECT 56.38 2.865 56.415 3.354 ;
      RECT 56.37 2.879 56.38 3.37 ;
      RECT 56.35 2.889 56.37 3.38 ;
      RECT 56.345 2.898 56.35 3.388 ;
      RECT 56.335 2.905 56.345 3.395 ;
      RECT 56.325 2.912 56.335 3.403 ;
      RECT 56.31 2.922 56.325 3.411 ;
      RECT 56.3 2.936 56.31 3.421 ;
      RECT 56.29 2.948 56.3 3.433 ;
      RECT 56.275 2.97 56.29 3.446 ;
      RECT 56.265 2.992 56.275 3.457 ;
      RECT 56.255 3.012 56.265 3.466 ;
      RECT 56.25 3.027 56.255 3.473 ;
      RECT 56.22 3.06 56.25 3.487 ;
      RECT 56.21 3.095 56.22 3.502 ;
      RECT 56.205 3.102 56.21 3.508 ;
      RECT 56.185 3.117 56.205 3.515 ;
      RECT 56.18 3.132 56.185 3.523 ;
      RECT 56.175 3.141 56.18 3.528 ;
      RECT 56.16 3.147 56.175 3.535 ;
      RECT 56.155 3.153 56.16 3.543 ;
      RECT 56.15 3.157 56.155 3.55 ;
      RECT 56.145 3.161 56.15 3.56 ;
      RECT 56.135 3.166 56.145 3.57 ;
      RECT 56.115 3.177 56.135 3.598 ;
      RECT 56.1 3.189 56.115 3.625 ;
      RECT 56.08 3.202 56.1 3.65 ;
      RECT 56.06 3.217 56.08 3.674 ;
      RECT 56.045 3.232 56.06 3.689 ;
      RECT 56.04 3.243 56.045 3.698 ;
      RECT 55.975 3.288 56.04 3.708 ;
      RECT 55.94 3.347 55.975 3.721 ;
      RECT 55.935 3.37 55.94 3.727 ;
      RECT 55.93 3.377 55.935 3.729 ;
      RECT 55.915 3.387 55.93 3.732 ;
      RECT 55.885 3.412 55.915 3.736 ;
      RECT 55.88 3.43 55.885 3.74 ;
      RECT 55.875 3.437 55.88 3.741 ;
      RECT 55.855 3.445 55.875 3.745 ;
      RECT 55.845 3.452 55.855 3.749 ;
      RECT 55.801 3.463 55.845 3.756 ;
      RECT 55.715 3.491 55.801 3.772 ;
      RECT 55.655 3.515 55.715 3.79 ;
      RECT 55.61 3.525 55.655 3.804 ;
      RECT 55.551 3.533 55.61 3.818 ;
      RECT 55.465 3.54 55.551 3.837 ;
      RECT 55.44 3.545 55.465 3.852 ;
      RECT 55.36 3.548 55.44 3.855 ;
      RECT 55.28 3.552 55.36 3.842 ;
      RECT 55.271 3.555 55.28 3.827 ;
      RECT 55.185 3.555 55.271 3.812 ;
      RECT 55.125 3.557 55.185 3.789 ;
      RECT 55.121 3.56 55.125 3.779 ;
      RECT 55.035 3.56 55.121 3.764 ;
      RECT 54.96 3.56 55.035 3.74 ;
      RECT 56.275 2.569 56.285 2.745 ;
      RECT 56.23 2.536 56.275 2.745 ;
      RECT 56.185 2.487 56.23 2.745 ;
      RECT 56.155 2.457 56.185 2.746 ;
      RECT 56.15 2.44 56.155 2.747 ;
      RECT 56.125 2.42 56.15 2.748 ;
      RECT 56.11 2.395 56.125 2.749 ;
      RECT 56.105 2.382 56.11 2.75 ;
      RECT 56.1 2.376 56.105 2.748 ;
      RECT 56.095 2.368 56.1 2.742 ;
      RECT 56.07 2.36 56.095 2.722 ;
      RECT 56.05 2.349 56.07 2.693 ;
      RECT 56.02 2.334 56.05 2.664 ;
      RECT 56 2.32 56.02 2.636 ;
      RECT 55.99 2.314 56 2.615 ;
      RECT 55.985 2.311 55.99 2.598 ;
      RECT 55.98 2.308 55.985 2.583 ;
      RECT 55.965 2.303 55.98 2.548 ;
      RECT 55.96 2.299 55.965 2.515 ;
      RECT 55.94 2.294 55.96 2.491 ;
      RECT 55.91 2.286 55.94 2.456 ;
      RECT 55.895 2.28 55.91 2.433 ;
      RECT 55.855 2.273 55.895 2.418 ;
      RECT 55.83 2.265 55.855 2.398 ;
      RECT 55.81 2.26 55.83 2.388 ;
      RECT 55.775 2.254 55.81 2.383 ;
      RECT 55.73 2.245 55.775 2.382 ;
      RECT 55.7 2.241 55.73 2.384 ;
      RECT 55.615 2.249 55.7 2.388 ;
      RECT 55.545 2.26 55.615 2.41 ;
      RECT 55.532 2.266 55.545 2.433 ;
      RECT 55.446 2.273 55.532 2.455 ;
      RECT 55.36 2.285 55.446 2.492 ;
      RECT 55.36 2.662 55.37 2.9 ;
      RECT 55.355 2.291 55.36 2.515 ;
      RECT 55.35 2.547 55.36 2.9 ;
      RECT 55.35 2.292 55.355 2.52 ;
      RECT 55.345 2.293 55.35 2.9 ;
      RECT 55.321 2.295 55.345 2.901 ;
      RECT 55.235 2.303 55.321 2.903 ;
      RECT 55.215 2.317 55.235 2.906 ;
      RECT 55.21 2.345 55.215 2.907 ;
      RECT 55.205 2.357 55.21 2.908 ;
      RECT 55.2 2.372 55.205 2.909 ;
      RECT 55.19 2.402 55.2 2.91 ;
      RECT 55.185 2.44 55.19 2.908 ;
      RECT 55.18 2.46 55.185 2.903 ;
      RECT 55.165 2.495 55.18 2.888 ;
      RECT 55.155 2.547 55.165 2.868 ;
      RECT 55.15 2.577 55.155 2.856 ;
      RECT 55.135 2.59 55.15 2.839 ;
      RECT 55.11 2.594 55.135 2.806 ;
      RECT 55.095 2.592 55.11 2.783 ;
      RECT 55.08 2.591 55.095 2.78 ;
      RECT 55.02 2.589 55.08 2.778 ;
      RECT 55.01 2.587 55.02 2.773 ;
      RECT 54.97 2.586 55.01 2.77 ;
      RECT 54.9 2.583 54.97 2.768 ;
      RECT 54.845 2.581 54.9 2.763 ;
      RECT 54.775 2.575 54.845 2.758 ;
      RECT 54.766 2.575 54.775 2.755 ;
      RECT 54.68 2.575 54.766 2.75 ;
      RECT 54.675 2.575 54.68 2.745 ;
      RECT 55.98 1.81 56.155 2.16 ;
      RECT 55.98 1.825 56.165 2.158 ;
      RECT 55.955 1.775 56.1 2.155 ;
      RECT 55.935 1.776 56.1 2.148 ;
      RECT 55.925 1.777 56.11 2.143 ;
      RECT 55.895 1.778 56.11 2.13 ;
      RECT 55.845 1.779 56.11 2.106 ;
      RECT 55.84 1.781 56.11 2.091 ;
      RECT 55.84 1.847 56.17 2.085 ;
      RECT 55.82 1.788 56.125 2.065 ;
      RECT 55.81 1.797 56.135 1.92 ;
      RECT 55.82 1.792 56.135 2.065 ;
      RECT 55.84 1.782 56.125 2.091 ;
      RECT 55.425 3.107 55.595 3.395 ;
      RECT 55.42 3.125 55.605 3.39 ;
      RECT 55.385 3.133 55.67 3.31 ;
      RECT 55.385 3.133 55.756 3.3 ;
      RECT 55.385 3.133 55.81 3.246 ;
      RECT 55.67 3.03 55.84 3.214 ;
      RECT 55.385 3.185 55.845 3.202 ;
      RECT 55.37 3.155 55.84 3.198 ;
      RECT 55.63 3.037 55.67 3.349 ;
      RECT 55.51 3.074 55.84 3.214 ;
      RECT 55.605 3.049 55.63 3.375 ;
      RECT 55.595 3.056 55.84 3.214 ;
      RECT 55.726 2.52 55.795 2.779 ;
      RECT 55.726 2.575 55.8 2.778 ;
      RECT 55.64 2.575 55.8 2.777 ;
      RECT 55.635 2.575 55.805 2.77 ;
      RECT 55.625 2.52 55.795 2.765 ;
      RECT 55.005 1.819 55.18 2.12 ;
      RECT 54.99 1.807 55.005 2.105 ;
      RECT 54.96 1.806 54.99 2.058 ;
      RECT 54.96 1.824 55.185 2.053 ;
      RECT 54.945 1.808 55.005 2.018 ;
      RECT 54.94 1.83 55.195 1.918 ;
      RECT 54.94 1.813 55.091 1.918 ;
      RECT 54.94 1.815 55.095 1.918 ;
      RECT 54.945 1.811 55.091 2.018 ;
      RECT 55.05 3.047 55.055 3.395 ;
      RECT 55.04 3.037 55.05 3.401 ;
      RECT 55.005 3.027 55.04 3.403 ;
      RECT 54.967 3.022 55.005 3.407 ;
      RECT 54.881 3.015 54.967 3.414 ;
      RECT 54.795 3.005 54.881 3.424 ;
      RECT 54.75 3 54.795 3.432 ;
      RECT 54.746 3 54.75 3.436 ;
      RECT 54.66 3 54.746 3.443 ;
      RECT 54.645 3 54.66 3.443 ;
      RECT 54.635 2.998 54.645 3.415 ;
      RECT 54.625 2.994 54.635 3.358 ;
      RECT 54.605 2.988 54.625 3.29 ;
      RECT 54.6 2.984 54.605 3.238 ;
      RECT 54.59 2.983 54.6 3.205 ;
      RECT 54.54 2.981 54.59 3.19 ;
      RECT 54.515 2.979 54.54 3.185 ;
      RECT 54.472 2.977 54.515 3.181 ;
      RECT 54.386 2.973 54.472 3.169 ;
      RECT 54.3 2.968 54.386 3.153 ;
      RECT 54.27 2.965 54.3 3.14 ;
      RECT 54.245 2.964 54.27 3.128 ;
      RECT 54.24 2.964 54.245 3.118 ;
      RECT 54.2 2.963 54.24 3.11 ;
      RECT 54.185 2.962 54.2 3.103 ;
      RECT 54.135 2.961 54.185 3.095 ;
      RECT 54.133 2.96 54.135 3.09 ;
      RECT 54.047 2.958 54.133 3.09 ;
      RECT 53.961 2.953 54.047 3.09 ;
      RECT 53.875 2.949 53.961 3.09 ;
      RECT 53.826 2.945 53.875 3.088 ;
      RECT 53.74 2.942 53.826 3.083 ;
      RECT 53.717 2.939 53.74 3.079 ;
      RECT 53.631 2.936 53.717 3.074 ;
      RECT 53.545 2.932 53.631 3.065 ;
      RECT 53.52 2.925 53.545 3.06 ;
      RECT 53.46 2.89 53.52 3.057 ;
      RECT 53.44 2.815 53.46 3.054 ;
      RECT 53.435 2.757 53.44 3.053 ;
      RECT 53.41 2.697 53.435 3.052 ;
      RECT 53.335 2.575 53.41 3.048 ;
      RECT 53.325 2.575 53.335 3.04 ;
      RECT 53.31 2.575 53.325 3.03 ;
      RECT 53.295 2.575 53.31 3 ;
      RECT 53.28 2.575 53.295 2.945 ;
      RECT 53.265 2.575 53.28 2.883 ;
      RECT 53.24 2.575 53.265 2.808 ;
      RECT 53.235 2.575 53.24 2.758 ;
      RECT 54.58 2.12 54.6 2.429 ;
      RECT 54.566 2.122 54.615 2.426 ;
      RECT 54.566 2.127 54.635 2.417 ;
      RECT 54.48 2.125 54.615 2.411 ;
      RECT 54.48 2.133 54.67 2.394 ;
      RECT 54.445 2.135 54.67 2.393 ;
      RECT 54.415 2.143 54.67 2.384 ;
      RECT 54.405 2.148 54.69 2.37 ;
      RECT 54.445 2.138 54.69 2.37 ;
      RECT 54.445 2.141 54.7 2.358 ;
      RECT 54.415 2.143 54.71 2.345 ;
      RECT 54.415 2.147 54.72 2.288 ;
      RECT 54.405 2.152 54.725 2.203 ;
      RECT 54.566 2.12 54.6 2.426 ;
      RECT 54.445 7.855 54.615 8.305 ;
      RECT 54.5 6.075 54.67 8.025 ;
      RECT 54.445 5.015 54.615 6.245 ;
      RECT 54.005 2.223 54.01 2.435 ;
      RECT 53.88 2.22 53.895 2.435 ;
      RECT 53.345 2.25 53.415 2.435 ;
      RECT 53.23 2.25 53.265 2.43 ;
      RECT 54.351 2.552 54.37 2.746 ;
      RECT 54.265 2.507 54.351 2.747 ;
      RECT 54.255 2.46 54.265 2.749 ;
      RECT 54.25 2.44 54.255 2.75 ;
      RECT 54.23 2.405 54.25 2.751 ;
      RECT 54.215 2.355 54.23 2.752 ;
      RECT 54.195 2.292 54.215 2.753 ;
      RECT 54.185 2.255 54.195 2.754 ;
      RECT 54.17 2.244 54.185 2.755 ;
      RECT 54.165 2.236 54.17 2.753 ;
      RECT 54.155 2.235 54.165 2.745 ;
      RECT 54.125 2.232 54.155 2.724 ;
      RECT 54.05 2.227 54.125 2.669 ;
      RECT 54.035 2.223 54.05 2.615 ;
      RECT 54.025 2.223 54.035 2.51 ;
      RECT 54.01 2.223 54.025 2.443 ;
      RECT 53.995 2.223 54.005 2.433 ;
      RECT 53.94 2.222 53.995 2.43 ;
      RECT 53.895 2.22 53.94 2.433 ;
      RECT 53.867 2.22 53.88 2.436 ;
      RECT 53.781 2.224 53.867 2.438 ;
      RECT 53.695 2.23 53.781 2.443 ;
      RECT 53.675 2.234 53.695 2.445 ;
      RECT 53.673 2.235 53.675 2.444 ;
      RECT 53.587 2.237 53.673 2.443 ;
      RECT 53.501 2.242 53.587 2.44 ;
      RECT 53.415 2.247 53.501 2.437 ;
      RECT 53.265 2.25 53.345 2.433 ;
      RECT 53.925 5.015 54.095 8.305 ;
      RECT 53.925 7.315 54.33 7.645 ;
      RECT 53.925 6.475 54.33 6.805 ;
      RECT 54.041 3.225 54.09 3.559 ;
      RECT 54.041 3.225 54.095 3.558 ;
      RECT 53.955 3.225 54.095 3.557 ;
      RECT 53.73 3.333 54.1 3.555 ;
      RECT 53.955 3.225 54.125 3.548 ;
      RECT 53.925 3.237 54.13 3.539 ;
      RECT 53.91 3.255 54.135 3.536 ;
      RECT 53.725 3.339 54.135 3.463 ;
      RECT 53.72 3.346 54.135 3.423 ;
      RECT 53.735 3.312 54.135 3.536 ;
      RECT 53.896 3.258 54.1 3.555 ;
      RECT 53.81 3.278 54.135 3.536 ;
      RECT 53.91 3.252 54.13 3.539 ;
      RECT 53.68 2.576 53.87 2.77 ;
      RECT 53.675 2.578 53.87 2.769 ;
      RECT 53.67 2.582 53.885 2.766 ;
      RECT 53.685 2.575 53.885 2.766 ;
      RECT 53.67 2.685 53.89 2.761 ;
      RECT 52.965 3.185 53.056 3.483 ;
      RECT 52.96 3.187 53.135 3.478 ;
      RECT 52.965 3.185 53.135 3.478 ;
      RECT 52.96 3.191 53.155 3.476 ;
      RECT 52.96 3.246 53.195 3.475 ;
      RECT 52.96 3.281 53.21 3.469 ;
      RECT 52.96 3.315 53.22 3.459 ;
      RECT 52.95 3.195 53.155 3.31 ;
      RECT 52.95 3.215 53.17 3.31 ;
      RECT 52.95 3.198 53.16 3.31 ;
      RECT 53.175 1.966 53.18 2.028 ;
      RECT 53.17 1.888 53.175 2.051 ;
      RECT 53.165 1.845 53.17 2.062 ;
      RECT 53.16 1.835 53.165 2.074 ;
      RECT 53.155 1.835 53.16 2.083 ;
      RECT 53.13 1.835 53.155 2.115 ;
      RECT 53.125 1.835 53.13 2.148 ;
      RECT 53.11 1.835 53.125 2.173 ;
      RECT 53.1 1.835 53.11 2.2 ;
      RECT 53.095 1.835 53.1 2.213 ;
      RECT 53.09 1.835 53.095 2.228 ;
      RECT 53.08 1.835 53.09 2.243 ;
      RECT 53.075 1.835 53.08 2.263 ;
      RECT 53.05 1.835 53.075 2.298 ;
      RECT 53.005 1.835 53.05 2.343 ;
      RECT 52.995 1.835 53.005 2.356 ;
      RECT 52.91 1.92 52.995 2.363 ;
      RECT 52.875 2.042 52.91 2.372 ;
      RECT 52.87 2.082 52.875 2.376 ;
      RECT 52.85 2.105 52.87 2.378 ;
      RECT 52.845 2.135 52.85 2.381 ;
      RECT 52.835 2.147 52.845 2.382 ;
      RECT 52.79 2.17 52.835 2.387 ;
      RECT 52.75 2.2 52.79 2.395 ;
      RECT 52.715 2.212 52.75 2.401 ;
      RECT 52.71 2.217 52.715 2.405 ;
      RECT 52.64 2.227 52.71 2.412 ;
      RECT 52.6 2.237 52.64 2.422 ;
      RECT 52.58 2.242 52.6 2.428 ;
      RECT 52.57 2.246 52.58 2.433 ;
      RECT 52.565 2.249 52.57 2.436 ;
      RECT 52.555 2.25 52.565 2.437 ;
      RECT 52.53 2.252 52.555 2.441 ;
      RECT 52.52 2.257 52.53 2.444 ;
      RECT 52.475 2.265 52.52 2.445 ;
      RECT 52.35 2.27 52.475 2.445 ;
      RECT 52.905 2.567 52.925 2.749 ;
      RECT 52.856 2.552 52.905 2.748 ;
      RECT 52.77 2.567 52.925 2.746 ;
      RECT 52.755 2.567 52.925 2.745 ;
      RECT 52.72 2.545 52.89 2.73 ;
      RECT 52.79 3.565 52.805 3.774 ;
      RECT 52.79 3.573 52.81 3.773 ;
      RECT 52.735 3.573 52.81 3.772 ;
      RECT 52.715 3.577 52.815 3.77 ;
      RECT 52.695 3.527 52.735 3.769 ;
      RECT 52.64 3.585 52.82 3.767 ;
      RECT 52.605 3.542 52.735 3.765 ;
      RECT 52.601 3.545 52.79 3.764 ;
      RECT 52.515 3.553 52.79 3.762 ;
      RECT 52.515 3.597 52.825 3.755 ;
      RECT 52.505 3.69 52.825 3.753 ;
      RECT 52.515 3.609 52.83 3.738 ;
      RECT 52.515 3.63 52.845 3.708 ;
      RECT 52.515 3.657 52.85 3.678 ;
      RECT 52.64 3.535 52.735 3.767 ;
      RECT 52.27 2.58 52.275 3.118 ;
      RECT 52.075 2.91 52.08 3.105 ;
      RECT 50.375 2.575 50.39 2.955 ;
      RECT 52.44 2.575 52.445 2.745 ;
      RECT 52.435 2.575 52.44 2.755 ;
      RECT 52.43 2.575 52.435 2.768 ;
      RECT 52.405 2.575 52.43 2.81 ;
      RECT 52.38 2.575 52.405 2.883 ;
      RECT 52.365 2.575 52.38 2.935 ;
      RECT 52.36 2.575 52.365 2.965 ;
      RECT 52.335 2.575 52.36 3.005 ;
      RECT 52.32 2.575 52.335 3.06 ;
      RECT 52.315 2.575 52.32 3.093 ;
      RECT 52.29 2.575 52.315 3.113 ;
      RECT 52.275 2.575 52.29 3.119 ;
      RECT 52.205 2.61 52.27 3.115 ;
      RECT 52.155 2.665 52.205 3.11 ;
      RECT 52.145 2.697 52.155 3.108 ;
      RECT 52.14 2.722 52.145 3.108 ;
      RECT 52.12 2.795 52.14 3.108 ;
      RECT 52.11 2.875 52.12 3.107 ;
      RECT 52.095 2.905 52.11 3.107 ;
      RECT 52.08 2.91 52.095 3.106 ;
      RECT 52.02 2.912 52.075 3.103 ;
      RECT 51.99 2.917 52.02 3.099 ;
      RECT 51.988 2.92 51.99 3.098 ;
      RECT 51.902 2.922 51.988 3.095 ;
      RECT 51.816 2.928 51.902 3.089 ;
      RECT 51.73 2.933 51.816 3.083 ;
      RECT 51.657 2.938 51.73 3.084 ;
      RECT 51.571 2.944 51.657 3.092 ;
      RECT 51.485 2.95 51.571 3.101 ;
      RECT 51.465 2.954 51.485 3.106 ;
      RECT 51.418 2.956 51.465 3.109 ;
      RECT 51.332 2.961 51.418 3.115 ;
      RECT 51.246 2.966 51.332 3.124 ;
      RECT 51.16 2.972 51.246 3.132 ;
      RECT 51.075 2.97 51.16 3.141 ;
      RECT 51.071 2.965 51.075 3.145 ;
      RECT 50.985 2.96 51.071 3.137 ;
      RECT 50.921 2.951 50.985 3.125 ;
      RECT 50.835 2.942 50.921 3.112 ;
      RECT 50.811 2.935 50.835 3.103 ;
      RECT 50.725 2.929 50.811 3.09 ;
      RECT 50.685 2.922 50.725 3.076 ;
      RECT 50.68 2.912 50.685 3.072 ;
      RECT 50.67 2.9 50.68 3.071 ;
      RECT 50.65 2.87 50.67 3.068 ;
      RECT 50.595 2.79 50.65 3.062 ;
      RECT 50.575 2.709 50.595 3.057 ;
      RECT 50.555 2.667 50.575 3.053 ;
      RECT 50.53 2.62 50.555 3.047 ;
      RECT 50.525 2.595 50.53 3.044 ;
      RECT 50.49 2.575 50.525 3.039 ;
      RECT 50.481 2.575 50.49 3.032 ;
      RECT 50.395 2.575 50.481 3.002 ;
      RECT 50.39 2.575 50.395 2.965 ;
      RECT 50.355 2.575 50.375 2.887 ;
      RECT 50.35 2.617 50.355 2.852 ;
      RECT 50.345 2.692 50.35 2.808 ;
      RECT 51.795 2.497 51.97 2.745 ;
      RECT 51.795 2.497 51.975 2.743 ;
      RECT 51.79 2.529 51.975 2.703 ;
      RECT 51.82 2.47 51.99 2.69 ;
      RECT 51.785 2.547 51.99 2.623 ;
      RECT 51.095 2.01 51.265 2.185 ;
      RECT 51.095 2.01 51.437 2.177 ;
      RECT 51.095 2.01 51.52 2.171 ;
      RECT 51.095 2.01 51.555 2.167 ;
      RECT 51.095 2.01 51.575 2.166 ;
      RECT 51.095 2.01 51.661 2.162 ;
      RECT 51.555 1.835 51.725 2.157 ;
      RECT 51.13 1.942 51.755 2.155 ;
      RECT 51.12 1.997 51.76 2.153 ;
      RECT 51.095 2.033 51.77 2.148 ;
      RECT 51.095 2.06 51.775 2.078 ;
      RECT 51.16 1.885 51.735 2.155 ;
      RECT 51.351 1.87 51.735 2.155 ;
      RECT 51.185 1.873 51.735 2.155 ;
      RECT 51.265 1.871 51.351 2.182 ;
      RECT 51.351 1.868 51.73 2.155 ;
      RECT 51.535 1.845 51.73 2.155 ;
      RECT 51.437 1.866 51.73 2.155 ;
      RECT 51.52 1.86 51.535 2.168 ;
      RECT 51.67 3.225 51.675 3.425 ;
      RECT 51.135 3.29 51.18 3.425 ;
      RECT 51.705 3.225 51.725 3.398 ;
      RECT 51.675 3.225 51.705 3.413 ;
      RECT 51.61 3.225 51.67 3.45 ;
      RECT 51.595 3.225 51.61 3.48 ;
      RECT 51.58 3.225 51.595 3.493 ;
      RECT 51.56 3.225 51.58 3.508 ;
      RECT 51.555 3.225 51.56 3.517 ;
      RECT 51.545 3.229 51.555 3.522 ;
      RECT 51.53 3.239 51.545 3.533 ;
      RECT 51.505 3.255 51.53 3.543 ;
      RECT 51.495 3.269 51.505 3.545 ;
      RECT 51.475 3.281 51.495 3.542 ;
      RECT 51.445 3.302 51.475 3.536 ;
      RECT 51.435 3.314 51.445 3.531 ;
      RECT 51.425 3.312 51.435 3.528 ;
      RECT 51.41 3.311 51.425 3.523 ;
      RECT 51.405 3.31 51.41 3.518 ;
      RECT 51.37 3.308 51.405 3.508 ;
      RECT 51.35 3.305 51.37 3.49 ;
      RECT 51.34 3.303 51.35 3.485 ;
      RECT 51.33 3.302 51.34 3.48 ;
      RECT 51.295 3.3 51.33 3.468 ;
      RECT 51.24 3.296 51.295 3.448 ;
      RECT 51.23 3.294 51.24 3.433 ;
      RECT 51.225 3.294 51.23 3.428 ;
      RECT 51.18 3.292 51.225 3.425 ;
      RECT 51.085 3.29 51.135 3.429 ;
      RECT 51.075 3.291 51.085 3.434 ;
      RECT 51.015 3.298 51.075 3.448 ;
      RECT 50.99 3.306 51.015 3.468 ;
      RECT 50.98 3.31 50.99 3.48 ;
      RECT 50.975 3.311 50.98 3.485 ;
      RECT 50.96 3.313 50.975 3.488 ;
      RECT 50.945 3.315 50.96 3.493 ;
      RECT 50.94 3.315 50.945 3.496 ;
      RECT 50.895 3.32 50.94 3.507 ;
      RECT 50.89 3.324 50.895 3.519 ;
      RECT 50.865 3.32 50.89 3.523 ;
      RECT 50.855 3.316 50.865 3.527 ;
      RECT 50.845 3.315 50.855 3.531 ;
      RECT 50.83 3.305 50.845 3.537 ;
      RECT 50.825 3.293 50.83 3.541 ;
      RECT 50.82 3.29 50.825 3.542 ;
      RECT 50.815 3.287 50.82 3.544 ;
      RECT 50.8 3.275 50.815 3.543 ;
      RECT 50.785 3.257 50.8 3.54 ;
      RECT 50.765 3.236 50.785 3.533 ;
      RECT 50.7 3.225 50.765 3.505 ;
      RECT 50.696 3.225 50.7 3.484 ;
      RECT 50.61 3.225 50.696 3.454 ;
      RECT 50.595 3.225 50.61 3.41 ;
      RECT 51.17 2.325 51.175 2.56 ;
      RECT 50.3 2.241 50.305 2.445 ;
      RECT 50.88 2.27 50.885 2.425 ;
      RECT 50.8 2.25 50.805 2.425 ;
      RECT 51.47 2.392 51.485 2.745 ;
      RECT 51.396 2.377 51.47 2.745 ;
      RECT 51.31 2.36 51.396 2.745 ;
      RECT 51.3 2.35 51.31 2.743 ;
      RECT 51.295 2.348 51.3 2.738 ;
      RECT 51.28 2.346 51.295 2.724 ;
      RECT 51.21 2.338 51.28 2.664 ;
      RECT 51.19 2.329 51.21 2.598 ;
      RECT 51.185 2.326 51.19 2.578 ;
      RECT 51.175 2.325 51.185 2.568 ;
      RECT 51.165 2.325 51.17 2.552 ;
      RECT 51.155 2.324 51.165 2.542 ;
      RECT 51.145 2.322 51.155 2.53 ;
      RECT 51.13 2.319 51.145 2.51 ;
      RECT 51.12 2.317 51.13 2.495 ;
      RECT 51.1 2.314 51.12 2.483 ;
      RECT 51.095 2.312 51.1 2.473 ;
      RECT 51.07 2.31 51.095 2.46 ;
      RECT 51.04 2.305 51.07 2.445 ;
      RECT 50.96 2.296 51.04 2.436 ;
      RECT 50.915 2.285 50.96 2.429 ;
      RECT 50.895 2.276 50.915 2.426 ;
      RECT 50.885 2.271 50.895 2.425 ;
      RECT 50.84 2.265 50.88 2.425 ;
      RECT 50.825 2.257 50.84 2.425 ;
      RECT 50.805 2.252 50.825 2.425 ;
      RECT 50.785 2.249 50.8 2.425 ;
      RECT 50.702 2.248 50.785 2.424 ;
      RECT 50.616 2.247 50.702 2.42 ;
      RECT 50.53 2.245 50.616 2.417 ;
      RECT 50.477 2.244 50.53 2.419 ;
      RECT 50.391 2.243 50.477 2.428 ;
      RECT 50.305 2.242 50.391 2.44 ;
      RECT 50.285 2.241 50.3 2.448 ;
      RECT 50.205 2.24 50.285 2.46 ;
      RECT 50.18 2.24 50.205 2.473 ;
      RECT 50.155 2.24 50.18 2.488 ;
      RECT 50.15 2.24 50.155 2.51 ;
      RECT 50.145 2.24 50.15 2.528 ;
      RECT 50.14 2.24 50.145 2.545 ;
      RECT 50.135 2.24 50.14 2.558 ;
      RECT 50.13 2.24 50.135 2.568 ;
      RECT 50.09 2.24 50.13 2.653 ;
      RECT 50.075 2.24 50.09 2.738 ;
      RECT 50.065 2.241 50.075 2.75 ;
      RECT 50.03 2.246 50.065 2.755 ;
      RECT 49.99 2.255 50.03 2.755 ;
      RECT 49.975 2.265 49.99 2.755 ;
      RECT 49.97 2.275 49.975 2.755 ;
      RECT 49.95 2.302 49.97 2.755 ;
      RECT 49.9 2.385 49.95 2.755 ;
      RECT 49.895 2.447 49.9 2.755 ;
      RECT 49.885 2.46 49.895 2.755 ;
      RECT 49.875 2.482 49.885 2.755 ;
      RECT 49.865 2.507 49.875 2.75 ;
      RECT 49.86 2.545 49.865 2.743 ;
      RECT 49.85 2.655 49.86 2.738 ;
      RECT 51.245 3.576 51.26 3.835 ;
      RECT 51.245 3.591 51.265 3.834 ;
      RECT 51.161 3.591 51.265 3.832 ;
      RECT 51.161 3.605 51.27 3.831 ;
      RECT 51.075 3.647 51.275 3.828 ;
      RECT 51.07 3.59 51.26 3.823 ;
      RECT 51.07 3.661 51.28 3.82 ;
      RECT 51.065 3.692 51.28 3.818 ;
      RECT 51.07 3.689 51.295 3.808 ;
      RECT 51.065 3.735 51.31 3.793 ;
      RECT 51.065 3.763 51.315 3.778 ;
      RECT 51.075 3.565 51.245 3.828 ;
      RECT 50.835 2.575 51.005 2.745 ;
      RECT 50.8 2.575 51.005 2.74 ;
      RECT 50.79 2.575 51.005 2.733 ;
      RECT 50.785 2.56 50.955 2.73 ;
      RECT 49.615 3.097 49.88 3.54 ;
      RECT 49.61 3.068 49.825 3.538 ;
      RECT 49.605 3.222 49.885 3.533 ;
      RECT 49.61 3.117 49.885 3.533 ;
      RECT 49.61 3.128 49.895 3.52 ;
      RECT 49.61 3.075 49.855 3.538 ;
      RECT 49.615 3.062 49.825 3.54 ;
      RECT 49.615 3.06 49.775 3.54 ;
      RECT 49.716 3.052 49.775 3.54 ;
      RECT 49.63 3.053 49.775 3.54 ;
      RECT 49.716 3.051 49.765 3.54 ;
      RECT 49.52 1.866 49.695 2.165 ;
      RECT 49.57 1.828 49.695 2.165 ;
      RECT 49.555 1.83 49.781 2.157 ;
      RECT 49.555 1.833 49.82 2.144 ;
      RECT 49.555 1.834 49.83 2.13 ;
      RECT 49.51 1.885 49.83 2.12 ;
      RECT 49.555 1.835 49.835 2.115 ;
      RECT 49.51 2.045 49.84 2.105 ;
      RECT 49.495 1.905 49.835 2.045 ;
      RECT 49.49 1.921 49.835 1.985 ;
      RECT 49.535 1.845 49.835 2.115 ;
      RECT 49.57 1.826 49.656 2.165 ;
      RECT 48.03 5.02 48.2 6.49 ;
      RECT 48.03 6.315 48.205 6.485 ;
      RECT 47.66 1.74 47.83 2.93 ;
      RECT 47.66 1.74 48.13 1.91 ;
      RECT 47.66 6.97 48.13 7.14 ;
      RECT 47.66 5.95 47.83 7.14 ;
      RECT 46.67 1.74 46.84 2.93 ;
      RECT 46.67 1.74 47.14 1.91 ;
      RECT 46.67 6.97 47.14 7.14 ;
      RECT 46.67 5.95 46.84 7.14 ;
      RECT 44.82 2.635 44.99 3.865 ;
      RECT 44.875 0.855 45.045 2.805 ;
      RECT 44.82 0.575 44.99 1.025 ;
      RECT 44.82 7.855 44.99 8.305 ;
      RECT 44.875 6.075 45.045 8.025 ;
      RECT 44.82 5.015 44.99 6.245 ;
      RECT 44.3 0.575 44.47 3.865 ;
      RECT 44.3 2.075 44.705 2.405 ;
      RECT 44.3 1.235 44.705 1.565 ;
      RECT 44.3 5.015 44.47 8.305 ;
      RECT 44.3 7.315 44.705 7.645 ;
      RECT 44.3 6.475 44.705 6.805 ;
      RECT 42.225 3.126 42.23 3.298 ;
      RECT 42.22 3.119 42.225 3.388 ;
      RECT 42.215 3.113 42.22 3.407 ;
      RECT 42.195 3.107 42.215 3.417 ;
      RECT 42.18 3.102 42.195 3.425 ;
      RECT 42.143 3.096 42.18 3.423 ;
      RECT 42.057 3.082 42.143 3.419 ;
      RECT 41.971 3.064 42.057 3.414 ;
      RECT 41.885 3.045 41.971 3.408 ;
      RECT 41.855 3.033 41.885 3.404 ;
      RECT 41.835 3.027 41.855 3.403 ;
      RECT 41.77 3.025 41.835 3.401 ;
      RECT 41.755 3.025 41.77 3.393 ;
      RECT 41.74 3.025 41.755 3.38 ;
      RECT 41.735 3.025 41.74 3.37 ;
      RECT 41.72 3.025 41.735 3.348 ;
      RECT 41.705 3.025 41.72 3.315 ;
      RECT 41.7 3.025 41.705 3.293 ;
      RECT 41.69 3.025 41.7 3.275 ;
      RECT 41.675 3.025 41.69 3.253 ;
      RECT 41.655 3.025 41.675 3.215 ;
      RECT 42.005 2.31 42.04 2.749 ;
      RECT 42.005 2.31 42.045 2.748 ;
      RECT 41.95 2.37 42.045 2.747 ;
      RECT 41.815 2.542 42.045 2.746 ;
      RECT 41.925 2.42 42.045 2.746 ;
      RECT 41.815 2.542 42.07 2.736 ;
      RECT 41.87 2.487 42.15 2.653 ;
      RECT 42.045 2.281 42.05 2.744 ;
      RECT 41.9 2.457 42.19 2.53 ;
      RECT 41.915 2.44 42.045 2.746 ;
      RECT 42.05 2.28 42.22 2.468 ;
      RECT 42.04 2.283 42.22 2.468 ;
      RECT 41.545 2.16 41.715 2.47 ;
      RECT 41.545 2.16 41.72 2.443 ;
      RECT 41.545 2.16 41.725 2.42 ;
      RECT 41.545 2.16 41.735 2.37 ;
      RECT 41.54 2.265 41.735 2.34 ;
      RECT 41.575 1.835 41.745 2.313 ;
      RECT 41.575 1.835 41.76 2.234 ;
      RECT 41.565 2.045 41.76 2.234 ;
      RECT 41.575 1.845 41.77 2.149 ;
      RECT 41.505 2.587 41.51 2.79 ;
      RECT 41.495 2.575 41.505 2.9 ;
      RECT 41.47 2.575 41.495 2.94 ;
      RECT 41.39 2.575 41.47 3.025 ;
      RECT 41.38 2.575 41.39 3.095 ;
      RECT 41.355 2.575 41.38 3.118 ;
      RECT 41.335 2.575 41.355 3.153 ;
      RECT 41.29 2.585 41.335 3.196 ;
      RECT 41.28 2.597 41.29 3.233 ;
      RECT 41.26 2.611 41.28 3.253 ;
      RECT 41.25 2.629 41.26 3.269 ;
      RECT 41.235 2.655 41.25 3.279 ;
      RECT 41.22 2.696 41.235 3.293 ;
      RECT 41.21 2.731 41.22 3.303 ;
      RECT 41.205 2.747 41.21 3.308 ;
      RECT 41.195 2.762 41.205 3.313 ;
      RECT 41.175 2.805 41.195 3.323 ;
      RECT 41.155 2.842 41.175 3.336 ;
      RECT 41.12 2.865 41.155 3.354 ;
      RECT 41.11 2.879 41.12 3.37 ;
      RECT 41.09 2.889 41.11 3.38 ;
      RECT 41.085 2.898 41.09 3.388 ;
      RECT 41.075 2.905 41.085 3.395 ;
      RECT 41.065 2.912 41.075 3.403 ;
      RECT 41.05 2.922 41.065 3.411 ;
      RECT 41.04 2.936 41.05 3.421 ;
      RECT 41.03 2.948 41.04 3.433 ;
      RECT 41.015 2.97 41.03 3.446 ;
      RECT 41.005 2.992 41.015 3.457 ;
      RECT 40.995 3.012 41.005 3.466 ;
      RECT 40.99 3.027 40.995 3.473 ;
      RECT 40.96 3.06 40.99 3.487 ;
      RECT 40.95 3.095 40.96 3.502 ;
      RECT 40.945 3.102 40.95 3.508 ;
      RECT 40.925 3.117 40.945 3.515 ;
      RECT 40.92 3.132 40.925 3.523 ;
      RECT 40.915 3.141 40.92 3.528 ;
      RECT 40.9 3.147 40.915 3.535 ;
      RECT 40.895 3.153 40.9 3.543 ;
      RECT 40.89 3.157 40.895 3.55 ;
      RECT 40.885 3.161 40.89 3.56 ;
      RECT 40.875 3.166 40.885 3.57 ;
      RECT 40.855 3.177 40.875 3.598 ;
      RECT 40.84 3.189 40.855 3.625 ;
      RECT 40.82 3.202 40.84 3.65 ;
      RECT 40.8 3.217 40.82 3.674 ;
      RECT 40.785 3.232 40.8 3.689 ;
      RECT 40.78 3.243 40.785 3.698 ;
      RECT 40.715 3.288 40.78 3.708 ;
      RECT 40.68 3.347 40.715 3.721 ;
      RECT 40.675 3.37 40.68 3.727 ;
      RECT 40.67 3.377 40.675 3.729 ;
      RECT 40.655 3.387 40.67 3.732 ;
      RECT 40.625 3.412 40.655 3.736 ;
      RECT 40.62 3.43 40.625 3.74 ;
      RECT 40.615 3.437 40.62 3.741 ;
      RECT 40.595 3.445 40.615 3.745 ;
      RECT 40.585 3.452 40.595 3.749 ;
      RECT 40.541 3.463 40.585 3.756 ;
      RECT 40.455 3.491 40.541 3.772 ;
      RECT 40.395 3.515 40.455 3.79 ;
      RECT 40.35 3.525 40.395 3.804 ;
      RECT 40.291 3.533 40.35 3.818 ;
      RECT 40.205 3.54 40.291 3.837 ;
      RECT 40.18 3.545 40.205 3.852 ;
      RECT 40.1 3.548 40.18 3.855 ;
      RECT 40.02 3.552 40.1 3.842 ;
      RECT 40.011 3.555 40.02 3.827 ;
      RECT 39.925 3.555 40.011 3.812 ;
      RECT 39.865 3.557 39.925 3.789 ;
      RECT 39.861 3.56 39.865 3.779 ;
      RECT 39.775 3.56 39.861 3.764 ;
      RECT 39.7 3.56 39.775 3.74 ;
      RECT 41.015 2.569 41.025 2.745 ;
      RECT 40.97 2.536 41.015 2.745 ;
      RECT 40.925 2.487 40.97 2.745 ;
      RECT 40.895 2.457 40.925 2.746 ;
      RECT 40.89 2.44 40.895 2.747 ;
      RECT 40.865 2.42 40.89 2.748 ;
      RECT 40.85 2.395 40.865 2.749 ;
      RECT 40.845 2.382 40.85 2.75 ;
      RECT 40.84 2.376 40.845 2.748 ;
      RECT 40.835 2.368 40.84 2.742 ;
      RECT 40.81 2.36 40.835 2.722 ;
      RECT 40.79 2.349 40.81 2.693 ;
      RECT 40.76 2.334 40.79 2.664 ;
      RECT 40.74 2.32 40.76 2.636 ;
      RECT 40.73 2.314 40.74 2.615 ;
      RECT 40.725 2.311 40.73 2.598 ;
      RECT 40.72 2.308 40.725 2.583 ;
      RECT 40.705 2.303 40.72 2.548 ;
      RECT 40.7 2.299 40.705 2.515 ;
      RECT 40.68 2.294 40.7 2.491 ;
      RECT 40.65 2.286 40.68 2.456 ;
      RECT 40.635 2.28 40.65 2.433 ;
      RECT 40.595 2.273 40.635 2.418 ;
      RECT 40.57 2.265 40.595 2.398 ;
      RECT 40.55 2.26 40.57 2.388 ;
      RECT 40.515 2.254 40.55 2.383 ;
      RECT 40.47 2.245 40.515 2.382 ;
      RECT 40.44 2.241 40.47 2.384 ;
      RECT 40.355 2.249 40.44 2.388 ;
      RECT 40.285 2.26 40.355 2.41 ;
      RECT 40.272 2.266 40.285 2.433 ;
      RECT 40.186 2.273 40.272 2.455 ;
      RECT 40.1 2.285 40.186 2.492 ;
      RECT 40.1 2.662 40.11 2.9 ;
      RECT 40.095 2.291 40.1 2.515 ;
      RECT 40.09 2.547 40.1 2.9 ;
      RECT 40.09 2.292 40.095 2.52 ;
      RECT 40.085 2.293 40.09 2.9 ;
      RECT 40.061 2.295 40.085 2.901 ;
      RECT 39.975 2.303 40.061 2.903 ;
      RECT 39.955 2.317 39.975 2.906 ;
      RECT 39.95 2.345 39.955 2.907 ;
      RECT 39.945 2.357 39.95 2.908 ;
      RECT 39.94 2.372 39.945 2.909 ;
      RECT 39.93 2.402 39.94 2.91 ;
      RECT 39.925 2.44 39.93 2.908 ;
      RECT 39.92 2.46 39.925 2.903 ;
      RECT 39.905 2.495 39.92 2.888 ;
      RECT 39.895 2.547 39.905 2.868 ;
      RECT 39.89 2.577 39.895 2.856 ;
      RECT 39.875 2.59 39.89 2.839 ;
      RECT 39.85 2.594 39.875 2.806 ;
      RECT 39.835 2.592 39.85 2.783 ;
      RECT 39.82 2.591 39.835 2.78 ;
      RECT 39.76 2.589 39.82 2.778 ;
      RECT 39.75 2.587 39.76 2.773 ;
      RECT 39.71 2.586 39.75 2.77 ;
      RECT 39.64 2.583 39.71 2.768 ;
      RECT 39.585 2.581 39.64 2.763 ;
      RECT 39.515 2.575 39.585 2.758 ;
      RECT 39.506 2.575 39.515 2.755 ;
      RECT 39.42 2.575 39.506 2.75 ;
      RECT 39.415 2.575 39.42 2.745 ;
      RECT 40.72 1.81 40.895 2.16 ;
      RECT 40.72 1.825 40.905 2.158 ;
      RECT 40.695 1.775 40.84 2.155 ;
      RECT 40.675 1.776 40.84 2.148 ;
      RECT 40.665 1.777 40.85 2.143 ;
      RECT 40.635 1.778 40.85 2.13 ;
      RECT 40.585 1.779 40.85 2.106 ;
      RECT 40.58 1.781 40.85 2.091 ;
      RECT 40.58 1.847 40.91 2.085 ;
      RECT 40.56 1.788 40.865 2.065 ;
      RECT 40.55 1.797 40.875 1.92 ;
      RECT 40.56 1.792 40.875 2.065 ;
      RECT 40.58 1.782 40.865 2.091 ;
      RECT 40.165 3.107 40.335 3.395 ;
      RECT 40.16 3.125 40.345 3.39 ;
      RECT 40.125 3.133 40.41 3.31 ;
      RECT 40.125 3.133 40.496 3.3 ;
      RECT 40.125 3.133 40.55 3.246 ;
      RECT 40.41 3.03 40.58 3.214 ;
      RECT 40.125 3.185 40.585 3.202 ;
      RECT 40.11 3.155 40.58 3.198 ;
      RECT 40.37 3.037 40.41 3.349 ;
      RECT 40.25 3.074 40.58 3.214 ;
      RECT 40.345 3.049 40.37 3.375 ;
      RECT 40.335 3.056 40.58 3.214 ;
      RECT 40.466 2.52 40.535 2.779 ;
      RECT 40.466 2.575 40.54 2.778 ;
      RECT 40.38 2.575 40.54 2.777 ;
      RECT 40.375 2.575 40.545 2.77 ;
      RECT 40.365 2.52 40.535 2.765 ;
      RECT 39.745 1.819 39.92 2.12 ;
      RECT 39.73 1.807 39.745 2.105 ;
      RECT 39.7 1.806 39.73 2.058 ;
      RECT 39.7 1.824 39.925 2.053 ;
      RECT 39.685 1.808 39.745 2.018 ;
      RECT 39.68 1.83 39.935 1.918 ;
      RECT 39.68 1.813 39.831 1.918 ;
      RECT 39.68 1.815 39.835 1.918 ;
      RECT 39.685 1.811 39.831 2.018 ;
      RECT 39.79 3.047 39.795 3.395 ;
      RECT 39.78 3.037 39.79 3.401 ;
      RECT 39.745 3.027 39.78 3.403 ;
      RECT 39.707 3.022 39.745 3.407 ;
      RECT 39.621 3.015 39.707 3.414 ;
      RECT 39.535 3.005 39.621 3.424 ;
      RECT 39.49 3 39.535 3.432 ;
      RECT 39.486 3 39.49 3.436 ;
      RECT 39.4 3 39.486 3.443 ;
      RECT 39.385 3 39.4 3.443 ;
      RECT 39.375 2.998 39.385 3.415 ;
      RECT 39.365 2.994 39.375 3.358 ;
      RECT 39.345 2.988 39.365 3.29 ;
      RECT 39.34 2.984 39.345 3.238 ;
      RECT 39.33 2.983 39.34 3.205 ;
      RECT 39.28 2.981 39.33 3.19 ;
      RECT 39.255 2.979 39.28 3.185 ;
      RECT 39.212 2.977 39.255 3.181 ;
      RECT 39.126 2.973 39.212 3.169 ;
      RECT 39.04 2.968 39.126 3.153 ;
      RECT 39.01 2.965 39.04 3.14 ;
      RECT 38.985 2.964 39.01 3.128 ;
      RECT 38.98 2.964 38.985 3.118 ;
      RECT 38.94 2.963 38.98 3.11 ;
      RECT 38.925 2.962 38.94 3.103 ;
      RECT 38.875 2.961 38.925 3.095 ;
      RECT 38.873 2.96 38.875 3.09 ;
      RECT 38.787 2.958 38.873 3.09 ;
      RECT 38.701 2.953 38.787 3.09 ;
      RECT 38.615 2.949 38.701 3.09 ;
      RECT 38.566 2.945 38.615 3.088 ;
      RECT 38.48 2.942 38.566 3.083 ;
      RECT 38.457 2.939 38.48 3.079 ;
      RECT 38.371 2.936 38.457 3.074 ;
      RECT 38.285 2.932 38.371 3.065 ;
      RECT 38.26 2.925 38.285 3.06 ;
      RECT 38.2 2.89 38.26 3.057 ;
      RECT 38.18 2.815 38.2 3.054 ;
      RECT 38.175 2.757 38.18 3.053 ;
      RECT 38.15 2.697 38.175 3.052 ;
      RECT 38.075 2.575 38.15 3.048 ;
      RECT 38.065 2.575 38.075 3.04 ;
      RECT 38.05 2.575 38.065 3.03 ;
      RECT 38.035 2.575 38.05 3 ;
      RECT 38.02 2.575 38.035 2.945 ;
      RECT 38.005 2.575 38.02 2.883 ;
      RECT 37.98 2.575 38.005 2.808 ;
      RECT 37.975 2.575 37.98 2.758 ;
      RECT 39.32 2.12 39.34 2.429 ;
      RECT 39.306 2.122 39.355 2.426 ;
      RECT 39.306 2.127 39.375 2.417 ;
      RECT 39.22 2.125 39.355 2.411 ;
      RECT 39.22 2.133 39.41 2.394 ;
      RECT 39.185 2.135 39.41 2.393 ;
      RECT 39.155 2.143 39.41 2.384 ;
      RECT 39.145 2.148 39.43 2.37 ;
      RECT 39.185 2.138 39.43 2.37 ;
      RECT 39.185 2.141 39.44 2.358 ;
      RECT 39.155 2.143 39.45 2.345 ;
      RECT 39.155 2.147 39.46 2.288 ;
      RECT 39.145 2.152 39.465 2.203 ;
      RECT 39.306 2.12 39.34 2.426 ;
      RECT 39.185 7.855 39.355 8.305 ;
      RECT 39.24 6.075 39.41 8.025 ;
      RECT 39.185 5.015 39.355 6.245 ;
      RECT 38.745 2.223 38.75 2.435 ;
      RECT 38.62 2.22 38.635 2.435 ;
      RECT 38.085 2.25 38.155 2.435 ;
      RECT 37.97 2.25 38.005 2.43 ;
      RECT 39.091 2.552 39.11 2.746 ;
      RECT 39.005 2.507 39.091 2.747 ;
      RECT 38.995 2.46 39.005 2.749 ;
      RECT 38.99 2.44 38.995 2.75 ;
      RECT 38.97 2.405 38.99 2.751 ;
      RECT 38.955 2.355 38.97 2.752 ;
      RECT 38.935 2.292 38.955 2.753 ;
      RECT 38.925 2.255 38.935 2.754 ;
      RECT 38.91 2.244 38.925 2.755 ;
      RECT 38.905 2.236 38.91 2.753 ;
      RECT 38.895 2.235 38.905 2.745 ;
      RECT 38.865 2.232 38.895 2.724 ;
      RECT 38.79 2.227 38.865 2.669 ;
      RECT 38.775 2.223 38.79 2.615 ;
      RECT 38.765 2.223 38.775 2.51 ;
      RECT 38.75 2.223 38.765 2.443 ;
      RECT 38.735 2.223 38.745 2.433 ;
      RECT 38.68 2.222 38.735 2.43 ;
      RECT 38.635 2.22 38.68 2.433 ;
      RECT 38.607 2.22 38.62 2.436 ;
      RECT 38.521 2.224 38.607 2.438 ;
      RECT 38.435 2.23 38.521 2.443 ;
      RECT 38.415 2.234 38.435 2.445 ;
      RECT 38.413 2.235 38.415 2.444 ;
      RECT 38.327 2.237 38.413 2.443 ;
      RECT 38.241 2.242 38.327 2.44 ;
      RECT 38.155 2.247 38.241 2.437 ;
      RECT 38.005 2.25 38.085 2.433 ;
      RECT 38.665 5.015 38.835 8.305 ;
      RECT 38.665 7.315 39.07 7.645 ;
      RECT 38.665 6.475 39.07 6.805 ;
      RECT 38.781 3.225 38.83 3.559 ;
      RECT 38.781 3.225 38.835 3.558 ;
      RECT 38.695 3.225 38.835 3.557 ;
      RECT 38.47 3.333 38.84 3.555 ;
      RECT 38.695 3.225 38.865 3.548 ;
      RECT 38.665 3.237 38.87 3.539 ;
      RECT 38.65 3.255 38.875 3.536 ;
      RECT 38.465 3.339 38.875 3.463 ;
      RECT 38.46 3.346 38.875 3.423 ;
      RECT 38.475 3.312 38.875 3.536 ;
      RECT 38.636 3.258 38.84 3.555 ;
      RECT 38.55 3.278 38.875 3.536 ;
      RECT 38.65 3.252 38.87 3.539 ;
      RECT 38.42 2.576 38.61 2.77 ;
      RECT 38.415 2.578 38.61 2.769 ;
      RECT 38.41 2.582 38.625 2.766 ;
      RECT 38.425 2.575 38.625 2.766 ;
      RECT 38.41 2.685 38.63 2.761 ;
      RECT 37.705 3.185 37.796 3.483 ;
      RECT 37.7 3.187 37.875 3.478 ;
      RECT 37.705 3.185 37.875 3.478 ;
      RECT 37.7 3.191 37.895 3.476 ;
      RECT 37.7 3.246 37.935 3.475 ;
      RECT 37.7 3.281 37.95 3.469 ;
      RECT 37.7 3.315 37.96 3.459 ;
      RECT 37.69 3.195 37.895 3.31 ;
      RECT 37.69 3.215 37.91 3.31 ;
      RECT 37.69 3.198 37.9 3.31 ;
      RECT 37.915 1.966 37.92 2.028 ;
      RECT 37.91 1.888 37.915 2.051 ;
      RECT 37.905 1.845 37.91 2.062 ;
      RECT 37.9 1.835 37.905 2.074 ;
      RECT 37.895 1.835 37.9 2.083 ;
      RECT 37.87 1.835 37.895 2.115 ;
      RECT 37.865 1.835 37.87 2.148 ;
      RECT 37.85 1.835 37.865 2.173 ;
      RECT 37.84 1.835 37.85 2.2 ;
      RECT 37.835 1.835 37.84 2.213 ;
      RECT 37.83 1.835 37.835 2.228 ;
      RECT 37.82 1.835 37.83 2.243 ;
      RECT 37.815 1.835 37.82 2.263 ;
      RECT 37.79 1.835 37.815 2.298 ;
      RECT 37.745 1.835 37.79 2.343 ;
      RECT 37.735 1.835 37.745 2.356 ;
      RECT 37.65 1.92 37.735 2.363 ;
      RECT 37.615 2.042 37.65 2.372 ;
      RECT 37.61 2.082 37.615 2.376 ;
      RECT 37.59 2.105 37.61 2.378 ;
      RECT 37.585 2.135 37.59 2.381 ;
      RECT 37.575 2.147 37.585 2.382 ;
      RECT 37.53 2.17 37.575 2.387 ;
      RECT 37.49 2.2 37.53 2.395 ;
      RECT 37.455 2.212 37.49 2.401 ;
      RECT 37.45 2.217 37.455 2.405 ;
      RECT 37.38 2.227 37.45 2.412 ;
      RECT 37.34 2.237 37.38 2.422 ;
      RECT 37.32 2.242 37.34 2.428 ;
      RECT 37.31 2.246 37.32 2.433 ;
      RECT 37.305 2.249 37.31 2.436 ;
      RECT 37.295 2.25 37.305 2.437 ;
      RECT 37.27 2.252 37.295 2.441 ;
      RECT 37.26 2.257 37.27 2.444 ;
      RECT 37.215 2.265 37.26 2.445 ;
      RECT 37.09 2.27 37.215 2.445 ;
      RECT 37.645 2.567 37.665 2.749 ;
      RECT 37.596 2.552 37.645 2.748 ;
      RECT 37.51 2.567 37.665 2.746 ;
      RECT 37.495 2.567 37.665 2.745 ;
      RECT 37.46 2.545 37.63 2.73 ;
      RECT 37.53 3.565 37.545 3.774 ;
      RECT 37.53 3.573 37.55 3.773 ;
      RECT 37.475 3.573 37.55 3.772 ;
      RECT 37.455 3.577 37.555 3.77 ;
      RECT 37.435 3.527 37.475 3.769 ;
      RECT 37.38 3.585 37.56 3.767 ;
      RECT 37.345 3.542 37.475 3.765 ;
      RECT 37.341 3.545 37.53 3.764 ;
      RECT 37.255 3.553 37.53 3.762 ;
      RECT 37.255 3.597 37.565 3.755 ;
      RECT 37.245 3.69 37.565 3.753 ;
      RECT 37.255 3.609 37.57 3.738 ;
      RECT 37.255 3.63 37.585 3.708 ;
      RECT 37.255 3.657 37.59 3.678 ;
      RECT 37.38 3.535 37.475 3.767 ;
      RECT 37.01 2.58 37.015 3.118 ;
      RECT 36.815 2.91 36.82 3.105 ;
      RECT 35.115 2.575 35.13 2.955 ;
      RECT 37.18 2.575 37.185 2.745 ;
      RECT 37.175 2.575 37.18 2.755 ;
      RECT 37.17 2.575 37.175 2.768 ;
      RECT 37.145 2.575 37.17 2.81 ;
      RECT 37.12 2.575 37.145 2.883 ;
      RECT 37.105 2.575 37.12 2.935 ;
      RECT 37.1 2.575 37.105 2.965 ;
      RECT 37.075 2.575 37.1 3.005 ;
      RECT 37.06 2.575 37.075 3.06 ;
      RECT 37.055 2.575 37.06 3.093 ;
      RECT 37.03 2.575 37.055 3.113 ;
      RECT 37.015 2.575 37.03 3.119 ;
      RECT 36.945 2.61 37.01 3.115 ;
      RECT 36.895 2.665 36.945 3.11 ;
      RECT 36.885 2.697 36.895 3.108 ;
      RECT 36.88 2.722 36.885 3.108 ;
      RECT 36.86 2.795 36.88 3.108 ;
      RECT 36.85 2.875 36.86 3.107 ;
      RECT 36.835 2.905 36.85 3.107 ;
      RECT 36.82 2.91 36.835 3.106 ;
      RECT 36.76 2.912 36.815 3.103 ;
      RECT 36.73 2.917 36.76 3.099 ;
      RECT 36.728 2.92 36.73 3.098 ;
      RECT 36.642 2.922 36.728 3.095 ;
      RECT 36.556 2.928 36.642 3.089 ;
      RECT 36.47 2.933 36.556 3.083 ;
      RECT 36.397 2.938 36.47 3.084 ;
      RECT 36.311 2.944 36.397 3.092 ;
      RECT 36.225 2.95 36.311 3.101 ;
      RECT 36.205 2.954 36.225 3.106 ;
      RECT 36.158 2.956 36.205 3.109 ;
      RECT 36.072 2.961 36.158 3.115 ;
      RECT 35.986 2.966 36.072 3.124 ;
      RECT 35.9 2.972 35.986 3.132 ;
      RECT 35.815 2.97 35.9 3.141 ;
      RECT 35.811 2.965 35.815 3.145 ;
      RECT 35.725 2.96 35.811 3.137 ;
      RECT 35.661 2.951 35.725 3.125 ;
      RECT 35.575 2.942 35.661 3.112 ;
      RECT 35.551 2.935 35.575 3.103 ;
      RECT 35.465 2.929 35.551 3.09 ;
      RECT 35.425 2.922 35.465 3.076 ;
      RECT 35.42 2.912 35.425 3.072 ;
      RECT 35.41 2.9 35.42 3.071 ;
      RECT 35.39 2.87 35.41 3.068 ;
      RECT 35.335 2.79 35.39 3.062 ;
      RECT 35.315 2.709 35.335 3.057 ;
      RECT 35.295 2.667 35.315 3.053 ;
      RECT 35.27 2.62 35.295 3.047 ;
      RECT 35.265 2.595 35.27 3.044 ;
      RECT 35.23 2.575 35.265 3.039 ;
      RECT 35.221 2.575 35.23 3.032 ;
      RECT 35.135 2.575 35.221 3.002 ;
      RECT 35.13 2.575 35.135 2.965 ;
      RECT 35.095 2.575 35.115 2.887 ;
      RECT 35.09 2.617 35.095 2.852 ;
      RECT 35.085 2.692 35.09 2.808 ;
      RECT 36.535 2.497 36.71 2.745 ;
      RECT 36.535 2.497 36.715 2.743 ;
      RECT 36.53 2.529 36.715 2.703 ;
      RECT 36.56 2.47 36.73 2.69 ;
      RECT 36.525 2.547 36.73 2.623 ;
      RECT 35.835 2.01 36.005 2.185 ;
      RECT 35.835 2.01 36.177 2.177 ;
      RECT 35.835 2.01 36.26 2.171 ;
      RECT 35.835 2.01 36.295 2.167 ;
      RECT 35.835 2.01 36.315 2.166 ;
      RECT 35.835 2.01 36.401 2.162 ;
      RECT 36.295 1.835 36.465 2.157 ;
      RECT 35.87 1.942 36.495 2.155 ;
      RECT 35.86 1.997 36.5 2.153 ;
      RECT 35.835 2.033 36.51 2.148 ;
      RECT 35.835 2.06 36.515 2.078 ;
      RECT 35.9 1.885 36.475 2.155 ;
      RECT 36.091 1.87 36.475 2.155 ;
      RECT 35.925 1.873 36.475 2.155 ;
      RECT 36.005 1.871 36.091 2.182 ;
      RECT 36.091 1.868 36.47 2.155 ;
      RECT 36.275 1.845 36.47 2.155 ;
      RECT 36.177 1.866 36.47 2.155 ;
      RECT 36.26 1.86 36.275 2.168 ;
      RECT 36.41 3.225 36.415 3.425 ;
      RECT 35.875 3.29 35.92 3.425 ;
      RECT 36.445 3.225 36.465 3.398 ;
      RECT 36.415 3.225 36.445 3.413 ;
      RECT 36.35 3.225 36.41 3.45 ;
      RECT 36.335 3.225 36.35 3.48 ;
      RECT 36.32 3.225 36.335 3.493 ;
      RECT 36.3 3.225 36.32 3.508 ;
      RECT 36.295 3.225 36.3 3.517 ;
      RECT 36.285 3.229 36.295 3.522 ;
      RECT 36.27 3.239 36.285 3.533 ;
      RECT 36.245 3.255 36.27 3.543 ;
      RECT 36.235 3.269 36.245 3.545 ;
      RECT 36.215 3.281 36.235 3.542 ;
      RECT 36.185 3.302 36.215 3.536 ;
      RECT 36.175 3.314 36.185 3.531 ;
      RECT 36.165 3.312 36.175 3.528 ;
      RECT 36.15 3.311 36.165 3.523 ;
      RECT 36.145 3.31 36.15 3.518 ;
      RECT 36.11 3.308 36.145 3.508 ;
      RECT 36.09 3.305 36.11 3.49 ;
      RECT 36.08 3.303 36.09 3.485 ;
      RECT 36.07 3.302 36.08 3.48 ;
      RECT 36.035 3.3 36.07 3.468 ;
      RECT 35.98 3.296 36.035 3.448 ;
      RECT 35.97 3.294 35.98 3.433 ;
      RECT 35.965 3.294 35.97 3.428 ;
      RECT 35.92 3.292 35.965 3.425 ;
      RECT 35.825 3.29 35.875 3.429 ;
      RECT 35.815 3.291 35.825 3.434 ;
      RECT 35.755 3.298 35.815 3.448 ;
      RECT 35.73 3.306 35.755 3.468 ;
      RECT 35.72 3.31 35.73 3.48 ;
      RECT 35.715 3.311 35.72 3.485 ;
      RECT 35.7 3.313 35.715 3.488 ;
      RECT 35.685 3.315 35.7 3.493 ;
      RECT 35.68 3.315 35.685 3.496 ;
      RECT 35.635 3.32 35.68 3.507 ;
      RECT 35.63 3.324 35.635 3.519 ;
      RECT 35.605 3.32 35.63 3.523 ;
      RECT 35.595 3.316 35.605 3.527 ;
      RECT 35.585 3.315 35.595 3.531 ;
      RECT 35.57 3.305 35.585 3.537 ;
      RECT 35.565 3.293 35.57 3.541 ;
      RECT 35.56 3.29 35.565 3.542 ;
      RECT 35.555 3.287 35.56 3.544 ;
      RECT 35.54 3.275 35.555 3.543 ;
      RECT 35.525 3.257 35.54 3.54 ;
      RECT 35.505 3.236 35.525 3.533 ;
      RECT 35.44 3.225 35.505 3.505 ;
      RECT 35.436 3.225 35.44 3.484 ;
      RECT 35.35 3.225 35.436 3.454 ;
      RECT 35.335 3.225 35.35 3.41 ;
      RECT 35.91 2.325 35.915 2.56 ;
      RECT 35.04 2.241 35.045 2.445 ;
      RECT 35.62 2.27 35.625 2.425 ;
      RECT 35.54 2.25 35.545 2.425 ;
      RECT 36.21 2.392 36.225 2.745 ;
      RECT 36.136 2.377 36.21 2.745 ;
      RECT 36.05 2.36 36.136 2.745 ;
      RECT 36.04 2.35 36.05 2.743 ;
      RECT 36.035 2.348 36.04 2.738 ;
      RECT 36.02 2.346 36.035 2.724 ;
      RECT 35.95 2.338 36.02 2.664 ;
      RECT 35.93 2.329 35.95 2.598 ;
      RECT 35.925 2.326 35.93 2.578 ;
      RECT 35.915 2.325 35.925 2.568 ;
      RECT 35.905 2.325 35.91 2.552 ;
      RECT 35.895 2.324 35.905 2.542 ;
      RECT 35.885 2.322 35.895 2.53 ;
      RECT 35.87 2.319 35.885 2.51 ;
      RECT 35.86 2.317 35.87 2.495 ;
      RECT 35.84 2.314 35.86 2.483 ;
      RECT 35.835 2.312 35.84 2.473 ;
      RECT 35.81 2.31 35.835 2.46 ;
      RECT 35.78 2.305 35.81 2.445 ;
      RECT 35.7 2.296 35.78 2.436 ;
      RECT 35.655 2.285 35.7 2.429 ;
      RECT 35.635 2.276 35.655 2.426 ;
      RECT 35.625 2.271 35.635 2.425 ;
      RECT 35.58 2.265 35.62 2.425 ;
      RECT 35.565 2.257 35.58 2.425 ;
      RECT 35.545 2.252 35.565 2.425 ;
      RECT 35.525 2.249 35.54 2.425 ;
      RECT 35.442 2.248 35.525 2.424 ;
      RECT 35.356 2.247 35.442 2.42 ;
      RECT 35.27 2.245 35.356 2.417 ;
      RECT 35.217 2.244 35.27 2.419 ;
      RECT 35.131 2.243 35.217 2.428 ;
      RECT 35.045 2.242 35.131 2.44 ;
      RECT 35.025 2.241 35.04 2.448 ;
      RECT 34.945 2.24 35.025 2.46 ;
      RECT 34.92 2.24 34.945 2.473 ;
      RECT 34.895 2.24 34.92 2.488 ;
      RECT 34.89 2.24 34.895 2.51 ;
      RECT 34.885 2.24 34.89 2.528 ;
      RECT 34.88 2.24 34.885 2.545 ;
      RECT 34.875 2.24 34.88 2.558 ;
      RECT 34.87 2.24 34.875 2.568 ;
      RECT 34.83 2.24 34.87 2.653 ;
      RECT 34.815 2.24 34.83 2.738 ;
      RECT 34.805 2.241 34.815 2.75 ;
      RECT 34.77 2.246 34.805 2.755 ;
      RECT 34.73 2.255 34.77 2.755 ;
      RECT 34.715 2.265 34.73 2.755 ;
      RECT 34.71 2.275 34.715 2.755 ;
      RECT 34.69 2.302 34.71 2.755 ;
      RECT 34.64 2.385 34.69 2.755 ;
      RECT 34.635 2.447 34.64 2.755 ;
      RECT 34.625 2.46 34.635 2.755 ;
      RECT 34.615 2.482 34.625 2.755 ;
      RECT 34.605 2.507 34.615 2.75 ;
      RECT 34.6 2.545 34.605 2.743 ;
      RECT 34.59 2.655 34.6 2.738 ;
      RECT 35.985 3.576 36 3.835 ;
      RECT 35.985 3.591 36.005 3.834 ;
      RECT 35.901 3.591 36.005 3.832 ;
      RECT 35.901 3.605 36.01 3.831 ;
      RECT 35.815 3.647 36.015 3.828 ;
      RECT 35.81 3.59 36 3.823 ;
      RECT 35.81 3.661 36.02 3.82 ;
      RECT 35.805 3.692 36.02 3.818 ;
      RECT 35.81 3.689 36.035 3.808 ;
      RECT 35.805 3.735 36.05 3.793 ;
      RECT 35.805 3.763 36.055 3.778 ;
      RECT 35.815 3.565 35.985 3.828 ;
      RECT 35.575 2.575 35.745 2.745 ;
      RECT 35.54 2.575 35.745 2.74 ;
      RECT 35.53 2.575 35.745 2.733 ;
      RECT 35.525 2.56 35.695 2.73 ;
      RECT 34.355 3.097 34.62 3.54 ;
      RECT 34.35 3.068 34.565 3.538 ;
      RECT 34.345 3.222 34.625 3.533 ;
      RECT 34.35 3.117 34.625 3.533 ;
      RECT 34.35 3.128 34.635 3.52 ;
      RECT 34.35 3.075 34.595 3.538 ;
      RECT 34.355 3.062 34.565 3.54 ;
      RECT 34.355 3.06 34.515 3.54 ;
      RECT 34.456 3.052 34.515 3.54 ;
      RECT 34.37 3.053 34.515 3.54 ;
      RECT 34.456 3.051 34.505 3.54 ;
      RECT 34.26 1.866 34.435 2.165 ;
      RECT 34.31 1.828 34.435 2.165 ;
      RECT 34.295 1.83 34.521 2.157 ;
      RECT 34.295 1.833 34.56 2.144 ;
      RECT 34.295 1.834 34.57 2.13 ;
      RECT 34.25 1.885 34.57 2.12 ;
      RECT 34.295 1.835 34.575 2.115 ;
      RECT 34.25 2.045 34.58 2.105 ;
      RECT 34.235 1.905 34.575 2.045 ;
      RECT 34.23 1.921 34.575 1.985 ;
      RECT 34.275 1.845 34.575 2.115 ;
      RECT 34.31 1.826 34.396 2.165 ;
      RECT 32.77 5.02 32.94 6.49 ;
      RECT 32.77 6.315 32.945 6.485 ;
      RECT 32.4 1.74 32.57 2.93 ;
      RECT 32.4 1.74 32.87 1.91 ;
      RECT 32.4 6.97 32.87 7.14 ;
      RECT 32.4 5.95 32.57 7.14 ;
      RECT 31.41 1.74 31.58 2.93 ;
      RECT 31.41 1.74 31.88 1.91 ;
      RECT 31.41 6.97 31.88 7.14 ;
      RECT 31.41 5.95 31.58 7.14 ;
      RECT 29.56 2.635 29.73 3.865 ;
      RECT 29.615 0.855 29.785 2.805 ;
      RECT 29.56 0.575 29.73 1.025 ;
      RECT 29.56 7.855 29.73 8.305 ;
      RECT 29.615 6.075 29.785 8.025 ;
      RECT 29.56 5.015 29.73 6.245 ;
      RECT 29.04 0.575 29.21 3.865 ;
      RECT 29.04 2.075 29.445 2.405 ;
      RECT 29.04 1.235 29.445 1.565 ;
      RECT 29.04 5.015 29.21 8.305 ;
      RECT 29.04 7.315 29.445 7.645 ;
      RECT 29.04 6.475 29.445 6.805 ;
      RECT 26.965 3.126 26.97 3.298 ;
      RECT 26.96 3.119 26.965 3.388 ;
      RECT 26.955 3.113 26.96 3.407 ;
      RECT 26.935 3.107 26.955 3.417 ;
      RECT 26.92 3.102 26.935 3.425 ;
      RECT 26.883 3.096 26.92 3.423 ;
      RECT 26.797 3.082 26.883 3.419 ;
      RECT 26.711 3.064 26.797 3.414 ;
      RECT 26.625 3.045 26.711 3.408 ;
      RECT 26.595 3.033 26.625 3.404 ;
      RECT 26.575 3.027 26.595 3.403 ;
      RECT 26.51 3.025 26.575 3.401 ;
      RECT 26.495 3.025 26.51 3.393 ;
      RECT 26.48 3.025 26.495 3.38 ;
      RECT 26.475 3.025 26.48 3.37 ;
      RECT 26.46 3.025 26.475 3.348 ;
      RECT 26.445 3.025 26.46 3.315 ;
      RECT 26.44 3.025 26.445 3.293 ;
      RECT 26.43 3.025 26.44 3.275 ;
      RECT 26.415 3.025 26.43 3.253 ;
      RECT 26.395 3.025 26.415 3.215 ;
      RECT 26.745 2.31 26.78 2.749 ;
      RECT 26.745 2.31 26.785 2.748 ;
      RECT 26.69 2.37 26.785 2.747 ;
      RECT 26.555 2.542 26.785 2.746 ;
      RECT 26.665 2.42 26.785 2.746 ;
      RECT 26.555 2.542 26.81 2.736 ;
      RECT 26.61 2.487 26.89 2.653 ;
      RECT 26.785 2.281 26.79 2.744 ;
      RECT 26.64 2.457 26.93 2.53 ;
      RECT 26.655 2.44 26.785 2.746 ;
      RECT 26.79 2.28 26.96 2.468 ;
      RECT 26.78 2.283 26.96 2.468 ;
      RECT 26.285 2.16 26.455 2.47 ;
      RECT 26.285 2.16 26.46 2.443 ;
      RECT 26.285 2.16 26.465 2.42 ;
      RECT 26.285 2.16 26.475 2.37 ;
      RECT 26.28 2.265 26.475 2.34 ;
      RECT 26.315 1.835 26.485 2.313 ;
      RECT 26.315 1.835 26.5 2.234 ;
      RECT 26.305 2.045 26.5 2.234 ;
      RECT 26.315 1.845 26.51 2.149 ;
      RECT 26.245 2.587 26.25 2.79 ;
      RECT 26.235 2.575 26.245 2.9 ;
      RECT 26.21 2.575 26.235 2.94 ;
      RECT 26.13 2.575 26.21 3.025 ;
      RECT 26.12 2.575 26.13 3.095 ;
      RECT 26.095 2.575 26.12 3.118 ;
      RECT 26.075 2.575 26.095 3.153 ;
      RECT 26.03 2.585 26.075 3.196 ;
      RECT 26.02 2.597 26.03 3.233 ;
      RECT 26 2.611 26.02 3.253 ;
      RECT 25.99 2.629 26 3.269 ;
      RECT 25.975 2.655 25.99 3.279 ;
      RECT 25.96 2.696 25.975 3.293 ;
      RECT 25.95 2.731 25.96 3.303 ;
      RECT 25.945 2.747 25.95 3.308 ;
      RECT 25.935 2.762 25.945 3.313 ;
      RECT 25.915 2.805 25.935 3.323 ;
      RECT 25.895 2.842 25.915 3.336 ;
      RECT 25.86 2.865 25.895 3.354 ;
      RECT 25.85 2.879 25.86 3.37 ;
      RECT 25.83 2.889 25.85 3.38 ;
      RECT 25.825 2.898 25.83 3.388 ;
      RECT 25.815 2.905 25.825 3.395 ;
      RECT 25.805 2.912 25.815 3.403 ;
      RECT 25.79 2.922 25.805 3.411 ;
      RECT 25.78 2.936 25.79 3.421 ;
      RECT 25.77 2.948 25.78 3.433 ;
      RECT 25.755 2.97 25.77 3.446 ;
      RECT 25.745 2.992 25.755 3.457 ;
      RECT 25.735 3.012 25.745 3.466 ;
      RECT 25.73 3.027 25.735 3.473 ;
      RECT 25.7 3.06 25.73 3.487 ;
      RECT 25.69 3.095 25.7 3.502 ;
      RECT 25.685 3.102 25.69 3.508 ;
      RECT 25.665 3.117 25.685 3.515 ;
      RECT 25.66 3.132 25.665 3.523 ;
      RECT 25.655 3.141 25.66 3.528 ;
      RECT 25.64 3.147 25.655 3.535 ;
      RECT 25.635 3.153 25.64 3.543 ;
      RECT 25.63 3.157 25.635 3.55 ;
      RECT 25.625 3.161 25.63 3.56 ;
      RECT 25.615 3.166 25.625 3.57 ;
      RECT 25.595 3.177 25.615 3.598 ;
      RECT 25.58 3.189 25.595 3.625 ;
      RECT 25.56 3.202 25.58 3.65 ;
      RECT 25.54 3.217 25.56 3.674 ;
      RECT 25.525 3.232 25.54 3.689 ;
      RECT 25.52 3.243 25.525 3.698 ;
      RECT 25.455 3.288 25.52 3.708 ;
      RECT 25.42 3.347 25.455 3.721 ;
      RECT 25.415 3.37 25.42 3.727 ;
      RECT 25.41 3.377 25.415 3.729 ;
      RECT 25.395 3.387 25.41 3.732 ;
      RECT 25.365 3.412 25.395 3.736 ;
      RECT 25.36 3.43 25.365 3.74 ;
      RECT 25.355 3.437 25.36 3.741 ;
      RECT 25.335 3.445 25.355 3.745 ;
      RECT 25.325 3.452 25.335 3.749 ;
      RECT 25.281 3.463 25.325 3.756 ;
      RECT 25.195 3.491 25.281 3.772 ;
      RECT 25.135 3.515 25.195 3.79 ;
      RECT 25.09 3.525 25.135 3.804 ;
      RECT 25.031 3.533 25.09 3.818 ;
      RECT 24.945 3.54 25.031 3.837 ;
      RECT 24.92 3.545 24.945 3.852 ;
      RECT 24.84 3.548 24.92 3.855 ;
      RECT 24.76 3.552 24.84 3.842 ;
      RECT 24.751 3.555 24.76 3.827 ;
      RECT 24.665 3.555 24.751 3.812 ;
      RECT 24.605 3.557 24.665 3.789 ;
      RECT 24.601 3.56 24.605 3.779 ;
      RECT 24.515 3.56 24.601 3.764 ;
      RECT 24.44 3.56 24.515 3.74 ;
      RECT 25.755 2.569 25.765 2.745 ;
      RECT 25.71 2.536 25.755 2.745 ;
      RECT 25.665 2.487 25.71 2.745 ;
      RECT 25.635 2.457 25.665 2.746 ;
      RECT 25.63 2.44 25.635 2.747 ;
      RECT 25.605 2.42 25.63 2.748 ;
      RECT 25.59 2.395 25.605 2.749 ;
      RECT 25.585 2.382 25.59 2.75 ;
      RECT 25.58 2.376 25.585 2.748 ;
      RECT 25.575 2.368 25.58 2.742 ;
      RECT 25.55 2.36 25.575 2.722 ;
      RECT 25.53 2.349 25.55 2.693 ;
      RECT 25.5 2.334 25.53 2.664 ;
      RECT 25.48 2.32 25.5 2.636 ;
      RECT 25.47 2.314 25.48 2.615 ;
      RECT 25.465 2.311 25.47 2.598 ;
      RECT 25.46 2.308 25.465 2.583 ;
      RECT 25.445 2.303 25.46 2.548 ;
      RECT 25.44 2.299 25.445 2.515 ;
      RECT 25.42 2.294 25.44 2.491 ;
      RECT 25.39 2.286 25.42 2.456 ;
      RECT 25.375 2.28 25.39 2.433 ;
      RECT 25.335 2.273 25.375 2.418 ;
      RECT 25.31 2.265 25.335 2.398 ;
      RECT 25.29 2.26 25.31 2.388 ;
      RECT 25.255 2.254 25.29 2.383 ;
      RECT 25.21 2.245 25.255 2.382 ;
      RECT 25.18 2.241 25.21 2.384 ;
      RECT 25.095 2.249 25.18 2.388 ;
      RECT 25.025 2.26 25.095 2.41 ;
      RECT 25.012 2.266 25.025 2.433 ;
      RECT 24.926 2.273 25.012 2.455 ;
      RECT 24.84 2.285 24.926 2.492 ;
      RECT 24.84 2.662 24.85 2.9 ;
      RECT 24.835 2.291 24.84 2.515 ;
      RECT 24.83 2.547 24.84 2.9 ;
      RECT 24.83 2.292 24.835 2.52 ;
      RECT 24.825 2.293 24.83 2.9 ;
      RECT 24.801 2.295 24.825 2.901 ;
      RECT 24.715 2.303 24.801 2.903 ;
      RECT 24.695 2.317 24.715 2.906 ;
      RECT 24.69 2.345 24.695 2.907 ;
      RECT 24.685 2.357 24.69 2.908 ;
      RECT 24.68 2.372 24.685 2.909 ;
      RECT 24.67 2.402 24.68 2.91 ;
      RECT 24.665 2.44 24.67 2.908 ;
      RECT 24.66 2.46 24.665 2.903 ;
      RECT 24.645 2.495 24.66 2.888 ;
      RECT 24.635 2.547 24.645 2.868 ;
      RECT 24.63 2.577 24.635 2.856 ;
      RECT 24.615 2.59 24.63 2.839 ;
      RECT 24.59 2.594 24.615 2.806 ;
      RECT 24.575 2.592 24.59 2.783 ;
      RECT 24.56 2.591 24.575 2.78 ;
      RECT 24.5 2.589 24.56 2.778 ;
      RECT 24.49 2.587 24.5 2.773 ;
      RECT 24.45 2.586 24.49 2.77 ;
      RECT 24.38 2.583 24.45 2.768 ;
      RECT 24.325 2.581 24.38 2.763 ;
      RECT 24.255 2.575 24.325 2.758 ;
      RECT 24.246 2.575 24.255 2.755 ;
      RECT 24.16 2.575 24.246 2.75 ;
      RECT 24.155 2.575 24.16 2.745 ;
      RECT 25.46 1.81 25.635 2.16 ;
      RECT 25.46 1.825 25.645 2.158 ;
      RECT 25.435 1.775 25.58 2.155 ;
      RECT 25.415 1.776 25.58 2.148 ;
      RECT 25.405 1.777 25.59 2.143 ;
      RECT 25.375 1.778 25.59 2.13 ;
      RECT 25.325 1.779 25.59 2.106 ;
      RECT 25.32 1.781 25.59 2.091 ;
      RECT 25.32 1.847 25.65 2.085 ;
      RECT 25.3 1.788 25.605 2.065 ;
      RECT 25.29 1.797 25.615 1.92 ;
      RECT 25.3 1.792 25.615 2.065 ;
      RECT 25.32 1.782 25.605 2.091 ;
      RECT 24.905 3.107 25.075 3.395 ;
      RECT 24.9 3.125 25.085 3.39 ;
      RECT 24.865 3.133 25.15 3.31 ;
      RECT 24.865 3.133 25.236 3.3 ;
      RECT 24.865 3.133 25.29 3.246 ;
      RECT 25.15 3.03 25.32 3.214 ;
      RECT 24.865 3.185 25.325 3.202 ;
      RECT 24.85 3.155 25.32 3.198 ;
      RECT 25.11 3.037 25.15 3.349 ;
      RECT 24.99 3.074 25.32 3.214 ;
      RECT 25.085 3.049 25.11 3.375 ;
      RECT 25.075 3.056 25.32 3.214 ;
      RECT 25.206 2.52 25.275 2.779 ;
      RECT 25.206 2.575 25.28 2.778 ;
      RECT 25.12 2.575 25.28 2.777 ;
      RECT 25.115 2.575 25.285 2.77 ;
      RECT 25.105 2.52 25.275 2.765 ;
      RECT 24.485 1.819 24.66 2.12 ;
      RECT 24.47 1.807 24.485 2.105 ;
      RECT 24.44 1.806 24.47 2.058 ;
      RECT 24.44 1.824 24.665 2.053 ;
      RECT 24.425 1.808 24.485 2.018 ;
      RECT 24.42 1.83 24.675 1.918 ;
      RECT 24.42 1.813 24.571 1.918 ;
      RECT 24.42 1.815 24.575 1.918 ;
      RECT 24.425 1.811 24.571 2.018 ;
      RECT 24.53 3.047 24.535 3.395 ;
      RECT 24.52 3.037 24.53 3.401 ;
      RECT 24.485 3.027 24.52 3.403 ;
      RECT 24.447 3.022 24.485 3.407 ;
      RECT 24.361 3.015 24.447 3.414 ;
      RECT 24.275 3.005 24.361 3.424 ;
      RECT 24.23 3 24.275 3.432 ;
      RECT 24.226 3 24.23 3.436 ;
      RECT 24.14 3 24.226 3.443 ;
      RECT 24.125 3 24.14 3.443 ;
      RECT 24.115 2.998 24.125 3.415 ;
      RECT 24.105 2.994 24.115 3.358 ;
      RECT 24.085 2.988 24.105 3.29 ;
      RECT 24.08 2.984 24.085 3.238 ;
      RECT 24.07 2.983 24.08 3.205 ;
      RECT 24.02 2.981 24.07 3.19 ;
      RECT 23.995 2.979 24.02 3.185 ;
      RECT 23.952 2.977 23.995 3.181 ;
      RECT 23.866 2.973 23.952 3.169 ;
      RECT 23.78 2.968 23.866 3.153 ;
      RECT 23.75 2.965 23.78 3.14 ;
      RECT 23.725 2.964 23.75 3.128 ;
      RECT 23.72 2.964 23.725 3.118 ;
      RECT 23.68 2.963 23.72 3.11 ;
      RECT 23.665 2.962 23.68 3.103 ;
      RECT 23.615 2.961 23.665 3.095 ;
      RECT 23.613 2.96 23.615 3.09 ;
      RECT 23.527 2.958 23.613 3.09 ;
      RECT 23.441 2.953 23.527 3.09 ;
      RECT 23.355 2.949 23.441 3.09 ;
      RECT 23.306 2.945 23.355 3.088 ;
      RECT 23.22 2.942 23.306 3.083 ;
      RECT 23.197 2.939 23.22 3.079 ;
      RECT 23.111 2.936 23.197 3.074 ;
      RECT 23.025 2.932 23.111 3.065 ;
      RECT 23 2.925 23.025 3.06 ;
      RECT 22.94 2.89 23 3.057 ;
      RECT 22.92 2.815 22.94 3.054 ;
      RECT 22.915 2.757 22.92 3.053 ;
      RECT 22.89 2.697 22.915 3.052 ;
      RECT 22.815 2.575 22.89 3.048 ;
      RECT 22.805 2.575 22.815 3.04 ;
      RECT 22.79 2.575 22.805 3.03 ;
      RECT 22.775 2.575 22.79 3 ;
      RECT 22.76 2.575 22.775 2.945 ;
      RECT 22.745 2.575 22.76 2.883 ;
      RECT 22.72 2.575 22.745 2.808 ;
      RECT 22.715 2.575 22.72 2.758 ;
      RECT 24.06 2.12 24.08 2.429 ;
      RECT 24.046 2.122 24.095 2.426 ;
      RECT 24.046 2.127 24.115 2.417 ;
      RECT 23.96 2.125 24.095 2.411 ;
      RECT 23.96 2.133 24.15 2.394 ;
      RECT 23.925 2.135 24.15 2.393 ;
      RECT 23.895 2.143 24.15 2.384 ;
      RECT 23.885 2.148 24.17 2.37 ;
      RECT 23.925 2.138 24.17 2.37 ;
      RECT 23.925 2.141 24.18 2.358 ;
      RECT 23.895 2.143 24.19 2.345 ;
      RECT 23.895 2.147 24.2 2.288 ;
      RECT 23.885 2.152 24.205 2.203 ;
      RECT 24.046 2.12 24.08 2.426 ;
      RECT 23.925 7.855 24.095 8.305 ;
      RECT 23.98 6.075 24.15 8.025 ;
      RECT 23.925 5.015 24.095 6.245 ;
      RECT 23.485 2.223 23.49 2.435 ;
      RECT 23.36 2.22 23.375 2.435 ;
      RECT 22.825 2.25 22.895 2.435 ;
      RECT 22.71 2.25 22.745 2.43 ;
      RECT 23.831 2.552 23.85 2.746 ;
      RECT 23.745 2.507 23.831 2.747 ;
      RECT 23.735 2.46 23.745 2.749 ;
      RECT 23.73 2.44 23.735 2.75 ;
      RECT 23.71 2.405 23.73 2.751 ;
      RECT 23.695 2.355 23.71 2.752 ;
      RECT 23.675 2.292 23.695 2.753 ;
      RECT 23.665 2.255 23.675 2.754 ;
      RECT 23.65 2.244 23.665 2.755 ;
      RECT 23.645 2.236 23.65 2.753 ;
      RECT 23.635 2.235 23.645 2.745 ;
      RECT 23.605 2.232 23.635 2.724 ;
      RECT 23.53 2.227 23.605 2.669 ;
      RECT 23.515 2.223 23.53 2.615 ;
      RECT 23.505 2.223 23.515 2.51 ;
      RECT 23.49 2.223 23.505 2.443 ;
      RECT 23.475 2.223 23.485 2.433 ;
      RECT 23.42 2.222 23.475 2.43 ;
      RECT 23.375 2.22 23.42 2.433 ;
      RECT 23.347 2.22 23.36 2.436 ;
      RECT 23.261 2.224 23.347 2.438 ;
      RECT 23.175 2.23 23.261 2.443 ;
      RECT 23.155 2.234 23.175 2.445 ;
      RECT 23.153 2.235 23.155 2.444 ;
      RECT 23.067 2.237 23.153 2.443 ;
      RECT 22.981 2.242 23.067 2.44 ;
      RECT 22.895 2.247 22.981 2.437 ;
      RECT 22.745 2.25 22.825 2.433 ;
      RECT 23.405 5.015 23.575 8.305 ;
      RECT 23.405 7.315 23.81 7.645 ;
      RECT 23.405 6.475 23.81 6.805 ;
      RECT 23.521 3.225 23.57 3.559 ;
      RECT 23.521 3.225 23.575 3.558 ;
      RECT 23.435 3.225 23.575 3.557 ;
      RECT 23.21 3.333 23.58 3.555 ;
      RECT 23.435 3.225 23.605 3.548 ;
      RECT 23.405 3.237 23.61 3.539 ;
      RECT 23.39 3.255 23.615 3.536 ;
      RECT 23.205 3.339 23.615 3.463 ;
      RECT 23.2 3.346 23.615 3.423 ;
      RECT 23.215 3.312 23.615 3.536 ;
      RECT 23.376 3.258 23.58 3.555 ;
      RECT 23.29 3.278 23.615 3.536 ;
      RECT 23.39 3.252 23.61 3.539 ;
      RECT 23.16 2.576 23.35 2.77 ;
      RECT 23.155 2.578 23.35 2.769 ;
      RECT 23.15 2.582 23.365 2.766 ;
      RECT 23.165 2.575 23.365 2.766 ;
      RECT 23.15 2.685 23.37 2.761 ;
      RECT 22.445 3.185 22.536 3.483 ;
      RECT 22.44 3.187 22.615 3.478 ;
      RECT 22.445 3.185 22.615 3.478 ;
      RECT 22.44 3.191 22.635 3.476 ;
      RECT 22.44 3.246 22.675 3.475 ;
      RECT 22.44 3.281 22.69 3.469 ;
      RECT 22.44 3.315 22.7 3.459 ;
      RECT 22.43 3.195 22.635 3.31 ;
      RECT 22.43 3.215 22.65 3.31 ;
      RECT 22.43 3.198 22.64 3.31 ;
      RECT 22.655 1.966 22.66 2.028 ;
      RECT 22.65 1.888 22.655 2.051 ;
      RECT 22.645 1.845 22.65 2.062 ;
      RECT 22.64 1.835 22.645 2.074 ;
      RECT 22.635 1.835 22.64 2.083 ;
      RECT 22.61 1.835 22.635 2.115 ;
      RECT 22.605 1.835 22.61 2.148 ;
      RECT 22.59 1.835 22.605 2.173 ;
      RECT 22.58 1.835 22.59 2.2 ;
      RECT 22.575 1.835 22.58 2.213 ;
      RECT 22.57 1.835 22.575 2.228 ;
      RECT 22.56 1.835 22.57 2.243 ;
      RECT 22.555 1.835 22.56 2.263 ;
      RECT 22.53 1.835 22.555 2.298 ;
      RECT 22.485 1.835 22.53 2.343 ;
      RECT 22.475 1.835 22.485 2.356 ;
      RECT 22.39 1.92 22.475 2.363 ;
      RECT 22.355 2.042 22.39 2.372 ;
      RECT 22.35 2.082 22.355 2.376 ;
      RECT 22.33 2.105 22.35 2.378 ;
      RECT 22.325 2.135 22.33 2.381 ;
      RECT 22.315 2.147 22.325 2.382 ;
      RECT 22.27 2.17 22.315 2.387 ;
      RECT 22.23 2.2 22.27 2.395 ;
      RECT 22.195 2.212 22.23 2.401 ;
      RECT 22.19 2.217 22.195 2.405 ;
      RECT 22.12 2.227 22.19 2.412 ;
      RECT 22.08 2.237 22.12 2.422 ;
      RECT 22.06 2.242 22.08 2.428 ;
      RECT 22.05 2.246 22.06 2.433 ;
      RECT 22.045 2.249 22.05 2.436 ;
      RECT 22.035 2.25 22.045 2.437 ;
      RECT 22.01 2.252 22.035 2.441 ;
      RECT 22 2.257 22.01 2.444 ;
      RECT 21.955 2.265 22 2.445 ;
      RECT 21.83 2.27 21.955 2.445 ;
      RECT 22.385 2.567 22.405 2.749 ;
      RECT 22.336 2.552 22.385 2.748 ;
      RECT 22.25 2.567 22.405 2.746 ;
      RECT 22.235 2.567 22.405 2.745 ;
      RECT 22.2 2.545 22.37 2.73 ;
      RECT 22.27 3.565 22.285 3.774 ;
      RECT 22.27 3.573 22.29 3.773 ;
      RECT 22.215 3.573 22.29 3.772 ;
      RECT 22.195 3.577 22.295 3.77 ;
      RECT 22.175 3.527 22.215 3.769 ;
      RECT 22.12 3.585 22.3 3.767 ;
      RECT 22.085 3.542 22.215 3.765 ;
      RECT 22.081 3.545 22.27 3.764 ;
      RECT 21.995 3.553 22.27 3.762 ;
      RECT 21.995 3.597 22.305 3.755 ;
      RECT 21.985 3.69 22.305 3.753 ;
      RECT 21.995 3.609 22.31 3.738 ;
      RECT 21.995 3.63 22.325 3.708 ;
      RECT 21.995 3.657 22.33 3.678 ;
      RECT 22.12 3.535 22.215 3.767 ;
      RECT 21.75 2.58 21.755 3.118 ;
      RECT 21.555 2.91 21.56 3.105 ;
      RECT 19.855 2.575 19.87 2.955 ;
      RECT 21.92 2.575 21.925 2.745 ;
      RECT 21.915 2.575 21.92 2.755 ;
      RECT 21.91 2.575 21.915 2.768 ;
      RECT 21.885 2.575 21.91 2.81 ;
      RECT 21.86 2.575 21.885 2.883 ;
      RECT 21.845 2.575 21.86 2.935 ;
      RECT 21.84 2.575 21.845 2.965 ;
      RECT 21.815 2.575 21.84 3.005 ;
      RECT 21.8 2.575 21.815 3.06 ;
      RECT 21.795 2.575 21.8 3.093 ;
      RECT 21.77 2.575 21.795 3.113 ;
      RECT 21.755 2.575 21.77 3.119 ;
      RECT 21.685 2.61 21.75 3.115 ;
      RECT 21.635 2.665 21.685 3.11 ;
      RECT 21.625 2.697 21.635 3.108 ;
      RECT 21.62 2.722 21.625 3.108 ;
      RECT 21.6 2.795 21.62 3.108 ;
      RECT 21.59 2.875 21.6 3.107 ;
      RECT 21.575 2.905 21.59 3.107 ;
      RECT 21.56 2.91 21.575 3.106 ;
      RECT 21.5 2.912 21.555 3.103 ;
      RECT 21.47 2.917 21.5 3.099 ;
      RECT 21.468 2.92 21.47 3.098 ;
      RECT 21.382 2.922 21.468 3.095 ;
      RECT 21.296 2.928 21.382 3.089 ;
      RECT 21.21 2.933 21.296 3.083 ;
      RECT 21.137 2.938 21.21 3.084 ;
      RECT 21.051 2.944 21.137 3.092 ;
      RECT 20.965 2.95 21.051 3.101 ;
      RECT 20.945 2.954 20.965 3.106 ;
      RECT 20.898 2.956 20.945 3.109 ;
      RECT 20.812 2.961 20.898 3.115 ;
      RECT 20.726 2.966 20.812 3.124 ;
      RECT 20.64 2.972 20.726 3.132 ;
      RECT 20.555 2.97 20.64 3.141 ;
      RECT 20.551 2.965 20.555 3.145 ;
      RECT 20.465 2.96 20.551 3.137 ;
      RECT 20.401 2.951 20.465 3.125 ;
      RECT 20.315 2.942 20.401 3.112 ;
      RECT 20.291 2.935 20.315 3.103 ;
      RECT 20.205 2.929 20.291 3.09 ;
      RECT 20.165 2.922 20.205 3.076 ;
      RECT 20.16 2.912 20.165 3.072 ;
      RECT 20.15 2.9 20.16 3.071 ;
      RECT 20.13 2.87 20.15 3.068 ;
      RECT 20.075 2.79 20.13 3.062 ;
      RECT 20.055 2.709 20.075 3.057 ;
      RECT 20.035 2.667 20.055 3.053 ;
      RECT 20.01 2.62 20.035 3.047 ;
      RECT 20.005 2.595 20.01 3.044 ;
      RECT 19.97 2.575 20.005 3.039 ;
      RECT 19.961 2.575 19.97 3.032 ;
      RECT 19.875 2.575 19.961 3.002 ;
      RECT 19.87 2.575 19.875 2.965 ;
      RECT 19.835 2.575 19.855 2.887 ;
      RECT 19.83 2.617 19.835 2.852 ;
      RECT 19.825 2.692 19.83 2.808 ;
      RECT 21.275 2.497 21.45 2.745 ;
      RECT 21.275 2.497 21.455 2.743 ;
      RECT 21.27 2.529 21.455 2.703 ;
      RECT 21.3 2.47 21.47 2.69 ;
      RECT 21.265 2.547 21.47 2.623 ;
      RECT 20.575 2.01 20.745 2.185 ;
      RECT 20.575 2.01 20.917 2.177 ;
      RECT 20.575 2.01 21 2.171 ;
      RECT 20.575 2.01 21.035 2.167 ;
      RECT 20.575 2.01 21.055 2.166 ;
      RECT 20.575 2.01 21.141 2.162 ;
      RECT 21.035 1.835 21.205 2.157 ;
      RECT 20.61 1.942 21.235 2.155 ;
      RECT 20.6 1.997 21.24 2.153 ;
      RECT 20.575 2.033 21.25 2.148 ;
      RECT 20.575 2.06 21.255 2.078 ;
      RECT 20.64 1.885 21.215 2.155 ;
      RECT 20.831 1.87 21.215 2.155 ;
      RECT 20.665 1.873 21.215 2.155 ;
      RECT 20.745 1.871 20.831 2.182 ;
      RECT 20.831 1.868 21.21 2.155 ;
      RECT 21.015 1.845 21.21 2.155 ;
      RECT 20.917 1.866 21.21 2.155 ;
      RECT 21 1.86 21.015 2.168 ;
      RECT 21.15 3.225 21.155 3.425 ;
      RECT 20.615 3.29 20.66 3.425 ;
      RECT 21.185 3.225 21.205 3.398 ;
      RECT 21.155 3.225 21.185 3.413 ;
      RECT 21.09 3.225 21.15 3.45 ;
      RECT 21.075 3.225 21.09 3.48 ;
      RECT 21.06 3.225 21.075 3.493 ;
      RECT 21.04 3.225 21.06 3.508 ;
      RECT 21.035 3.225 21.04 3.517 ;
      RECT 21.025 3.229 21.035 3.522 ;
      RECT 21.01 3.239 21.025 3.533 ;
      RECT 20.985 3.255 21.01 3.543 ;
      RECT 20.975 3.269 20.985 3.545 ;
      RECT 20.955 3.281 20.975 3.542 ;
      RECT 20.925 3.302 20.955 3.536 ;
      RECT 20.915 3.314 20.925 3.531 ;
      RECT 20.905 3.312 20.915 3.528 ;
      RECT 20.89 3.311 20.905 3.523 ;
      RECT 20.885 3.31 20.89 3.518 ;
      RECT 20.85 3.308 20.885 3.508 ;
      RECT 20.83 3.305 20.85 3.49 ;
      RECT 20.82 3.303 20.83 3.485 ;
      RECT 20.81 3.302 20.82 3.48 ;
      RECT 20.775 3.3 20.81 3.468 ;
      RECT 20.72 3.296 20.775 3.448 ;
      RECT 20.71 3.294 20.72 3.433 ;
      RECT 20.705 3.294 20.71 3.428 ;
      RECT 20.66 3.292 20.705 3.425 ;
      RECT 20.565 3.29 20.615 3.429 ;
      RECT 20.555 3.291 20.565 3.434 ;
      RECT 20.495 3.298 20.555 3.448 ;
      RECT 20.47 3.306 20.495 3.468 ;
      RECT 20.46 3.31 20.47 3.48 ;
      RECT 20.455 3.311 20.46 3.485 ;
      RECT 20.44 3.313 20.455 3.488 ;
      RECT 20.425 3.315 20.44 3.493 ;
      RECT 20.42 3.315 20.425 3.496 ;
      RECT 20.375 3.32 20.42 3.507 ;
      RECT 20.37 3.324 20.375 3.519 ;
      RECT 20.345 3.32 20.37 3.523 ;
      RECT 20.335 3.316 20.345 3.527 ;
      RECT 20.325 3.315 20.335 3.531 ;
      RECT 20.31 3.305 20.325 3.537 ;
      RECT 20.305 3.293 20.31 3.541 ;
      RECT 20.3 3.29 20.305 3.542 ;
      RECT 20.295 3.287 20.3 3.544 ;
      RECT 20.28 3.275 20.295 3.543 ;
      RECT 20.265 3.257 20.28 3.54 ;
      RECT 20.245 3.236 20.265 3.533 ;
      RECT 20.18 3.225 20.245 3.505 ;
      RECT 20.176 3.225 20.18 3.484 ;
      RECT 20.09 3.225 20.176 3.454 ;
      RECT 20.075 3.225 20.09 3.41 ;
      RECT 20.65 2.325 20.655 2.56 ;
      RECT 19.78 2.241 19.785 2.445 ;
      RECT 20.36 2.27 20.365 2.425 ;
      RECT 20.28 2.25 20.285 2.425 ;
      RECT 20.95 2.392 20.965 2.745 ;
      RECT 20.876 2.377 20.95 2.745 ;
      RECT 20.79 2.36 20.876 2.745 ;
      RECT 20.78 2.35 20.79 2.743 ;
      RECT 20.775 2.348 20.78 2.738 ;
      RECT 20.76 2.346 20.775 2.724 ;
      RECT 20.69 2.338 20.76 2.664 ;
      RECT 20.67 2.329 20.69 2.598 ;
      RECT 20.665 2.326 20.67 2.578 ;
      RECT 20.655 2.325 20.665 2.568 ;
      RECT 20.645 2.325 20.65 2.552 ;
      RECT 20.635 2.324 20.645 2.542 ;
      RECT 20.625 2.322 20.635 2.53 ;
      RECT 20.61 2.319 20.625 2.51 ;
      RECT 20.6 2.317 20.61 2.495 ;
      RECT 20.58 2.314 20.6 2.483 ;
      RECT 20.575 2.312 20.58 2.473 ;
      RECT 20.55 2.31 20.575 2.46 ;
      RECT 20.52 2.305 20.55 2.445 ;
      RECT 20.44 2.296 20.52 2.436 ;
      RECT 20.395 2.285 20.44 2.429 ;
      RECT 20.375 2.276 20.395 2.426 ;
      RECT 20.365 2.271 20.375 2.425 ;
      RECT 20.32 2.265 20.36 2.425 ;
      RECT 20.305 2.257 20.32 2.425 ;
      RECT 20.285 2.252 20.305 2.425 ;
      RECT 20.265 2.249 20.28 2.425 ;
      RECT 20.182 2.248 20.265 2.424 ;
      RECT 20.096 2.247 20.182 2.42 ;
      RECT 20.01 2.245 20.096 2.417 ;
      RECT 19.957 2.244 20.01 2.419 ;
      RECT 19.871 2.243 19.957 2.428 ;
      RECT 19.785 2.242 19.871 2.44 ;
      RECT 19.765 2.241 19.78 2.448 ;
      RECT 19.685 2.24 19.765 2.46 ;
      RECT 19.66 2.24 19.685 2.473 ;
      RECT 19.635 2.24 19.66 2.488 ;
      RECT 19.63 2.24 19.635 2.51 ;
      RECT 19.625 2.24 19.63 2.528 ;
      RECT 19.62 2.24 19.625 2.545 ;
      RECT 19.615 2.24 19.62 2.558 ;
      RECT 19.61 2.24 19.615 2.568 ;
      RECT 19.57 2.24 19.61 2.653 ;
      RECT 19.555 2.24 19.57 2.738 ;
      RECT 19.545 2.241 19.555 2.75 ;
      RECT 19.51 2.246 19.545 2.755 ;
      RECT 19.47 2.255 19.51 2.755 ;
      RECT 19.455 2.265 19.47 2.755 ;
      RECT 19.45 2.275 19.455 2.755 ;
      RECT 19.43 2.302 19.45 2.755 ;
      RECT 19.38 2.385 19.43 2.755 ;
      RECT 19.375 2.447 19.38 2.755 ;
      RECT 19.365 2.46 19.375 2.755 ;
      RECT 19.355 2.482 19.365 2.755 ;
      RECT 19.345 2.507 19.355 2.75 ;
      RECT 19.34 2.545 19.345 2.743 ;
      RECT 19.33 2.655 19.34 2.738 ;
      RECT 20.725 3.576 20.74 3.835 ;
      RECT 20.725 3.591 20.745 3.834 ;
      RECT 20.641 3.591 20.745 3.832 ;
      RECT 20.641 3.605 20.75 3.831 ;
      RECT 20.555 3.647 20.755 3.828 ;
      RECT 20.55 3.59 20.74 3.823 ;
      RECT 20.55 3.661 20.76 3.82 ;
      RECT 20.545 3.692 20.76 3.818 ;
      RECT 20.55 3.689 20.775 3.808 ;
      RECT 20.545 3.735 20.79 3.793 ;
      RECT 20.545 3.763 20.795 3.778 ;
      RECT 20.555 3.565 20.725 3.828 ;
      RECT 20.315 2.575 20.485 2.745 ;
      RECT 20.28 2.575 20.485 2.74 ;
      RECT 20.27 2.575 20.485 2.733 ;
      RECT 20.265 2.56 20.435 2.73 ;
      RECT 19.095 3.097 19.36 3.54 ;
      RECT 19.09 3.068 19.305 3.538 ;
      RECT 19.085 3.222 19.365 3.533 ;
      RECT 19.09 3.117 19.365 3.533 ;
      RECT 19.09 3.128 19.375 3.52 ;
      RECT 19.09 3.075 19.335 3.538 ;
      RECT 19.095 3.062 19.305 3.54 ;
      RECT 19.095 3.06 19.255 3.54 ;
      RECT 19.196 3.052 19.255 3.54 ;
      RECT 19.11 3.053 19.255 3.54 ;
      RECT 19.196 3.051 19.245 3.54 ;
      RECT 19 1.866 19.175 2.165 ;
      RECT 19.05 1.828 19.175 2.165 ;
      RECT 19.035 1.83 19.261 2.157 ;
      RECT 19.035 1.833 19.3 2.144 ;
      RECT 19.035 1.834 19.31 2.13 ;
      RECT 18.99 1.885 19.31 2.12 ;
      RECT 19.035 1.835 19.315 2.115 ;
      RECT 18.99 2.045 19.32 2.105 ;
      RECT 18.975 1.905 19.315 2.045 ;
      RECT 18.97 1.921 19.315 1.985 ;
      RECT 19.015 1.845 19.315 2.115 ;
      RECT 19.05 1.826 19.136 2.165 ;
      RECT 17.51 5.02 17.68 6.49 ;
      RECT 17.51 6.315 17.685 6.485 ;
      RECT 17.14 1.74 17.31 2.93 ;
      RECT 17.14 1.74 17.61 1.91 ;
      RECT 17.14 6.97 17.61 7.14 ;
      RECT 17.14 5.95 17.31 7.14 ;
      RECT 16.15 1.74 16.32 2.93 ;
      RECT 16.15 1.74 16.62 1.91 ;
      RECT 16.15 6.97 16.62 7.14 ;
      RECT 16.15 5.95 16.32 7.14 ;
      RECT 14.3 2.635 14.47 3.865 ;
      RECT 14.355 0.855 14.525 2.805 ;
      RECT 14.3 0.575 14.47 1.025 ;
      RECT 14.3 7.855 14.47 8.305 ;
      RECT 14.355 6.075 14.525 8.025 ;
      RECT 14.3 5.015 14.47 6.245 ;
      RECT 13.78 0.575 13.95 3.865 ;
      RECT 13.78 2.075 14.185 2.405 ;
      RECT 13.78 1.235 14.185 1.565 ;
      RECT 13.78 5.015 13.95 8.305 ;
      RECT 13.78 7.315 14.185 7.645 ;
      RECT 13.78 6.475 14.185 6.805 ;
      RECT 11.705 3.126 11.71 3.298 ;
      RECT 11.7 3.119 11.705 3.388 ;
      RECT 11.695 3.113 11.7 3.407 ;
      RECT 11.675 3.107 11.695 3.417 ;
      RECT 11.66 3.102 11.675 3.425 ;
      RECT 11.623 3.096 11.66 3.423 ;
      RECT 11.537 3.082 11.623 3.419 ;
      RECT 11.451 3.064 11.537 3.414 ;
      RECT 11.365 3.045 11.451 3.408 ;
      RECT 11.335 3.033 11.365 3.404 ;
      RECT 11.315 3.027 11.335 3.403 ;
      RECT 11.25 3.025 11.315 3.401 ;
      RECT 11.235 3.025 11.25 3.393 ;
      RECT 11.22 3.025 11.235 3.38 ;
      RECT 11.215 3.025 11.22 3.37 ;
      RECT 11.2 3.025 11.215 3.348 ;
      RECT 11.185 3.025 11.2 3.315 ;
      RECT 11.18 3.025 11.185 3.293 ;
      RECT 11.17 3.025 11.18 3.275 ;
      RECT 11.155 3.025 11.17 3.253 ;
      RECT 11.135 3.025 11.155 3.215 ;
      RECT 11.485 2.31 11.52 2.749 ;
      RECT 11.485 2.31 11.525 2.748 ;
      RECT 11.43 2.37 11.525 2.747 ;
      RECT 11.295 2.542 11.525 2.746 ;
      RECT 11.405 2.42 11.525 2.746 ;
      RECT 11.295 2.542 11.55 2.736 ;
      RECT 11.35 2.487 11.63 2.653 ;
      RECT 11.525 2.281 11.53 2.744 ;
      RECT 11.38 2.457 11.67 2.53 ;
      RECT 11.395 2.44 11.525 2.746 ;
      RECT 11.53 2.28 11.7 2.468 ;
      RECT 11.52 2.283 11.7 2.468 ;
      RECT 11.025 2.16 11.195 2.47 ;
      RECT 11.025 2.16 11.2 2.443 ;
      RECT 11.025 2.16 11.205 2.42 ;
      RECT 11.025 2.16 11.215 2.37 ;
      RECT 11.02 2.265 11.215 2.34 ;
      RECT 11.055 1.835 11.225 2.313 ;
      RECT 11.055 1.835 11.24 2.234 ;
      RECT 11.045 2.045 11.24 2.234 ;
      RECT 11.055 1.845 11.25 2.149 ;
      RECT 10.985 2.587 10.99 2.79 ;
      RECT 10.975 2.575 10.985 2.9 ;
      RECT 10.95 2.575 10.975 2.94 ;
      RECT 10.87 2.575 10.95 3.025 ;
      RECT 10.86 2.575 10.87 3.095 ;
      RECT 10.835 2.575 10.86 3.118 ;
      RECT 10.815 2.575 10.835 3.153 ;
      RECT 10.77 2.585 10.815 3.196 ;
      RECT 10.76 2.597 10.77 3.233 ;
      RECT 10.74 2.611 10.76 3.253 ;
      RECT 10.73 2.629 10.74 3.269 ;
      RECT 10.715 2.655 10.73 3.279 ;
      RECT 10.7 2.696 10.715 3.293 ;
      RECT 10.69 2.731 10.7 3.303 ;
      RECT 10.685 2.747 10.69 3.308 ;
      RECT 10.675 2.762 10.685 3.313 ;
      RECT 10.655 2.805 10.675 3.323 ;
      RECT 10.635 2.842 10.655 3.336 ;
      RECT 10.6 2.865 10.635 3.354 ;
      RECT 10.59 2.879 10.6 3.37 ;
      RECT 10.57 2.889 10.59 3.38 ;
      RECT 10.565 2.898 10.57 3.388 ;
      RECT 10.555 2.905 10.565 3.395 ;
      RECT 10.545 2.912 10.555 3.403 ;
      RECT 10.53 2.922 10.545 3.411 ;
      RECT 10.52 2.936 10.53 3.421 ;
      RECT 10.51 2.948 10.52 3.433 ;
      RECT 10.495 2.97 10.51 3.446 ;
      RECT 10.485 2.992 10.495 3.457 ;
      RECT 10.475 3.012 10.485 3.466 ;
      RECT 10.47 3.027 10.475 3.473 ;
      RECT 10.44 3.06 10.47 3.487 ;
      RECT 10.43 3.095 10.44 3.502 ;
      RECT 10.425 3.102 10.43 3.508 ;
      RECT 10.405 3.117 10.425 3.515 ;
      RECT 10.4 3.132 10.405 3.523 ;
      RECT 10.395 3.141 10.4 3.528 ;
      RECT 10.38 3.147 10.395 3.535 ;
      RECT 10.375 3.153 10.38 3.543 ;
      RECT 10.37 3.157 10.375 3.55 ;
      RECT 10.365 3.161 10.37 3.56 ;
      RECT 10.355 3.166 10.365 3.57 ;
      RECT 10.335 3.177 10.355 3.598 ;
      RECT 10.32 3.189 10.335 3.625 ;
      RECT 10.3 3.202 10.32 3.65 ;
      RECT 10.28 3.217 10.3 3.674 ;
      RECT 10.265 3.232 10.28 3.689 ;
      RECT 10.26 3.243 10.265 3.698 ;
      RECT 10.195 3.288 10.26 3.708 ;
      RECT 10.16 3.347 10.195 3.721 ;
      RECT 10.155 3.37 10.16 3.727 ;
      RECT 10.15 3.377 10.155 3.729 ;
      RECT 10.135 3.387 10.15 3.732 ;
      RECT 10.105 3.412 10.135 3.736 ;
      RECT 10.1 3.43 10.105 3.74 ;
      RECT 10.095 3.437 10.1 3.741 ;
      RECT 10.075 3.445 10.095 3.745 ;
      RECT 10.065 3.452 10.075 3.749 ;
      RECT 10.021 3.463 10.065 3.756 ;
      RECT 9.935 3.491 10.021 3.772 ;
      RECT 9.875 3.515 9.935 3.79 ;
      RECT 9.83 3.525 9.875 3.804 ;
      RECT 9.771 3.533 9.83 3.818 ;
      RECT 9.685 3.54 9.771 3.837 ;
      RECT 9.66 3.545 9.685 3.852 ;
      RECT 9.58 3.548 9.66 3.855 ;
      RECT 9.5 3.552 9.58 3.842 ;
      RECT 9.491 3.555 9.5 3.827 ;
      RECT 9.405 3.555 9.491 3.812 ;
      RECT 9.345 3.557 9.405 3.789 ;
      RECT 9.341 3.56 9.345 3.779 ;
      RECT 9.255 3.56 9.341 3.764 ;
      RECT 9.18 3.56 9.255 3.74 ;
      RECT 10.495 2.569 10.505 2.745 ;
      RECT 10.45 2.536 10.495 2.745 ;
      RECT 10.405 2.487 10.45 2.745 ;
      RECT 10.375 2.457 10.405 2.746 ;
      RECT 10.37 2.44 10.375 2.747 ;
      RECT 10.345 2.42 10.37 2.748 ;
      RECT 10.33 2.395 10.345 2.749 ;
      RECT 10.325 2.382 10.33 2.75 ;
      RECT 10.32 2.376 10.325 2.748 ;
      RECT 10.315 2.368 10.32 2.742 ;
      RECT 10.29 2.36 10.315 2.722 ;
      RECT 10.27 2.349 10.29 2.693 ;
      RECT 10.24 2.334 10.27 2.664 ;
      RECT 10.22 2.32 10.24 2.636 ;
      RECT 10.21 2.314 10.22 2.615 ;
      RECT 10.205 2.311 10.21 2.598 ;
      RECT 10.2 2.308 10.205 2.583 ;
      RECT 10.185 2.303 10.2 2.548 ;
      RECT 10.18 2.299 10.185 2.515 ;
      RECT 10.16 2.294 10.18 2.491 ;
      RECT 10.13 2.286 10.16 2.456 ;
      RECT 10.115 2.28 10.13 2.433 ;
      RECT 10.075 2.273 10.115 2.418 ;
      RECT 10.05 2.265 10.075 2.398 ;
      RECT 10.03 2.26 10.05 2.388 ;
      RECT 9.995 2.254 10.03 2.383 ;
      RECT 9.95 2.245 9.995 2.382 ;
      RECT 9.92 2.241 9.95 2.384 ;
      RECT 9.835 2.249 9.92 2.388 ;
      RECT 9.765 2.26 9.835 2.41 ;
      RECT 9.752 2.266 9.765 2.433 ;
      RECT 9.666 2.273 9.752 2.455 ;
      RECT 9.58 2.285 9.666 2.492 ;
      RECT 9.58 2.662 9.59 2.9 ;
      RECT 9.575 2.291 9.58 2.515 ;
      RECT 9.57 2.547 9.58 2.9 ;
      RECT 9.57 2.292 9.575 2.52 ;
      RECT 9.565 2.293 9.57 2.9 ;
      RECT 9.541 2.295 9.565 2.901 ;
      RECT 9.455 2.303 9.541 2.903 ;
      RECT 9.435 2.317 9.455 2.906 ;
      RECT 9.43 2.345 9.435 2.907 ;
      RECT 9.425 2.357 9.43 2.908 ;
      RECT 9.42 2.372 9.425 2.909 ;
      RECT 9.41 2.402 9.42 2.91 ;
      RECT 9.405 2.44 9.41 2.908 ;
      RECT 9.4 2.46 9.405 2.903 ;
      RECT 9.385 2.495 9.4 2.888 ;
      RECT 9.375 2.547 9.385 2.868 ;
      RECT 9.37 2.577 9.375 2.856 ;
      RECT 9.355 2.59 9.37 2.839 ;
      RECT 9.33 2.594 9.355 2.806 ;
      RECT 9.315 2.592 9.33 2.783 ;
      RECT 9.3 2.591 9.315 2.78 ;
      RECT 9.24 2.589 9.3 2.778 ;
      RECT 9.23 2.587 9.24 2.773 ;
      RECT 9.19 2.586 9.23 2.77 ;
      RECT 9.12 2.583 9.19 2.768 ;
      RECT 9.065 2.581 9.12 2.763 ;
      RECT 8.995 2.575 9.065 2.758 ;
      RECT 8.986 2.575 8.995 2.755 ;
      RECT 8.9 2.575 8.986 2.75 ;
      RECT 8.895 2.575 8.9 2.745 ;
      RECT 10.2 1.81 10.375 2.16 ;
      RECT 10.2 1.825 10.385 2.158 ;
      RECT 10.175 1.775 10.32 2.155 ;
      RECT 10.155 1.776 10.32 2.148 ;
      RECT 10.145 1.777 10.33 2.143 ;
      RECT 10.115 1.778 10.33 2.13 ;
      RECT 10.065 1.779 10.33 2.106 ;
      RECT 10.06 1.781 10.33 2.091 ;
      RECT 10.06 1.847 10.39 2.085 ;
      RECT 10.04 1.788 10.345 2.065 ;
      RECT 10.03 1.797 10.355 1.92 ;
      RECT 10.04 1.792 10.355 2.065 ;
      RECT 10.06 1.782 10.345 2.091 ;
      RECT 9.645 3.107 9.815 3.395 ;
      RECT 9.64 3.125 9.825 3.39 ;
      RECT 9.605 3.133 9.89 3.31 ;
      RECT 9.605 3.133 9.976 3.3 ;
      RECT 9.605 3.133 10.03 3.246 ;
      RECT 9.89 3.03 10.06 3.214 ;
      RECT 9.605 3.185 10.065 3.202 ;
      RECT 9.59 3.155 10.06 3.198 ;
      RECT 9.85 3.037 9.89 3.349 ;
      RECT 9.73 3.074 10.06 3.214 ;
      RECT 9.825 3.049 9.85 3.375 ;
      RECT 9.815 3.056 10.06 3.214 ;
      RECT 9.946 2.52 10.015 2.779 ;
      RECT 9.946 2.575 10.02 2.778 ;
      RECT 9.86 2.575 10.02 2.777 ;
      RECT 9.855 2.575 10.025 2.77 ;
      RECT 9.845 2.52 10.015 2.765 ;
      RECT 9.225 1.819 9.4 2.12 ;
      RECT 9.21 1.807 9.225 2.105 ;
      RECT 9.18 1.806 9.21 2.058 ;
      RECT 9.18 1.824 9.405 2.053 ;
      RECT 9.165 1.808 9.225 2.018 ;
      RECT 9.16 1.83 9.415 1.918 ;
      RECT 9.16 1.813 9.311 1.918 ;
      RECT 9.16 1.815 9.315 1.918 ;
      RECT 9.165 1.811 9.311 2.018 ;
      RECT 9.27 3.047 9.275 3.395 ;
      RECT 9.26 3.037 9.27 3.401 ;
      RECT 9.225 3.027 9.26 3.403 ;
      RECT 9.187 3.022 9.225 3.407 ;
      RECT 9.101 3.015 9.187 3.414 ;
      RECT 9.015 3.005 9.101 3.424 ;
      RECT 8.97 3 9.015 3.432 ;
      RECT 8.966 3 8.97 3.436 ;
      RECT 8.88 3 8.966 3.443 ;
      RECT 8.865 3 8.88 3.443 ;
      RECT 8.855 2.998 8.865 3.415 ;
      RECT 8.845 2.994 8.855 3.358 ;
      RECT 8.825 2.988 8.845 3.29 ;
      RECT 8.82 2.984 8.825 3.238 ;
      RECT 8.81 2.983 8.82 3.205 ;
      RECT 8.76 2.981 8.81 3.19 ;
      RECT 8.735 2.979 8.76 3.185 ;
      RECT 8.692 2.977 8.735 3.181 ;
      RECT 8.606 2.973 8.692 3.169 ;
      RECT 8.52 2.968 8.606 3.153 ;
      RECT 8.49 2.965 8.52 3.14 ;
      RECT 8.465 2.964 8.49 3.128 ;
      RECT 8.46 2.964 8.465 3.118 ;
      RECT 8.42 2.963 8.46 3.11 ;
      RECT 8.405 2.962 8.42 3.103 ;
      RECT 8.355 2.961 8.405 3.095 ;
      RECT 8.353 2.96 8.355 3.09 ;
      RECT 8.267 2.958 8.353 3.09 ;
      RECT 8.181 2.953 8.267 3.09 ;
      RECT 8.095 2.949 8.181 3.09 ;
      RECT 8.046 2.945 8.095 3.088 ;
      RECT 7.96 2.942 8.046 3.083 ;
      RECT 7.937 2.939 7.96 3.079 ;
      RECT 7.851 2.936 7.937 3.074 ;
      RECT 7.765 2.932 7.851 3.065 ;
      RECT 7.74 2.925 7.765 3.06 ;
      RECT 7.68 2.89 7.74 3.057 ;
      RECT 7.66 2.815 7.68 3.054 ;
      RECT 7.655 2.757 7.66 3.053 ;
      RECT 7.63 2.697 7.655 3.052 ;
      RECT 7.555 2.575 7.63 3.048 ;
      RECT 7.545 2.575 7.555 3.04 ;
      RECT 7.53 2.575 7.545 3.03 ;
      RECT 7.515 2.575 7.53 3 ;
      RECT 7.5 2.575 7.515 2.945 ;
      RECT 7.485 2.575 7.5 2.883 ;
      RECT 7.46 2.575 7.485 2.808 ;
      RECT 7.455 2.575 7.46 2.758 ;
      RECT 8.8 2.12 8.82 2.429 ;
      RECT 8.786 2.122 8.835 2.426 ;
      RECT 8.786 2.127 8.855 2.417 ;
      RECT 8.7 2.125 8.835 2.411 ;
      RECT 8.7 2.133 8.89 2.394 ;
      RECT 8.665 2.135 8.89 2.393 ;
      RECT 8.635 2.143 8.89 2.384 ;
      RECT 8.625 2.148 8.91 2.37 ;
      RECT 8.665 2.138 8.91 2.37 ;
      RECT 8.665 2.141 8.92 2.358 ;
      RECT 8.635 2.143 8.93 2.345 ;
      RECT 8.635 2.147 8.94 2.288 ;
      RECT 8.625 2.152 8.945 2.203 ;
      RECT 8.786 2.12 8.82 2.426 ;
      RECT 8.665 7.855 8.835 8.305 ;
      RECT 8.72 6.075 8.89 8.025 ;
      RECT 8.665 5.015 8.835 6.245 ;
      RECT 8.225 2.223 8.23 2.435 ;
      RECT 8.1 2.22 8.115 2.435 ;
      RECT 7.565 2.25 7.635 2.435 ;
      RECT 7.45 2.25 7.485 2.43 ;
      RECT 8.571 2.552 8.59 2.746 ;
      RECT 8.485 2.507 8.571 2.747 ;
      RECT 8.475 2.46 8.485 2.749 ;
      RECT 8.47 2.44 8.475 2.75 ;
      RECT 8.45 2.405 8.47 2.751 ;
      RECT 8.435 2.355 8.45 2.752 ;
      RECT 8.415 2.292 8.435 2.753 ;
      RECT 8.405 2.255 8.415 2.754 ;
      RECT 8.39 2.244 8.405 2.755 ;
      RECT 8.385 2.236 8.39 2.753 ;
      RECT 8.375 2.235 8.385 2.745 ;
      RECT 8.345 2.232 8.375 2.724 ;
      RECT 8.27 2.227 8.345 2.669 ;
      RECT 8.255 2.223 8.27 2.615 ;
      RECT 8.245 2.223 8.255 2.51 ;
      RECT 8.23 2.223 8.245 2.443 ;
      RECT 8.215 2.223 8.225 2.433 ;
      RECT 8.16 2.222 8.215 2.43 ;
      RECT 8.115 2.22 8.16 2.433 ;
      RECT 8.087 2.22 8.1 2.436 ;
      RECT 8.001 2.224 8.087 2.438 ;
      RECT 7.915 2.23 8.001 2.443 ;
      RECT 7.895 2.234 7.915 2.445 ;
      RECT 7.893 2.235 7.895 2.444 ;
      RECT 7.807 2.237 7.893 2.443 ;
      RECT 7.721 2.242 7.807 2.44 ;
      RECT 7.635 2.247 7.721 2.437 ;
      RECT 7.485 2.25 7.565 2.433 ;
      RECT 8.145 5.015 8.315 8.305 ;
      RECT 8.145 7.315 8.55 7.645 ;
      RECT 8.145 6.475 8.55 6.805 ;
      RECT 8.261 3.225 8.31 3.559 ;
      RECT 8.261 3.225 8.315 3.558 ;
      RECT 8.175 3.225 8.315 3.557 ;
      RECT 7.95 3.333 8.32 3.555 ;
      RECT 8.175 3.225 8.345 3.548 ;
      RECT 8.145 3.237 8.35 3.539 ;
      RECT 8.13 3.255 8.355 3.536 ;
      RECT 7.945 3.339 8.355 3.463 ;
      RECT 7.94 3.346 8.355 3.423 ;
      RECT 7.955 3.312 8.355 3.536 ;
      RECT 8.116 3.258 8.32 3.555 ;
      RECT 8.03 3.278 8.355 3.536 ;
      RECT 8.13 3.252 8.35 3.539 ;
      RECT 7.9 2.576 8.09 2.77 ;
      RECT 7.895 2.578 8.09 2.769 ;
      RECT 7.89 2.582 8.105 2.766 ;
      RECT 7.905 2.575 8.105 2.766 ;
      RECT 7.89 2.685 8.11 2.761 ;
      RECT 7.185 3.185 7.276 3.483 ;
      RECT 7.18 3.187 7.355 3.478 ;
      RECT 7.185 3.185 7.355 3.478 ;
      RECT 7.18 3.191 7.375 3.476 ;
      RECT 7.18 3.246 7.415 3.475 ;
      RECT 7.18 3.281 7.43 3.469 ;
      RECT 7.18 3.315 7.44 3.459 ;
      RECT 7.17 3.195 7.375 3.31 ;
      RECT 7.17 3.215 7.39 3.31 ;
      RECT 7.17 3.198 7.38 3.31 ;
      RECT 7.395 1.966 7.4 2.028 ;
      RECT 7.39 1.888 7.395 2.051 ;
      RECT 7.385 1.845 7.39 2.062 ;
      RECT 7.38 1.835 7.385 2.074 ;
      RECT 7.375 1.835 7.38 2.083 ;
      RECT 7.35 1.835 7.375 2.115 ;
      RECT 7.345 1.835 7.35 2.148 ;
      RECT 7.33 1.835 7.345 2.173 ;
      RECT 7.32 1.835 7.33 2.2 ;
      RECT 7.315 1.835 7.32 2.213 ;
      RECT 7.31 1.835 7.315 2.228 ;
      RECT 7.3 1.835 7.31 2.243 ;
      RECT 7.295 1.835 7.3 2.263 ;
      RECT 7.27 1.835 7.295 2.298 ;
      RECT 7.225 1.835 7.27 2.343 ;
      RECT 7.215 1.835 7.225 2.356 ;
      RECT 7.13 1.92 7.215 2.363 ;
      RECT 7.095 2.042 7.13 2.372 ;
      RECT 7.09 2.082 7.095 2.376 ;
      RECT 7.07 2.105 7.09 2.378 ;
      RECT 7.065 2.135 7.07 2.381 ;
      RECT 7.055 2.147 7.065 2.382 ;
      RECT 7.01 2.17 7.055 2.387 ;
      RECT 6.97 2.2 7.01 2.395 ;
      RECT 6.935 2.212 6.97 2.401 ;
      RECT 6.93 2.217 6.935 2.405 ;
      RECT 6.86 2.227 6.93 2.412 ;
      RECT 6.82 2.237 6.86 2.422 ;
      RECT 6.8 2.242 6.82 2.428 ;
      RECT 6.79 2.246 6.8 2.433 ;
      RECT 6.785 2.249 6.79 2.436 ;
      RECT 6.775 2.25 6.785 2.437 ;
      RECT 6.75 2.252 6.775 2.441 ;
      RECT 6.74 2.257 6.75 2.444 ;
      RECT 6.695 2.265 6.74 2.445 ;
      RECT 6.57 2.27 6.695 2.445 ;
      RECT 7.125 2.567 7.145 2.749 ;
      RECT 7.076 2.552 7.125 2.748 ;
      RECT 6.99 2.567 7.145 2.746 ;
      RECT 6.975 2.567 7.145 2.745 ;
      RECT 6.94 2.545 7.11 2.73 ;
      RECT 7.01 3.565 7.025 3.774 ;
      RECT 7.01 3.573 7.03 3.773 ;
      RECT 6.955 3.573 7.03 3.772 ;
      RECT 6.935 3.577 7.035 3.77 ;
      RECT 6.915 3.527 6.955 3.769 ;
      RECT 6.86 3.585 7.04 3.767 ;
      RECT 6.825 3.542 6.955 3.765 ;
      RECT 6.821 3.545 7.01 3.764 ;
      RECT 6.735 3.553 7.01 3.762 ;
      RECT 6.735 3.597 7.045 3.755 ;
      RECT 6.725 3.69 7.045 3.753 ;
      RECT 6.735 3.609 7.05 3.738 ;
      RECT 6.735 3.63 7.065 3.708 ;
      RECT 6.735 3.657 7.07 3.678 ;
      RECT 6.86 3.535 6.955 3.767 ;
      RECT 6.49 2.58 6.495 3.118 ;
      RECT 6.295 2.91 6.3 3.105 ;
      RECT 4.595 2.575 4.61 2.955 ;
      RECT 6.66 2.575 6.665 2.745 ;
      RECT 6.655 2.575 6.66 2.755 ;
      RECT 6.65 2.575 6.655 2.768 ;
      RECT 6.625 2.575 6.65 2.81 ;
      RECT 6.6 2.575 6.625 2.883 ;
      RECT 6.585 2.575 6.6 2.935 ;
      RECT 6.58 2.575 6.585 2.965 ;
      RECT 6.555 2.575 6.58 3.005 ;
      RECT 6.54 2.575 6.555 3.06 ;
      RECT 6.535 2.575 6.54 3.093 ;
      RECT 6.51 2.575 6.535 3.113 ;
      RECT 6.495 2.575 6.51 3.119 ;
      RECT 6.425 2.61 6.49 3.115 ;
      RECT 6.375 2.665 6.425 3.11 ;
      RECT 6.365 2.697 6.375 3.108 ;
      RECT 6.36 2.722 6.365 3.108 ;
      RECT 6.34 2.795 6.36 3.108 ;
      RECT 6.33 2.875 6.34 3.107 ;
      RECT 6.315 2.905 6.33 3.107 ;
      RECT 6.3 2.91 6.315 3.106 ;
      RECT 6.24 2.912 6.295 3.103 ;
      RECT 6.21 2.917 6.24 3.099 ;
      RECT 6.208 2.92 6.21 3.098 ;
      RECT 6.122 2.922 6.208 3.095 ;
      RECT 6.036 2.928 6.122 3.089 ;
      RECT 5.95 2.933 6.036 3.083 ;
      RECT 5.877 2.938 5.95 3.084 ;
      RECT 5.791 2.944 5.877 3.092 ;
      RECT 5.705 2.95 5.791 3.101 ;
      RECT 5.685 2.954 5.705 3.106 ;
      RECT 5.638 2.956 5.685 3.109 ;
      RECT 5.552 2.961 5.638 3.115 ;
      RECT 5.466 2.966 5.552 3.124 ;
      RECT 5.38 2.972 5.466 3.132 ;
      RECT 5.295 2.97 5.38 3.141 ;
      RECT 5.291 2.965 5.295 3.145 ;
      RECT 5.205 2.96 5.291 3.137 ;
      RECT 5.141 2.951 5.205 3.125 ;
      RECT 5.055 2.942 5.141 3.112 ;
      RECT 5.031 2.935 5.055 3.103 ;
      RECT 4.945 2.929 5.031 3.09 ;
      RECT 4.905 2.922 4.945 3.076 ;
      RECT 4.9 2.912 4.905 3.072 ;
      RECT 4.89 2.9 4.9 3.071 ;
      RECT 4.87 2.87 4.89 3.068 ;
      RECT 4.815 2.79 4.87 3.062 ;
      RECT 4.795 2.709 4.815 3.057 ;
      RECT 4.775 2.667 4.795 3.053 ;
      RECT 4.75 2.62 4.775 3.047 ;
      RECT 4.745 2.595 4.75 3.044 ;
      RECT 4.71 2.575 4.745 3.039 ;
      RECT 4.701 2.575 4.71 3.032 ;
      RECT 4.615 2.575 4.701 3.002 ;
      RECT 4.61 2.575 4.615 2.965 ;
      RECT 4.575 2.575 4.595 2.887 ;
      RECT 4.57 2.617 4.575 2.852 ;
      RECT 4.565 2.692 4.57 2.808 ;
      RECT 6.015 2.497 6.19 2.745 ;
      RECT 6.015 2.497 6.195 2.743 ;
      RECT 6.01 2.529 6.195 2.703 ;
      RECT 6.04 2.47 6.21 2.69 ;
      RECT 6.005 2.547 6.21 2.623 ;
      RECT 5.315 2.01 5.485 2.185 ;
      RECT 5.315 2.01 5.657 2.177 ;
      RECT 5.315 2.01 5.74 2.171 ;
      RECT 5.315 2.01 5.775 2.167 ;
      RECT 5.315 2.01 5.795 2.166 ;
      RECT 5.315 2.01 5.881 2.162 ;
      RECT 5.775 1.835 5.945 2.157 ;
      RECT 5.35 1.942 5.975 2.155 ;
      RECT 5.34 1.997 5.98 2.153 ;
      RECT 5.315 2.033 5.99 2.148 ;
      RECT 5.315 2.06 5.995 2.078 ;
      RECT 5.38 1.885 5.955 2.155 ;
      RECT 5.571 1.87 5.955 2.155 ;
      RECT 5.405 1.873 5.955 2.155 ;
      RECT 5.485 1.871 5.571 2.182 ;
      RECT 5.571 1.868 5.95 2.155 ;
      RECT 5.755 1.845 5.95 2.155 ;
      RECT 5.657 1.866 5.95 2.155 ;
      RECT 5.74 1.86 5.755 2.168 ;
      RECT 5.89 3.225 5.895 3.425 ;
      RECT 5.355 3.29 5.4 3.425 ;
      RECT 5.925 3.225 5.945 3.398 ;
      RECT 5.895 3.225 5.925 3.413 ;
      RECT 5.83 3.225 5.89 3.45 ;
      RECT 5.815 3.225 5.83 3.48 ;
      RECT 5.8 3.225 5.815 3.493 ;
      RECT 5.78 3.225 5.8 3.508 ;
      RECT 5.775 3.225 5.78 3.517 ;
      RECT 5.765 3.229 5.775 3.522 ;
      RECT 5.75 3.239 5.765 3.533 ;
      RECT 5.725 3.255 5.75 3.543 ;
      RECT 5.715 3.269 5.725 3.545 ;
      RECT 5.695 3.281 5.715 3.542 ;
      RECT 5.665 3.302 5.695 3.536 ;
      RECT 5.655 3.314 5.665 3.531 ;
      RECT 5.645 3.312 5.655 3.528 ;
      RECT 5.63 3.311 5.645 3.523 ;
      RECT 5.625 3.31 5.63 3.518 ;
      RECT 5.59 3.308 5.625 3.508 ;
      RECT 5.57 3.305 5.59 3.49 ;
      RECT 5.56 3.303 5.57 3.485 ;
      RECT 5.55 3.302 5.56 3.48 ;
      RECT 5.515 3.3 5.55 3.468 ;
      RECT 5.46 3.296 5.515 3.448 ;
      RECT 5.45 3.294 5.46 3.433 ;
      RECT 5.445 3.294 5.45 3.428 ;
      RECT 5.4 3.292 5.445 3.425 ;
      RECT 5.305 3.29 5.355 3.429 ;
      RECT 5.295 3.291 5.305 3.434 ;
      RECT 5.235 3.298 5.295 3.448 ;
      RECT 5.21 3.306 5.235 3.468 ;
      RECT 5.2 3.31 5.21 3.48 ;
      RECT 5.195 3.311 5.2 3.485 ;
      RECT 5.18 3.313 5.195 3.488 ;
      RECT 5.165 3.315 5.18 3.493 ;
      RECT 5.16 3.315 5.165 3.496 ;
      RECT 5.115 3.32 5.16 3.507 ;
      RECT 5.11 3.324 5.115 3.519 ;
      RECT 5.085 3.32 5.11 3.523 ;
      RECT 5.075 3.316 5.085 3.527 ;
      RECT 5.065 3.315 5.075 3.531 ;
      RECT 5.05 3.305 5.065 3.537 ;
      RECT 5.045 3.293 5.05 3.541 ;
      RECT 5.04 3.29 5.045 3.542 ;
      RECT 5.035 3.287 5.04 3.544 ;
      RECT 5.02 3.275 5.035 3.543 ;
      RECT 5.005 3.257 5.02 3.54 ;
      RECT 4.985 3.236 5.005 3.533 ;
      RECT 4.92 3.225 4.985 3.505 ;
      RECT 4.916 3.225 4.92 3.484 ;
      RECT 4.83 3.225 4.916 3.454 ;
      RECT 4.815 3.225 4.83 3.41 ;
      RECT 5.39 2.325 5.395 2.56 ;
      RECT 4.52 2.241 4.525 2.445 ;
      RECT 5.1 2.27 5.105 2.425 ;
      RECT 5.02 2.25 5.025 2.425 ;
      RECT 5.69 2.392 5.705 2.745 ;
      RECT 5.616 2.377 5.69 2.745 ;
      RECT 5.53 2.36 5.616 2.745 ;
      RECT 5.52 2.35 5.53 2.743 ;
      RECT 5.515 2.348 5.52 2.738 ;
      RECT 5.5 2.346 5.515 2.724 ;
      RECT 5.43 2.338 5.5 2.664 ;
      RECT 5.41 2.329 5.43 2.598 ;
      RECT 5.405 2.326 5.41 2.578 ;
      RECT 5.395 2.325 5.405 2.568 ;
      RECT 5.385 2.325 5.39 2.552 ;
      RECT 5.375 2.324 5.385 2.542 ;
      RECT 5.365 2.322 5.375 2.53 ;
      RECT 5.35 2.319 5.365 2.51 ;
      RECT 5.34 2.317 5.35 2.495 ;
      RECT 5.32 2.314 5.34 2.483 ;
      RECT 5.315 2.312 5.32 2.473 ;
      RECT 5.29 2.31 5.315 2.46 ;
      RECT 5.26 2.305 5.29 2.445 ;
      RECT 5.18 2.296 5.26 2.436 ;
      RECT 5.135 2.285 5.18 2.429 ;
      RECT 5.115 2.276 5.135 2.426 ;
      RECT 5.105 2.271 5.115 2.425 ;
      RECT 5.06 2.265 5.1 2.425 ;
      RECT 5.045 2.257 5.06 2.425 ;
      RECT 5.025 2.252 5.045 2.425 ;
      RECT 5.005 2.249 5.02 2.425 ;
      RECT 4.922 2.248 5.005 2.424 ;
      RECT 4.836 2.247 4.922 2.42 ;
      RECT 4.75 2.245 4.836 2.417 ;
      RECT 4.697 2.244 4.75 2.419 ;
      RECT 4.611 2.243 4.697 2.428 ;
      RECT 4.525 2.242 4.611 2.44 ;
      RECT 4.505 2.241 4.52 2.448 ;
      RECT 4.425 2.24 4.505 2.46 ;
      RECT 4.4 2.24 4.425 2.473 ;
      RECT 4.375 2.24 4.4 2.488 ;
      RECT 4.37 2.24 4.375 2.51 ;
      RECT 4.365 2.24 4.37 2.528 ;
      RECT 4.36 2.24 4.365 2.545 ;
      RECT 4.355 2.24 4.36 2.558 ;
      RECT 4.35 2.24 4.355 2.568 ;
      RECT 4.31 2.24 4.35 2.653 ;
      RECT 4.295 2.24 4.31 2.738 ;
      RECT 4.285 2.241 4.295 2.75 ;
      RECT 4.25 2.246 4.285 2.755 ;
      RECT 4.21 2.255 4.25 2.755 ;
      RECT 4.195 2.265 4.21 2.755 ;
      RECT 4.19 2.275 4.195 2.755 ;
      RECT 4.17 2.302 4.19 2.755 ;
      RECT 4.12 2.385 4.17 2.755 ;
      RECT 4.115 2.447 4.12 2.755 ;
      RECT 4.105 2.46 4.115 2.755 ;
      RECT 4.095 2.482 4.105 2.755 ;
      RECT 4.085 2.507 4.095 2.75 ;
      RECT 4.08 2.545 4.085 2.743 ;
      RECT 4.07 2.655 4.08 2.738 ;
      RECT 5.465 3.576 5.48 3.835 ;
      RECT 5.465 3.591 5.485 3.834 ;
      RECT 5.381 3.591 5.485 3.832 ;
      RECT 5.381 3.605 5.49 3.831 ;
      RECT 5.295 3.647 5.495 3.828 ;
      RECT 5.29 3.59 5.48 3.823 ;
      RECT 5.29 3.661 5.5 3.82 ;
      RECT 5.285 3.692 5.5 3.818 ;
      RECT 5.29 3.689 5.515 3.808 ;
      RECT 5.285 3.735 5.53 3.793 ;
      RECT 5.285 3.763 5.535 3.778 ;
      RECT 5.295 3.565 5.465 3.828 ;
      RECT 5.055 2.575 5.225 2.745 ;
      RECT 5.02 2.575 5.225 2.74 ;
      RECT 5.01 2.575 5.225 2.733 ;
      RECT 5.005 2.56 5.175 2.73 ;
      RECT 3.835 3.097 4.1 3.54 ;
      RECT 3.83 3.068 4.045 3.538 ;
      RECT 3.825 3.222 4.105 3.533 ;
      RECT 3.83 3.117 4.105 3.533 ;
      RECT 3.83 3.128 4.115 3.52 ;
      RECT 3.83 3.075 4.075 3.538 ;
      RECT 3.835 3.062 4.045 3.54 ;
      RECT 3.835 3.06 3.995 3.54 ;
      RECT 3.936 3.052 3.995 3.54 ;
      RECT 3.85 3.053 3.995 3.54 ;
      RECT 3.936 3.051 3.985 3.54 ;
      RECT 3.74 1.866 3.915 2.165 ;
      RECT 3.79 1.828 3.915 2.165 ;
      RECT 3.775 1.83 4.001 2.157 ;
      RECT 3.775 1.833 4.04 2.144 ;
      RECT 3.775 1.834 4.05 2.13 ;
      RECT 3.73 1.885 4.05 2.12 ;
      RECT 3.775 1.835 4.055 2.115 ;
      RECT 3.73 2.045 4.06 2.105 ;
      RECT 3.715 1.905 4.055 2.045 ;
      RECT 3.71 1.921 4.055 1.985 ;
      RECT 3.755 1.845 4.055 2.115 ;
      RECT 3.79 1.826 3.876 2.165 ;
      RECT 1.17 7.855 1.34 8.305 ;
      RECT 1.225 6.075 1.395 8.025 ;
      RECT 1.17 5.015 1.34 6.245 ;
      RECT 0.65 5.015 0.82 8.305 ;
      RECT 0.65 7.315 1.055 7.645 ;
      RECT 0.65 6.475 1.055 6.805 ;
      RECT 78.55 7.8 78.72 8.31 ;
      RECT 77.56 0.57 77.73 1.08 ;
      RECT 77.56 2.39 77.73 3.86 ;
      RECT 77.56 5.02 77.73 6.49 ;
      RECT 77.56 7.8 77.73 8.31 ;
      RECT 76.2 0.575 76.37 3.865 ;
      RECT 76.2 5.015 76.37 8.305 ;
      RECT 75.77 0.575 75.94 1.085 ;
      RECT 75.77 1.655 75.94 3.865 ;
      RECT 75.77 5.015 75.94 7.225 ;
      RECT 75.77 7.795 75.94 8.305 ;
      RECT 70.565 5.015 70.735 8.305 ;
      RECT 70.135 5.015 70.305 7.225 ;
      RECT 70.135 7.795 70.305 8.305 ;
      RECT 63.29 7.8 63.46 8.31 ;
      RECT 62.3 0.57 62.47 1.08 ;
      RECT 62.3 2.39 62.47 3.86 ;
      RECT 62.3 5.02 62.47 6.49 ;
      RECT 62.3 7.8 62.47 8.31 ;
      RECT 60.94 0.575 61.11 3.865 ;
      RECT 60.94 5.015 61.11 8.305 ;
      RECT 60.51 0.575 60.68 1.085 ;
      RECT 60.51 1.655 60.68 3.865 ;
      RECT 60.51 5.015 60.68 7.225 ;
      RECT 60.51 7.795 60.68 8.305 ;
      RECT 55.305 5.015 55.475 8.305 ;
      RECT 54.875 5.015 55.045 7.225 ;
      RECT 54.875 7.795 55.045 8.305 ;
      RECT 48.03 7.8 48.2 8.31 ;
      RECT 47.04 0.57 47.21 1.08 ;
      RECT 47.04 2.39 47.21 3.86 ;
      RECT 47.04 5.02 47.21 6.49 ;
      RECT 47.04 7.8 47.21 8.31 ;
      RECT 45.68 0.575 45.85 3.865 ;
      RECT 45.68 5.015 45.85 8.305 ;
      RECT 45.25 0.575 45.42 1.085 ;
      RECT 45.25 1.655 45.42 3.865 ;
      RECT 45.25 5.015 45.42 7.225 ;
      RECT 45.25 7.795 45.42 8.305 ;
      RECT 40.045 5.015 40.215 8.305 ;
      RECT 39.615 5.015 39.785 7.225 ;
      RECT 39.615 7.795 39.785 8.305 ;
      RECT 32.77 7.8 32.94 8.31 ;
      RECT 31.78 0.57 31.95 1.08 ;
      RECT 31.78 2.39 31.95 3.86 ;
      RECT 31.78 5.02 31.95 6.49 ;
      RECT 31.78 7.8 31.95 8.31 ;
      RECT 30.42 0.575 30.59 3.865 ;
      RECT 30.42 5.015 30.59 8.305 ;
      RECT 29.99 0.575 30.16 1.085 ;
      RECT 29.99 1.655 30.16 3.865 ;
      RECT 29.99 5.015 30.16 7.225 ;
      RECT 29.99 7.795 30.16 8.305 ;
      RECT 24.785 5.015 24.955 8.305 ;
      RECT 24.355 5.015 24.525 7.225 ;
      RECT 24.355 7.795 24.525 8.305 ;
      RECT 17.51 7.8 17.68 8.31 ;
      RECT 16.52 0.57 16.69 1.08 ;
      RECT 16.52 2.39 16.69 3.86 ;
      RECT 16.52 5.02 16.69 6.49 ;
      RECT 16.52 7.8 16.69 8.31 ;
      RECT 15.16 0.575 15.33 3.865 ;
      RECT 15.16 5.015 15.33 8.305 ;
      RECT 14.73 0.575 14.9 1.085 ;
      RECT 14.73 1.655 14.9 3.865 ;
      RECT 14.73 5.015 14.9 7.225 ;
      RECT 14.73 7.795 14.9 8.305 ;
      RECT 9.525 5.015 9.695 8.305 ;
      RECT 9.095 5.015 9.265 7.225 ;
      RECT 9.095 7.795 9.265 8.305 ;
      RECT 1.6 5.015 1.77 7.225 ;
      RECT 1.6 7.795 1.77 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8_b0r2 ;
  SIZE 79.095 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 17.515 0.915 17.685 1.085 ;
        RECT 17.51 0.91 17.68 1.08 ;
        RECT 17.51 2.39 17.68 2.56 ;
      LAYER li1 ;
        RECT 17.515 0.915 17.685 1.085 ;
        RECT 17.51 0.57 17.68 1.08 ;
        RECT 17.51 2.39 17.68 3.86 ;
      LAYER met1 ;
        RECT 17.45 2.36 17.74 2.59 ;
        RECT 17.45 0.88 17.74 1.11 ;
        RECT 17.51 0.88 17.68 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 32.775 0.915 32.945 1.085 ;
        RECT 32.77 0.91 32.94 1.08 ;
        RECT 32.77 2.39 32.94 2.56 ;
      LAYER li1 ;
        RECT 32.775 0.915 32.945 1.085 ;
        RECT 32.77 0.57 32.94 1.08 ;
        RECT 32.77 2.39 32.94 3.86 ;
      LAYER met1 ;
        RECT 32.71 2.36 33 2.59 ;
        RECT 32.71 0.88 33 1.11 ;
        RECT 32.77 0.88 32.94 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 48.035 0.915 48.205 1.085 ;
        RECT 48.03 0.91 48.2 1.08 ;
        RECT 48.03 2.39 48.2 2.56 ;
      LAYER li1 ;
        RECT 48.035 0.915 48.205 1.085 ;
        RECT 48.03 0.57 48.2 1.08 ;
        RECT 48.03 2.39 48.2 3.86 ;
      LAYER met1 ;
        RECT 47.97 2.36 48.26 2.59 ;
        RECT 47.97 0.88 48.26 1.11 ;
        RECT 48.03 0.88 48.2 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 63.295 0.915 63.465 1.085 ;
        RECT 63.29 0.91 63.46 1.08 ;
        RECT 63.29 2.39 63.46 2.56 ;
      LAYER li1 ;
        RECT 63.295 0.915 63.465 1.085 ;
        RECT 63.29 0.57 63.46 1.08 ;
        RECT 63.29 2.39 63.46 3.86 ;
      LAYER met1 ;
        RECT 63.23 2.36 63.52 2.59 ;
        RECT 63.23 0.88 63.52 1.11 ;
        RECT 63.29 0.88 63.46 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 78.555 0.915 78.725 1.085 ;
        RECT 78.55 0.91 78.72 1.08 ;
        RECT 78.55 2.39 78.72 2.56 ;
      LAYER li1 ;
        RECT 78.555 0.915 78.725 1.085 ;
        RECT 78.55 0.57 78.72 1.08 ;
        RECT 78.55 2.39 78.72 3.86 ;
      LAYER met1 ;
        RECT 78.49 2.36 78.78 2.59 ;
        RECT 78.49 0.88 78.78 1.11 ;
        RECT 78.55 0.88 78.72 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 13.28 2.705 13.62 3.055 ;
        RECT 13.275 5.86 13.615 6.21 ;
        RECT 13.355 2.705 13.53 6.21 ;
      LAYER li1 ;
        RECT 13.36 1.66 13.53 2.935 ;
        RECT 13.36 5.945 13.53 7.22 ;
        RECT 7.725 5.945 7.895 7.22 ;
      LAYER met1 ;
        RECT 13.28 2.765 13.76 2.935 ;
        RECT 13.28 2.705 13.62 3.055 ;
        RECT 7.665 5.945 13.76 6.115 ;
        RECT 13.275 5.86 13.615 6.21 ;
        RECT 7.665 5.915 7.955 6.145 ;
      LAYER mcon ;
        RECT 7.725 5.945 7.895 6.115 ;
        RECT 13.36 5.945 13.53 6.115 ;
        RECT 13.36 2.765 13.53 2.935 ;
      LAYER via1 ;
        RECT 13.375 5.96 13.525 6.11 ;
        RECT 13.38 2.805 13.53 2.955 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 28.54 2.705 28.88 3.055 ;
        RECT 28.535 5.86 28.875 6.21 ;
        RECT 28.615 2.705 28.79 6.21 ;
      LAYER li1 ;
        RECT 28.62 1.66 28.79 2.935 ;
        RECT 28.62 5.945 28.79 7.22 ;
        RECT 22.985 5.945 23.155 7.22 ;
      LAYER met1 ;
        RECT 28.54 2.765 29.02 2.935 ;
        RECT 28.54 2.705 28.88 3.055 ;
        RECT 22.925 5.945 29.02 6.115 ;
        RECT 28.535 5.86 28.875 6.21 ;
        RECT 22.925 5.915 23.215 6.145 ;
      LAYER mcon ;
        RECT 22.985 5.945 23.155 6.115 ;
        RECT 28.62 5.945 28.79 6.115 ;
        RECT 28.62 2.765 28.79 2.935 ;
      LAYER via1 ;
        RECT 28.635 5.96 28.785 6.11 ;
        RECT 28.64 2.805 28.79 2.955 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 43.8 2.705 44.14 3.055 ;
        RECT 43.795 5.86 44.135 6.21 ;
        RECT 43.875 2.705 44.05 6.21 ;
      LAYER li1 ;
        RECT 43.88 1.66 44.05 2.935 ;
        RECT 43.88 5.945 44.05 7.22 ;
        RECT 38.245 5.945 38.415 7.22 ;
      LAYER met1 ;
        RECT 43.8 2.765 44.28 2.935 ;
        RECT 43.8 2.705 44.14 3.055 ;
        RECT 38.185 5.945 44.28 6.115 ;
        RECT 43.795 5.86 44.135 6.21 ;
        RECT 38.185 5.915 38.475 6.145 ;
      LAYER mcon ;
        RECT 38.245 5.945 38.415 6.115 ;
        RECT 43.88 5.945 44.05 6.115 ;
        RECT 43.88 2.765 44.05 2.935 ;
      LAYER via1 ;
        RECT 43.895 5.96 44.045 6.11 ;
        RECT 43.9 2.805 44.05 2.955 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 59.06 2.705 59.4 3.055 ;
        RECT 59.055 5.86 59.395 6.21 ;
        RECT 59.135 2.705 59.31 6.21 ;
      LAYER li1 ;
        RECT 59.14 1.66 59.31 2.935 ;
        RECT 59.14 5.945 59.31 7.22 ;
        RECT 53.505 5.945 53.675 7.22 ;
      LAYER met1 ;
        RECT 59.06 2.765 59.54 2.935 ;
        RECT 59.06 2.705 59.4 3.055 ;
        RECT 53.445 5.945 59.54 6.115 ;
        RECT 59.055 5.86 59.395 6.21 ;
        RECT 53.445 5.915 53.735 6.145 ;
      LAYER mcon ;
        RECT 53.505 5.945 53.675 6.115 ;
        RECT 59.14 5.945 59.31 6.115 ;
        RECT 59.14 2.765 59.31 2.935 ;
      LAYER via1 ;
        RECT 59.155 5.96 59.305 6.11 ;
        RECT 59.16 2.805 59.31 2.955 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 74.32 2.705 74.66 3.055 ;
        RECT 74.315 5.86 74.655 6.21 ;
        RECT 74.395 2.705 74.57 6.21 ;
      LAYER li1 ;
        RECT 74.4 1.66 74.57 2.935 ;
        RECT 74.4 5.945 74.57 7.22 ;
        RECT 68.765 5.945 68.935 7.22 ;
      LAYER met1 ;
        RECT 74.32 2.765 74.8 2.935 ;
        RECT 74.32 2.705 74.66 3.055 ;
        RECT 68.705 5.945 74.8 6.115 ;
        RECT 74.315 5.86 74.655 6.21 ;
        RECT 68.705 5.915 68.995 6.145 ;
      LAYER mcon ;
        RECT 68.765 5.945 68.935 6.115 ;
        RECT 74.4 5.945 74.57 6.115 ;
        RECT 74.4 2.765 74.57 2.935 ;
      LAYER via1 ;
        RECT 74.415 5.96 74.565 6.11 ;
        RECT 74.42 2.805 74.57 2.955 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 5.945 0.4 7.22 ;
      LAYER met1 ;
        RECT 0.17 5.945 0.63 6.115 ;
        RECT 0.17 5.915 0.46 6.145 ;
      LAYER mcon ;
        RECT 0.23 5.945 0.4 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 1.61 4.255 2.415 4.635 ;
      LAYER met2 ;
        RECT 1.8 4.255 2.18 4.635 ;
      LAYER li1 ;
        RECT 0 4.44 79.095 4.745 ;
        RECT 64.585 4.135 79.095 4.745 ;
        RECT 76.96 4.13 78.94 4.75 ;
        RECT 78.12 3.4 78.29 5.48 ;
        RECT 77.13 3.4 77.3 5.48 ;
        RECT 74.39 3.405 74.56 5.475 ;
        RECT 71.615 3.635 71.785 4.745 ;
        RECT 69.695 3.635 69.865 4.745 ;
        RECT 68.755 3.635 68.925 5.475 ;
        RECT 67.295 3.635 67.465 4.745 ;
        RECT 65.375 3.635 65.545 4.745 ;
        RECT 2.075 4.14 79.095 4.745 ;
        RECT 49.325 4.135 63.835 4.745 ;
        RECT 61.7 4.13 63.68 4.75 ;
        RECT 62.86 3.4 63.03 5.48 ;
        RECT 61.87 3.4 62.04 5.48 ;
        RECT 59.13 3.405 59.3 5.475 ;
        RECT 56.355 3.635 56.525 4.745 ;
        RECT 54.435 3.635 54.605 4.745 ;
        RECT 53.495 3.635 53.665 5.475 ;
        RECT 52.035 3.635 52.205 4.745 ;
        RECT 50.115 3.635 50.285 4.745 ;
        RECT 34.065 4.135 48.575 4.745 ;
        RECT 46.44 4.13 48.42 4.75 ;
        RECT 47.6 3.4 47.77 5.48 ;
        RECT 46.61 3.4 46.78 5.48 ;
        RECT 43.87 3.405 44.04 5.475 ;
        RECT 41.095 3.635 41.265 4.745 ;
        RECT 39.175 3.635 39.345 4.745 ;
        RECT 38.235 3.635 38.405 5.475 ;
        RECT 36.775 3.635 36.945 4.745 ;
        RECT 34.855 3.635 35.025 4.745 ;
        RECT 18.805 4.135 33.315 4.745 ;
        RECT 31.18 4.13 33.16 4.75 ;
        RECT 32.34 3.4 32.51 5.48 ;
        RECT 31.35 3.4 31.52 5.48 ;
        RECT 28.61 3.405 28.78 5.475 ;
        RECT 25.835 3.635 26.005 4.745 ;
        RECT 23.915 3.635 24.085 4.745 ;
        RECT 22.975 3.635 23.145 5.475 ;
        RECT 21.515 3.635 21.685 4.745 ;
        RECT 19.595 3.635 19.765 4.745 ;
        RECT 3.545 4.135 18.055 4.745 ;
        RECT 15.92 4.13 17.9 4.75 ;
        RECT 17.08 3.4 17.25 5.48 ;
        RECT 16.09 3.4 16.26 5.48 ;
        RECT 13.35 3.405 13.52 5.475 ;
        RECT 10.575 3.635 10.745 4.745 ;
        RECT 8.655 3.635 8.825 4.745 ;
        RECT 7.715 3.635 7.885 5.475 ;
        RECT 6.255 3.635 6.425 4.745 ;
        RECT 4.335 3.635 4.505 4.745 ;
        RECT 2.03 4.44 2.2 8.305 ;
        RECT 0 4.14 79.095 4.39 ;
        RECT 0 4.14 1.905 4.745 ;
        RECT 0.22 4.14 0.39 5.475 ;
      LAYER met1 ;
        RECT 0 4.14 79.095 4.745 ;
        RECT 64.585 4.135 79.095 4.745 ;
        RECT 76.96 4.13 78.94 4.75 ;
        RECT 64.585 3.98 73.325 4.745 ;
        RECT 49.325 4.135 63.835 4.745 ;
        RECT 61.7 4.13 63.68 4.75 ;
        RECT 49.325 3.98 58.065 4.745 ;
        RECT 34.065 4.135 48.575 4.745 ;
        RECT 46.44 4.13 48.42 4.75 ;
        RECT 34.065 3.98 42.805 4.745 ;
        RECT 18.805 4.135 33.315 4.745 ;
        RECT 31.18 4.13 33.16 4.75 ;
        RECT 18.805 3.98 27.545 4.745 ;
        RECT 3.545 4.135 18.055 4.745 ;
        RECT 15.92 4.13 17.9 4.75 ;
        RECT 3.545 3.98 12.285 4.745 ;
        RECT 1.97 6.655 2.26 6.885 ;
        RECT 1.8 6.685 2.26 6.855 ;
      LAYER via2 ;
        RECT 1.89 4.345 2.09 4.545 ;
      LAYER mcon ;
        RECT 2.03 6.685 2.2 6.855 ;
        RECT 2.34 4.545 2.51 4.715 ;
        RECT 3.69 4.135 3.86 4.305 ;
        RECT 4.15 4.135 4.32 4.305 ;
        RECT 4.61 4.135 4.78 4.305 ;
        RECT 5.07 4.135 5.24 4.305 ;
        RECT 5.53 4.135 5.7 4.305 ;
        RECT 5.99 4.135 6.16 4.305 ;
        RECT 6.45 4.135 6.62 4.305 ;
        RECT 6.91 4.135 7.08 4.305 ;
        RECT 7.37 4.135 7.54 4.305 ;
        RECT 7.83 4.135 8 4.305 ;
        RECT 8.29 4.135 8.46 4.305 ;
        RECT 8.75 4.135 8.92 4.305 ;
        RECT 9.21 4.135 9.38 4.305 ;
        RECT 9.67 4.135 9.84 4.305 ;
        RECT 9.835 4.545 10.005 4.715 ;
        RECT 10.13 4.135 10.3 4.305 ;
        RECT 10.59 4.135 10.76 4.305 ;
        RECT 11.05 4.135 11.22 4.305 ;
        RECT 11.51 4.135 11.68 4.305 ;
        RECT 11.97 4.135 12.14 4.305 ;
        RECT 15.47 4.545 15.64 4.715 ;
        RECT 15.47 4.165 15.64 4.335 ;
        RECT 16.17 4.55 16.34 4.72 ;
        RECT 16.17 4.16 16.34 4.33 ;
        RECT 17.16 4.55 17.33 4.72 ;
        RECT 17.16 4.16 17.33 4.33 ;
        RECT 18.95 4.135 19.12 4.305 ;
        RECT 19.41 4.135 19.58 4.305 ;
        RECT 19.87 4.135 20.04 4.305 ;
        RECT 20.33 4.135 20.5 4.305 ;
        RECT 20.79 4.135 20.96 4.305 ;
        RECT 21.25 4.135 21.42 4.305 ;
        RECT 21.71 4.135 21.88 4.305 ;
        RECT 22.17 4.135 22.34 4.305 ;
        RECT 22.63 4.135 22.8 4.305 ;
        RECT 23.09 4.135 23.26 4.305 ;
        RECT 23.55 4.135 23.72 4.305 ;
        RECT 24.01 4.135 24.18 4.305 ;
        RECT 24.47 4.135 24.64 4.305 ;
        RECT 24.93 4.135 25.1 4.305 ;
        RECT 25.095 4.545 25.265 4.715 ;
        RECT 25.39 4.135 25.56 4.305 ;
        RECT 25.85 4.135 26.02 4.305 ;
        RECT 26.31 4.135 26.48 4.305 ;
        RECT 26.77 4.135 26.94 4.305 ;
        RECT 27.23 4.135 27.4 4.305 ;
        RECT 30.73 4.545 30.9 4.715 ;
        RECT 30.73 4.165 30.9 4.335 ;
        RECT 31.43 4.55 31.6 4.72 ;
        RECT 31.43 4.16 31.6 4.33 ;
        RECT 32.42 4.55 32.59 4.72 ;
        RECT 32.42 4.16 32.59 4.33 ;
        RECT 34.21 4.135 34.38 4.305 ;
        RECT 34.67 4.135 34.84 4.305 ;
        RECT 35.13 4.135 35.3 4.305 ;
        RECT 35.59 4.135 35.76 4.305 ;
        RECT 36.05 4.135 36.22 4.305 ;
        RECT 36.51 4.135 36.68 4.305 ;
        RECT 36.97 4.135 37.14 4.305 ;
        RECT 37.43 4.135 37.6 4.305 ;
        RECT 37.89 4.135 38.06 4.305 ;
        RECT 38.35 4.135 38.52 4.305 ;
        RECT 38.81 4.135 38.98 4.305 ;
        RECT 39.27 4.135 39.44 4.305 ;
        RECT 39.73 4.135 39.9 4.305 ;
        RECT 40.19 4.135 40.36 4.305 ;
        RECT 40.355 4.545 40.525 4.715 ;
        RECT 40.65 4.135 40.82 4.305 ;
        RECT 41.11 4.135 41.28 4.305 ;
        RECT 41.57 4.135 41.74 4.305 ;
        RECT 42.03 4.135 42.2 4.305 ;
        RECT 42.49 4.135 42.66 4.305 ;
        RECT 45.99 4.545 46.16 4.715 ;
        RECT 45.99 4.165 46.16 4.335 ;
        RECT 46.69 4.55 46.86 4.72 ;
        RECT 46.69 4.16 46.86 4.33 ;
        RECT 47.68 4.55 47.85 4.72 ;
        RECT 47.68 4.16 47.85 4.33 ;
        RECT 49.47 4.135 49.64 4.305 ;
        RECT 49.93 4.135 50.1 4.305 ;
        RECT 50.39 4.135 50.56 4.305 ;
        RECT 50.85 4.135 51.02 4.305 ;
        RECT 51.31 4.135 51.48 4.305 ;
        RECT 51.77 4.135 51.94 4.305 ;
        RECT 52.23 4.135 52.4 4.305 ;
        RECT 52.69 4.135 52.86 4.305 ;
        RECT 53.15 4.135 53.32 4.305 ;
        RECT 53.61 4.135 53.78 4.305 ;
        RECT 54.07 4.135 54.24 4.305 ;
        RECT 54.53 4.135 54.7 4.305 ;
        RECT 54.99 4.135 55.16 4.305 ;
        RECT 55.45 4.135 55.62 4.305 ;
        RECT 55.615 4.545 55.785 4.715 ;
        RECT 55.91 4.135 56.08 4.305 ;
        RECT 56.37 4.135 56.54 4.305 ;
        RECT 56.83 4.135 57 4.305 ;
        RECT 57.29 4.135 57.46 4.305 ;
        RECT 57.75 4.135 57.92 4.305 ;
        RECT 61.25 4.545 61.42 4.715 ;
        RECT 61.25 4.165 61.42 4.335 ;
        RECT 61.95 4.55 62.12 4.72 ;
        RECT 61.95 4.16 62.12 4.33 ;
        RECT 62.94 4.55 63.11 4.72 ;
        RECT 62.94 4.16 63.11 4.33 ;
        RECT 64.73 4.135 64.9 4.305 ;
        RECT 65.19 4.135 65.36 4.305 ;
        RECT 65.65 4.135 65.82 4.305 ;
        RECT 66.11 4.135 66.28 4.305 ;
        RECT 66.57 4.135 66.74 4.305 ;
        RECT 67.03 4.135 67.2 4.305 ;
        RECT 67.49 4.135 67.66 4.305 ;
        RECT 67.95 4.135 68.12 4.305 ;
        RECT 68.41 4.135 68.58 4.305 ;
        RECT 68.87 4.135 69.04 4.305 ;
        RECT 69.33 4.135 69.5 4.305 ;
        RECT 69.79 4.135 69.96 4.305 ;
        RECT 70.25 4.135 70.42 4.305 ;
        RECT 70.71 4.135 70.88 4.305 ;
        RECT 70.875 4.545 71.045 4.715 ;
        RECT 71.17 4.135 71.34 4.305 ;
        RECT 71.63 4.135 71.8 4.305 ;
        RECT 72.09 4.135 72.26 4.305 ;
        RECT 72.55 4.135 72.72 4.305 ;
        RECT 73.01 4.135 73.18 4.305 ;
        RECT 76.51 4.545 76.68 4.715 ;
        RECT 76.51 4.165 76.68 4.335 ;
        RECT 77.21 4.55 77.38 4.72 ;
        RECT 77.21 4.16 77.38 4.33 ;
        RECT 78.2 4.55 78.37 4.72 ;
        RECT 78.2 4.16 78.37 4.33 ;
      LAYER via1 ;
        RECT 1.915 4.37 2.065 4.52 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 73.705 0.95 74.035 3.055 ;
      RECT 73.705 2.735 74.05 3.025 ;
      RECT 67.695 0.95 68.025 2.585 ;
      RECT 67.695 0.95 74.035 1.28 ;
      RECT 70.035 7.055 70.405 7.425 ;
      RECT 70.07 4.27 70.37 7.425 ;
      RECT 65.88 4.27 70.37 4.57 ;
      RECT 69.06 1.855 69.36 4.57 ;
      RECT 65.88 2.435 66.18 4.57 ;
      RECT 69.015 2.76 69.36 3.49 ;
      RECT 65.775 2.015 66.105 2.745 ;
      RECT 68.655 1.855 69.385 2.185 ;
      RECT 58.445 0.95 58.775 3.055 ;
      RECT 58.445 2.735 58.79 3.025 ;
      RECT 52.435 0.95 52.765 2.585 ;
      RECT 52.435 0.95 58.775 1.28 ;
      RECT 54.775 7.055 55.145 7.425 ;
      RECT 54.81 4.27 55.11 7.425 ;
      RECT 50.62 4.27 55.11 4.57 ;
      RECT 53.8 1.855 54.1 4.57 ;
      RECT 50.62 2.435 50.92 4.57 ;
      RECT 53.755 2.76 54.1 3.49 ;
      RECT 50.515 2.015 50.845 2.745 ;
      RECT 53.395 1.855 54.125 2.185 ;
      RECT 43.185 0.95 43.515 3.055 ;
      RECT 43.185 2.735 43.53 3.025 ;
      RECT 37.175 0.95 37.505 2.585 ;
      RECT 37.175 0.95 43.515 1.28 ;
      RECT 39.515 7.055 39.885 7.425 ;
      RECT 39.55 4.27 39.85 7.425 ;
      RECT 35.36 4.27 39.85 4.57 ;
      RECT 38.54 1.855 38.84 4.57 ;
      RECT 35.36 2.435 35.66 4.57 ;
      RECT 38.495 2.76 38.84 3.49 ;
      RECT 35.255 2.015 35.585 2.745 ;
      RECT 38.135 1.855 38.865 2.185 ;
      RECT 27.925 0.95 28.255 3.055 ;
      RECT 27.925 2.735 28.27 3.025 ;
      RECT 21.915 0.95 22.245 2.585 ;
      RECT 21.915 0.95 28.255 1.28 ;
      RECT 24.255 7.055 24.625 7.425 ;
      RECT 24.29 4.27 24.59 7.425 ;
      RECT 20.1 4.27 24.59 4.57 ;
      RECT 23.28 1.855 23.58 4.57 ;
      RECT 20.1 2.435 20.4 4.57 ;
      RECT 23.235 2.76 23.58 3.49 ;
      RECT 19.995 2.015 20.325 2.745 ;
      RECT 22.875 1.855 23.605 2.185 ;
      RECT 12.665 0.95 12.995 3.055 ;
      RECT 12.665 2.735 13.01 3.025 ;
      RECT 6.655 0.95 6.985 2.585 ;
      RECT 6.655 0.95 12.995 1.28 ;
      RECT 8.995 7.055 9.365 7.425 ;
      RECT 9.03 4.27 9.33 7.425 ;
      RECT 4.84 4.27 9.33 4.57 ;
      RECT 8.02 1.855 8.32 4.57 ;
      RECT 4.84 2.435 5.14 4.57 ;
      RECT 7.975 2.76 8.32 3.49 ;
      RECT 4.735 2.015 5.065 2.745 ;
      RECT 7.615 1.855 8.345 2.185 ;
      RECT 72.135 2.015 72.465 2.745 ;
      RECT 70.935 2.88 71.265 3.61 ;
      RECT 70.095 1.855 70.825 2.185 ;
      RECT 66.495 2.015 66.825 2.745 ;
      RECT 56.875 2.015 57.205 2.745 ;
      RECT 55.675 2.88 56.005 3.61 ;
      RECT 54.835 1.855 55.565 2.185 ;
      RECT 51.235 2.015 51.565 2.745 ;
      RECT 41.615 2.015 41.945 2.745 ;
      RECT 40.415 2.88 40.745 3.61 ;
      RECT 39.575 1.855 40.305 2.185 ;
      RECT 35.975 2.015 36.305 2.745 ;
      RECT 26.355 2.015 26.685 2.745 ;
      RECT 25.155 2.88 25.485 3.61 ;
      RECT 24.315 1.855 25.045 2.185 ;
      RECT 20.715 2.015 21.045 2.745 ;
      RECT 11.095 2.015 11.425 2.745 ;
      RECT 9.895 2.88 10.225 3.61 ;
      RECT 9.055 1.855 9.785 2.185 ;
      RECT 5.455 2.015 5.785 2.745 ;
      RECT 0.005 8.5 0.81 8.88 ;
    LAYER via2 ;
      RECT 73.805 2.78 74.005 2.98 ;
      RECT 72.2 2.48 72.4 2.68 ;
      RECT 71 3.04 71.2 3.24 ;
      RECT 70.16 1.92 70.36 2.12 ;
      RECT 70.12 7.14 70.32 7.34 ;
      RECT 69.08 2.825 69.28 3.025 ;
      RECT 68.72 1.92 68.92 2.12 ;
      RECT 67.76 1.92 67.96 2.12 ;
      RECT 66.56 2.48 66.76 2.68 ;
      RECT 65.84 2.48 66.04 2.68 ;
      RECT 58.545 2.78 58.745 2.98 ;
      RECT 56.94 2.48 57.14 2.68 ;
      RECT 55.74 3.04 55.94 3.24 ;
      RECT 54.9 1.92 55.1 2.12 ;
      RECT 54.86 7.14 55.06 7.34 ;
      RECT 53.82 2.825 54.02 3.025 ;
      RECT 53.46 1.92 53.66 2.12 ;
      RECT 52.5 1.92 52.7 2.12 ;
      RECT 51.3 2.48 51.5 2.68 ;
      RECT 50.58 2.48 50.78 2.68 ;
      RECT 43.285 2.78 43.485 2.98 ;
      RECT 41.68 2.48 41.88 2.68 ;
      RECT 40.48 3.04 40.68 3.24 ;
      RECT 39.64 1.92 39.84 2.12 ;
      RECT 39.6 7.14 39.8 7.34 ;
      RECT 38.56 2.825 38.76 3.025 ;
      RECT 38.2 1.92 38.4 2.12 ;
      RECT 37.24 1.92 37.44 2.12 ;
      RECT 36.04 2.48 36.24 2.68 ;
      RECT 35.32 2.48 35.52 2.68 ;
      RECT 28.025 2.78 28.225 2.98 ;
      RECT 26.42 2.48 26.62 2.68 ;
      RECT 25.22 3.04 25.42 3.24 ;
      RECT 24.38 1.92 24.58 2.12 ;
      RECT 24.34 7.14 24.54 7.34 ;
      RECT 23.3 2.825 23.5 3.025 ;
      RECT 22.94 1.92 23.14 2.12 ;
      RECT 21.98 1.92 22.18 2.12 ;
      RECT 20.78 2.48 20.98 2.68 ;
      RECT 20.06 2.48 20.26 2.68 ;
      RECT 12.765 2.78 12.965 2.98 ;
      RECT 11.16 2.48 11.36 2.68 ;
      RECT 9.96 3.04 10.16 3.24 ;
      RECT 9.12 1.92 9.32 2.12 ;
      RECT 9.08 7.14 9.28 7.34 ;
      RECT 8.04 2.825 8.24 3.025 ;
      RECT 7.68 1.92 7.88 2.12 ;
      RECT 6.72 1.92 6.92 2.12 ;
      RECT 5.52 2.48 5.72 2.68 ;
      RECT 4.8 2.48 5 2.68 ;
      RECT 0.285 8.59 0.485 8.79 ;
    LAYER met2 ;
      RECT 1.225 8.4 78.725 8.57 ;
      RECT 78.555 7.275 78.725 8.57 ;
      RECT 1.225 6.255 1.395 8.57 ;
      RECT 78.525 7.275 78.875 7.625 ;
      RECT 1.165 6.255 1.455 6.605 ;
      RECT 75.365 6.22 75.685 6.545 ;
      RECT 75.395 5.695 75.565 6.545 ;
      RECT 75.395 5.695 75.57 6.045 ;
      RECT 75.395 5.695 76.37 5.87 ;
      RECT 76.195 1.965 76.37 5.87 ;
      RECT 76.14 1.965 76.49 2.315 ;
      RECT 76.165 6.655 76.49 6.98 ;
      RECT 75.05 6.745 76.49 6.915 ;
      RECT 75.05 2.395 75.21 6.915 ;
      RECT 75.365 2.365 75.685 2.685 ;
      RECT 75.05 2.395 75.685 2.565 ;
      RECT 73.715 2.705 74.1 3.055 ;
      RECT 73.705 2.77 74.1 2.97 ;
      RECT 73.85 2.7 74.02 3.055 ;
      RECT 72.16 2.44 72.44 2.72 ;
      RECT 72.155 2.44 72.44 2.673 ;
      RECT 72.135 2.44 72.44 2.65 ;
      RECT 72.125 2.44 72.44 2.63 ;
      RECT 72.115 2.44 72.44 2.615 ;
      RECT 72.09 2.44 72.44 2.588 ;
      RECT 72.08 2.44 72.44 2.563 ;
      RECT 72.035 2.295 72.315 2.555 ;
      RECT 72.035 2.39 72.415 2.555 ;
      RECT 72.035 2.335 72.36 2.555 ;
      RECT 72.035 2.327 72.355 2.555 ;
      RECT 72.035 2.317 72.35 2.555 ;
      RECT 72.035 2.305 72.345 2.555 ;
      RECT 70.96 3 71.24 3.28 ;
      RECT 70.96 3 71.275 3.26 ;
      RECT 63.24 6.655 63.59 7.005 ;
      RECT 70.705 6.61 71.055 6.96 ;
      RECT 63.24 6.685 71.055 6.885 ;
      RECT 70.995 2.42 71.045 2.68 ;
      RECT 70.785 2.42 70.79 2.68 ;
      RECT 69.98 1.975 70.01 2.235 ;
      RECT 69.75 1.975 69.825 2.235 ;
      RECT 70.97 2.37 70.995 2.68 ;
      RECT 70.965 2.327 70.97 2.68 ;
      RECT 70.96 2.31 70.965 2.68 ;
      RECT 70.955 2.297 70.96 2.68 ;
      RECT 70.88 2.18 70.955 2.68 ;
      RECT 70.835 1.997 70.88 2.68 ;
      RECT 70.83 1.925 70.835 2.68 ;
      RECT 70.815 1.9 70.83 2.68 ;
      RECT 70.79 1.862 70.815 2.68 ;
      RECT 70.78 1.842 70.79 2.402 ;
      RECT 70.765 1.834 70.78 2.357 ;
      RECT 70.76 1.826 70.765 2.328 ;
      RECT 70.755 1.823 70.76 2.308 ;
      RECT 70.75 1.82 70.755 2.288 ;
      RECT 70.745 1.817 70.75 2.268 ;
      RECT 70.715 1.806 70.745 2.205 ;
      RECT 70.695 1.791 70.715 2.12 ;
      RECT 70.69 1.783 70.695 2.083 ;
      RECT 70.68 1.777 70.69 2.05 ;
      RECT 70.665 1.769 70.68 2.01 ;
      RECT 70.66 1.762 70.665 1.97 ;
      RECT 70.655 1.759 70.66 1.948 ;
      RECT 70.65 1.756 70.655 1.935 ;
      RECT 70.645 1.755 70.65 1.925 ;
      RECT 70.63 1.749 70.645 1.915 ;
      RECT 70.605 1.736 70.63 1.9 ;
      RECT 70.555 1.711 70.605 1.871 ;
      RECT 70.54 1.69 70.555 1.846 ;
      RECT 70.53 1.683 70.54 1.835 ;
      RECT 70.475 1.664 70.53 1.808 ;
      RECT 70.45 1.642 70.475 1.781 ;
      RECT 70.445 1.635 70.45 1.776 ;
      RECT 70.43 1.635 70.445 1.774 ;
      RECT 70.405 1.627 70.43 1.77 ;
      RECT 70.39 1.625 70.405 1.766 ;
      RECT 70.36 1.625 70.39 1.763 ;
      RECT 70.35 1.625 70.36 1.758 ;
      RECT 70.305 1.625 70.35 1.756 ;
      RECT 70.276 1.625 70.305 1.757 ;
      RECT 70.19 1.625 70.276 1.759 ;
      RECT 70.176 1.626 70.19 1.761 ;
      RECT 70.09 1.627 70.176 1.763 ;
      RECT 70.075 1.628 70.09 1.773 ;
      RECT 70.07 1.629 70.075 1.782 ;
      RECT 70.05 1.632 70.07 1.792 ;
      RECT 70.035 1.64 70.05 1.807 ;
      RECT 70.015 1.658 70.035 1.822 ;
      RECT 70.005 1.67 70.015 1.845 ;
      RECT 69.995 1.679 70.005 1.875 ;
      RECT 69.98 1.691 69.995 1.92 ;
      RECT 69.925 1.724 69.98 2.235 ;
      RECT 69.92 1.752 69.925 2.235 ;
      RECT 69.9 1.767 69.92 2.235 ;
      RECT 69.865 1.827 69.9 2.235 ;
      RECT 69.863 1.877 69.865 2.235 ;
      RECT 69.86 1.885 69.863 2.235 ;
      RECT 69.85 1.9 69.86 2.235 ;
      RECT 69.845 1.912 69.85 2.235 ;
      RECT 69.835 1.937 69.845 2.235 ;
      RECT 69.825 1.965 69.835 2.235 ;
      RECT 67.73 3.47 67.78 3.73 ;
      RECT 70.64 3.02 70.7 3.28 ;
      RECT 70.625 3.02 70.64 3.29 ;
      RECT 70.606 3.02 70.625 3.323 ;
      RECT 70.52 3.02 70.606 3.448 ;
      RECT 70.44 3.02 70.52 3.63 ;
      RECT 70.435 3.257 70.44 3.715 ;
      RECT 70.41 3.327 70.435 3.743 ;
      RECT 70.405 3.397 70.41 3.77 ;
      RECT 70.385 3.469 70.405 3.792 ;
      RECT 70.38 3.536 70.385 3.815 ;
      RECT 70.37 3.565 70.38 3.83 ;
      RECT 70.36 3.587 70.37 3.847 ;
      RECT 70.355 3.597 70.36 3.858 ;
      RECT 70.35 3.605 70.355 3.866 ;
      RECT 70.34 3.613 70.35 3.878 ;
      RECT 70.335 3.625 70.34 3.888 ;
      RECT 70.33 3.633 70.335 3.893 ;
      RECT 70.31 3.651 70.33 3.903 ;
      RECT 70.305 3.668 70.31 3.91 ;
      RECT 70.3 3.676 70.305 3.911 ;
      RECT 70.295 3.687 70.3 3.913 ;
      RECT 70.255 3.725 70.295 3.923 ;
      RECT 70.25 3.76 70.255 3.934 ;
      RECT 70.245 3.765 70.25 3.937 ;
      RECT 70.22 3.775 70.245 3.944 ;
      RECT 70.21 3.789 70.22 3.953 ;
      RECT 70.19 3.801 70.21 3.956 ;
      RECT 70.14 3.82 70.19 3.96 ;
      RECT 70.095 3.835 70.14 3.965 ;
      RECT 70.03 3.838 70.095 3.971 ;
      RECT 70.015 3.836 70.03 3.978 ;
      RECT 69.985 3.835 70.015 3.978 ;
      RECT 69.946 3.834 69.985 3.974 ;
      RECT 69.86 3.831 69.946 3.97 ;
      RECT 69.843 3.829 69.86 3.967 ;
      RECT 69.757 3.827 69.843 3.964 ;
      RECT 69.671 3.824 69.757 3.958 ;
      RECT 69.585 3.82 69.671 3.953 ;
      RECT 69.507 3.817 69.585 3.949 ;
      RECT 69.421 3.814 69.507 3.947 ;
      RECT 69.335 3.811 69.421 3.944 ;
      RECT 69.277 3.809 69.335 3.941 ;
      RECT 69.191 3.806 69.277 3.939 ;
      RECT 69.105 3.802 69.191 3.937 ;
      RECT 69.019 3.799 69.105 3.934 ;
      RECT 68.933 3.795 69.019 3.932 ;
      RECT 68.847 3.791 68.933 3.929 ;
      RECT 68.761 3.788 68.847 3.927 ;
      RECT 68.675 3.784 68.761 3.924 ;
      RECT 68.589 3.781 68.675 3.922 ;
      RECT 68.503 3.777 68.589 3.919 ;
      RECT 68.417 3.774 68.503 3.917 ;
      RECT 68.331 3.77 68.417 3.914 ;
      RECT 68.245 3.767 68.331 3.912 ;
      RECT 68.235 3.765 68.245 3.908 ;
      RECT 68.23 3.765 68.235 3.906 ;
      RECT 68.19 3.76 68.23 3.9 ;
      RECT 68.176 3.751 68.19 3.893 ;
      RECT 68.09 3.721 68.176 3.878 ;
      RECT 68.07 3.687 68.09 3.863 ;
      RECT 68 3.656 68.07 3.85 ;
      RECT 67.995 3.631 68 3.839 ;
      RECT 67.99 3.625 67.995 3.837 ;
      RECT 67.921 3.47 67.99 3.825 ;
      RECT 67.835 3.47 67.921 3.799 ;
      RECT 67.81 3.47 67.835 3.778 ;
      RECT 67.805 3.47 67.81 3.768 ;
      RECT 67.8 3.47 67.805 3.76 ;
      RECT 67.78 3.47 67.8 3.743 ;
      RECT 70.2 2.04 70.46 2.3 ;
      RECT 70.185 2.04 70.46 2.203 ;
      RECT 70.155 2.04 70.46 2.178 ;
      RECT 70.12 1.88 70.4 2.16 ;
      RECT 70.09 3.37 70.15 3.63 ;
      RECT 69.115 2.06 69.17 2.32 ;
      RECT 70.05 3.327 70.09 3.63 ;
      RECT 70.021 3.248 70.05 3.63 ;
      RECT 69.935 3.12 70.021 3.63 ;
      RECT 69.915 3 69.935 3.63 ;
      RECT 69.89 2.951 69.915 3.63 ;
      RECT 69.885 2.916 69.89 3.48 ;
      RECT 69.855 2.876 69.885 3.418 ;
      RECT 69.83 2.813 69.855 3.333 ;
      RECT 69.82 2.775 69.83 3.27 ;
      RECT 69.805 2.75 69.82 3.231 ;
      RECT 69.762 2.708 69.805 3.137 ;
      RECT 69.76 2.681 69.762 3.064 ;
      RECT 69.755 2.676 69.76 3.055 ;
      RECT 69.75 2.669 69.755 3.03 ;
      RECT 69.745 2.663 69.75 3.015 ;
      RECT 69.74 2.657 69.745 3.003 ;
      RECT 69.73 2.648 69.74 2.985 ;
      RECT 69.725 2.639 69.73 2.963 ;
      RECT 69.7 2.62 69.725 2.913 ;
      RECT 69.695 2.601 69.7 2.863 ;
      RECT 69.68 2.587 69.695 2.823 ;
      RECT 69.675 2.573 69.68 2.79 ;
      RECT 69.67 2.566 69.675 2.783 ;
      RECT 69.655 2.553 69.67 2.775 ;
      RECT 69.61 2.515 69.655 2.748 ;
      RECT 69.58 2.468 69.61 2.713 ;
      RECT 69.56 2.437 69.58 2.69 ;
      RECT 69.48 2.37 69.56 2.643 ;
      RECT 69.45 2.3 69.48 2.59 ;
      RECT 69.445 2.277 69.45 2.573 ;
      RECT 69.415 2.255 69.445 2.558 ;
      RECT 69.385 2.214 69.415 2.53 ;
      RECT 69.38 2.189 69.385 2.515 ;
      RECT 69.375 2.183 69.38 2.508 ;
      RECT 69.365 2.06 69.375 2.5 ;
      RECT 69.355 2.06 69.365 2.493 ;
      RECT 69.35 2.06 69.355 2.485 ;
      RECT 69.33 2.06 69.35 2.473 ;
      RECT 69.28 2.06 69.33 2.443 ;
      RECT 69.225 2.06 69.28 2.393 ;
      RECT 69.195 2.06 69.225 2.353 ;
      RECT 69.17 2.06 69.195 2.33 ;
      RECT 69.04 2.785 69.32 3.065 ;
      RECT 69.005 2.7 69.265 2.96 ;
      RECT 69.005 2.782 69.275 2.96 ;
      RECT 67.205 2.155 67.21 2.64 ;
      RECT 67.095 2.34 67.1 2.64 ;
      RECT 67.005 2.38 67.07 2.64 ;
      RECT 68.68 1.88 68.77 2.51 ;
      RECT 68.645 1.93 68.65 2.51 ;
      RECT 68.59 1.955 68.6 2.51 ;
      RECT 68.545 1.955 68.555 2.51 ;
      RECT 68.915 1.88 68.96 2.16 ;
      RECT 67.765 1.61 67.965 1.75 ;
      RECT 68.881 1.88 68.915 2.172 ;
      RECT 68.795 1.88 68.881 2.212 ;
      RECT 68.78 1.88 68.795 2.253 ;
      RECT 68.775 1.88 68.78 2.273 ;
      RECT 68.77 1.88 68.775 2.293 ;
      RECT 68.65 1.922 68.68 2.51 ;
      RECT 68.6 1.942 68.645 2.51 ;
      RECT 68.585 1.957 68.59 2.51 ;
      RECT 68.555 1.957 68.585 2.51 ;
      RECT 68.51 1.942 68.545 2.51 ;
      RECT 68.505 1.93 68.51 2.29 ;
      RECT 68.5 1.927 68.505 2.27 ;
      RECT 68.485 1.917 68.5 2.223 ;
      RECT 68.48 1.91 68.485 2.186 ;
      RECT 68.475 1.907 68.48 2.169 ;
      RECT 68.46 1.897 68.475 2.125 ;
      RECT 68.455 1.888 68.46 2.085 ;
      RECT 68.45 1.884 68.455 2.07 ;
      RECT 68.44 1.878 68.45 2.053 ;
      RECT 68.4 1.859 68.44 2.028 ;
      RECT 68.395 1.841 68.4 2.008 ;
      RECT 68.385 1.835 68.395 2.003 ;
      RECT 68.355 1.819 68.385 1.99 ;
      RECT 68.34 1.801 68.355 1.973 ;
      RECT 68.325 1.789 68.34 1.96 ;
      RECT 68.32 1.781 68.325 1.953 ;
      RECT 68.29 1.767 68.32 1.94 ;
      RECT 68.285 1.752 68.29 1.928 ;
      RECT 68.275 1.746 68.285 1.92 ;
      RECT 68.255 1.734 68.275 1.908 ;
      RECT 68.245 1.722 68.255 1.895 ;
      RECT 68.215 1.706 68.245 1.88 ;
      RECT 68.195 1.686 68.215 1.863 ;
      RECT 68.19 1.676 68.195 1.853 ;
      RECT 68.165 1.664 68.19 1.84 ;
      RECT 68.16 1.652 68.165 1.828 ;
      RECT 68.155 1.647 68.16 1.824 ;
      RECT 68.14 1.64 68.155 1.816 ;
      RECT 68.13 1.627 68.14 1.806 ;
      RECT 68.125 1.625 68.13 1.8 ;
      RECT 68.1 1.618 68.125 1.789 ;
      RECT 68.095 1.611 68.1 1.778 ;
      RECT 68.07 1.61 68.095 1.765 ;
      RECT 68.051 1.61 68.07 1.755 ;
      RECT 67.965 1.61 68.051 1.752 ;
      RECT 67.735 1.61 67.765 1.755 ;
      RECT 67.695 1.617 67.735 1.768 ;
      RECT 67.67 1.627 67.695 1.781 ;
      RECT 67.655 1.636 67.67 1.791 ;
      RECT 67.625 1.641 67.655 1.81 ;
      RECT 67.62 1.647 67.625 1.828 ;
      RECT 67.6 1.657 67.62 1.843 ;
      RECT 67.59 1.67 67.6 1.863 ;
      RECT 67.575 1.682 67.59 1.88 ;
      RECT 67.57 1.692 67.575 1.89 ;
      RECT 67.565 1.697 67.57 1.895 ;
      RECT 67.555 1.705 67.565 1.908 ;
      RECT 67.505 1.737 67.555 1.945 ;
      RECT 67.49 1.772 67.505 1.986 ;
      RECT 67.485 1.782 67.49 2.001 ;
      RECT 67.48 1.787 67.485 2.008 ;
      RECT 67.455 1.803 67.48 2.028 ;
      RECT 67.44 1.824 67.455 2.053 ;
      RECT 67.415 1.845 67.44 2.078 ;
      RECT 67.405 1.864 67.415 2.101 ;
      RECT 67.38 1.882 67.405 2.124 ;
      RECT 67.365 1.902 67.38 2.148 ;
      RECT 67.36 1.912 67.365 2.16 ;
      RECT 67.345 1.924 67.36 2.18 ;
      RECT 67.335 1.939 67.345 2.22 ;
      RECT 67.33 1.947 67.335 2.248 ;
      RECT 67.32 1.957 67.33 2.268 ;
      RECT 67.315 1.97 67.32 2.293 ;
      RECT 67.31 1.983 67.315 2.313 ;
      RECT 67.305 1.989 67.31 2.335 ;
      RECT 67.295 1.998 67.305 2.355 ;
      RECT 67.29 2.018 67.295 2.378 ;
      RECT 67.285 2.024 67.29 2.398 ;
      RECT 67.28 2.031 67.285 2.42 ;
      RECT 67.275 2.042 67.28 2.433 ;
      RECT 67.265 2.052 67.275 2.458 ;
      RECT 67.245 2.077 67.265 2.64 ;
      RECT 67.215 2.117 67.245 2.64 ;
      RECT 67.21 2.147 67.215 2.64 ;
      RECT 67.185 2.175 67.205 2.64 ;
      RECT 67.155 2.22 67.185 2.64 ;
      RECT 67.15 2.247 67.155 2.64 ;
      RECT 67.13 2.265 67.15 2.64 ;
      RECT 67.12 2.29 67.13 2.64 ;
      RECT 67.115 2.302 67.12 2.64 ;
      RECT 67.1 2.325 67.115 2.64 ;
      RECT 67.08 2.352 67.095 2.64 ;
      RECT 67.07 2.375 67.08 2.64 ;
      RECT 68.86 3.26 68.94 3.52 ;
      RECT 68.095 2.48 68.165 2.74 ;
      RECT 68.826 3.227 68.86 3.52 ;
      RECT 68.74 3.13 68.826 3.52 ;
      RECT 68.72 3.042 68.74 3.52 ;
      RECT 68.71 3.012 68.72 3.52 ;
      RECT 68.7 2.992 68.71 3.52 ;
      RECT 68.68 2.979 68.7 3.52 ;
      RECT 68.665 2.969 68.68 3.348 ;
      RECT 68.66 2.962 68.665 3.303 ;
      RECT 68.65 2.956 68.66 3.293 ;
      RECT 68.64 2.948 68.65 3.275 ;
      RECT 68.635 2.942 68.64 3.263 ;
      RECT 68.625 2.937 68.635 3.25 ;
      RECT 68.605 2.927 68.625 3.223 ;
      RECT 68.565 2.906 68.605 3.175 ;
      RECT 68.55 2.887 68.565 3.133 ;
      RECT 68.525 2.873 68.55 3.103 ;
      RECT 68.515 2.861 68.525 3.07 ;
      RECT 68.51 2.856 68.515 3.06 ;
      RECT 68.48 2.842 68.51 3.04 ;
      RECT 68.47 2.826 68.48 3.013 ;
      RECT 68.465 2.821 68.47 3.003 ;
      RECT 68.44 2.812 68.465 2.983 ;
      RECT 68.43 2.8 68.44 2.963 ;
      RECT 68.36 2.768 68.43 2.938 ;
      RECT 68.355 2.737 68.36 2.915 ;
      RECT 68.306 2.48 68.355 2.898 ;
      RECT 68.22 2.48 68.306 2.857 ;
      RECT 68.165 2.48 68.22 2.785 ;
      RECT 68.255 3.265 68.415 3.525 ;
      RECT 67.78 1.88 67.83 2.565 ;
      RECT 67.57 2.305 67.605 2.565 ;
      RECT 67.885 1.88 67.89 2.34 ;
      RECT 67.975 1.88 68 2.16 ;
      RECT 68.25 3.262 68.255 3.525 ;
      RECT 68.215 3.25 68.25 3.525 ;
      RECT 68.155 3.223 68.215 3.525 ;
      RECT 68.15 3.206 68.155 3.379 ;
      RECT 68.145 3.203 68.15 3.366 ;
      RECT 68.125 3.196 68.145 3.353 ;
      RECT 68.09 3.179 68.125 3.335 ;
      RECT 68.05 3.158 68.09 3.315 ;
      RECT 68.045 3.146 68.05 3.303 ;
      RECT 68.005 3.132 68.045 3.289 ;
      RECT 67.985 3.115 68.005 3.271 ;
      RECT 67.975 3.107 67.985 3.263 ;
      RECT 67.96 1.88 67.975 2.178 ;
      RECT 67.945 3.097 67.975 3.25 ;
      RECT 67.93 1.88 67.96 2.223 ;
      RECT 67.935 3.087 67.945 3.237 ;
      RECT 67.905 3.072 67.935 3.224 ;
      RECT 67.89 1.88 67.93 2.29 ;
      RECT 67.89 3.04 67.905 3.21 ;
      RECT 67.885 3.012 67.89 3.204 ;
      RECT 67.88 1.88 67.885 2.345 ;
      RECT 67.87 2.982 67.885 3.198 ;
      RECT 67.875 1.88 67.88 2.358 ;
      RECT 67.865 1.88 67.875 2.378 ;
      RECT 67.83 2.895 67.87 3.183 ;
      RECT 67.83 1.88 67.865 2.418 ;
      RECT 67.825 2.827 67.83 3.171 ;
      RECT 67.81 2.782 67.825 3.166 ;
      RECT 67.805 2.72 67.81 3.161 ;
      RECT 67.78 2.627 67.805 3.154 ;
      RECT 67.775 1.88 67.78 3.146 ;
      RECT 67.76 1.88 67.775 3.133 ;
      RECT 67.74 1.88 67.76 3.09 ;
      RECT 67.73 1.88 67.74 3.04 ;
      RECT 67.725 1.88 67.73 3.013 ;
      RECT 67.72 1.88 67.725 2.991 ;
      RECT 67.715 2.106 67.72 2.974 ;
      RECT 67.71 2.128 67.715 2.952 ;
      RECT 67.705 2.17 67.71 2.935 ;
      RECT 67.675 2.22 67.705 2.879 ;
      RECT 67.67 2.247 67.675 2.821 ;
      RECT 67.655 2.265 67.67 2.785 ;
      RECT 67.65 2.283 67.655 2.749 ;
      RECT 67.644 2.29 67.65 2.73 ;
      RECT 67.64 2.297 67.644 2.713 ;
      RECT 67.635 2.302 67.64 2.682 ;
      RECT 67.625 2.305 67.635 2.657 ;
      RECT 67.615 2.305 67.625 2.623 ;
      RECT 67.61 2.305 67.615 2.6 ;
      RECT 67.605 2.305 67.61 2.58 ;
      RECT 66.52 2.44 66.8 2.72 ;
      RECT 66.52 2.44 66.82 2.615 ;
      RECT 66.61 2.33 66.87 2.59 ;
      RECT 66.575 2.425 66.87 2.59 ;
      RECT 66.7 0.945 66.865 2.59 ;
      RECT 66.6 0.945 66.97 1.315 ;
      RECT 66.225 3.47 66.485 3.73 ;
      RECT 66.245 3.397 66.425 3.73 ;
      RECT 66.245 3.14 66.42 3.73 ;
      RECT 66.245 2.932 66.41 3.73 ;
      RECT 66.25 2.85 66.41 3.73 ;
      RECT 66.25 2.615 66.4 3.73 ;
      RECT 66.25 2.462 66.395 3.73 ;
      RECT 66.255 2.447 66.395 3.73 ;
      RECT 66.305 2.162 66.395 3.73 ;
      RECT 66.26 2.397 66.395 3.73 ;
      RECT 66.29 2.215 66.395 3.73 ;
      RECT 66.275 2.327 66.395 3.73 ;
      RECT 66.28 2.285 66.395 3.73 ;
      RECT 66.275 2.327 66.41 2.39 ;
      RECT 66.31 1.915 66.415 2.335 ;
      RECT 66.31 1.915 66.43 2.318 ;
      RECT 66.31 1.915 66.465 2.28 ;
      RECT 66.305 2.162 66.515 2.213 ;
      RECT 66.31 1.915 66.57 2.175 ;
      RECT 65.57 2.62 65.83 2.88 ;
      RECT 65.57 2.62 65.84 2.838 ;
      RECT 65.57 2.62 65.926 2.809 ;
      RECT 65.57 2.62 65.995 2.761 ;
      RECT 65.57 2.62 66.03 2.73 ;
      RECT 65.8 2.44 66.08 2.72 ;
      RECT 65.635 2.605 66.08 2.72 ;
      RECT 65.725 2.482 65.83 2.88 ;
      RECT 65.655 2.545 66.08 2.72 ;
      RECT 60.105 6.22 60.425 6.545 ;
      RECT 60.135 5.695 60.305 6.545 ;
      RECT 60.135 5.695 60.31 6.045 ;
      RECT 60.135 5.695 61.11 5.87 ;
      RECT 60.935 1.965 61.11 5.87 ;
      RECT 60.88 1.965 61.23 2.315 ;
      RECT 60.905 6.655 61.23 6.98 ;
      RECT 59.79 6.745 61.23 6.915 ;
      RECT 59.79 2.395 59.95 6.915 ;
      RECT 60.105 2.365 60.425 2.685 ;
      RECT 59.79 2.395 60.425 2.565 ;
      RECT 58.455 2.705 58.84 3.055 ;
      RECT 58.445 2.77 58.84 2.97 ;
      RECT 58.59 2.7 58.76 3.055 ;
      RECT 56.9 2.44 57.18 2.72 ;
      RECT 56.895 2.44 57.18 2.673 ;
      RECT 56.875 2.44 57.18 2.65 ;
      RECT 56.865 2.44 57.18 2.63 ;
      RECT 56.855 2.44 57.18 2.615 ;
      RECT 56.83 2.44 57.18 2.588 ;
      RECT 56.82 2.44 57.18 2.563 ;
      RECT 56.775 2.295 57.055 2.555 ;
      RECT 56.775 2.39 57.155 2.555 ;
      RECT 56.775 2.335 57.1 2.555 ;
      RECT 56.775 2.327 57.095 2.555 ;
      RECT 56.775 2.317 57.09 2.555 ;
      RECT 56.775 2.305 57.085 2.555 ;
      RECT 55.7 3 55.98 3.28 ;
      RECT 55.7 3 56.015 3.26 ;
      RECT 47.98 6.655 48.33 7.005 ;
      RECT 55.445 6.61 55.795 6.96 ;
      RECT 47.98 6.685 55.795 6.885 ;
      RECT 55.735 2.42 55.785 2.68 ;
      RECT 55.525 2.42 55.53 2.68 ;
      RECT 54.72 1.975 54.75 2.235 ;
      RECT 54.49 1.975 54.565 2.235 ;
      RECT 55.71 2.37 55.735 2.68 ;
      RECT 55.705 2.327 55.71 2.68 ;
      RECT 55.7 2.31 55.705 2.68 ;
      RECT 55.695 2.297 55.7 2.68 ;
      RECT 55.62 2.18 55.695 2.68 ;
      RECT 55.575 1.997 55.62 2.68 ;
      RECT 55.57 1.925 55.575 2.68 ;
      RECT 55.555 1.9 55.57 2.68 ;
      RECT 55.53 1.862 55.555 2.68 ;
      RECT 55.52 1.842 55.53 2.402 ;
      RECT 55.505 1.834 55.52 2.357 ;
      RECT 55.5 1.826 55.505 2.328 ;
      RECT 55.495 1.823 55.5 2.308 ;
      RECT 55.49 1.82 55.495 2.288 ;
      RECT 55.485 1.817 55.49 2.268 ;
      RECT 55.455 1.806 55.485 2.205 ;
      RECT 55.435 1.791 55.455 2.12 ;
      RECT 55.43 1.783 55.435 2.083 ;
      RECT 55.42 1.777 55.43 2.05 ;
      RECT 55.405 1.769 55.42 2.01 ;
      RECT 55.4 1.762 55.405 1.97 ;
      RECT 55.395 1.759 55.4 1.948 ;
      RECT 55.39 1.756 55.395 1.935 ;
      RECT 55.385 1.755 55.39 1.925 ;
      RECT 55.37 1.749 55.385 1.915 ;
      RECT 55.345 1.736 55.37 1.9 ;
      RECT 55.295 1.711 55.345 1.871 ;
      RECT 55.28 1.69 55.295 1.846 ;
      RECT 55.27 1.683 55.28 1.835 ;
      RECT 55.215 1.664 55.27 1.808 ;
      RECT 55.19 1.642 55.215 1.781 ;
      RECT 55.185 1.635 55.19 1.776 ;
      RECT 55.17 1.635 55.185 1.774 ;
      RECT 55.145 1.627 55.17 1.77 ;
      RECT 55.13 1.625 55.145 1.766 ;
      RECT 55.1 1.625 55.13 1.763 ;
      RECT 55.09 1.625 55.1 1.758 ;
      RECT 55.045 1.625 55.09 1.756 ;
      RECT 55.016 1.625 55.045 1.757 ;
      RECT 54.93 1.625 55.016 1.759 ;
      RECT 54.916 1.626 54.93 1.761 ;
      RECT 54.83 1.627 54.916 1.763 ;
      RECT 54.815 1.628 54.83 1.773 ;
      RECT 54.81 1.629 54.815 1.782 ;
      RECT 54.79 1.632 54.81 1.792 ;
      RECT 54.775 1.64 54.79 1.807 ;
      RECT 54.755 1.658 54.775 1.822 ;
      RECT 54.745 1.67 54.755 1.845 ;
      RECT 54.735 1.679 54.745 1.875 ;
      RECT 54.72 1.691 54.735 1.92 ;
      RECT 54.665 1.724 54.72 2.235 ;
      RECT 54.66 1.752 54.665 2.235 ;
      RECT 54.64 1.767 54.66 2.235 ;
      RECT 54.605 1.827 54.64 2.235 ;
      RECT 54.603 1.877 54.605 2.235 ;
      RECT 54.6 1.885 54.603 2.235 ;
      RECT 54.59 1.9 54.6 2.235 ;
      RECT 54.585 1.912 54.59 2.235 ;
      RECT 54.575 1.937 54.585 2.235 ;
      RECT 54.565 1.965 54.575 2.235 ;
      RECT 52.47 3.47 52.52 3.73 ;
      RECT 55.38 3.02 55.44 3.28 ;
      RECT 55.365 3.02 55.38 3.29 ;
      RECT 55.346 3.02 55.365 3.323 ;
      RECT 55.26 3.02 55.346 3.448 ;
      RECT 55.18 3.02 55.26 3.63 ;
      RECT 55.175 3.257 55.18 3.715 ;
      RECT 55.15 3.327 55.175 3.743 ;
      RECT 55.145 3.397 55.15 3.77 ;
      RECT 55.125 3.469 55.145 3.792 ;
      RECT 55.12 3.536 55.125 3.815 ;
      RECT 55.11 3.565 55.12 3.83 ;
      RECT 55.1 3.587 55.11 3.847 ;
      RECT 55.095 3.597 55.1 3.858 ;
      RECT 55.09 3.605 55.095 3.866 ;
      RECT 55.08 3.613 55.09 3.878 ;
      RECT 55.075 3.625 55.08 3.888 ;
      RECT 55.07 3.633 55.075 3.893 ;
      RECT 55.05 3.651 55.07 3.903 ;
      RECT 55.045 3.668 55.05 3.91 ;
      RECT 55.04 3.676 55.045 3.911 ;
      RECT 55.035 3.687 55.04 3.913 ;
      RECT 54.995 3.725 55.035 3.923 ;
      RECT 54.99 3.76 54.995 3.934 ;
      RECT 54.985 3.765 54.99 3.937 ;
      RECT 54.96 3.775 54.985 3.944 ;
      RECT 54.95 3.789 54.96 3.953 ;
      RECT 54.93 3.801 54.95 3.956 ;
      RECT 54.88 3.82 54.93 3.96 ;
      RECT 54.835 3.835 54.88 3.965 ;
      RECT 54.77 3.838 54.835 3.971 ;
      RECT 54.755 3.836 54.77 3.978 ;
      RECT 54.725 3.835 54.755 3.978 ;
      RECT 54.686 3.834 54.725 3.974 ;
      RECT 54.6 3.831 54.686 3.97 ;
      RECT 54.583 3.829 54.6 3.967 ;
      RECT 54.497 3.827 54.583 3.964 ;
      RECT 54.411 3.824 54.497 3.958 ;
      RECT 54.325 3.82 54.411 3.953 ;
      RECT 54.247 3.817 54.325 3.949 ;
      RECT 54.161 3.814 54.247 3.947 ;
      RECT 54.075 3.811 54.161 3.944 ;
      RECT 54.017 3.809 54.075 3.941 ;
      RECT 53.931 3.806 54.017 3.939 ;
      RECT 53.845 3.802 53.931 3.937 ;
      RECT 53.759 3.799 53.845 3.934 ;
      RECT 53.673 3.795 53.759 3.932 ;
      RECT 53.587 3.791 53.673 3.929 ;
      RECT 53.501 3.788 53.587 3.927 ;
      RECT 53.415 3.784 53.501 3.924 ;
      RECT 53.329 3.781 53.415 3.922 ;
      RECT 53.243 3.777 53.329 3.919 ;
      RECT 53.157 3.774 53.243 3.917 ;
      RECT 53.071 3.77 53.157 3.914 ;
      RECT 52.985 3.767 53.071 3.912 ;
      RECT 52.975 3.765 52.985 3.908 ;
      RECT 52.97 3.765 52.975 3.906 ;
      RECT 52.93 3.76 52.97 3.9 ;
      RECT 52.916 3.751 52.93 3.893 ;
      RECT 52.83 3.721 52.916 3.878 ;
      RECT 52.81 3.687 52.83 3.863 ;
      RECT 52.74 3.656 52.81 3.85 ;
      RECT 52.735 3.631 52.74 3.839 ;
      RECT 52.73 3.625 52.735 3.837 ;
      RECT 52.661 3.47 52.73 3.825 ;
      RECT 52.575 3.47 52.661 3.799 ;
      RECT 52.55 3.47 52.575 3.778 ;
      RECT 52.545 3.47 52.55 3.768 ;
      RECT 52.54 3.47 52.545 3.76 ;
      RECT 52.52 3.47 52.54 3.743 ;
      RECT 54.94 2.04 55.2 2.3 ;
      RECT 54.925 2.04 55.2 2.203 ;
      RECT 54.895 2.04 55.2 2.178 ;
      RECT 54.86 1.88 55.14 2.16 ;
      RECT 54.83 3.37 54.89 3.63 ;
      RECT 53.855 2.06 53.91 2.32 ;
      RECT 54.79 3.327 54.83 3.63 ;
      RECT 54.761 3.248 54.79 3.63 ;
      RECT 54.675 3.12 54.761 3.63 ;
      RECT 54.655 3 54.675 3.63 ;
      RECT 54.63 2.951 54.655 3.63 ;
      RECT 54.625 2.916 54.63 3.48 ;
      RECT 54.595 2.876 54.625 3.418 ;
      RECT 54.57 2.813 54.595 3.333 ;
      RECT 54.56 2.775 54.57 3.27 ;
      RECT 54.545 2.75 54.56 3.231 ;
      RECT 54.502 2.708 54.545 3.137 ;
      RECT 54.5 2.681 54.502 3.064 ;
      RECT 54.495 2.676 54.5 3.055 ;
      RECT 54.49 2.669 54.495 3.03 ;
      RECT 54.485 2.663 54.49 3.015 ;
      RECT 54.48 2.657 54.485 3.003 ;
      RECT 54.47 2.648 54.48 2.985 ;
      RECT 54.465 2.639 54.47 2.963 ;
      RECT 54.44 2.62 54.465 2.913 ;
      RECT 54.435 2.601 54.44 2.863 ;
      RECT 54.42 2.587 54.435 2.823 ;
      RECT 54.415 2.573 54.42 2.79 ;
      RECT 54.41 2.566 54.415 2.783 ;
      RECT 54.395 2.553 54.41 2.775 ;
      RECT 54.35 2.515 54.395 2.748 ;
      RECT 54.32 2.468 54.35 2.713 ;
      RECT 54.3 2.437 54.32 2.69 ;
      RECT 54.22 2.37 54.3 2.643 ;
      RECT 54.19 2.3 54.22 2.59 ;
      RECT 54.185 2.277 54.19 2.573 ;
      RECT 54.155 2.255 54.185 2.558 ;
      RECT 54.125 2.214 54.155 2.53 ;
      RECT 54.12 2.189 54.125 2.515 ;
      RECT 54.115 2.183 54.12 2.508 ;
      RECT 54.105 2.06 54.115 2.5 ;
      RECT 54.095 2.06 54.105 2.493 ;
      RECT 54.09 2.06 54.095 2.485 ;
      RECT 54.07 2.06 54.09 2.473 ;
      RECT 54.02 2.06 54.07 2.443 ;
      RECT 53.965 2.06 54.02 2.393 ;
      RECT 53.935 2.06 53.965 2.353 ;
      RECT 53.91 2.06 53.935 2.33 ;
      RECT 53.78 2.785 54.06 3.065 ;
      RECT 53.745 2.7 54.005 2.96 ;
      RECT 53.745 2.782 54.015 2.96 ;
      RECT 51.945 2.155 51.95 2.64 ;
      RECT 51.835 2.34 51.84 2.64 ;
      RECT 51.745 2.38 51.81 2.64 ;
      RECT 53.42 1.88 53.51 2.51 ;
      RECT 53.385 1.93 53.39 2.51 ;
      RECT 53.33 1.955 53.34 2.51 ;
      RECT 53.285 1.955 53.295 2.51 ;
      RECT 53.655 1.88 53.7 2.16 ;
      RECT 52.505 1.61 52.705 1.75 ;
      RECT 53.621 1.88 53.655 2.172 ;
      RECT 53.535 1.88 53.621 2.212 ;
      RECT 53.52 1.88 53.535 2.253 ;
      RECT 53.515 1.88 53.52 2.273 ;
      RECT 53.51 1.88 53.515 2.293 ;
      RECT 53.39 1.922 53.42 2.51 ;
      RECT 53.34 1.942 53.385 2.51 ;
      RECT 53.325 1.957 53.33 2.51 ;
      RECT 53.295 1.957 53.325 2.51 ;
      RECT 53.25 1.942 53.285 2.51 ;
      RECT 53.245 1.93 53.25 2.29 ;
      RECT 53.24 1.927 53.245 2.27 ;
      RECT 53.225 1.917 53.24 2.223 ;
      RECT 53.22 1.91 53.225 2.186 ;
      RECT 53.215 1.907 53.22 2.169 ;
      RECT 53.2 1.897 53.215 2.125 ;
      RECT 53.195 1.888 53.2 2.085 ;
      RECT 53.19 1.884 53.195 2.07 ;
      RECT 53.18 1.878 53.19 2.053 ;
      RECT 53.14 1.859 53.18 2.028 ;
      RECT 53.135 1.841 53.14 2.008 ;
      RECT 53.125 1.835 53.135 2.003 ;
      RECT 53.095 1.819 53.125 1.99 ;
      RECT 53.08 1.801 53.095 1.973 ;
      RECT 53.065 1.789 53.08 1.96 ;
      RECT 53.06 1.781 53.065 1.953 ;
      RECT 53.03 1.767 53.06 1.94 ;
      RECT 53.025 1.752 53.03 1.928 ;
      RECT 53.015 1.746 53.025 1.92 ;
      RECT 52.995 1.734 53.015 1.908 ;
      RECT 52.985 1.722 52.995 1.895 ;
      RECT 52.955 1.706 52.985 1.88 ;
      RECT 52.935 1.686 52.955 1.863 ;
      RECT 52.93 1.676 52.935 1.853 ;
      RECT 52.905 1.664 52.93 1.84 ;
      RECT 52.9 1.652 52.905 1.828 ;
      RECT 52.895 1.647 52.9 1.824 ;
      RECT 52.88 1.64 52.895 1.816 ;
      RECT 52.87 1.627 52.88 1.806 ;
      RECT 52.865 1.625 52.87 1.8 ;
      RECT 52.84 1.618 52.865 1.789 ;
      RECT 52.835 1.611 52.84 1.778 ;
      RECT 52.81 1.61 52.835 1.765 ;
      RECT 52.791 1.61 52.81 1.755 ;
      RECT 52.705 1.61 52.791 1.752 ;
      RECT 52.475 1.61 52.505 1.755 ;
      RECT 52.435 1.617 52.475 1.768 ;
      RECT 52.41 1.627 52.435 1.781 ;
      RECT 52.395 1.636 52.41 1.791 ;
      RECT 52.365 1.641 52.395 1.81 ;
      RECT 52.36 1.647 52.365 1.828 ;
      RECT 52.34 1.657 52.36 1.843 ;
      RECT 52.33 1.67 52.34 1.863 ;
      RECT 52.315 1.682 52.33 1.88 ;
      RECT 52.31 1.692 52.315 1.89 ;
      RECT 52.305 1.697 52.31 1.895 ;
      RECT 52.295 1.705 52.305 1.908 ;
      RECT 52.245 1.737 52.295 1.945 ;
      RECT 52.23 1.772 52.245 1.986 ;
      RECT 52.225 1.782 52.23 2.001 ;
      RECT 52.22 1.787 52.225 2.008 ;
      RECT 52.195 1.803 52.22 2.028 ;
      RECT 52.18 1.824 52.195 2.053 ;
      RECT 52.155 1.845 52.18 2.078 ;
      RECT 52.145 1.864 52.155 2.101 ;
      RECT 52.12 1.882 52.145 2.124 ;
      RECT 52.105 1.902 52.12 2.148 ;
      RECT 52.1 1.912 52.105 2.16 ;
      RECT 52.085 1.924 52.1 2.18 ;
      RECT 52.075 1.939 52.085 2.22 ;
      RECT 52.07 1.947 52.075 2.248 ;
      RECT 52.06 1.957 52.07 2.268 ;
      RECT 52.055 1.97 52.06 2.293 ;
      RECT 52.05 1.983 52.055 2.313 ;
      RECT 52.045 1.989 52.05 2.335 ;
      RECT 52.035 1.998 52.045 2.355 ;
      RECT 52.03 2.018 52.035 2.378 ;
      RECT 52.025 2.024 52.03 2.398 ;
      RECT 52.02 2.031 52.025 2.42 ;
      RECT 52.015 2.042 52.02 2.433 ;
      RECT 52.005 2.052 52.015 2.458 ;
      RECT 51.985 2.077 52.005 2.64 ;
      RECT 51.955 2.117 51.985 2.64 ;
      RECT 51.95 2.147 51.955 2.64 ;
      RECT 51.925 2.175 51.945 2.64 ;
      RECT 51.895 2.22 51.925 2.64 ;
      RECT 51.89 2.247 51.895 2.64 ;
      RECT 51.87 2.265 51.89 2.64 ;
      RECT 51.86 2.29 51.87 2.64 ;
      RECT 51.855 2.302 51.86 2.64 ;
      RECT 51.84 2.325 51.855 2.64 ;
      RECT 51.82 2.352 51.835 2.64 ;
      RECT 51.81 2.375 51.82 2.64 ;
      RECT 53.6 3.26 53.68 3.52 ;
      RECT 52.835 2.48 52.905 2.74 ;
      RECT 53.566 3.227 53.6 3.52 ;
      RECT 53.48 3.13 53.566 3.52 ;
      RECT 53.46 3.042 53.48 3.52 ;
      RECT 53.45 3.012 53.46 3.52 ;
      RECT 53.44 2.992 53.45 3.52 ;
      RECT 53.42 2.979 53.44 3.52 ;
      RECT 53.405 2.969 53.42 3.348 ;
      RECT 53.4 2.962 53.405 3.303 ;
      RECT 53.39 2.956 53.4 3.293 ;
      RECT 53.38 2.948 53.39 3.275 ;
      RECT 53.375 2.942 53.38 3.263 ;
      RECT 53.365 2.937 53.375 3.25 ;
      RECT 53.345 2.927 53.365 3.223 ;
      RECT 53.305 2.906 53.345 3.175 ;
      RECT 53.29 2.887 53.305 3.133 ;
      RECT 53.265 2.873 53.29 3.103 ;
      RECT 53.255 2.861 53.265 3.07 ;
      RECT 53.25 2.856 53.255 3.06 ;
      RECT 53.22 2.842 53.25 3.04 ;
      RECT 53.21 2.826 53.22 3.013 ;
      RECT 53.205 2.821 53.21 3.003 ;
      RECT 53.18 2.812 53.205 2.983 ;
      RECT 53.17 2.8 53.18 2.963 ;
      RECT 53.1 2.768 53.17 2.938 ;
      RECT 53.095 2.737 53.1 2.915 ;
      RECT 53.046 2.48 53.095 2.898 ;
      RECT 52.96 2.48 53.046 2.857 ;
      RECT 52.905 2.48 52.96 2.785 ;
      RECT 52.995 3.265 53.155 3.525 ;
      RECT 52.52 1.88 52.57 2.565 ;
      RECT 52.31 2.305 52.345 2.565 ;
      RECT 52.625 1.88 52.63 2.34 ;
      RECT 52.715 1.88 52.74 2.16 ;
      RECT 52.99 3.262 52.995 3.525 ;
      RECT 52.955 3.25 52.99 3.525 ;
      RECT 52.895 3.223 52.955 3.525 ;
      RECT 52.89 3.206 52.895 3.379 ;
      RECT 52.885 3.203 52.89 3.366 ;
      RECT 52.865 3.196 52.885 3.353 ;
      RECT 52.83 3.179 52.865 3.335 ;
      RECT 52.79 3.158 52.83 3.315 ;
      RECT 52.785 3.146 52.79 3.303 ;
      RECT 52.745 3.132 52.785 3.289 ;
      RECT 52.725 3.115 52.745 3.271 ;
      RECT 52.715 3.107 52.725 3.263 ;
      RECT 52.7 1.88 52.715 2.178 ;
      RECT 52.685 3.097 52.715 3.25 ;
      RECT 52.67 1.88 52.7 2.223 ;
      RECT 52.675 3.087 52.685 3.237 ;
      RECT 52.645 3.072 52.675 3.224 ;
      RECT 52.63 1.88 52.67 2.29 ;
      RECT 52.63 3.04 52.645 3.21 ;
      RECT 52.625 3.012 52.63 3.204 ;
      RECT 52.62 1.88 52.625 2.345 ;
      RECT 52.61 2.982 52.625 3.198 ;
      RECT 52.615 1.88 52.62 2.358 ;
      RECT 52.605 1.88 52.615 2.378 ;
      RECT 52.57 2.895 52.61 3.183 ;
      RECT 52.57 1.88 52.605 2.418 ;
      RECT 52.565 2.827 52.57 3.171 ;
      RECT 52.55 2.782 52.565 3.166 ;
      RECT 52.545 2.72 52.55 3.161 ;
      RECT 52.52 2.627 52.545 3.154 ;
      RECT 52.515 1.88 52.52 3.146 ;
      RECT 52.5 1.88 52.515 3.133 ;
      RECT 52.48 1.88 52.5 3.09 ;
      RECT 52.47 1.88 52.48 3.04 ;
      RECT 52.465 1.88 52.47 3.013 ;
      RECT 52.46 1.88 52.465 2.991 ;
      RECT 52.455 2.106 52.46 2.974 ;
      RECT 52.45 2.128 52.455 2.952 ;
      RECT 52.445 2.17 52.45 2.935 ;
      RECT 52.415 2.22 52.445 2.879 ;
      RECT 52.41 2.247 52.415 2.821 ;
      RECT 52.395 2.265 52.41 2.785 ;
      RECT 52.39 2.283 52.395 2.749 ;
      RECT 52.384 2.29 52.39 2.73 ;
      RECT 52.38 2.297 52.384 2.713 ;
      RECT 52.375 2.302 52.38 2.682 ;
      RECT 52.365 2.305 52.375 2.657 ;
      RECT 52.355 2.305 52.365 2.623 ;
      RECT 52.35 2.305 52.355 2.6 ;
      RECT 52.345 2.305 52.35 2.58 ;
      RECT 51.26 2.44 51.54 2.72 ;
      RECT 51.26 2.44 51.56 2.615 ;
      RECT 51.35 2.33 51.61 2.59 ;
      RECT 51.315 2.425 51.61 2.59 ;
      RECT 51.44 0.945 51.605 2.59 ;
      RECT 51.34 0.945 51.71 1.315 ;
      RECT 50.965 3.47 51.225 3.73 ;
      RECT 50.985 3.397 51.165 3.73 ;
      RECT 50.985 3.14 51.16 3.73 ;
      RECT 50.985 2.932 51.15 3.73 ;
      RECT 50.99 2.85 51.15 3.73 ;
      RECT 50.99 2.615 51.14 3.73 ;
      RECT 50.99 2.462 51.135 3.73 ;
      RECT 50.995 2.447 51.135 3.73 ;
      RECT 51.045 2.162 51.135 3.73 ;
      RECT 51 2.397 51.135 3.73 ;
      RECT 51.03 2.215 51.135 3.73 ;
      RECT 51.015 2.327 51.135 3.73 ;
      RECT 51.02 2.285 51.135 3.73 ;
      RECT 51.015 2.327 51.15 2.39 ;
      RECT 51.05 1.915 51.155 2.335 ;
      RECT 51.05 1.915 51.17 2.318 ;
      RECT 51.05 1.915 51.205 2.28 ;
      RECT 51.045 2.162 51.255 2.213 ;
      RECT 51.05 1.915 51.31 2.175 ;
      RECT 50.31 2.62 50.57 2.88 ;
      RECT 50.31 2.62 50.58 2.838 ;
      RECT 50.31 2.62 50.666 2.809 ;
      RECT 50.31 2.62 50.735 2.761 ;
      RECT 50.31 2.62 50.77 2.73 ;
      RECT 50.54 2.44 50.82 2.72 ;
      RECT 50.375 2.605 50.82 2.72 ;
      RECT 50.465 2.482 50.57 2.88 ;
      RECT 50.395 2.545 50.82 2.72 ;
      RECT 44.845 6.22 45.165 6.545 ;
      RECT 44.875 5.695 45.045 6.545 ;
      RECT 44.875 5.695 45.05 6.045 ;
      RECT 44.875 5.695 45.85 5.87 ;
      RECT 45.675 1.965 45.85 5.87 ;
      RECT 45.62 1.965 45.97 2.315 ;
      RECT 45.645 6.655 45.97 6.98 ;
      RECT 44.53 6.745 45.97 6.915 ;
      RECT 44.53 2.395 44.69 6.915 ;
      RECT 44.845 2.365 45.165 2.685 ;
      RECT 44.53 2.395 45.165 2.565 ;
      RECT 43.195 2.705 43.58 3.055 ;
      RECT 43.185 2.77 43.58 2.97 ;
      RECT 43.33 2.7 43.5 3.055 ;
      RECT 41.64 2.44 41.92 2.72 ;
      RECT 41.635 2.44 41.92 2.673 ;
      RECT 41.615 2.44 41.92 2.65 ;
      RECT 41.605 2.44 41.92 2.63 ;
      RECT 41.595 2.44 41.92 2.615 ;
      RECT 41.57 2.44 41.92 2.588 ;
      RECT 41.56 2.44 41.92 2.563 ;
      RECT 41.515 2.295 41.795 2.555 ;
      RECT 41.515 2.39 41.895 2.555 ;
      RECT 41.515 2.335 41.84 2.555 ;
      RECT 41.515 2.327 41.835 2.555 ;
      RECT 41.515 2.317 41.83 2.555 ;
      RECT 41.515 2.305 41.825 2.555 ;
      RECT 40.44 3 40.72 3.28 ;
      RECT 40.44 3 40.755 3.26 ;
      RECT 32.765 6.66 33.115 7.01 ;
      RECT 40.185 6.615 40.535 6.965 ;
      RECT 32.765 6.69 40.535 6.89 ;
      RECT 40.475 2.42 40.525 2.68 ;
      RECT 40.265 2.42 40.27 2.68 ;
      RECT 39.46 1.975 39.49 2.235 ;
      RECT 39.23 1.975 39.305 2.235 ;
      RECT 40.45 2.37 40.475 2.68 ;
      RECT 40.445 2.327 40.45 2.68 ;
      RECT 40.44 2.31 40.445 2.68 ;
      RECT 40.435 2.297 40.44 2.68 ;
      RECT 40.36 2.18 40.435 2.68 ;
      RECT 40.315 1.997 40.36 2.68 ;
      RECT 40.31 1.925 40.315 2.68 ;
      RECT 40.295 1.9 40.31 2.68 ;
      RECT 40.27 1.862 40.295 2.68 ;
      RECT 40.26 1.842 40.27 2.402 ;
      RECT 40.245 1.834 40.26 2.357 ;
      RECT 40.24 1.826 40.245 2.328 ;
      RECT 40.235 1.823 40.24 2.308 ;
      RECT 40.23 1.82 40.235 2.288 ;
      RECT 40.225 1.817 40.23 2.268 ;
      RECT 40.195 1.806 40.225 2.205 ;
      RECT 40.175 1.791 40.195 2.12 ;
      RECT 40.17 1.783 40.175 2.083 ;
      RECT 40.16 1.777 40.17 2.05 ;
      RECT 40.145 1.769 40.16 2.01 ;
      RECT 40.14 1.762 40.145 1.97 ;
      RECT 40.135 1.759 40.14 1.948 ;
      RECT 40.13 1.756 40.135 1.935 ;
      RECT 40.125 1.755 40.13 1.925 ;
      RECT 40.11 1.749 40.125 1.915 ;
      RECT 40.085 1.736 40.11 1.9 ;
      RECT 40.035 1.711 40.085 1.871 ;
      RECT 40.02 1.69 40.035 1.846 ;
      RECT 40.01 1.683 40.02 1.835 ;
      RECT 39.955 1.664 40.01 1.808 ;
      RECT 39.93 1.642 39.955 1.781 ;
      RECT 39.925 1.635 39.93 1.776 ;
      RECT 39.91 1.635 39.925 1.774 ;
      RECT 39.885 1.627 39.91 1.77 ;
      RECT 39.87 1.625 39.885 1.766 ;
      RECT 39.84 1.625 39.87 1.763 ;
      RECT 39.83 1.625 39.84 1.758 ;
      RECT 39.785 1.625 39.83 1.756 ;
      RECT 39.756 1.625 39.785 1.757 ;
      RECT 39.67 1.625 39.756 1.759 ;
      RECT 39.656 1.626 39.67 1.761 ;
      RECT 39.57 1.627 39.656 1.763 ;
      RECT 39.555 1.628 39.57 1.773 ;
      RECT 39.55 1.629 39.555 1.782 ;
      RECT 39.53 1.632 39.55 1.792 ;
      RECT 39.515 1.64 39.53 1.807 ;
      RECT 39.495 1.658 39.515 1.822 ;
      RECT 39.485 1.67 39.495 1.845 ;
      RECT 39.475 1.679 39.485 1.875 ;
      RECT 39.46 1.691 39.475 1.92 ;
      RECT 39.405 1.724 39.46 2.235 ;
      RECT 39.4 1.752 39.405 2.235 ;
      RECT 39.38 1.767 39.4 2.235 ;
      RECT 39.345 1.827 39.38 2.235 ;
      RECT 39.343 1.877 39.345 2.235 ;
      RECT 39.34 1.885 39.343 2.235 ;
      RECT 39.33 1.9 39.34 2.235 ;
      RECT 39.325 1.912 39.33 2.235 ;
      RECT 39.315 1.937 39.325 2.235 ;
      RECT 39.305 1.965 39.315 2.235 ;
      RECT 37.21 3.47 37.26 3.73 ;
      RECT 40.12 3.02 40.18 3.28 ;
      RECT 40.105 3.02 40.12 3.29 ;
      RECT 40.086 3.02 40.105 3.323 ;
      RECT 40 3.02 40.086 3.448 ;
      RECT 39.92 3.02 40 3.63 ;
      RECT 39.915 3.257 39.92 3.715 ;
      RECT 39.89 3.327 39.915 3.743 ;
      RECT 39.885 3.397 39.89 3.77 ;
      RECT 39.865 3.469 39.885 3.792 ;
      RECT 39.86 3.536 39.865 3.815 ;
      RECT 39.85 3.565 39.86 3.83 ;
      RECT 39.84 3.587 39.85 3.847 ;
      RECT 39.835 3.597 39.84 3.858 ;
      RECT 39.83 3.605 39.835 3.866 ;
      RECT 39.82 3.613 39.83 3.878 ;
      RECT 39.815 3.625 39.82 3.888 ;
      RECT 39.81 3.633 39.815 3.893 ;
      RECT 39.79 3.651 39.81 3.903 ;
      RECT 39.785 3.668 39.79 3.91 ;
      RECT 39.78 3.676 39.785 3.911 ;
      RECT 39.775 3.687 39.78 3.913 ;
      RECT 39.735 3.725 39.775 3.923 ;
      RECT 39.73 3.76 39.735 3.934 ;
      RECT 39.725 3.765 39.73 3.937 ;
      RECT 39.7 3.775 39.725 3.944 ;
      RECT 39.69 3.789 39.7 3.953 ;
      RECT 39.67 3.801 39.69 3.956 ;
      RECT 39.62 3.82 39.67 3.96 ;
      RECT 39.575 3.835 39.62 3.965 ;
      RECT 39.51 3.838 39.575 3.971 ;
      RECT 39.495 3.836 39.51 3.978 ;
      RECT 39.465 3.835 39.495 3.978 ;
      RECT 39.426 3.834 39.465 3.974 ;
      RECT 39.34 3.831 39.426 3.97 ;
      RECT 39.323 3.829 39.34 3.967 ;
      RECT 39.237 3.827 39.323 3.964 ;
      RECT 39.151 3.824 39.237 3.958 ;
      RECT 39.065 3.82 39.151 3.953 ;
      RECT 38.987 3.817 39.065 3.949 ;
      RECT 38.901 3.814 38.987 3.947 ;
      RECT 38.815 3.811 38.901 3.944 ;
      RECT 38.757 3.809 38.815 3.941 ;
      RECT 38.671 3.806 38.757 3.939 ;
      RECT 38.585 3.802 38.671 3.937 ;
      RECT 38.499 3.799 38.585 3.934 ;
      RECT 38.413 3.795 38.499 3.932 ;
      RECT 38.327 3.791 38.413 3.929 ;
      RECT 38.241 3.788 38.327 3.927 ;
      RECT 38.155 3.784 38.241 3.924 ;
      RECT 38.069 3.781 38.155 3.922 ;
      RECT 37.983 3.777 38.069 3.919 ;
      RECT 37.897 3.774 37.983 3.917 ;
      RECT 37.811 3.77 37.897 3.914 ;
      RECT 37.725 3.767 37.811 3.912 ;
      RECT 37.715 3.765 37.725 3.908 ;
      RECT 37.71 3.765 37.715 3.906 ;
      RECT 37.67 3.76 37.71 3.9 ;
      RECT 37.656 3.751 37.67 3.893 ;
      RECT 37.57 3.721 37.656 3.878 ;
      RECT 37.55 3.687 37.57 3.863 ;
      RECT 37.48 3.656 37.55 3.85 ;
      RECT 37.475 3.631 37.48 3.839 ;
      RECT 37.47 3.625 37.475 3.837 ;
      RECT 37.401 3.47 37.47 3.825 ;
      RECT 37.315 3.47 37.401 3.799 ;
      RECT 37.29 3.47 37.315 3.778 ;
      RECT 37.285 3.47 37.29 3.768 ;
      RECT 37.28 3.47 37.285 3.76 ;
      RECT 37.26 3.47 37.28 3.743 ;
      RECT 39.68 2.04 39.94 2.3 ;
      RECT 39.665 2.04 39.94 2.203 ;
      RECT 39.635 2.04 39.94 2.178 ;
      RECT 39.6 1.88 39.88 2.16 ;
      RECT 39.57 3.37 39.63 3.63 ;
      RECT 38.595 2.06 38.65 2.32 ;
      RECT 39.53 3.327 39.57 3.63 ;
      RECT 39.501 3.248 39.53 3.63 ;
      RECT 39.415 3.12 39.501 3.63 ;
      RECT 39.395 3 39.415 3.63 ;
      RECT 39.37 2.951 39.395 3.63 ;
      RECT 39.365 2.916 39.37 3.48 ;
      RECT 39.335 2.876 39.365 3.418 ;
      RECT 39.31 2.813 39.335 3.333 ;
      RECT 39.3 2.775 39.31 3.27 ;
      RECT 39.285 2.75 39.3 3.231 ;
      RECT 39.242 2.708 39.285 3.137 ;
      RECT 39.24 2.681 39.242 3.064 ;
      RECT 39.235 2.676 39.24 3.055 ;
      RECT 39.23 2.669 39.235 3.03 ;
      RECT 39.225 2.663 39.23 3.015 ;
      RECT 39.22 2.657 39.225 3.003 ;
      RECT 39.21 2.648 39.22 2.985 ;
      RECT 39.205 2.639 39.21 2.963 ;
      RECT 39.18 2.62 39.205 2.913 ;
      RECT 39.175 2.601 39.18 2.863 ;
      RECT 39.16 2.587 39.175 2.823 ;
      RECT 39.155 2.573 39.16 2.79 ;
      RECT 39.15 2.566 39.155 2.783 ;
      RECT 39.135 2.553 39.15 2.775 ;
      RECT 39.09 2.515 39.135 2.748 ;
      RECT 39.06 2.468 39.09 2.713 ;
      RECT 39.04 2.437 39.06 2.69 ;
      RECT 38.96 2.37 39.04 2.643 ;
      RECT 38.93 2.3 38.96 2.59 ;
      RECT 38.925 2.277 38.93 2.573 ;
      RECT 38.895 2.255 38.925 2.558 ;
      RECT 38.865 2.214 38.895 2.53 ;
      RECT 38.86 2.189 38.865 2.515 ;
      RECT 38.855 2.183 38.86 2.508 ;
      RECT 38.845 2.06 38.855 2.5 ;
      RECT 38.835 2.06 38.845 2.493 ;
      RECT 38.83 2.06 38.835 2.485 ;
      RECT 38.81 2.06 38.83 2.473 ;
      RECT 38.76 2.06 38.81 2.443 ;
      RECT 38.705 2.06 38.76 2.393 ;
      RECT 38.675 2.06 38.705 2.353 ;
      RECT 38.65 2.06 38.675 2.33 ;
      RECT 38.52 2.785 38.8 3.065 ;
      RECT 38.485 2.7 38.745 2.96 ;
      RECT 38.485 2.782 38.755 2.96 ;
      RECT 36.685 2.155 36.69 2.64 ;
      RECT 36.575 2.34 36.58 2.64 ;
      RECT 36.485 2.38 36.55 2.64 ;
      RECT 38.16 1.88 38.25 2.51 ;
      RECT 38.125 1.93 38.13 2.51 ;
      RECT 38.07 1.955 38.08 2.51 ;
      RECT 38.025 1.955 38.035 2.51 ;
      RECT 38.395 1.88 38.44 2.16 ;
      RECT 37.245 1.61 37.445 1.75 ;
      RECT 38.361 1.88 38.395 2.172 ;
      RECT 38.275 1.88 38.361 2.212 ;
      RECT 38.26 1.88 38.275 2.253 ;
      RECT 38.255 1.88 38.26 2.273 ;
      RECT 38.25 1.88 38.255 2.293 ;
      RECT 38.13 1.922 38.16 2.51 ;
      RECT 38.08 1.942 38.125 2.51 ;
      RECT 38.065 1.957 38.07 2.51 ;
      RECT 38.035 1.957 38.065 2.51 ;
      RECT 37.99 1.942 38.025 2.51 ;
      RECT 37.985 1.93 37.99 2.29 ;
      RECT 37.98 1.927 37.985 2.27 ;
      RECT 37.965 1.917 37.98 2.223 ;
      RECT 37.96 1.91 37.965 2.186 ;
      RECT 37.955 1.907 37.96 2.169 ;
      RECT 37.94 1.897 37.955 2.125 ;
      RECT 37.935 1.888 37.94 2.085 ;
      RECT 37.93 1.884 37.935 2.07 ;
      RECT 37.92 1.878 37.93 2.053 ;
      RECT 37.88 1.859 37.92 2.028 ;
      RECT 37.875 1.841 37.88 2.008 ;
      RECT 37.865 1.835 37.875 2.003 ;
      RECT 37.835 1.819 37.865 1.99 ;
      RECT 37.82 1.801 37.835 1.973 ;
      RECT 37.805 1.789 37.82 1.96 ;
      RECT 37.8 1.781 37.805 1.953 ;
      RECT 37.77 1.767 37.8 1.94 ;
      RECT 37.765 1.752 37.77 1.928 ;
      RECT 37.755 1.746 37.765 1.92 ;
      RECT 37.735 1.734 37.755 1.908 ;
      RECT 37.725 1.722 37.735 1.895 ;
      RECT 37.695 1.706 37.725 1.88 ;
      RECT 37.675 1.686 37.695 1.863 ;
      RECT 37.67 1.676 37.675 1.853 ;
      RECT 37.645 1.664 37.67 1.84 ;
      RECT 37.64 1.652 37.645 1.828 ;
      RECT 37.635 1.647 37.64 1.824 ;
      RECT 37.62 1.64 37.635 1.816 ;
      RECT 37.61 1.627 37.62 1.806 ;
      RECT 37.605 1.625 37.61 1.8 ;
      RECT 37.58 1.618 37.605 1.789 ;
      RECT 37.575 1.611 37.58 1.778 ;
      RECT 37.55 1.61 37.575 1.765 ;
      RECT 37.531 1.61 37.55 1.755 ;
      RECT 37.445 1.61 37.531 1.752 ;
      RECT 37.215 1.61 37.245 1.755 ;
      RECT 37.175 1.617 37.215 1.768 ;
      RECT 37.15 1.627 37.175 1.781 ;
      RECT 37.135 1.636 37.15 1.791 ;
      RECT 37.105 1.641 37.135 1.81 ;
      RECT 37.1 1.647 37.105 1.828 ;
      RECT 37.08 1.657 37.1 1.843 ;
      RECT 37.07 1.67 37.08 1.863 ;
      RECT 37.055 1.682 37.07 1.88 ;
      RECT 37.05 1.692 37.055 1.89 ;
      RECT 37.045 1.697 37.05 1.895 ;
      RECT 37.035 1.705 37.045 1.908 ;
      RECT 36.985 1.737 37.035 1.945 ;
      RECT 36.97 1.772 36.985 1.986 ;
      RECT 36.965 1.782 36.97 2.001 ;
      RECT 36.96 1.787 36.965 2.008 ;
      RECT 36.935 1.803 36.96 2.028 ;
      RECT 36.92 1.824 36.935 2.053 ;
      RECT 36.895 1.845 36.92 2.078 ;
      RECT 36.885 1.864 36.895 2.101 ;
      RECT 36.86 1.882 36.885 2.124 ;
      RECT 36.845 1.902 36.86 2.148 ;
      RECT 36.84 1.912 36.845 2.16 ;
      RECT 36.825 1.924 36.84 2.18 ;
      RECT 36.815 1.939 36.825 2.22 ;
      RECT 36.81 1.947 36.815 2.248 ;
      RECT 36.8 1.957 36.81 2.268 ;
      RECT 36.795 1.97 36.8 2.293 ;
      RECT 36.79 1.983 36.795 2.313 ;
      RECT 36.785 1.989 36.79 2.335 ;
      RECT 36.775 1.998 36.785 2.355 ;
      RECT 36.77 2.018 36.775 2.378 ;
      RECT 36.765 2.024 36.77 2.398 ;
      RECT 36.76 2.031 36.765 2.42 ;
      RECT 36.755 2.042 36.76 2.433 ;
      RECT 36.745 2.052 36.755 2.458 ;
      RECT 36.725 2.077 36.745 2.64 ;
      RECT 36.695 2.117 36.725 2.64 ;
      RECT 36.69 2.147 36.695 2.64 ;
      RECT 36.665 2.175 36.685 2.64 ;
      RECT 36.635 2.22 36.665 2.64 ;
      RECT 36.63 2.247 36.635 2.64 ;
      RECT 36.61 2.265 36.63 2.64 ;
      RECT 36.6 2.29 36.61 2.64 ;
      RECT 36.595 2.302 36.6 2.64 ;
      RECT 36.58 2.325 36.595 2.64 ;
      RECT 36.56 2.352 36.575 2.64 ;
      RECT 36.55 2.375 36.56 2.64 ;
      RECT 38.34 3.26 38.42 3.52 ;
      RECT 37.575 2.48 37.645 2.74 ;
      RECT 38.306 3.227 38.34 3.52 ;
      RECT 38.22 3.13 38.306 3.52 ;
      RECT 38.2 3.042 38.22 3.52 ;
      RECT 38.19 3.012 38.2 3.52 ;
      RECT 38.18 2.992 38.19 3.52 ;
      RECT 38.16 2.979 38.18 3.52 ;
      RECT 38.145 2.969 38.16 3.348 ;
      RECT 38.14 2.962 38.145 3.303 ;
      RECT 38.13 2.956 38.14 3.293 ;
      RECT 38.12 2.948 38.13 3.275 ;
      RECT 38.115 2.942 38.12 3.263 ;
      RECT 38.105 2.937 38.115 3.25 ;
      RECT 38.085 2.927 38.105 3.223 ;
      RECT 38.045 2.906 38.085 3.175 ;
      RECT 38.03 2.887 38.045 3.133 ;
      RECT 38.005 2.873 38.03 3.103 ;
      RECT 37.995 2.861 38.005 3.07 ;
      RECT 37.99 2.856 37.995 3.06 ;
      RECT 37.96 2.842 37.99 3.04 ;
      RECT 37.95 2.826 37.96 3.013 ;
      RECT 37.945 2.821 37.95 3.003 ;
      RECT 37.92 2.812 37.945 2.983 ;
      RECT 37.91 2.8 37.92 2.963 ;
      RECT 37.84 2.768 37.91 2.938 ;
      RECT 37.835 2.737 37.84 2.915 ;
      RECT 37.786 2.48 37.835 2.898 ;
      RECT 37.7 2.48 37.786 2.857 ;
      RECT 37.645 2.48 37.7 2.785 ;
      RECT 37.735 3.265 37.895 3.525 ;
      RECT 37.26 1.88 37.31 2.565 ;
      RECT 37.05 2.305 37.085 2.565 ;
      RECT 37.365 1.88 37.37 2.34 ;
      RECT 37.455 1.88 37.48 2.16 ;
      RECT 37.73 3.262 37.735 3.525 ;
      RECT 37.695 3.25 37.73 3.525 ;
      RECT 37.635 3.223 37.695 3.525 ;
      RECT 37.63 3.206 37.635 3.379 ;
      RECT 37.625 3.203 37.63 3.366 ;
      RECT 37.605 3.196 37.625 3.353 ;
      RECT 37.57 3.179 37.605 3.335 ;
      RECT 37.53 3.158 37.57 3.315 ;
      RECT 37.525 3.146 37.53 3.303 ;
      RECT 37.485 3.132 37.525 3.289 ;
      RECT 37.465 3.115 37.485 3.271 ;
      RECT 37.455 3.107 37.465 3.263 ;
      RECT 37.44 1.88 37.455 2.178 ;
      RECT 37.425 3.097 37.455 3.25 ;
      RECT 37.41 1.88 37.44 2.223 ;
      RECT 37.415 3.087 37.425 3.237 ;
      RECT 37.385 3.072 37.415 3.224 ;
      RECT 37.37 1.88 37.41 2.29 ;
      RECT 37.37 3.04 37.385 3.21 ;
      RECT 37.365 3.012 37.37 3.204 ;
      RECT 37.36 1.88 37.365 2.345 ;
      RECT 37.35 2.982 37.365 3.198 ;
      RECT 37.355 1.88 37.36 2.358 ;
      RECT 37.345 1.88 37.355 2.378 ;
      RECT 37.31 2.895 37.35 3.183 ;
      RECT 37.31 1.88 37.345 2.418 ;
      RECT 37.305 2.827 37.31 3.171 ;
      RECT 37.29 2.782 37.305 3.166 ;
      RECT 37.285 2.72 37.29 3.161 ;
      RECT 37.26 2.627 37.285 3.154 ;
      RECT 37.255 1.88 37.26 3.146 ;
      RECT 37.24 1.88 37.255 3.133 ;
      RECT 37.22 1.88 37.24 3.09 ;
      RECT 37.21 1.88 37.22 3.04 ;
      RECT 37.205 1.88 37.21 3.013 ;
      RECT 37.2 1.88 37.205 2.991 ;
      RECT 37.195 2.106 37.2 2.974 ;
      RECT 37.19 2.128 37.195 2.952 ;
      RECT 37.185 2.17 37.19 2.935 ;
      RECT 37.155 2.22 37.185 2.879 ;
      RECT 37.15 2.247 37.155 2.821 ;
      RECT 37.135 2.265 37.15 2.785 ;
      RECT 37.13 2.283 37.135 2.749 ;
      RECT 37.124 2.29 37.13 2.73 ;
      RECT 37.12 2.297 37.124 2.713 ;
      RECT 37.115 2.302 37.12 2.682 ;
      RECT 37.105 2.305 37.115 2.657 ;
      RECT 37.095 2.305 37.105 2.623 ;
      RECT 37.09 2.305 37.095 2.6 ;
      RECT 37.085 2.305 37.09 2.58 ;
      RECT 36 2.44 36.28 2.72 ;
      RECT 36 2.44 36.3 2.615 ;
      RECT 36.09 2.33 36.35 2.59 ;
      RECT 36.055 2.425 36.35 2.59 ;
      RECT 36.18 0.945 36.345 2.59 ;
      RECT 36.08 0.945 36.45 1.315 ;
      RECT 35.705 3.47 35.965 3.73 ;
      RECT 35.725 3.397 35.905 3.73 ;
      RECT 35.725 3.14 35.9 3.73 ;
      RECT 35.725 2.932 35.89 3.73 ;
      RECT 35.73 2.85 35.89 3.73 ;
      RECT 35.73 2.615 35.88 3.73 ;
      RECT 35.73 2.462 35.875 3.73 ;
      RECT 35.735 2.447 35.875 3.73 ;
      RECT 35.785 2.162 35.875 3.73 ;
      RECT 35.74 2.397 35.875 3.73 ;
      RECT 35.77 2.215 35.875 3.73 ;
      RECT 35.755 2.327 35.875 3.73 ;
      RECT 35.76 2.285 35.875 3.73 ;
      RECT 35.755 2.327 35.89 2.39 ;
      RECT 35.79 1.915 35.895 2.335 ;
      RECT 35.79 1.915 35.91 2.318 ;
      RECT 35.79 1.915 35.945 2.28 ;
      RECT 35.785 2.162 35.995 2.213 ;
      RECT 35.79 1.915 36.05 2.175 ;
      RECT 35.05 2.62 35.31 2.88 ;
      RECT 35.05 2.62 35.32 2.838 ;
      RECT 35.05 2.62 35.406 2.809 ;
      RECT 35.05 2.62 35.475 2.761 ;
      RECT 35.05 2.62 35.51 2.73 ;
      RECT 35.28 2.44 35.56 2.72 ;
      RECT 35.115 2.605 35.56 2.72 ;
      RECT 35.205 2.482 35.31 2.88 ;
      RECT 35.135 2.545 35.56 2.72 ;
      RECT 29.585 6.22 29.905 6.545 ;
      RECT 29.615 5.695 29.785 6.545 ;
      RECT 29.615 5.695 29.79 6.045 ;
      RECT 29.615 5.695 30.59 5.87 ;
      RECT 30.415 1.965 30.59 5.87 ;
      RECT 30.36 1.965 30.71 2.315 ;
      RECT 30.385 6.655 30.71 6.98 ;
      RECT 29.27 6.745 30.71 6.915 ;
      RECT 29.27 2.395 29.43 6.915 ;
      RECT 29.585 2.365 29.905 2.685 ;
      RECT 29.27 2.395 29.905 2.565 ;
      RECT 27.935 2.705 28.32 3.055 ;
      RECT 27.925 2.77 28.32 2.97 ;
      RECT 28.07 2.7 28.24 3.055 ;
      RECT 26.38 2.44 26.66 2.72 ;
      RECT 26.375 2.44 26.66 2.673 ;
      RECT 26.355 2.44 26.66 2.65 ;
      RECT 26.345 2.44 26.66 2.63 ;
      RECT 26.335 2.44 26.66 2.615 ;
      RECT 26.31 2.44 26.66 2.588 ;
      RECT 26.3 2.44 26.66 2.563 ;
      RECT 26.255 2.295 26.535 2.555 ;
      RECT 26.255 2.39 26.635 2.555 ;
      RECT 26.255 2.335 26.58 2.555 ;
      RECT 26.255 2.327 26.575 2.555 ;
      RECT 26.255 2.317 26.57 2.555 ;
      RECT 26.255 2.305 26.565 2.555 ;
      RECT 25.18 3 25.46 3.28 ;
      RECT 25.18 3 25.495 3.26 ;
      RECT 17.505 6.655 17.855 7.005 ;
      RECT 24.925 6.61 25.275 6.96 ;
      RECT 17.505 6.685 25.275 6.885 ;
      RECT 25.215 2.42 25.265 2.68 ;
      RECT 25.005 2.42 25.01 2.68 ;
      RECT 24.2 1.975 24.23 2.235 ;
      RECT 23.97 1.975 24.045 2.235 ;
      RECT 25.19 2.37 25.215 2.68 ;
      RECT 25.185 2.327 25.19 2.68 ;
      RECT 25.18 2.31 25.185 2.68 ;
      RECT 25.175 2.297 25.18 2.68 ;
      RECT 25.1 2.18 25.175 2.68 ;
      RECT 25.055 1.997 25.1 2.68 ;
      RECT 25.05 1.925 25.055 2.68 ;
      RECT 25.035 1.9 25.05 2.68 ;
      RECT 25.01 1.862 25.035 2.68 ;
      RECT 25 1.842 25.01 2.402 ;
      RECT 24.985 1.834 25 2.357 ;
      RECT 24.98 1.826 24.985 2.328 ;
      RECT 24.975 1.823 24.98 2.308 ;
      RECT 24.97 1.82 24.975 2.288 ;
      RECT 24.965 1.817 24.97 2.268 ;
      RECT 24.935 1.806 24.965 2.205 ;
      RECT 24.915 1.791 24.935 2.12 ;
      RECT 24.91 1.783 24.915 2.083 ;
      RECT 24.9 1.777 24.91 2.05 ;
      RECT 24.885 1.769 24.9 2.01 ;
      RECT 24.88 1.762 24.885 1.97 ;
      RECT 24.875 1.759 24.88 1.948 ;
      RECT 24.87 1.756 24.875 1.935 ;
      RECT 24.865 1.755 24.87 1.925 ;
      RECT 24.85 1.749 24.865 1.915 ;
      RECT 24.825 1.736 24.85 1.9 ;
      RECT 24.775 1.711 24.825 1.871 ;
      RECT 24.76 1.69 24.775 1.846 ;
      RECT 24.75 1.683 24.76 1.835 ;
      RECT 24.695 1.664 24.75 1.808 ;
      RECT 24.67 1.642 24.695 1.781 ;
      RECT 24.665 1.635 24.67 1.776 ;
      RECT 24.65 1.635 24.665 1.774 ;
      RECT 24.625 1.627 24.65 1.77 ;
      RECT 24.61 1.625 24.625 1.766 ;
      RECT 24.58 1.625 24.61 1.763 ;
      RECT 24.57 1.625 24.58 1.758 ;
      RECT 24.525 1.625 24.57 1.756 ;
      RECT 24.496 1.625 24.525 1.757 ;
      RECT 24.41 1.625 24.496 1.759 ;
      RECT 24.396 1.626 24.41 1.761 ;
      RECT 24.31 1.627 24.396 1.763 ;
      RECT 24.295 1.628 24.31 1.773 ;
      RECT 24.29 1.629 24.295 1.782 ;
      RECT 24.27 1.632 24.29 1.792 ;
      RECT 24.255 1.64 24.27 1.807 ;
      RECT 24.235 1.658 24.255 1.822 ;
      RECT 24.225 1.67 24.235 1.845 ;
      RECT 24.215 1.679 24.225 1.875 ;
      RECT 24.2 1.691 24.215 1.92 ;
      RECT 24.145 1.724 24.2 2.235 ;
      RECT 24.14 1.752 24.145 2.235 ;
      RECT 24.12 1.767 24.14 2.235 ;
      RECT 24.085 1.827 24.12 2.235 ;
      RECT 24.083 1.877 24.085 2.235 ;
      RECT 24.08 1.885 24.083 2.235 ;
      RECT 24.07 1.9 24.08 2.235 ;
      RECT 24.065 1.912 24.07 2.235 ;
      RECT 24.055 1.937 24.065 2.235 ;
      RECT 24.045 1.965 24.055 2.235 ;
      RECT 21.95 3.47 22 3.73 ;
      RECT 24.86 3.02 24.92 3.28 ;
      RECT 24.845 3.02 24.86 3.29 ;
      RECT 24.826 3.02 24.845 3.323 ;
      RECT 24.74 3.02 24.826 3.448 ;
      RECT 24.66 3.02 24.74 3.63 ;
      RECT 24.655 3.257 24.66 3.715 ;
      RECT 24.63 3.327 24.655 3.743 ;
      RECT 24.625 3.397 24.63 3.77 ;
      RECT 24.605 3.469 24.625 3.792 ;
      RECT 24.6 3.536 24.605 3.815 ;
      RECT 24.59 3.565 24.6 3.83 ;
      RECT 24.58 3.587 24.59 3.847 ;
      RECT 24.575 3.597 24.58 3.858 ;
      RECT 24.57 3.605 24.575 3.866 ;
      RECT 24.56 3.613 24.57 3.878 ;
      RECT 24.555 3.625 24.56 3.888 ;
      RECT 24.55 3.633 24.555 3.893 ;
      RECT 24.53 3.651 24.55 3.903 ;
      RECT 24.525 3.668 24.53 3.91 ;
      RECT 24.52 3.676 24.525 3.911 ;
      RECT 24.515 3.687 24.52 3.913 ;
      RECT 24.475 3.725 24.515 3.923 ;
      RECT 24.47 3.76 24.475 3.934 ;
      RECT 24.465 3.765 24.47 3.937 ;
      RECT 24.44 3.775 24.465 3.944 ;
      RECT 24.43 3.789 24.44 3.953 ;
      RECT 24.41 3.801 24.43 3.956 ;
      RECT 24.36 3.82 24.41 3.96 ;
      RECT 24.315 3.835 24.36 3.965 ;
      RECT 24.25 3.838 24.315 3.971 ;
      RECT 24.235 3.836 24.25 3.978 ;
      RECT 24.205 3.835 24.235 3.978 ;
      RECT 24.166 3.834 24.205 3.974 ;
      RECT 24.08 3.831 24.166 3.97 ;
      RECT 24.063 3.829 24.08 3.967 ;
      RECT 23.977 3.827 24.063 3.964 ;
      RECT 23.891 3.824 23.977 3.958 ;
      RECT 23.805 3.82 23.891 3.953 ;
      RECT 23.727 3.817 23.805 3.949 ;
      RECT 23.641 3.814 23.727 3.947 ;
      RECT 23.555 3.811 23.641 3.944 ;
      RECT 23.497 3.809 23.555 3.941 ;
      RECT 23.411 3.806 23.497 3.939 ;
      RECT 23.325 3.802 23.411 3.937 ;
      RECT 23.239 3.799 23.325 3.934 ;
      RECT 23.153 3.795 23.239 3.932 ;
      RECT 23.067 3.791 23.153 3.929 ;
      RECT 22.981 3.788 23.067 3.927 ;
      RECT 22.895 3.784 22.981 3.924 ;
      RECT 22.809 3.781 22.895 3.922 ;
      RECT 22.723 3.777 22.809 3.919 ;
      RECT 22.637 3.774 22.723 3.917 ;
      RECT 22.551 3.77 22.637 3.914 ;
      RECT 22.465 3.767 22.551 3.912 ;
      RECT 22.455 3.765 22.465 3.908 ;
      RECT 22.45 3.765 22.455 3.906 ;
      RECT 22.41 3.76 22.45 3.9 ;
      RECT 22.396 3.751 22.41 3.893 ;
      RECT 22.31 3.721 22.396 3.878 ;
      RECT 22.29 3.687 22.31 3.863 ;
      RECT 22.22 3.656 22.29 3.85 ;
      RECT 22.215 3.631 22.22 3.839 ;
      RECT 22.21 3.625 22.215 3.837 ;
      RECT 22.141 3.47 22.21 3.825 ;
      RECT 22.055 3.47 22.141 3.799 ;
      RECT 22.03 3.47 22.055 3.778 ;
      RECT 22.025 3.47 22.03 3.768 ;
      RECT 22.02 3.47 22.025 3.76 ;
      RECT 22 3.47 22.02 3.743 ;
      RECT 24.42 2.04 24.68 2.3 ;
      RECT 24.405 2.04 24.68 2.203 ;
      RECT 24.375 2.04 24.68 2.178 ;
      RECT 24.34 1.88 24.62 2.16 ;
      RECT 24.31 3.37 24.37 3.63 ;
      RECT 23.335 2.06 23.39 2.32 ;
      RECT 24.27 3.327 24.31 3.63 ;
      RECT 24.241 3.248 24.27 3.63 ;
      RECT 24.155 3.12 24.241 3.63 ;
      RECT 24.135 3 24.155 3.63 ;
      RECT 24.11 2.951 24.135 3.63 ;
      RECT 24.105 2.916 24.11 3.48 ;
      RECT 24.075 2.876 24.105 3.418 ;
      RECT 24.05 2.813 24.075 3.333 ;
      RECT 24.04 2.775 24.05 3.27 ;
      RECT 24.025 2.75 24.04 3.231 ;
      RECT 23.982 2.708 24.025 3.137 ;
      RECT 23.98 2.681 23.982 3.064 ;
      RECT 23.975 2.676 23.98 3.055 ;
      RECT 23.97 2.669 23.975 3.03 ;
      RECT 23.965 2.663 23.97 3.015 ;
      RECT 23.96 2.657 23.965 3.003 ;
      RECT 23.95 2.648 23.96 2.985 ;
      RECT 23.945 2.639 23.95 2.963 ;
      RECT 23.92 2.62 23.945 2.913 ;
      RECT 23.915 2.601 23.92 2.863 ;
      RECT 23.9 2.587 23.915 2.823 ;
      RECT 23.895 2.573 23.9 2.79 ;
      RECT 23.89 2.566 23.895 2.783 ;
      RECT 23.875 2.553 23.89 2.775 ;
      RECT 23.83 2.515 23.875 2.748 ;
      RECT 23.8 2.468 23.83 2.713 ;
      RECT 23.78 2.437 23.8 2.69 ;
      RECT 23.7 2.37 23.78 2.643 ;
      RECT 23.67 2.3 23.7 2.59 ;
      RECT 23.665 2.277 23.67 2.573 ;
      RECT 23.635 2.255 23.665 2.558 ;
      RECT 23.605 2.214 23.635 2.53 ;
      RECT 23.6 2.189 23.605 2.515 ;
      RECT 23.595 2.183 23.6 2.508 ;
      RECT 23.585 2.06 23.595 2.5 ;
      RECT 23.575 2.06 23.585 2.493 ;
      RECT 23.57 2.06 23.575 2.485 ;
      RECT 23.55 2.06 23.57 2.473 ;
      RECT 23.5 2.06 23.55 2.443 ;
      RECT 23.445 2.06 23.5 2.393 ;
      RECT 23.415 2.06 23.445 2.353 ;
      RECT 23.39 2.06 23.415 2.33 ;
      RECT 23.26 2.785 23.54 3.065 ;
      RECT 23.225 2.7 23.485 2.96 ;
      RECT 23.225 2.782 23.495 2.96 ;
      RECT 21.425 2.155 21.43 2.64 ;
      RECT 21.315 2.34 21.32 2.64 ;
      RECT 21.225 2.38 21.29 2.64 ;
      RECT 22.9 1.88 22.99 2.51 ;
      RECT 22.865 1.93 22.87 2.51 ;
      RECT 22.81 1.955 22.82 2.51 ;
      RECT 22.765 1.955 22.775 2.51 ;
      RECT 23.135 1.88 23.18 2.16 ;
      RECT 21.985 1.61 22.185 1.75 ;
      RECT 23.101 1.88 23.135 2.172 ;
      RECT 23.015 1.88 23.101 2.212 ;
      RECT 23 1.88 23.015 2.253 ;
      RECT 22.995 1.88 23 2.273 ;
      RECT 22.99 1.88 22.995 2.293 ;
      RECT 22.87 1.922 22.9 2.51 ;
      RECT 22.82 1.942 22.865 2.51 ;
      RECT 22.805 1.957 22.81 2.51 ;
      RECT 22.775 1.957 22.805 2.51 ;
      RECT 22.73 1.942 22.765 2.51 ;
      RECT 22.725 1.93 22.73 2.29 ;
      RECT 22.72 1.927 22.725 2.27 ;
      RECT 22.705 1.917 22.72 2.223 ;
      RECT 22.7 1.91 22.705 2.186 ;
      RECT 22.695 1.907 22.7 2.169 ;
      RECT 22.68 1.897 22.695 2.125 ;
      RECT 22.675 1.888 22.68 2.085 ;
      RECT 22.67 1.884 22.675 2.07 ;
      RECT 22.66 1.878 22.67 2.053 ;
      RECT 22.62 1.859 22.66 2.028 ;
      RECT 22.615 1.841 22.62 2.008 ;
      RECT 22.605 1.835 22.615 2.003 ;
      RECT 22.575 1.819 22.605 1.99 ;
      RECT 22.56 1.801 22.575 1.973 ;
      RECT 22.545 1.789 22.56 1.96 ;
      RECT 22.54 1.781 22.545 1.953 ;
      RECT 22.51 1.767 22.54 1.94 ;
      RECT 22.505 1.752 22.51 1.928 ;
      RECT 22.495 1.746 22.505 1.92 ;
      RECT 22.475 1.734 22.495 1.908 ;
      RECT 22.465 1.722 22.475 1.895 ;
      RECT 22.435 1.706 22.465 1.88 ;
      RECT 22.415 1.686 22.435 1.863 ;
      RECT 22.41 1.676 22.415 1.853 ;
      RECT 22.385 1.664 22.41 1.84 ;
      RECT 22.38 1.652 22.385 1.828 ;
      RECT 22.375 1.647 22.38 1.824 ;
      RECT 22.36 1.64 22.375 1.816 ;
      RECT 22.35 1.627 22.36 1.806 ;
      RECT 22.345 1.625 22.35 1.8 ;
      RECT 22.32 1.618 22.345 1.789 ;
      RECT 22.315 1.611 22.32 1.778 ;
      RECT 22.29 1.61 22.315 1.765 ;
      RECT 22.271 1.61 22.29 1.755 ;
      RECT 22.185 1.61 22.271 1.752 ;
      RECT 21.955 1.61 21.985 1.755 ;
      RECT 21.915 1.617 21.955 1.768 ;
      RECT 21.89 1.627 21.915 1.781 ;
      RECT 21.875 1.636 21.89 1.791 ;
      RECT 21.845 1.641 21.875 1.81 ;
      RECT 21.84 1.647 21.845 1.828 ;
      RECT 21.82 1.657 21.84 1.843 ;
      RECT 21.81 1.67 21.82 1.863 ;
      RECT 21.795 1.682 21.81 1.88 ;
      RECT 21.79 1.692 21.795 1.89 ;
      RECT 21.785 1.697 21.79 1.895 ;
      RECT 21.775 1.705 21.785 1.908 ;
      RECT 21.725 1.737 21.775 1.945 ;
      RECT 21.71 1.772 21.725 1.986 ;
      RECT 21.705 1.782 21.71 2.001 ;
      RECT 21.7 1.787 21.705 2.008 ;
      RECT 21.675 1.803 21.7 2.028 ;
      RECT 21.66 1.824 21.675 2.053 ;
      RECT 21.635 1.845 21.66 2.078 ;
      RECT 21.625 1.864 21.635 2.101 ;
      RECT 21.6 1.882 21.625 2.124 ;
      RECT 21.585 1.902 21.6 2.148 ;
      RECT 21.58 1.912 21.585 2.16 ;
      RECT 21.565 1.924 21.58 2.18 ;
      RECT 21.555 1.939 21.565 2.22 ;
      RECT 21.55 1.947 21.555 2.248 ;
      RECT 21.54 1.957 21.55 2.268 ;
      RECT 21.535 1.97 21.54 2.293 ;
      RECT 21.53 1.983 21.535 2.313 ;
      RECT 21.525 1.989 21.53 2.335 ;
      RECT 21.515 1.998 21.525 2.355 ;
      RECT 21.51 2.018 21.515 2.378 ;
      RECT 21.505 2.024 21.51 2.398 ;
      RECT 21.5 2.031 21.505 2.42 ;
      RECT 21.495 2.042 21.5 2.433 ;
      RECT 21.485 2.052 21.495 2.458 ;
      RECT 21.465 2.077 21.485 2.64 ;
      RECT 21.435 2.117 21.465 2.64 ;
      RECT 21.43 2.147 21.435 2.64 ;
      RECT 21.405 2.175 21.425 2.64 ;
      RECT 21.375 2.22 21.405 2.64 ;
      RECT 21.37 2.247 21.375 2.64 ;
      RECT 21.35 2.265 21.37 2.64 ;
      RECT 21.34 2.29 21.35 2.64 ;
      RECT 21.335 2.302 21.34 2.64 ;
      RECT 21.32 2.325 21.335 2.64 ;
      RECT 21.3 2.352 21.315 2.64 ;
      RECT 21.29 2.375 21.3 2.64 ;
      RECT 23.08 3.26 23.16 3.52 ;
      RECT 22.315 2.48 22.385 2.74 ;
      RECT 23.046 3.227 23.08 3.52 ;
      RECT 22.96 3.13 23.046 3.52 ;
      RECT 22.94 3.042 22.96 3.52 ;
      RECT 22.93 3.012 22.94 3.52 ;
      RECT 22.92 2.992 22.93 3.52 ;
      RECT 22.9 2.979 22.92 3.52 ;
      RECT 22.885 2.969 22.9 3.348 ;
      RECT 22.88 2.962 22.885 3.303 ;
      RECT 22.87 2.956 22.88 3.293 ;
      RECT 22.86 2.948 22.87 3.275 ;
      RECT 22.855 2.942 22.86 3.263 ;
      RECT 22.845 2.937 22.855 3.25 ;
      RECT 22.825 2.927 22.845 3.223 ;
      RECT 22.785 2.906 22.825 3.175 ;
      RECT 22.77 2.887 22.785 3.133 ;
      RECT 22.745 2.873 22.77 3.103 ;
      RECT 22.735 2.861 22.745 3.07 ;
      RECT 22.73 2.856 22.735 3.06 ;
      RECT 22.7 2.842 22.73 3.04 ;
      RECT 22.69 2.826 22.7 3.013 ;
      RECT 22.685 2.821 22.69 3.003 ;
      RECT 22.66 2.812 22.685 2.983 ;
      RECT 22.65 2.8 22.66 2.963 ;
      RECT 22.58 2.768 22.65 2.938 ;
      RECT 22.575 2.737 22.58 2.915 ;
      RECT 22.526 2.48 22.575 2.898 ;
      RECT 22.44 2.48 22.526 2.857 ;
      RECT 22.385 2.48 22.44 2.785 ;
      RECT 22.475 3.265 22.635 3.525 ;
      RECT 22 1.88 22.05 2.565 ;
      RECT 21.79 2.305 21.825 2.565 ;
      RECT 22.105 1.88 22.11 2.34 ;
      RECT 22.195 1.88 22.22 2.16 ;
      RECT 22.47 3.262 22.475 3.525 ;
      RECT 22.435 3.25 22.47 3.525 ;
      RECT 22.375 3.223 22.435 3.525 ;
      RECT 22.37 3.206 22.375 3.379 ;
      RECT 22.365 3.203 22.37 3.366 ;
      RECT 22.345 3.196 22.365 3.353 ;
      RECT 22.31 3.179 22.345 3.335 ;
      RECT 22.27 3.158 22.31 3.315 ;
      RECT 22.265 3.146 22.27 3.303 ;
      RECT 22.225 3.132 22.265 3.289 ;
      RECT 22.205 3.115 22.225 3.271 ;
      RECT 22.195 3.107 22.205 3.263 ;
      RECT 22.18 1.88 22.195 2.178 ;
      RECT 22.165 3.097 22.195 3.25 ;
      RECT 22.15 1.88 22.18 2.223 ;
      RECT 22.155 3.087 22.165 3.237 ;
      RECT 22.125 3.072 22.155 3.224 ;
      RECT 22.11 1.88 22.15 2.29 ;
      RECT 22.11 3.04 22.125 3.21 ;
      RECT 22.105 3.012 22.11 3.204 ;
      RECT 22.1 1.88 22.105 2.345 ;
      RECT 22.09 2.982 22.105 3.198 ;
      RECT 22.095 1.88 22.1 2.358 ;
      RECT 22.085 1.88 22.095 2.378 ;
      RECT 22.05 2.895 22.09 3.183 ;
      RECT 22.05 1.88 22.085 2.418 ;
      RECT 22.045 2.827 22.05 3.171 ;
      RECT 22.03 2.782 22.045 3.166 ;
      RECT 22.025 2.72 22.03 3.161 ;
      RECT 22 2.627 22.025 3.154 ;
      RECT 21.995 1.88 22 3.146 ;
      RECT 21.98 1.88 21.995 3.133 ;
      RECT 21.96 1.88 21.98 3.09 ;
      RECT 21.95 1.88 21.96 3.04 ;
      RECT 21.945 1.88 21.95 3.013 ;
      RECT 21.94 1.88 21.945 2.991 ;
      RECT 21.935 2.106 21.94 2.974 ;
      RECT 21.93 2.128 21.935 2.952 ;
      RECT 21.925 2.17 21.93 2.935 ;
      RECT 21.895 2.22 21.925 2.879 ;
      RECT 21.89 2.247 21.895 2.821 ;
      RECT 21.875 2.265 21.89 2.785 ;
      RECT 21.87 2.283 21.875 2.749 ;
      RECT 21.864 2.29 21.87 2.73 ;
      RECT 21.86 2.297 21.864 2.713 ;
      RECT 21.855 2.302 21.86 2.682 ;
      RECT 21.845 2.305 21.855 2.657 ;
      RECT 21.835 2.305 21.845 2.623 ;
      RECT 21.83 2.305 21.835 2.6 ;
      RECT 21.825 2.305 21.83 2.58 ;
      RECT 20.74 2.44 21.02 2.72 ;
      RECT 20.74 2.44 21.04 2.615 ;
      RECT 20.83 2.33 21.09 2.59 ;
      RECT 20.795 2.425 21.09 2.59 ;
      RECT 20.92 0.945 21.085 2.59 ;
      RECT 20.82 0.945 21.19 1.315 ;
      RECT 20.445 3.47 20.705 3.73 ;
      RECT 20.465 3.397 20.645 3.73 ;
      RECT 20.465 3.14 20.64 3.73 ;
      RECT 20.465 2.932 20.63 3.73 ;
      RECT 20.47 2.85 20.63 3.73 ;
      RECT 20.47 2.615 20.62 3.73 ;
      RECT 20.47 2.462 20.615 3.73 ;
      RECT 20.475 2.447 20.615 3.73 ;
      RECT 20.525 2.162 20.615 3.73 ;
      RECT 20.48 2.397 20.615 3.73 ;
      RECT 20.51 2.215 20.615 3.73 ;
      RECT 20.495 2.327 20.615 3.73 ;
      RECT 20.5 2.285 20.615 3.73 ;
      RECT 20.495 2.327 20.63 2.39 ;
      RECT 20.53 1.915 20.635 2.335 ;
      RECT 20.53 1.915 20.65 2.318 ;
      RECT 20.53 1.915 20.685 2.28 ;
      RECT 20.525 2.162 20.735 2.213 ;
      RECT 20.53 1.915 20.79 2.175 ;
      RECT 19.79 2.62 20.05 2.88 ;
      RECT 19.79 2.62 20.06 2.838 ;
      RECT 19.79 2.62 20.146 2.809 ;
      RECT 19.79 2.62 20.215 2.761 ;
      RECT 19.79 2.62 20.25 2.73 ;
      RECT 20.02 2.44 20.3 2.72 ;
      RECT 19.855 2.605 20.3 2.72 ;
      RECT 19.945 2.482 20.05 2.88 ;
      RECT 19.875 2.545 20.3 2.72 ;
      RECT 14.325 6.22 14.645 6.545 ;
      RECT 14.355 5.695 14.525 6.545 ;
      RECT 14.355 5.695 14.53 6.045 ;
      RECT 14.355 5.695 15.33 5.87 ;
      RECT 15.155 1.965 15.33 5.87 ;
      RECT 15.1 1.965 15.45 2.315 ;
      RECT 15.125 6.655 15.45 6.98 ;
      RECT 14.01 6.745 15.45 6.915 ;
      RECT 14.01 2.395 14.17 6.915 ;
      RECT 14.325 2.365 14.645 2.685 ;
      RECT 14.01 2.395 14.645 2.565 ;
      RECT 12.675 2.705 13.06 3.055 ;
      RECT 12.665 2.77 13.06 2.97 ;
      RECT 12.81 2.7 12.98 3.055 ;
      RECT 11.12 2.44 11.4 2.72 ;
      RECT 11.115 2.44 11.4 2.673 ;
      RECT 11.095 2.44 11.4 2.65 ;
      RECT 11.085 2.44 11.4 2.63 ;
      RECT 11.075 2.44 11.4 2.615 ;
      RECT 11.05 2.44 11.4 2.588 ;
      RECT 11.04 2.44 11.4 2.563 ;
      RECT 10.995 2.295 11.275 2.555 ;
      RECT 10.995 2.39 11.375 2.555 ;
      RECT 10.995 2.335 11.32 2.555 ;
      RECT 10.995 2.327 11.315 2.555 ;
      RECT 10.995 2.317 11.31 2.555 ;
      RECT 10.995 2.305 11.305 2.555 ;
      RECT 9.92 3 10.2 3.28 ;
      RECT 9.92 3 10.235 3.26 ;
      RECT 1.54 6.995 1.83 7.345 ;
      RECT 1.54 7.07 2.905 7.24 ;
      RECT 2.735 6.685 2.905 7.24 ;
      RECT 9.665 6.605 10.015 6.955 ;
      RECT 2.735 6.685 10.015 6.855 ;
      RECT 9.955 2.42 10.005 2.68 ;
      RECT 9.745 2.42 9.75 2.68 ;
      RECT 8.94 1.975 8.97 2.235 ;
      RECT 8.71 1.975 8.785 2.235 ;
      RECT 9.93 2.37 9.955 2.68 ;
      RECT 9.925 2.327 9.93 2.68 ;
      RECT 9.92 2.31 9.925 2.68 ;
      RECT 9.915 2.297 9.92 2.68 ;
      RECT 9.84 2.18 9.915 2.68 ;
      RECT 9.795 1.997 9.84 2.68 ;
      RECT 9.79 1.925 9.795 2.68 ;
      RECT 9.775 1.9 9.79 2.68 ;
      RECT 9.75 1.862 9.775 2.68 ;
      RECT 9.74 1.842 9.75 2.402 ;
      RECT 9.725 1.834 9.74 2.357 ;
      RECT 9.72 1.826 9.725 2.328 ;
      RECT 9.715 1.823 9.72 2.308 ;
      RECT 9.71 1.82 9.715 2.288 ;
      RECT 9.705 1.817 9.71 2.268 ;
      RECT 9.675 1.806 9.705 2.205 ;
      RECT 9.655 1.791 9.675 2.12 ;
      RECT 9.65 1.783 9.655 2.083 ;
      RECT 9.64 1.777 9.65 2.05 ;
      RECT 9.625 1.769 9.64 2.01 ;
      RECT 9.62 1.762 9.625 1.97 ;
      RECT 9.615 1.759 9.62 1.948 ;
      RECT 9.61 1.756 9.615 1.935 ;
      RECT 9.605 1.755 9.61 1.925 ;
      RECT 9.59 1.749 9.605 1.915 ;
      RECT 9.565 1.736 9.59 1.9 ;
      RECT 9.515 1.711 9.565 1.871 ;
      RECT 9.5 1.69 9.515 1.846 ;
      RECT 9.49 1.683 9.5 1.835 ;
      RECT 9.435 1.664 9.49 1.808 ;
      RECT 9.41 1.642 9.435 1.781 ;
      RECT 9.405 1.635 9.41 1.776 ;
      RECT 9.39 1.635 9.405 1.774 ;
      RECT 9.365 1.627 9.39 1.77 ;
      RECT 9.35 1.625 9.365 1.766 ;
      RECT 9.32 1.625 9.35 1.763 ;
      RECT 9.31 1.625 9.32 1.758 ;
      RECT 9.265 1.625 9.31 1.756 ;
      RECT 9.236 1.625 9.265 1.757 ;
      RECT 9.15 1.625 9.236 1.759 ;
      RECT 9.136 1.626 9.15 1.761 ;
      RECT 9.05 1.627 9.136 1.763 ;
      RECT 9.035 1.628 9.05 1.773 ;
      RECT 9.03 1.629 9.035 1.782 ;
      RECT 9.01 1.632 9.03 1.792 ;
      RECT 8.995 1.64 9.01 1.807 ;
      RECT 8.975 1.658 8.995 1.822 ;
      RECT 8.965 1.67 8.975 1.845 ;
      RECT 8.955 1.679 8.965 1.875 ;
      RECT 8.94 1.691 8.955 1.92 ;
      RECT 8.885 1.724 8.94 2.235 ;
      RECT 8.88 1.752 8.885 2.235 ;
      RECT 8.86 1.767 8.88 2.235 ;
      RECT 8.825 1.827 8.86 2.235 ;
      RECT 8.823 1.877 8.825 2.235 ;
      RECT 8.82 1.885 8.823 2.235 ;
      RECT 8.81 1.9 8.82 2.235 ;
      RECT 8.805 1.912 8.81 2.235 ;
      RECT 8.795 1.937 8.805 2.235 ;
      RECT 8.785 1.965 8.795 2.235 ;
      RECT 6.69 3.47 6.74 3.73 ;
      RECT 9.6 3.02 9.66 3.28 ;
      RECT 9.585 3.02 9.6 3.29 ;
      RECT 9.566 3.02 9.585 3.323 ;
      RECT 9.48 3.02 9.566 3.448 ;
      RECT 9.4 3.02 9.48 3.63 ;
      RECT 9.395 3.257 9.4 3.715 ;
      RECT 9.37 3.327 9.395 3.743 ;
      RECT 9.365 3.397 9.37 3.77 ;
      RECT 9.345 3.469 9.365 3.792 ;
      RECT 9.34 3.536 9.345 3.815 ;
      RECT 9.33 3.565 9.34 3.83 ;
      RECT 9.32 3.587 9.33 3.847 ;
      RECT 9.315 3.597 9.32 3.858 ;
      RECT 9.31 3.605 9.315 3.866 ;
      RECT 9.3 3.613 9.31 3.878 ;
      RECT 9.295 3.625 9.3 3.888 ;
      RECT 9.29 3.633 9.295 3.893 ;
      RECT 9.27 3.651 9.29 3.903 ;
      RECT 9.265 3.668 9.27 3.91 ;
      RECT 9.26 3.676 9.265 3.911 ;
      RECT 9.255 3.687 9.26 3.913 ;
      RECT 9.215 3.725 9.255 3.923 ;
      RECT 9.21 3.76 9.215 3.934 ;
      RECT 9.205 3.765 9.21 3.937 ;
      RECT 9.18 3.775 9.205 3.944 ;
      RECT 9.17 3.789 9.18 3.953 ;
      RECT 9.15 3.801 9.17 3.956 ;
      RECT 9.1 3.82 9.15 3.96 ;
      RECT 9.055 3.835 9.1 3.965 ;
      RECT 8.99 3.838 9.055 3.971 ;
      RECT 8.975 3.836 8.99 3.978 ;
      RECT 8.945 3.835 8.975 3.978 ;
      RECT 8.906 3.834 8.945 3.974 ;
      RECT 8.82 3.831 8.906 3.97 ;
      RECT 8.803 3.829 8.82 3.967 ;
      RECT 8.717 3.827 8.803 3.964 ;
      RECT 8.631 3.824 8.717 3.958 ;
      RECT 8.545 3.82 8.631 3.953 ;
      RECT 8.467 3.817 8.545 3.949 ;
      RECT 8.381 3.814 8.467 3.947 ;
      RECT 8.295 3.811 8.381 3.944 ;
      RECT 8.237 3.809 8.295 3.941 ;
      RECT 8.151 3.806 8.237 3.939 ;
      RECT 8.065 3.802 8.151 3.937 ;
      RECT 7.979 3.799 8.065 3.934 ;
      RECT 7.893 3.795 7.979 3.932 ;
      RECT 7.807 3.791 7.893 3.929 ;
      RECT 7.721 3.788 7.807 3.927 ;
      RECT 7.635 3.784 7.721 3.924 ;
      RECT 7.549 3.781 7.635 3.922 ;
      RECT 7.463 3.777 7.549 3.919 ;
      RECT 7.377 3.774 7.463 3.917 ;
      RECT 7.291 3.77 7.377 3.914 ;
      RECT 7.205 3.767 7.291 3.912 ;
      RECT 7.195 3.765 7.205 3.908 ;
      RECT 7.19 3.765 7.195 3.906 ;
      RECT 7.15 3.76 7.19 3.9 ;
      RECT 7.136 3.751 7.15 3.893 ;
      RECT 7.05 3.721 7.136 3.878 ;
      RECT 7.03 3.687 7.05 3.863 ;
      RECT 6.96 3.656 7.03 3.85 ;
      RECT 6.955 3.631 6.96 3.839 ;
      RECT 6.95 3.625 6.955 3.837 ;
      RECT 6.881 3.47 6.95 3.825 ;
      RECT 6.795 3.47 6.881 3.799 ;
      RECT 6.77 3.47 6.795 3.778 ;
      RECT 6.765 3.47 6.77 3.768 ;
      RECT 6.76 3.47 6.765 3.76 ;
      RECT 6.74 3.47 6.76 3.743 ;
      RECT 9.16 2.04 9.42 2.3 ;
      RECT 9.145 2.04 9.42 2.203 ;
      RECT 9.115 2.04 9.42 2.178 ;
      RECT 9.08 1.88 9.36 2.16 ;
      RECT 9.05 3.37 9.11 3.63 ;
      RECT 8.075 2.06 8.13 2.32 ;
      RECT 9.01 3.327 9.05 3.63 ;
      RECT 8.981 3.248 9.01 3.63 ;
      RECT 8.895 3.12 8.981 3.63 ;
      RECT 8.875 3 8.895 3.63 ;
      RECT 8.85 2.951 8.875 3.63 ;
      RECT 8.845 2.916 8.85 3.48 ;
      RECT 8.815 2.876 8.845 3.418 ;
      RECT 8.79 2.813 8.815 3.333 ;
      RECT 8.78 2.775 8.79 3.27 ;
      RECT 8.765 2.75 8.78 3.231 ;
      RECT 8.722 2.708 8.765 3.137 ;
      RECT 8.72 2.681 8.722 3.064 ;
      RECT 8.715 2.676 8.72 3.055 ;
      RECT 8.71 2.669 8.715 3.03 ;
      RECT 8.705 2.663 8.71 3.015 ;
      RECT 8.7 2.657 8.705 3.003 ;
      RECT 8.69 2.648 8.7 2.985 ;
      RECT 8.685 2.639 8.69 2.963 ;
      RECT 8.66 2.62 8.685 2.913 ;
      RECT 8.655 2.601 8.66 2.863 ;
      RECT 8.64 2.587 8.655 2.823 ;
      RECT 8.635 2.573 8.64 2.79 ;
      RECT 8.63 2.566 8.635 2.783 ;
      RECT 8.615 2.553 8.63 2.775 ;
      RECT 8.57 2.515 8.615 2.748 ;
      RECT 8.54 2.468 8.57 2.713 ;
      RECT 8.52 2.437 8.54 2.69 ;
      RECT 8.44 2.37 8.52 2.643 ;
      RECT 8.41 2.3 8.44 2.59 ;
      RECT 8.405 2.277 8.41 2.573 ;
      RECT 8.375 2.255 8.405 2.558 ;
      RECT 8.345 2.214 8.375 2.53 ;
      RECT 8.34 2.189 8.345 2.515 ;
      RECT 8.335 2.183 8.34 2.508 ;
      RECT 8.325 2.06 8.335 2.5 ;
      RECT 8.315 2.06 8.325 2.493 ;
      RECT 8.31 2.06 8.315 2.485 ;
      RECT 8.29 2.06 8.31 2.473 ;
      RECT 8.24 2.06 8.29 2.443 ;
      RECT 8.185 2.06 8.24 2.393 ;
      RECT 8.155 2.06 8.185 2.353 ;
      RECT 8.13 2.06 8.155 2.33 ;
      RECT 8 2.785 8.28 3.065 ;
      RECT 7.965 2.7 8.225 2.96 ;
      RECT 7.965 2.782 8.235 2.96 ;
      RECT 6.165 2.155 6.17 2.64 ;
      RECT 6.055 2.34 6.06 2.64 ;
      RECT 5.965 2.38 6.03 2.64 ;
      RECT 7.64 1.88 7.73 2.51 ;
      RECT 7.605 1.93 7.61 2.51 ;
      RECT 7.55 1.955 7.56 2.51 ;
      RECT 7.505 1.955 7.515 2.51 ;
      RECT 7.875 1.88 7.92 2.16 ;
      RECT 6.725 1.61 6.925 1.75 ;
      RECT 7.841 1.88 7.875 2.172 ;
      RECT 7.755 1.88 7.841 2.212 ;
      RECT 7.74 1.88 7.755 2.253 ;
      RECT 7.735 1.88 7.74 2.273 ;
      RECT 7.73 1.88 7.735 2.293 ;
      RECT 7.61 1.922 7.64 2.51 ;
      RECT 7.56 1.942 7.605 2.51 ;
      RECT 7.545 1.957 7.55 2.51 ;
      RECT 7.515 1.957 7.545 2.51 ;
      RECT 7.47 1.942 7.505 2.51 ;
      RECT 7.465 1.93 7.47 2.29 ;
      RECT 7.46 1.927 7.465 2.27 ;
      RECT 7.445 1.917 7.46 2.223 ;
      RECT 7.44 1.91 7.445 2.186 ;
      RECT 7.435 1.907 7.44 2.169 ;
      RECT 7.42 1.897 7.435 2.125 ;
      RECT 7.415 1.888 7.42 2.085 ;
      RECT 7.41 1.884 7.415 2.07 ;
      RECT 7.4 1.878 7.41 2.053 ;
      RECT 7.36 1.859 7.4 2.028 ;
      RECT 7.355 1.841 7.36 2.008 ;
      RECT 7.345 1.835 7.355 2.003 ;
      RECT 7.315 1.819 7.345 1.99 ;
      RECT 7.3 1.801 7.315 1.973 ;
      RECT 7.285 1.789 7.3 1.96 ;
      RECT 7.28 1.781 7.285 1.953 ;
      RECT 7.25 1.767 7.28 1.94 ;
      RECT 7.245 1.752 7.25 1.928 ;
      RECT 7.235 1.746 7.245 1.92 ;
      RECT 7.215 1.734 7.235 1.908 ;
      RECT 7.205 1.722 7.215 1.895 ;
      RECT 7.175 1.706 7.205 1.88 ;
      RECT 7.155 1.686 7.175 1.863 ;
      RECT 7.15 1.676 7.155 1.853 ;
      RECT 7.125 1.664 7.15 1.84 ;
      RECT 7.12 1.652 7.125 1.828 ;
      RECT 7.115 1.647 7.12 1.824 ;
      RECT 7.1 1.64 7.115 1.816 ;
      RECT 7.09 1.627 7.1 1.806 ;
      RECT 7.085 1.625 7.09 1.8 ;
      RECT 7.06 1.618 7.085 1.789 ;
      RECT 7.055 1.611 7.06 1.778 ;
      RECT 7.03 1.61 7.055 1.765 ;
      RECT 7.011 1.61 7.03 1.755 ;
      RECT 6.925 1.61 7.011 1.752 ;
      RECT 6.695 1.61 6.725 1.755 ;
      RECT 6.655 1.617 6.695 1.768 ;
      RECT 6.63 1.627 6.655 1.781 ;
      RECT 6.615 1.636 6.63 1.791 ;
      RECT 6.585 1.641 6.615 1.81 ;
      RECT 6.58 1.647 6.585 1.828 ;
      RECT 6.56 1.657 6.58 1.843 ;
      RECT 6.55 1.67 6.56 1.863 ;
      RECT 6.535 1.682 6.55 1.88 ;
      RECT 6.53 1.692 6.535 1.89 ;
      RECT 6.525 1.697 6.53 1.895 ;
      RECT 6.515 1.705 6.525 1.908 ;
      RECT 6.465 1.737 6.515 1.945 ;
      RECT 6.45 1.772 6.465 1.986 ;
      RECT 6.445 1.782 6.45 2.001 ;
      RECT 6.44 1.787 6.445 2.008 ;
      RECT 6.415 1.803 6.44 2.028 ;
      RECT 6.4 1.824 6.415 2.053 ;
      RECT 6.375 1.845 6.4 2.078 ;
      RECT 6.365 1.864 6.375 2.101 ;
      RECT 6.34 1.882 6.365 2.124 ;
      RECT 6.325 1.902 6.34 2.148 ;
      RECT 6.32 1.912 6.325 2.16 ;
      RECT 6.305 1.924 6.32 2.18 ;
      RECT 6.295 1.939 6.305 2.22 ;
      RECT 6.29 1.947 6.295 2.248 ;
      RECT 6.28 1.957 6.29 2.268 ;
      RECT 6.275 1.97 6.28 2.293 ;
      RECT 6.27 1.983 6.275 2.313 ;
      RECT 6.265 1.989 6.27 2.335 ;
      RECT 6.255 1.998 6.265 2.355 ;
      RECT 6.25 2.018 6.255 2.378 ;
      RECT 6.245 2.024 6.25 2.398 ;
      RECT 6.24 2.031 6.245 2.42 ;
      RECT 6.235 2.042 6.24 2.433 ;
      RECT 6.225 2.052 6.235 2.458 ;
      RECT 6.205 2.077 6.225 2.64 ;
      RECT 6.175 2.117 6.205 2.64 ;
      RECT 6.17 2.147 6.175 2.64 ;
      RECT 6.145 2.175 6.165 2.64 ;
      RECT 6.115 2.22 6.145 2.64 ;
      RECT 6.11 2.247 6.115 2.64 ;
      RECT 6.09 2.265 6.11 2.64 ;
      RECT 6.08 2.29 6.09 2.64 ;
      RECT 6.075 2.302 6.08 2.64 ;
      RECT 6.06 2.325 6.075 2.64 ;
      RECT 6.04 2.352 6.055 2.64 ;
      RECT 6.03 2.375 6.04 2.64 ;
      RECT 7.82 3.26 7.9 3.52 ;
      RECT 7.055 2.48 7.125 2.74 ;
      RECT 7.786 3.227 7.82 3.52 ;
      RECT 7.7 3.13 7.786 3.52 ;
      RECT 7.68 3.042 7.7 3.52 ;
      RECT 7.67 3.012 7.68 3.52 ;
      RECT 7.66 2.992 7.67 3.52 ;
      RECT 7.64 2.979 7.66 3.52 ;
      RECT 7.625 2.969 7.64 3.348 ;
      RECT 7.62 2.962 7.625 3.303 ;
      RECT 7.61 2.956 7.62 3.293 ;
      RECT 7.6 2.948 7.61 3.275 ;
      RECT 7.595 2.942 7.6 3.263 ;
      RECT 7.585 2.937 7.595 3.25 ;
      RECT 7.565 2.927 7.585 3.223 ;
      RECT 7.525 2.906 7.565 3.175 ;
      RECT 7.51 2.887 7.525 3.133 ;
      RECT 7.485 2.873 7.51 3.103 ;
      RECT 7.475 2.861 7.485 3.07 ;
      RECT 7.47 2.856 7.475 3.06 ;
      RECT 7.44 2.842 7.47 3.04 ;
      RECT 7.43 2.826 7.44 3.013 ;
      RECT 7.425 2.821 7.43 3.003 ;
      RECT 7.4 2.812 7.425 2.983 ;
      RECT 7.39 2.8 7.4 2.963 ;
      RECT 7.32 2.768 7.39 2.938 ;
      RECT 7.315 2.737 7.32 2.915 ;
      RECT 7.266 2.48 7.315 2.898 ;
      RECT 7.18 2.48 7.266 2.857 ;
      RECT 7.125 2.48 7.18 2.785 ;
      RECT 7.215 3.265 7.375 3.525 ;
      RECT 6.74 1.88 6.79 2.565 ;
      RECT 6.53 2.305 6.565 2.565 ;
      RECT 6.845 1.88 6.85 2.34 ;
      RECT 6.935 1.88 6.96 2.16 ;
      RECT 7.21 3.262 7.215 3.525 ;
      RECT 7.175 3.25 7.21 3.525 ;
      RECT 7.115 3.223 7.175 3.525 ;
      RECT 7.11 3.206 7.115 3.379 ;
      RECT 7.105 3.203 7.11 3.366 ;
      RECT 7.085 3.196 7.105 3.353 ;
      RECT 7.05 3.179 7.085 3.335 ;
      RECT 7.01 3.158 7.05 3.315 ;
      RECT 7.005 3.146 7.01 3.303 ;
      RECT 6.965 3.132 7.005 3.289 ;
      RECT 6.945 3.115 6.965 3.271 ;
      RECT 6.935 3.107 6.945 3.263 ;
      RECT 6.92 1.88 6.935 2.178 ;
      RECT 6.905 3.097 6.935 3.25 ;
      RECT 6.89 1.88 6.92 2.223 ;
      RECT 6.895 3.087 6.905 3.237 ;
      RECT 6.865 3.072 6.895 3.224 ;
      RECT 6.85 1.88 6.89 2.29 ;
      RECT 6.85 3.04 6.865 3.21 ;
      RECT 6.845 3.012 6.85 3.204 ;
      RECT 6.84 1.88 6.845 2.345 ;
      RECT 6.83 2.982 6.845 3.198 ;
      RECT 6.835 1.88 6.84 2.358 ;
      RECT 6.825 1.88 6.835 2.378 ;
      RECT 6.79 2.895 6.83 3.183 ;
      RECT 6.79 1.88 6.825 2.418 ;
      RECT 6.785 2.827 6.79 3.171 ;
      RECT 6.77 2.782 6.785 3.166 ;
      RECT 6.765 2.72 6.77 3.161 ;
      RECT 6.74 2.627 6.765 3.154 ;
      RECT 6.735 1.88 6.74 3.146 ;
      RECT 6.72 1.88 6.735 3.133 ;
      RECT 6.7 1.88 6.72 3.09 ;
      RECT 6.69 1.88 6.7 3.04 ;
      RECT 6.685 1.88 6.69 3.013 ;
      RECT 6.68 1.88 6.685 2.991 ;
      RECT 6.675 2.106 6.68 2.974 ;
      RECT 6.67 2.128 6.675 2.952 ;
      RECT 6.665 2.17 6.67 2.935 ;
      RECT 6.635 2.22 6.665 2.879 ;
      RECT 6.63 2.247 6.635 2.821 ;
      RECT 6.615 2.265 6.63 2.785 ;
      RECT 6.61 2.283 6.615 2.749 ;
      RECT 6.604 2.29 6.61 2.73 ;
      RECT 6.6 2.297 6.604 2.713 ;
      RECT 6.595 2.302 6.6 2.682 ;
      RECT 6.585 2.305 6.595 2.657 ;
      RECT 6.575 2.305 6.585 2.623 ;
      RECT 6.57 2.305 6.575 2.6 ;
      RECT 6.565 2.305 6.57 2.58 ;
      RECT 5.48 2.44 5.76 2.72 ;
      RECT 5.48 2.44 5.78 2.615 ;
      RECT 5.57 2.33 5.83 2.59 ;
      RECT 5.535 2.425 5.83 2.59 ;
      RECT 5.66 0.945 5.825 2.59 ;
      RECT 5.56 0.945 5.93 1.315 ;
      RECT 5.185 3.47 5.445 3.73 ;
      RECT 5.205 3.397 5.385 3.73 ;
      RECT 5.205 3.14 5.38 3.73 ;
      RECT 5.205 2.932 5.37 3.73 ;
      RECT 5.21 2.85 5.37 3.73 ;
      RECT 5.21 2.615 5.36 3.73 ;
      RECT 5.21 2.462 5.355 3.73 ;
      RECT 5.215 2.447 5.355 3.73 ;
      RECT 5.265 2.162 5.355 3.73 ;
      RECT 5.22 2.397 5.355 3.73 ;
      RECT 5.25 2.215 5.355 3.73 ;
      RECT 5.235 2.327 5.355 3.73 ;
      RECT 5.24 2.285 5.355 3.73 ;
      RECT 5.235 2.327 5.37 2.39 ;
      RECT 5.27 1.915 5.375 2.335 ;
      RECT 5.27 1.915 5.39 2.318 ;
      RECT 5.27 1.915 5.425 2.28 ;
      RECT 5.265 2.162 5.475 2.213 ;
      RECT 5.27 1.915 5.53 2.175 ;
      RECT 4.53 2.62 4.79 2.88 ;
      RECT 4.53 2.62 4.8 2.838 ;
      RECT 4.53 2.62 4.886 2.809 ;
      RECT 4.53 2.62 4.955 2.761 ;
      RECT 4.53 2.62 4.99 2.73 ;
      RECT 4.76 2.44 5.04 2.72 ;
      RECT 4.595 2.605 5.04 2.72 ;
      RECT 4.685 2.482 4.79 2.88 ;
      RECT 4.615 2.545 5.04 2.72 ;
      RECT 0.195 8.5 0.575 8.88 ;
      RECT 0.235 8.48 0.405 8.88 ;
      RECT 70.035 7.055 70.405 7.425 ;
      RECT 54.775 7.055 55.145 7.425 ;
      RECT 39.515 7.055 39.885 7.425 ;
      RECT 24.255 7.055 24.625 7.425 ;
      RECT 8.995 7.055 9.365 7.425 ;
    LAYER via1 ;
      RECT 78.625 7.375 78.775 7.525 ;
      RECT 76.255 6.74 76.405 6.89 ;
      RECT 76.24 2.065 76.39 2.215 ;
      RECT 75.45 2.45 75.6 2.6 ;
      RECT 75.45 6.325 75.6 6.475 ;
      RECT 73.86 2.805 74.01 2.955 ;
      RECT 72.09 2.35 72.24 2.5 ;
      RECT 71.07 3.055 71.22 3.205 ;
      RECT 70.84 2.475 70.99 2.625 ;
      RECT 70.805 6.71 70.955 6.86 ;
      RECT 70.495 3.075 70.645 3.225 ;
      RECT 70.255 2.095 70.405 2.245 ;
      RECT 70.145 7.165 70.295 7.315 ;
      RECT 69.945 3.425 70.095 3.575 ;
      RECT 69.805 2.03 69.955 2.18 ;
      RECT 69.17 2.115 69.32 2.265 ;
      RECT 69.06 2.755 69.21 2.905 ;
      RECT 68.735 3.315 68.885 3.465 ;
      RECT 68.565 2.305 68.715 2.455 ;
      RECT 68.21 3.32 68.36 3.47 ;
      RECT 68.15 2.535 68.3 2.685 ;
      RECT 67.785 3.525 67.935 3.675 ;
      RECT 67.625 2.36 67.775 2.51 ;
      RECT 67.06 2.435 67.21 2.585 ;
      RECT 66.71 1.055 66.86 1.205 ;
      RECT 66.665 2.385 66.815 2.535 ;
      RECT 66.365 1.97 66.515 2.12 ;
      RECT 66.28 3.525 66.43 3.675 ;
      RECT 65.625 2.675 65.775 2.825 ;
      RECT 63.34 6.755 63.49 6.905 ;
      RECT 60.995 6.74 61.145 6.89 ;
      RECT 60.98 2.065 61.13 2.215 ;
      RECT 60.19 2.45 60.34 2.6 ;
      RECT 60.19 6.325 60.34 6.475 ;
      RECT 58.6 2.805 58.75 2.955 ;
      RECT 56.83 2.35 56.98 2.5 ;
      RECT 55.81 3.055 55.96 3.205 ;
      RECT 55.58 2.475 55.73 2.625 ;
      RECT 55.545 6.71 55.695 6.86 ;
      RECT 55.235 3.075 55.385 3.225 ;
      RECT 54.995 2.095 55.145 2.245 ;
      RECT 54.885 7.165 55.035 7.315 ;
      RECT 54.685 3.425 54.835 3.575 ;
      RECT 54.545 2.03 54.695 2.18 ;
      RECT 53.91 2.115 54.06 2.265 ;
      RECT 53.8 2.755 53.95 2.905 ;
      RECT 53.475 3.315 53.625 3.465 ;
      RECT 53.305 2.305 53.455 2.455 ;
      RECT 52.95 3.32 53.1 3.47 ;
      RECT 52.89 2.535 53.04 2.685 ;
      RECT 52.525 3.525 52.675 3.675 ;
      RECT 52.365 2.36 52.515 2.51 ;
      RECT 51.8 2.435 51.95 2.585 ;
      RECT 51.45 1.055 51.6 1.205 ;
      RECT 51.405 2.385 51.555 2.535 ;
      RECT 51.105 1.97 51.255 2.12 ;
      RECT 51.02 3.525 51.17 3.675 ;
      RECT 50.365 2.675 50.515 2.825 ;
      RECT 48.08 6.755 48.23 6.905 ;
      RECT 45.735 6.74 45.885 6.89 ;
      RECT 45.72 2.065 45.87 2.215 ;
      RECT 44.93 2.45 45.08 2.6 ;
      RECT 44.93 6.325 45.08 6.475 ;
      RECT 43.34 2.805 43.49 2.955 ;
      RECT 41.57 2.35 41.72 2.5 ;
      RECT 40.55 3.055 40.7 3.205 ;
      RECT 40.32 2.475 40.47 2.625 ;
      RECT 40.285 6.715 40.435 6.865 ;
      RECT 39.975 3.075 40.125 3.225 ;
      RECT 39.735 2.095 39.885 2.245 ;
      RECT 39.625 7.165 39.775 7.315 ;
      RECT 39.425 3.425 39.575 3.575 ;
      RECT 39.285 2.03 39.435 2.18 ;
      RECT 38.65 2.115 38.8 2.265 ;
      RECT 38.54 2.755 38.69 2.905 ;
      RECT 38.215 3.315 38.365 3.465 ;
      RECT 38.045 2.305 38.195 2.455 ;
      RECT 37.69 3.32 37.84 3.47 ;
      RECT 37.63 2.535 37.78 2.685 ;
      RECT 37.265 3.525 37.415 3.675 ;
      RECT 37.105 2.36 37.255 2.51 ;
      RECT 36.54 2.435 36.69 2.585 ;
      RECT 36.19 1.055 36.34 1.205 ;
      RECT 36.145 2.385 36.295 2.535 ;
      RECT 35.845 1.97 35.995 2.12 ;
      RECT 35.76 3.525 35.91 3.675 ;
      RECT 35.105 2.675 35.255 2.825 ;
      RECT 32.865 6.76 33.015 6.91 ;
      RECT 30.475 6.74 30.625 6.89 ;
      RECT 30.46 2.065 30.61 2.215 ;
      RECT 29.67 2.45 29.82 2.6 ;
      RECT 29.67 6.325 29.82 6.475 ;
      RECT 28.08 2.805 28.23 2.955 ;
      RECT 26.31 2.35 26.46 2.5 ;
      RECT 25.29 3.055 25.44 3.205 ;
      RECT 25.06 2.475 25.21 2.625 ;
      RECT 25.025 6.71 25.175 6.86 ;
      RECT 24.715 3.075 24.865 3.225 ;
      RECT 24.475 2.095 24.625 2.245 ;
      RECT 24.365 7.165 24.515 7.315 ;
      RECT 24.165 3.425 24.315 3.575 ;
      RECT 24.025 2.03 24.175 2.18 ;
      RECT 23.39 2.115 23.54 2.265 ;
      RECT 23.28 2.755 23.43 2.905 ;
      RECT 22.955 3.315 23.105 3.465 ;
      RECT 22.785 2.305 22.935 2.455 ;
      RECT 22.43 3.32 22.58 3.47 ;
      RECT 22.37 2.535 22.52 2.685 ;
      RECT 22.005 3.525 22.155 3.675 ;
      RECT 21.845 2.36 21.995 2.51 ;
      RECT 21.28 2.435 21.43 2.585 ;
      RECT 20.93 1.055 21.08 1.205 ;
      RECT 20.885 2.385 21.035 2.535 ;
      RECT 20.585 1.97 20.735 2.12 ;
      RECT 20.5 3.525 20.65 3.675 ;
      RECT 19.845 2.675 19.995 2.825 ;
      RECT 17.605 6.755 17.755 6.905 ;
      RECT 15.215 6.74 15.365 6.89 ;
      RECT 15.2 2.065 15.35 2.215 ;
      RECT 14.41 2.45 14.56 2.6 ;
      RECT 14.41 6.325 14.56 6.475 ;
      RECT 12.82 2.805 12.97 2.955 ;
      RECT 11.05 2.35 11.2 2.5 ;
      RECT 10.03 3.055 10.18 3.205 ;
      RECT 9.8 2.475 9.95 2.625 ;
      RECT 9.765 6.705 9.915 6.855 ;
      RECT 9.455 3.075 9.605 3.225 ;
      RECT 9.215 2.095 9.365 2.245 ;
      RECT 9.105 7.165 9.255 7.315 ;
      RECT 8.905 3.425 9.055 3.575 ;
      RECT 8.765 2.03 8.915 2.18 ;
      RECT 8.13 2.115 8.28 2.265 ;
      RECT 8.02 2.755 8.17 2.905 ;
      RECT 7.695 3.315 7.845 3.465 ;
      RECT 7.525 2.305 7.675 2.455 ;
      RECT 7.17 3.32 7.32 3.47 ;
      RECT 7.11 2.535 7.26 2.685 ;
      RECT 6.745 3.525 6.895 3.675 ;
      RECT 6.585 2.36 6.735 2.51 ;
      RECT 6.02 2.435 6.17 2.585 ;
      RECT 5.67 1.055 5.82 1.205 ;
      RECT 5.625 2.385 5.775 2.535 ;
      RECT 5.325 1.97 5.475 2.12 ;
      RECT 5.24 3.525 5.39 3.675 ;
      RECT 4.585 2.675 4.735 2.825 ;
      RECT 1.61 7.095 1.76 7.245 ;
      RECT 1.235 6.355 1.385 6.505 ;
      RECT 0.31 8.615 0.46 8.765 ;
    LAYER met1 ;
      RECT 64.585 0 73.325 1.74 ;
      RECT 49.325 0 58.065 1.74 ;
      RECT 34.065 0 42.805 1.74 ;
      RECT 18.805 0 27.545 1.74 ;
      RECT 3.545 0 12.285 1.74 ;
      RECT 78.915 0 79.095 0.305 ;
      RECT 63.655 0 76.965 0.305 ;
      RECT 48.395 0 61.705 0.305 ;
      RECT 33.135 0 46.445 0.305 ;
      RECT 17.875 0 31.185 0.305 ;
      RECT 0 0 15.925 0.305 ;
      RECT 0 0 79.095 0.3 ;
      RECT 0 8.58 79.095 8.88 ;
      RECT 78.915 8.575 79.095 8.88 ;
      RECT 63.655 8.575 76.965 8.88 ;
      RECT 48.395 8.575 61.705 8.88 ;
      RECT 33.135 8.575 46.445 8.88 ;
      RECT 17.875 8.575 31.185 8.88 ;
      RECT 0 8.575 15.925 8.88 ;
      RECT 69.53 6.315 69.7 8.88 ;
      RECT 54.27 6.315 54.44 8.88 ;
      RECT 39.01 6.315 39.18 8.88 ;
      RECT 23.75 6.315 23.92 8.88 ;
      RECT 8.49 6.315 8.66 8.88 ;
      RECT 0.005 8.565 0.81 8.88 ;
      RECT 0.21 8.545 0.56 8.88 ;
      RECT 69.7 6.285 69.99 6.515 ;
      RECT 54.44 6.285 54.73 6.515 ;
      RECT 39.18 6.285 39.47 6.515 ;
      RECT 23.92 6.285 24.21 6.515 ;
      RECT 8.66 6.285 8.95 6.515 ;
      RECT 78.49 7.77 78.78 8 ;
      RECT 78.55 6.29 78.72 8 ;
      RECT 78.525 7.275 78.875 7.625 ;
      RECT 78.49 6.29 78.78 6.52 ;
      RECT 78.085 2.395 78.19 2.965 ;
      RECT 78.085 2.73 78.41 2.96 ;
      RECT 78.085 2.76 78.58 2.93 ;
      RECT 78.085 2.395 78.275 2.96 ;
      RECT 77.5 2.36 77.79 2.59 ;
      RECT 77.5 2.395 78.275 2.565 ;
      RECT 77.56 0.88 77.73 2.59 ;
      RECT 77.5 0.88 77.79 1.11 ;
      RECT 77.5 7.77 77.79 8 ;
      RECT 77.56 6.29 77.73 8 ;
      RECT 77.5 6.29 77.79 6.52 ;
      RECT 77.5 6.325 78.355 6.485 ;
      RECT 78.185 5.92 78.355 6.485 ;
      RECT 77.5 6.32 77.895 6.485 ;
      RECT 78.12 5.92 78.41 6.15 ;
      RECT 78.12 5.95 78.58 6.12 ;
      RECT 77.13 2.73 77.42 2.96 ;
      RECT 77.13 2.76 77.59 2.93 ;
      RECT 77.195 1.655 77.36 2.96 ;
      RECT 75.71 1.625 76 1.855 ;
      RECT 75.71 1.655 77.36 1.825 ;
      RECT 75.77 0.885 75.94 1.855 ;
      RECT 75.71 0.885 76 1.115 ;
      RECT 75.71 7.765 76 7.995 ;
      RECT 75.77 7.025 75.94 7.995 ;
      RECT 75.77 7.12 77.36 7.29 ;
      RECT 77.19 5.92 77.36 7.29 ;
      RECT 75.71 7.025 76 7.255 ;
      RECT 77.13 5.92 77.42 6.15 ;
      RECT 77.13 5.95 77.59 6.12 ;
      RECT 73.76 2.705 74.1 3.055 ;
      RECT 73.85 2.025 74.02 3.055 ;
      RECT 76.14 1.965 76.49 2.315 ;
      RECT 73.85 2.025 76.49 2.195 ;
      RECT 76.165 6.655 76.49 6.98 ;
      RECT 70.705 6.61 71.055 6.96 ;
      RECT 76.14 6.655 76.49 6.885 ;
      RECT 70.505 6.655 71.055 6.885 ;
      RECT 70.335 6.685 76.49 6.855 ;
      RECT 75.365 2.365 75.685 2.685 ;
      RECT 75.335 2.365 75.685 2.595 ;
      RECT 75.165 2.395 75.685 2.565 ;
      RECT 75.365 6.255 75.685 6.545 ;
      RECT 75.335 6.285 75.685 6.515 ;
      RECT 75.165 6.315 75.685 6.485 ;
      RECT 71.055 2.985 71.205 3.26 ;
      RECT 71.595 2.065 71.6 2.285 ;
      RECT 72.745 2.265 72.76 2.463 ;
      RECT 72.71 2.257 72.745 2.47 ;
      RECT 72.68 2.25 72.71 2.47 ;
      RECT 72.625 2.215 72.68 2.47 ;
      RECT 72.56 2.152 72.625 2.47 ;
      RECT 72.555 2.117 72.56 2.468 ;
      RECT 72.55 2.112 72.555 2.46 ;
      RECT 72.545 2.107 72.55 2.446 ;
      RECT 72.54 2.104 72.545 2.439 ;
      RECT 72.495 2.094 72.54 2.39 ;
      RECT 72.475 2.081 72.495 2.325 ;
      RECT 72.47 2.076 72.475 2.298 ;
      RECT 72.465 2.075 72.47 2.291 ;
      RECT 72.46 2.074 72.465 2.284 ;
      RECT 72.375 2.059 72.46 2.23 ;
      RECT 72.345 2.04 72.375 2.18 ;
      RECT 72.265 2.023 72.345 2.165 ;
      RECT 72.23 2.01 72.265 2.15 ;
      RECT 72.222 2.01 72.23 2.145 ;
      RECT 72.136 2.011 72.222 2.145 ;
      RECT 72.05 2.013 72.136 2.145 ;
      RECT 72.025 2.014 72.05 2.149 ;
      RECT 71.95 2.02 72.025 2.164 ;
      RECT 71.867 2.032 71.95 2.188 ;
      RECT 71.781 2.045 71.867 2.214 ;
      RECT 71.695 2.058 71.781 2.24 ;
      RECT 71.66 2.067 71.695 2.259 ;
      RECT 71.61 2.067 71.66 2.272 ;
      RECT 71.6 2.065 71.61 2.283 ;
      RECT 71.585 2.062 71.595 2.285 ;
      RECT 71.57 2.054 71.585 2.293 ;
      RECT 71.555 2.046 71.57 2.313 ;
      RECT 71.55 2.041 71.555 2.37 ;
      RECT 71.535 2.036 71.55 2.443 ;
      RECT 71.53 2.031 71.535 2.485 ;
      RECT 71.525 2.029 71.53 2.513 ;
      RECT 71.52 2.027 71.525 2.535 ;
      RECT 71.51 2.023 71.52 2.578 ;
      RECT 71.505 2.02 71.51 2.603 ;
      RECT 71.5 2.018 71.505 2.623 ;
      RECT 71.495 2.016 71.5 2.647 ;
      RECT 71.49 2.012 71.495 2.67 ;
      RECT 71.485 2.008 71.49 2.693 ;
      RECT 71.45 1.998 71.485 2.8 ;
      RECT 71.445 1.988 71.45 2.898 ;
      RECT 71.44 1.986 71.445 2.925 ;
      RECT 71.435 1.985 71.44 2.945 ;
      RECT 71.43 1.977 71.435 2.965 ;
      RECT 71.425 1.972 71.43 3 ;
      RECT 71.42 1.97 71.425 3.018 ;
      RECT 71.415 1.97 71.42 3.043 ;
      RECT 71.41 1.97 71.415 3.065 ;
      RECT 71.375 1.97 71.41 3.108 ;
      RECT 71.35 1.97 71.375 3.137 ;
      RECT 71.34 1.97 71.35 2.323 ;
      RECT 71.343 2.38 71.35 3.147 ;
      RECT 71.34 2.437 71.343 3.15 ;
      RECT 71.335 1.97 71.34 2.295 ;
      RECT 71.335 2.487 71.34 3.153 ;
      RECT 71.325 1.97 71.335 2.285 ;
      RECT 71.33 2.54 71.335 3.156 ;
      RECT 71.325 2.625 71.33 3.16 ;
      RECT 71.315 1.97 71.325 2.273 ;
      RECT 71.32 2.672 71.325 3.164 ;
      RECT 71.315 2.747 71.32 3.168 ;
      RECT 71.28 1.97 71.315 2.248 ;
      RECT 71.305 2.83 71.315 3.173 ;
      RECT 71.295 2.897 71.305 3.18 ;
      RECT 71.29 2.925 71.295 3.185 ;
      RECT 71.28 2.938 71.29 3.191 ;
      RECT 71.235 1.97 71.28 2.205 ;
      RECT 71.275 2.943 71.28 3.198 ;
      RECT 71.235 2.96 71.275 3.26 ;
      RECT 71.23 1.972 71.235 2.178 ;
      RECT 71.205 2.98 71.235 3.26 ;
      RECT 71.225 1.977 71.23 2.15 ;
      RECT 71.015 2.989 71.055 3.26 ;
      RECT 70.99 2.997 71.015 3.23 ;
      RECT 70.945 3.005 70.99 3.23 ;
      RECT 70.93 3.01 70.945 3.225 ;
      RECT 70.92 3.01 70.93 3.219 ;
      RECT 70.91 3.017 70.92 3.216 ;
      RECT 70.905 3.055 70.91 3.205 ;
      RECT 70.9 3.117 70.905 3.183 ;
      RECT 72.17 2.992 72.355 3.215 ;
      RECT 72.17 3.007 72.36 3.211 ;
      RECT 72.16 2.28 72.245 3.21 ;
      RECT 72.16 3.007 72.365 3.204 ;
      RECT 72.155 3.015 72.365 3.203 ;
      RECT 72.36 2.735 72.68 3.055 ;
      RECT 72.155 2.907 72.325 2.998 ;
      RECT 72.15 2.907 72.325 2.98 ;
      RECT 72.14 2.715 72.275 2.955 ;
      RECT 72.135 2.715 72.275 2.9 ;
      RECT 72.095 2.295 72.265 2.8 ;
      RECT 72.08 2.295 72.265 2.67 ;
      RECT 72.075 2.295 72.265 2.623 ;
      RECT 72.07 2.295 72.265 2.603 ;
      RECT 72.065 2.295 72.265 2.578 ;
      RECT 72.035 2.295 72.295 2.555 ;
      RECT 72.045 2.292 72.255 2.555 ;
      RECT 72.17 2.287 72.255 3.215 ;
      RECT 72.055 2.28 72.245 2.555 ;
      RECT 72.05 2.285 72.245 2.555 ;
      RECT 70.88 2.497 71.065 2.71 ;
      RECT 70.88 2.505 71.075 2.703 ;
      RECT 70.86 2.505 71.075 2.7 ;
      RECT 70.855 2.505 71.075 2.685 ;
      RECT 70.785 2.42 71.045 2.68 ;
      RECT 70.785 2.565 71.08 2.593 ;
      RECT 70.44 3.02 70.7 3.28 ;
      RECT 70.465 2.965 70.66 3.28 ;
      RECT 70.46 2.714 70.64 3.008 ;
      RECT 70.46 2.72 70.65 3.008 ;
      RECT 70.44 2.722 70.65 2.953 ;
      RECT 70.435 2.732 70.65 2.82 ;
      RECT 70.465 2.712 70.64 3.28 ;
      RECT 70.551 2.71 70.64 3.28 ;
      RECT 70.41 1.93 70.445 2.3 ;
      RECT 70.2 2.04 70.205 2.3 ;
      RECT 70.445 1.937 70.46 2.3 ;
      RECT 70.335 1.93 70.41 2.378 ;
      RECT 70.325 1.93 70.335 2.463 ;
      RECT 70.3 1.93 70.325 2.498 ;
      RECT 70.26 1.93 70.3 2.566 ;
      RECT 70.25 1.937 70.26 2.618 ;
      RECT 70.22 2.04 70.25 2.659 ;
      RECT 70.215 2.04 70.22 2.698 ;
      RECT 70.205 2.04 70.215 2.718 ;
      RECT 70.2 2.335 70.205 2.755 ;
      RECT 70.195 2.352 70.2 2.775 ;
      RECT 70.18 2.415 70.195 2.815 ;
      RECT 70.175 2.458 70.18 2.85 ;
      RECT 70.17 2.466 70.175 2.863 ;
      RECT 70.16 2.48 70.17 2.885 ;
      RECT 70.135 2.515 70.16 2.95 ;
      RECT 70.125 2.55 70.135 3.013 ;
      RECT 70.105 2.58 70.125 3.074 ;
      RECT 70.09 2.616 70.105 3.141 ;
      RECT 70.08 2.644 70.09 3.18 ;
      RECT 70.07 2.666 70.08 3.2 ;
      RECT 70.065 2.676 70.07 3.211 ;
      RECT 70.06 2.685 70.065 3.214 ;
      RECT 70.05 2.703 70.06 3.218 ;
      RECT 70.04 2.721 70.05 3.219 ;
      RECT 70.015 2.76 70.04 3.216 ;
      RECT 69.995 2.802 70.015 3.213 ;
      RECT 69.98 2.84 69.995 3.212 ;
      RECT 69.945 2.875 69.98 3.209 ;
      RECT 69.94 2.897 69.945 3.207 ;
      RECT 69.875 2.937 69.94 3.204 ;
      RECT 69.87 2.977 69.875 3.2 ;
      RECT 69.855 2.987 69.87 3.191 ;
      RECT 69.845 3.107 69.855 3.176 ;
      RECT 70.325 3.52 70.335 3.78 ;
      RECT 70.325 3.523 70.345 3.779 ;
      RECT 70.315 3.513 70.325 3.778 ;
      RECT 70.305 3.528 70.385 3.774 ;
      RECT 70.29 3.507 70.305 3.772 ;
      RECT 70.265 3.532 70.39 3.768 ;
      RECT 70.25 3.492 70.265 3.763 ;
      RECT 70.25 3.534 70.4 3.762 ;
      RECT 70.25 3.542 70.415 3.755 ;
      RECT 70.19 3.479 70.25 3.745 ;
      RECT 70.18 3.466 70.19 3.727 ;
      RECT 70.155 3.456 70.18 3.717 ;
      RECT 70.15 3.446 70.155 3.709 ;
      RECT 70.085 3.542 70.415 3.691 ;
      RECT 70 3.542 70.415 3.653 ;
      RECT 69.89 3.37 70.15 3.63 ;
      RECT 70.265 3.5 70.29 3.768 ;
      RECT 70.305 3.51 70.315 3.774 ;
      RECT 69.89 3.518 70.33 3.63 ;
      RECT 70.075 7.765 70.365 7.995 ;
      RECT 70.135 7.025 70.305 7.995 ;
      RECT 70.035 7.055 70.405 7.425 ;
      RECT 70.075 7.025 70.365 7.425 ;
      RECT 69.105 3.275 69.135 3.575 ;
      RECT 68.88 3.26 68.885 3.535 ;
      RECT 68.68 3.26 68.835 3.52 ;
      RECT 69.98 1.975 70.01 2.235 ;
      RECT 69.97 1.975 69.98 2.343 ;
      RECT 69.95 1.975 69.97 2.353 ;
      RECT 69.935 1.975 69.95 2.365 ;
      RECT 69.88 1.975 69.935 2.415 ;
      RECT 69.865 1.975 69.88 2.463 ;
      RECT 69.835 1.975 69.865 2.498 ;
      RECT 69.78 1.975 69.835 2.56 ;
      RECT 69.76 1.975 69.78 2.628 ;
      RECT 69.755 1.975 69.76 2.658 ;
      RECT 69.75 1.975 69.755 2.67 ;
      RECT 69.745 2.092 69.75 2.688 ;
      RECT 69.725 2.11 69.745 2.713 ;
      RECT 69.705 2.137 69.725 2.763 ;
      RECT 69.7 2.157 69.705 2.794 ;
      RECT 69.695 2.165 69.7 2.811 ;
      RECT 69.68 2.191 69.695 2.84 ;
      RECT 69.665 2.233 69.68 2.875 ;
      RECT 69.66 2.262 69.665 2.898 ;
      RECT 69.655 2.277 69.66 2.911 ;
      RECT 69.65 2.3 69.655 2.922 ;
      RECT 69.64 2.32 69.65 2.94 ;
      RECT 69.63 2.35 69.64 2.963 ;
      RECT 69.625 2.372 69.63 2.983 ;
      RECT 69.62 2.387 69.625 2.998 ;
      RECT 69.605 2.417 69.62 3.025 ;
      RECT 69.6 2.447 69.605 3.051 ;
      RECT 69.595 2.465 69.6 3.063 ;
      RECT 69.585 2.495 69.595 3.082 ;
      RECT 69.575 2.52 69.585 3.107 ;
      RECT 69.57 2.54 69.575 3.126 ;
      RECT 69.565 2.557 69.57 3.139 ;
      RECT 69.555 2.583 69.565 3.158 ;
      RECT 69.545 2.621 69.555 3.185 ;
      RECT 69.54 2.647 69.545 3.205 ;
      RECT 69.535 2.657 69.54 3.215 ;
      RECT 69.53 2.67 69.535 3.23 ;
      RECT 69.525 2.685 69.53 3.24 ;
      RECT 69.52 2.707 69.525 3.255 ;
      RECT 69.515 2.725 69.52 3.266 ;
      RECT 69.51 2.735 69.515 3.277 ;
      RECT 69.505 2.743 69.51 3.289 ;
      RECT 69.5 2.751 69.505 3.3 ;
      RECT 69.495 2.777 69.5 3.313 ;
      RECT 69.485 2.805 69.495 3.326 ;
      RECT 69.48 2.835 69.485 3.335 ;
      RECT 69.475 2.85 69.48 3.342 ;
      RECT 69.46 2.875 69.475 3.349 ;
      RECT 69.455 2.897 69.46 3.355 ;
      RECT 69.45 2.922 69.455 3.358 ;
      RECT 69.441 2.95 69.45 3.362 ;
      RECT 69.435 2.967 69.441 3.367 ;
      RECT 69.43 2.985 69.435 3.371 ;
      RECT 69.425 2.997 69.43 3.374 ;
      RECT 69.42 3.018 69.425 3.378 ;
      RECT 69.415 3.036 69.42 3.381 ;
      RECT 69.41 3.05 69.415 3.384 ;
      RECT 69.405 3.067 69.41 3.387 ;
      RECT 69.4 3.08 69.405 3.39 ;
      RECT 69.375 3.117 69.4 3.398 ;
      RECT 69.37 3.162 69.375 3.407 ;
      RECT 69.365 3.19 69.37 3.41 ;
      RECT 69.355 3.21 69.365 3.414 ;
      RECT 69.35 3.23 69.355 3.419 ;
      RECT 69.345 3.245 69.35 3.422 ;
      RECT 69.325 3.255 69.345 3.429 ;
      RECT 69.26 3.262 69.325 3.455 ;
      RECT 69.225 3.265 69.26 3.483 ;
      RECT 69.21 3.268 69.225 3.498 ;
      RECT 69.2 3.269 69.21 3.513 ;
      RECT 69.19 3.27 69.2 3.53 ;
      RECT 69.185 3.27 69.19 3.545 ;
      RECT 69.18 3.27 69.185 3.553 ;
      RECT 69.165 3.271 69.18 3.568 ;
      RECT 69.135 3.273 69.165 3.575 ;
      RECT 69.025 3.28 69.105 3.575 ;
      RECT 68.98 3.285 69.025 3.575 ;
      RECT 68.97 3.286 68.98 3.565 ;
      RECT 68.96 3.287 68.97 3.558 ;
      RECT 68.94 3.289 68.96 3.553 ;
      RECT 68.93 3.26 68.94 3.548 ;
      RECT 68.885 3.26 68.93 3.54 ;
      RECT 68.855 3.26 68.88 3.53 ;
      RECT 68.835 3.26 68.855 3.523 ;
      RECT 69.115 2.06 69.375 2.32 ;
      RECT 68.995 2.075 69.005 2.24 ;
      RECT 68.98 2.075 68.985 2.235 ;
      RECT 66.345 1.915 66.53 2.205 ;
      RECT 68.16 2.04 68.175 2.195 ;
      RECT 66.31 1.915 66.335 2.175 ;
      RECT 68.725 1.965 68.73 2.107 ;
      RECT 68.64 1.96 68.665 2.1 ;
      RECT 69.04 2.077 69.115 2.27 ;
      RECT 69.025 2.075 69.04 2.253 ;
      RECT 69.005 2.075 69.025 2.245 ;
      RECT 68.985 2.075 68.995 2.238 ;
      RECT 68.94 2.07 68.98 2.228 ;
      RECT 68.9 2.045 68.94 2.213 ;
      RECT 68.885 2.02 68.9 2.203 ;
      RECT 68.88 2.014 68.885 2.201 ;
      RECT 68.845 2.006 68.88 2.184 ;
      RECT 68.84 1.999 68.845 2.172 ;
      RECT 68.82 1.994 68.84 2.16 ;
      RECT 68.81 1.988 68.82 2.145 ;
      RECT 68.79 1.983 68.81 2.13 ;
      RECT 68.78 1.978 68.79 2.123 ;
      RECT 68.775 1.976 68.78 2.118 ;
      RECT 68.77 1.975 68.775 2.115 ;
      RECT 68.73 1.97 68.77 2.111 ;
      RECT 68.71 1.964 68.725 2.106 ;
      RECT 68.675 1.961 68.71 2.103 ;
      RECT 68.665 1.96 68.675 2.101 ;
      RECT 68.605 1.96 68.64 2.098 ;
      RECT 68.56 1.96 68.605 2.098 ;
      RECT 68.51 1.96 68.56 2.101 ;
      RECT 68.495 1.962 68.51 2.103 ;
      RECT 68.48 1.965 68.495 2.104 ;
      RECT 68.47 1.97 68.48 2.105 ;
      RECT 68.44 1.975 68.47 2.11 ;
      RECT 68.43 1.981 68.44 2.118 ;
      RECT 68.42 1.983 68.43 2.122 ;
      RECT 68.41 1.987 68.42 2.126 ;
      RECT 68.385 1.993 68.41 2.134 ;
      RECT 68.375 1.998 68.385 2.142 ;
      RECT 68.36 2.002 68.375 2.146 ;
      RECT 68.325 2.008 68.36 2.154 ;
      RECT 68.305 2.013 68.325 2.164 ;
      RECT 68.275 2.02 68.305 2.173 ;
      RECT 68.23 2.029 68.275 2.187 ;
      RECT 68.225 2.034 68.23 2.198 ;
      RECT 68.205 2.037 68.225 2.199 ;
      RECT 68.175 2.04 68.205 2.197 ;
      RECT 68.14 2.04 68.16 2.193 ;
      RECT 68.07 2.04 68.14 2.184 ;
      RECT 68.055 2.037 68.07 2.176 ;
      RECT 68.015 2.03 68.055 2.171 ;
      RECT 67.99 2.02 68.015 2.164 ;
      RECT 67.985 2.014 67.99 2.161 ;
      RECT 67.945 2.008 67.985 2.158 ;
      RECT 67.93 2.001 67.945 2.153 ;
      RECT 67.91 1.997 67.93 2.148 ;
      RECT 67.895 1.992 67.91 2.144 ;
      RECT 67.88 1.987 67.895 2.142 ;
      RECT 67.865 1.983 67.88 2.141 ;
      RECT 67.85 1.981 67.865 2.137 ;
      RECT 67.84 1.979 67.85 2.132 ;
      RECT 67.825 1.976 67.84 2.128 ;
      RECT 67.815 1.974 67.825 2.123 ;
      RECT 67.795 1.971 67.815 2.119 ;
      RECT 67.75 1.97 67.795 2.117 ;
      RECT 67.69 1.972 67.75 2.118 ;
      RECT 67.67 1.974 67.69 2.12 ;
      RECT 67.64 1.977 67.67 2.121 ;
      RECT 67.59 1.982 67.64 2.123 ;
      RECT 67.585 1.985 67.59 2.125 ;
      RECT 67.575 1.987 67.585 2.128 ;
      RECT 67.57 1.989 67.575 2.131 ;
      RECT 67.52 1.992 67.57 2.138 ;
      RECT 67.5 1.996 67.52 2.15 ;
      RECT 67.49 1.999 67.5 2.156 ;
      RECT 67.48 2 67.49 2.159 ;
      RECT 67.441 2.003 67.48 2.161 ;
      RECT 67.355 2.01 67.441 2.164 ;
      RECT 67.281 2.02 67.355 2.168 ;
      RECT 67.195 2.031 67.281 2.173 ;
      RECT 67.18 2.038 67.195 2.175 ;
      RECT 67.125 2.042 67.18 2.176 ;
      RECT 67.111 2.045 67.125 2.178 ;
      RECT 67.025 2.045 67.111 2.18 ;
      RECT 66.985 2.042 67.025 2.183 ;
      RECT 66.961 2.038 66.985 2.185 ;
      RECT 66.875 2.028 66.961 2.188 ;
      RECT 66.845 2.017 66.875 2.189 ;
      RECT 66.826 2.013 66.845 2.188 ;
      RECT 66.74 2.006 66.826 2.185 ;
      RECT 66.68 1.995 66.74 2.182 ;
      RECT 66.66 1.987 66.68 2.18 ;
      RECT 66.625 1.982 66.66 2.179 ;
      RECT 66.6 1.977 66.625 2.178 ;
      RECT 66.57 1.972 66.6 2.177 ;
      RECT 66.545 1.915 66.57 2.176 ;
      RECT 66.53 1.915 66.545 2.2 ;
      RECT 66.335 1.915 66.345 2.2 ;
      RECT 68.11 2.935 68.115 3.075 ;
      RECT 67.77 2.935 67.805 3.073 ;
      RECT 67.345 2.92 67.36 3.065 ;
      RECT 69.175 2.7 69.265 2.96 ;
      RECT 69.005 2.565 69.105 2.96 ;
      RECT 66.04 2.54 66.12 2.75 ;
      RECT 69.13 2.677 69.175 2.96 ;
      RECT 69.12 2.647 69.13 2.96 ;
      RECT 69.105 2.57 69.12 2.96 ;
      RECT 68.92 2.565 69.005 2.925 ;
      RECT 68.915 2.567 68.92 2.92 ;
      RECT 68.91 2.572 68.915 2.92 ;
      RECT 68.875 2.672 68.91 2.92 ;
      RECT 68.865 2.7 68.875 2.92 ;
      RECT 68.855 2.715 68.865 2.92 ;
      RECT 68.845 2.727 68.855 2.92 ;
      RECT 68.84 2.737 68.845 2.92 ;
      RECT 68.825 2.747 68.84 2.922 ;
      RECT 68.82 2.762 68.825 2.924 ;
      RECT 68.805 2.775 68.82 2.926 ;
      RECT 68.8 2.79 68.805 2.929 ;
      RECT 68.78 2.8 68.8 2.933 ;
      RECT 68.765 2.81 68.78 2.936 ;
      RECT 68.73 2.817 68.765 2.941 ;
      RECT 68.686 2.824 68.73 2.949 ;
      RECT 68.6 2.836 68.686 2.962 ;
      RECT 68.575 2.847 68.6 2.973 ;
      RECT 68.545 2.852 68.575 2.978 ;
      RECT 68.51 2.857 68.545 2.986 ;
      RECT 68.48 2.862 68.51 2.993 ;
      RECT 68.455 2.867 68.48 2.998 ;
      RECT 68.39 2.874 68.455 3.007 ;
      RECT 68.32 2.887 68.39 3.023 ;
      RECT 68.29 2.897 68.32 3.035 ;
      RECT 68.265 2.902 68.29 3.042 ;
      RECT 68.21 2.909 68.265 3.05 ;
      RECT 68.205 2.916 68.21 3.055 ;
      RECT 68.2 2.918 68.205 3.056 ;
      RECT 68.185 2.92 68.2 3.058 ;
      RECT 68.18 2.92 68.185 3.061 ;
      RECT 68.115 2.927 68.18 3.068 ;
      RECT 68.08 2.937 68.11 3.078 ;
      RECT 68.063 2.94 68.08 3.08 ;
      RECT 67.977 2.939 68.063 3.079 ;
      RECT 67.891 2.937 67.977 3.076 ;
      RECT 67.805 2.936 67.891 3.074 ;
      RECT 67.704 2.934 67.77 3.073 ;
      RECT 67.618 2.931 67.704 3.071 ;
      RECT 67.532 2.927 67.618 3.069 ;
      RECT 67.446 2.924 67.532 3.068 ;
      RECT 67.36 2.921 67.446 3.066 ;
      RECT 67.26 2.92 67.345 3.063 ;
      RECT 67.21 2.918 67.26 3.061 ;
      RECT 67.19 2.915 67.21 3.059 ;
      RECT 67.17 2.913 67.19 3.056 ;
      RECT 67.145 2.909 67.17 3.053 ;
      RECT 67.1 2.903 67.145 3.048 ;
      RECT 67.06 2.897 67.1 3.04 ;
      RECT 67.035 2.892 67.06 3.033 ;
      RECT 66.98 2.885 67.035 3.025 ;
      RECT 66.956 2.878 66.98 3.018 ;
      RECT 66.87 2.869 66.956 3.008 ;
      RECT 66.84 2.861 66.87 2.998 ;
      RECT 66.81 2.857 66.84 2.993 ;
      RECT 66.805 2.854 66.81 2.99 ;
      RECT 66.8 2.853 66.805 2.99 ;
      RECT 66.725 2.846 66.8 2.983 ;
      RECT 66.686 2.837 66.725 2.972 ;
      RECT 66.6 2.827 66.686 2.96 ;
      RECT 66.56 2.817 66.6 2.948 ;
      RECT 66.521 2.812 66.56 2.941 ;
      RECT 66.435 2.802 66.521 2.93 ;
      RECT 66.395 2.79 66.435 2.919 ;
      RECT 66.36 2.775 66.395 2.912 ;
      RECT 66.35 2.765 66.36 2.909 ;
      RECT 66.33 2.75 66.35 2.907 ;
      RECT 66.3 2.72 66.33 2.903 ;
      RECT 66.29 2.7 66.3 2.898 ;
      RECT 66.285 2.692 66.29 2.895 ;
      RECT 66.28 2.685 66.285 2.893 ;
      RECT 66.265 2.672 66.28 2.886 ;
      RECT 66.26 2.662 66.265 2.878 ;
      RECT 66.255 2.655 66.26 2.873 ;
      RECT 66.25 2.65 66.255 2.869 ;
      RECT 66.235 2.637 66.25 2.861 ;
      RECT 66.23 2.547 66.235 2.85 ;
      RECT 66.225 2.542 66.23 2.843 ;
      RECT 66.15 2.54 66.225 2.803 ;
      RECT 66.12 2.54 66.15 2.758 ;
      RECT 66.025 2.545 66.04 2.745 ;
      RECT 68.51 2.25 68.77 2.51 ;
      RECT 68.495 2.238 68.675 2.475 ;
      RECT 68.49 2.239 68.675 2.473 ;
      RECT 68.475 2.243 68.685 2.463 ;
      RECT 68.47 2.248 68.69 2.433 ;
      RECT 68.475 2.245 68.69 2.463 ;
      RECT 68.49 2.24 68.685 2.473 ;
      RECT 68.51 2.237 68.675 2.51 ;
      RECT 68.51 2.236 68.665 2.51 ;
      RECT 68.535 2.235 68.665 2.51 ;
      RECT 68.095 2.48 68.355 2.74 ;
      RECT 67.97 2.525 68.355 2.735 ;
      RECT 67.96 2.53 68.355 2.73 ;
      RECT 67.975 3.47 67.99 3.78 ;
      RECT 66.57 3.24 66.58 3.37 ;
      RECT 66.35 3.235 66.455 3.37 ;
      RECT 66.265 3.24 66.315 3.37 ;
      RECT 64.815 1.975 64.82 3.08 ;
      RECT 68.07 3.562 68.075 3.698 ;
      RECT 68.065 3.557 68.07 3.758 ;
      RECT 68.06 3.555 68.065 3.771 ;
      RECT 68.045 3.552 68.06 3.773 ;
      RECT 68.04 3.547 68.045 3.775 ;
      RECT 68.035 3.543 68.04 3.778 ;
      RECT 68.02 3.538 68.035 3.78 ;
      RECT 67.99 3.53 68.02 3.78 ;
      RECT 67.951 3.47 67.975 3.78 ;
      RECT 67.865 3.47 67.951 3.777 ;
      RECT 67.835 3.47 67.865 3.77 ;
      RECT 67.81 3.47 67.835 3.763 ;
      RECT 67.785 3.47 67.81 3.755 ;
      RECT 67.77 3.47 67.785 3.748 ;
      RECT 67.745 3.47 67.77 3.74 ;
      RECT 67.73 3.47 67.745 3.733 ;
      RECT 67.69 3.48 67.73 3.722 ;
      RECT 67.68 3.475 67.69 3.712 ;
      RECT 67.676 3.474 67.68 3.709 ;
      RECT 67.59 3.466 67.676 3.692 ;
      RECT 67.557 3.455 67.59 3.669 ;
      RECT 67.471 3.444 67.557 3.647 ;
      RECT 67.385 3.428 67.471 3.616 ;
      RECT 67.315 3.413 67.385 3.588 ;
      RECT 67.305 3.406 67.315 3.575 ;
      RECT 67.275 3.403 67.305 3.565 ;
      RECT 67.25 3.399 67.275 3.558 ;
      RECT 67.235 3.396 67.25 3.553 ;
      RECT 67.23 3.395 67.235 3.548 ;
      RECT 67.2 3.39 67.23 3.541 ;
      RECT 67.195 3.385 67.2 3.536 ;
      RECT 67.18 3.382 67.195 3.531 ;
      RECT 67.175 3.377 67.18 3.526 ;
      RECT 67.155 3.372 67.175 3.523 ;
      RECT 67.14 3.367 67.155 3.515 ;
      RECT 67.125 3.361 67.14 3.51 ;
      RECT 67.095 3.352 67.125 3.503 ;
      RECT 67.09 3.345 67.095 3.495 ;
      RECT 67.085 3.343 67.09 3.493 ;
      RECT 67.08 3.342 67.085 3.49 ;
      RECT 67.04 3.335 67.08 3.483 ;
      RECT 67.026 3.325 67.04 3.473 ;
      RECT 66.975 3.314 67.026 3.461 ;
      RECT 66.95 3.3 66.975 3.447 ;
      RECT 66.925 3.289 66.95 3.439 ;
      RECT 66.905 3.278 66.925 3.433 ;
      RECT 66.895 3.272 66.905 3.428 ;
      RECT 66.89 3.27 66.895 3.424 ;
      RECT 66.87 3.265 66.89 3.419 ;
      RECT 66.84 3.255 66.87 3.409 ;
      RECT 66.835 3.247 66.84 3.402 ;
      RECT 66.82 3.245 66.835 3.398 ;
      RECT 66.8 3.245 66.82 3.393 ;
      RECT 66.795 3.244 66.8 3.391 ;
      RECT 66.79 3.244 66.795 3.388 ;
      RECT 66.75 3.243 66.79 3.383 ;
      RECT 66.725 3.242 66.75 3.378 ;
      RECT 66.665 3.241 66.725 3.375 ;
      RECT 66.58 3.24 66.665 3.373 ;
      RECT 66.541 3.239 66.57 3.37 ;
      RECT 66.455 3.237 66.541 3.37 ;
      RECT 66.315 3.237 66.35 3.37 ;
      RECT 66.225 3.241 66.265 3.373 ;
      RECT 66.21 3.244 66.225 3.38 ;
      RECT 66.2 3.245 66.21 3.387 ;
      RECT 66.175 3.248 66.2 3.392 ;
      RECT 66.17 3.25 66.175 3.395 ;
      RECT 66.12 3.252 66.17 3.396 ;
      RECT 66.081 3.256 66.12 3.398 ;
      RECT 65.995 3.258 66.081 3.401 ;
      RECT 65.977 3.26 65.995 3.403 ;
      RECT 65.891 3.263 65.977 3.405 ;
      RECT 65.805 3.267 65.891 3.408 ;
      RECT 65.768 3.271 65.805 3.411 ;
      RECT 65.682 3.274 65.768 3.414 ;
      RECT 65.596 3.278 65.682 3.417 ;
      RECT 65.51 3.283 65.596 3.421 ;
      RECT 65.49 3.285 65.51 3.424 ;
      RECT 65.47 3.284 65.49 3.425 ;
      RECT 65.421 3.281 65.47 3.426 ;
      RECT 65.335 3.276 65.421 3.429 ;
      RECT 65.285 3.271 65.335 3.431 ;
      RECT 65.261 3.269 65.285 3.432 ;
      RECT 65.175 3.264 65.261 3.434 ;
      RECT 65.15 3.26 65.175 3.433 ;
      RECT 65.14 3.257 65.15 3.431 ;
      RECT 65.13 3.25 65.14 3.428 ;
      RECT 65.125 3.23 65.13 3.423 ;
      RECT 65.115 3.2 65.125 3.418 ;
      RECT 65.1 3.07 65.115 3.409 ;
      RECT 65.095 3.062 65.1 3.402 ;
      RECT 65.075 3.055 65.095 3.394 ;
      RECT 65.07 3.037 65.075 3.386 ;
      RECT 65.06 3.017 65.07 3.381 ;
      RECT 65.055 2.99 65.06 3.377 ;
      RECT 65.05 2.967 65.055 3.374 ;
      RECT 65.03 2.925 65.05 3.366 ;
      RECT 64.995 2.84 65.03 3.35 ;
      RECT 64.99 2.772 64.995 3.338 ;
      RECT 64.975 2.742 64.99 3.332 ;
      RECT 64.97 1.987 64.975 2.233 ;
      RECT 64.96 2.712 64.975 3.323 ;
      RECT 64.965 1.982 64.97 2.265 ;
      RECT 64.96 1.977 64.965 2.308 ;
      RECT 64.955 1.975 64.96 2.343 ;
      RECT 64.94 2.675 64.96 3.313 ;
      RECT 64.95 1.975 64.955 2.38 ;
      RECT 64.935 1.975 64.95 2.478 ;
      RECT 64.935 2.648 64.94 3.306 ;
      RECT 64.93 1.975 64.935 2.553 ;
      RECT 64.93 2.636 64.935 3.303 ;
      RECT 64.925 1.975 64.93 2.585 ;
      RECT 64.925 2.615 64.93 3.3 ;
      RECT 64.92 1.975 64.925 3.297 ;
      RECT 64.885 1.975 64.92 3.283 ;
      RECT 64.87 1.975 64.885 3.265 ;
      RECT 64.85 1.975 64.87 3.255 ;
      RECT 64.825 1.975 64.85 3.238 ;
      RECT 64.82 1.975 64.825 3.188 ;
      RECT 64.81 1.975 64.815 3.018 ;
      RECT 64.805 1.975 64.81 2.925 ;
      RECT 64.8 1.975 64.805 2.838 ;
      RECT 64.795 1.975 64.8 2.77 ;
      RECT 64.79 1.975 64.795 2.713 ;
      RECT 64.78 1.975 64.79 2.608 ;
      RECT 64.775 1.975 64.78 2.48 ;
      RECT 64.77 1.975 64.775 2.398 ;
      RECT 64.765 1.977 64.77 2.315 ;
      RECT 64.76 1.982 64.765 2.248 ;
      RECT 64.755 1.987 64.76 2.175 ;
      RECT 67.57 2.305 67.83 2.565 ;
      RECT 67.59 2.272 67.8 2.565 ;
      RECT 67.59 2.27 67.79 2.565 ;
      RECT 67.6 2.257 67.79 2.565 ;
      RECT 67.6 2.255 67.715 2.565 ;
      RECT 67.075 2.38 67.25 2.66 ;
      RECT 67.07 2.38 67.25 2.658 ;
      RECT 67.07 2.38 67.265 2.655 ;
      RECT 67.06 2.38 67.265 2.653 ;
      RECT 67.005 2.38 67.265 2.64 ;
      RECT 67.005 2.455 67.27 2.618 ;
      RECT 66.55 2.392 66.57 2.635 ;
      RECT 66.55 2.392 66.61 2.634 ;
      RECT 66.545 2.394 66.61 2.633 ;
      RECT 66.545 2.394 66.696 2.632 ;
      RECT 66.545 2.394 66.765 2.631 ;
      RECT 66.545 2.394 66.785 2.623 ;
      RECT 66.525 2.397 66.785 2.621 ;
      RECT 66.51 2.407 66.785 2.606 ;
      RECT 66.51 2.407 66.8 2.605 ;
      RECT 66.505 2.416 66.8 2.597 ;
      RECT 66.505 2.416 66.805 2.593 ;
      RECT 66.61 2.33 66.87 2.59 ;
      RECT 66.5 2.418 66.87 2.475 ;
      RECT 66.57 2.385 66.87 2.59 ;
      RECT 66.535 3.578 66.54 3.785 ;
      RECT 66.485 3.572 66.535 3.784 ;
      RECT 66.452 3.586 66.545 3.783 ;
      RECT 66.366 3.586 66.545 3.782 ;
      RECT 66.28 3.586 66.545 3.781 ;
      RECT 66.28 3.685 66.55 3.778 ;
      RECT 66.275 3.685 66.55 3.773 ;
      RECT 66.27 3.685 66.55 3.755 ;
      RECT 66.265 3.685 66.55 3.738 ;
      RECT 66.225 3.47 66.485 3.73 ;
      RECT 65.685 2.62 65.771 3.034 ;
      RECT 65.685 2.62 65.81 3.031 ;
      RECT 65.685 2.62 65.83 3.021 ;
      RECT 65.64 2.62 65.83 3.018 ;
      RECT 65.64 2.772 65.84 3.008 ;
      RECT 65.64 2.793 65.845 3.002 ;
      RECT 65.64 2.811 65.85 2.998 ;
      RECT 65.64 2.831 65.86 2.993 ;
      RECT 65.615 2.831 65.86 2.99 ;
      RECT 65.605 2.831 65.86 2.968 ;
      RECT 65.605 2.847 65.865 2.938 ;
      RECT 65.57 2.62 65.83 2.925 ;
      RECT 65.57 2.859 65.87 2.88 ;
      RECT 63.23 7.77 63.52 8 ;
      RECT 63.29 6.29 63.46 8 ;
      RECT 63.24 6.655 63.59 7.005 ;
      RECT 63.23 6.29 63.52 6.52 ;
      RECT 62.825 2.395 62.93 2.965 ;
      RECT 62.825 2.73 63.15 2.96 ;
      RECT 62.825 2.76 63.32 2.93 ;
      RECT 62.825 2.395 63.015 2.96 ;
      RECT 62.24 2.36 62.53 2.59 ;
      RECT 62.24 2.395 63.015 2.565 ;
      RECT 62.3 0.88 62.47 2.59 ;
      RECT 62.24 0.88 62.53 1.11 ;
      RECT 62.24 7.77 62.53 8 ;
      RECT 62.3 6.29 62.47 8 ;
      RECT 62.24 6.29 62.53 6.52 ;
      RECT 62.24 6.325 63.095 6.485 ;
      RECT 62.925 5.92 63.095 6.485 ;
      RECT 62.24 6.32 62.635 6.485 ;
      RECT 62.86 5.92 63.15 6.15 ;
      RECT 62.86 5.95 63.32 6.12 ;
      RECT 61.87 2.73 62.16 2.96 ;
      RECT 61.87 2.76 62.33 2.93 ;
      RECT 61.935 1.655 62.1 2.96 ;
      RECT 60.45 1.625 60.74 1.855 ;
      RECT 60.45 1.655 62.1 1.825 ;
      RECT 60.51 0.885 60.68 1.855 ;
      RECT 60.45 0.885 60.74 1.115 ;
      RECT 60.45 7.765 60.74 7.995 ;
      RECT 60.51 7.025 60.68 7.995 ;
      RECT 60.51 7.12 62.1 7.29 ;
      RECT 61.93 5.92 62.1 7.29 ;
      RECT 60.45 7.025 60.74 7.255 ;
      RECT 61.87 5.92 62.16 6.15 ;
      RECT 61.87 5.95 62.33 6.12 ;
      RECT 58.5 2.705 58.84 3.055 ;
      RECT 58.59 2.025 58.76 3.055 ;
      RECT 60.88 1.965 61.23 2.315 ;
      RECT 58.59 2.025 61.23 2.195 ;
      RECT 60.905 6.655 61.23 6.98 ;
      RECT 55.445 6.61 55.795 6.96 ;
      RECT 60.88 6.655 61.23 6.885 ;
      RECT 55.245 6.655 55.795 6.885 ;
      RECT 55.075 6.685 61.23 6.855 ;
      RECT 60.105 2.365 60.425 2.685 ;
      RECT 60.075 2.365 60.425 2.595 ;
      RECT 59.905 2.395 60.425 2.565 ;
      RECT 60.105 6.255 60.425 6.545 ;
      RECT 60.075 6.285 60.425 6.515 ;
      RECT 59.905 6.315 60.425 6.485 ;
      RECT 55.795 2.985 55.945 3.26 ;
      RECT 56.335 2.065 56.34 2.285 ;
      RECT 57.485 2.265 57.5 2.463 ;
      RECT 57.45 2.257 57.485 2.47 ;
      RECT 57.42 2.25 57.45 2.47 ;
      RECT 57.365 2.215 57.42 2.47 ;
      RECT 57.3 2.152 57.365 2.47 ;
      RECT 57.295 2.117 57.3 2.468 ;
      RECT 57.29 2.112 57.295 2.46 ;
      RECT 57.285 2.107 57.29 2.446 ;
      RECT 57.28 2.104 57.285 2.439 ;
      RECT 57.235 2.094 57.28 2.39 ;
      RECT 57.215 2.081 57.235 2.325 ;
      RECT 57.21 2.076 57.215 2.298 ;
      RECT 57.205 2.075 57.21 2.291 ;
      RECT 57.2 2.074 57.205 2.284 ;
      RECT 57.115 2.059 57.2 2.23 ;
      RECT 57.085 2.04 57.115 2.18 ;
      RECT 57.005 2.023 57.085 2.165 ;
      RECT 56.97 2.01 57.005 2.15 ;
      RECT 56.962 2.01 56.97 2.145 ;
      RECT 56.876 2.011 56.962 2.145 ;
      RECT 56.79 2.013 56.876 2.145 ;
      RECT 56.765 2.014 56.79 2.149 ;
      RECT 56.69 2.02 56.765 2.164 ;
      RECT 56.607 2.032 56.69 2.188 ;
      RECT 56.521 2.045 56.607 2.214 ;
      RECT 56.435 2.058 56.521 2.24 ;
      RECT 56.4 2.067 56.435 2.259 ;
      RECT 56.35 2.067 56.4 2.272 ;
      RECT 56.34 2.065 56.35 2.283 ;
      RECT 56.325 2.062 56.335 2.285 ;
      RECT 56.31 2.054 56.325 2.293 ;
      RECT 56.295 2.046 56.31 2.313 ;
      RECT 56.29 2.041 56.295 2.37 ;
      RECT 56.275 2.036 56.29 2.443 ;
      RECT 56.27 2.031 56.275 2.485 ;
      RECT 56.265 2.029 56.27 2.513 ;
      RECT 56.26 2.027 56.265 2.535 ;
      RECT 56.25 2.023 56.26 2.578 ;
      RECT 56.245 2.02 56.25 2.603 ;
      RECT 56.24 2.018 56.245 2.623 ;
      RECT 56.235 2.016 56.24 2.647 ;
      RECT 56.23 2.012 56.235 2.67 ;
      RECT 56.225 2.008 56.23 2.693 ;
      RECT 56.19 1.998 56.225 2.8 ;
      RECT 56.185 1.988 56.19 2.898 ;
      RECT 56.18 1.986 56.185 2.925 ;
      RECT 56.175 1.985 56.18 2.945 ;
      RECT 56.17 1.977 56.175 2.965 ;
      RECT 56.165 1.972 56.17 3 ;
      RECT 56.16 1.97 56.165 3.018 ;
      RECT 56.155 1.97 56.16 3.043 ;
      RECT 56.15 1.97 56.155 3.065 ;
      RECT 56.115 1.97 56.15 3.108 ;
      RECT 56.09 1.97 56.115 3.137 ;
      RECT 56.08 1.97 56.09 2.323 ;
      RECT 56.083 2.38 56.09 3.147 ;
      RECT 56.08 2.437 56.083 3.15 ;
      RECT 56.075 1.97 56.08 2.295 ;
      RECT 56.075 2.487 56.08 3.153 ;
      RECT 56.065 1.97 56.075 2.285 ;
      RECT 56.07 2.54 56.075 3.156 ;
      RECT 56.065 2.625 56.07 3.16 ;
      RECT 56.055 1.97 56.065 2.273 ;
      RECT 56.06 2.672 56.065 3.164 ;
      RECT 56.055 2.747 56.06 3.168 ;
      RECT 56.02 1.97 56.055 2.248 ;
      RECT 56.045 2.83 56.055 3.173 ;
      RECT 56.035 2.897 56.045 3.18 ;
      RECT 56.03 2.925 56.035 3.185 ;
      RECT 56.02 2.938 56.03 3.191 ;
      RECT 55.975 1.97 56.02 2.205 ;
      RECT 56.015 2.943 56.02 3.198 ;
      RECT 55.975 2.96 56.015 3.26 ;
      RECT 55.97 1.972 55.975 2.178 ;
      RECT 55.945 2.98 55.975 3.26 ;
      RECT 55.965 1.977 55.97 2.15 ;
      RECT 55.755 2.989 55.795 3.26 ;
      RECT 55.73 2.997 55.755 3.23 ;
      RECT 55.685 3.005 55.73 3.23 ;
      RECT 55.67 3.01 55.685 3.225 ;
      RECT 55.66 3.01 55.67 3.219 ;
      RECT 55.65 3.017 55.66 3.216 ;
      RECT 55.645 3.055 55.65 3.205 ;
      RECT 55.64 3.117 55.645 3.183 ;
      RECT 56.91 2.992 57.095 3.215 ;
      RECT 56.91 3.007 57.1 3.211 ;
      RECT 56.9 2.28 56.985 3.21 ;
      RECT 56.9 3.007 57.105 3.204 ;
      RECT 56.895 3.015 57.105 3.203 ;
      RECT 57.1 2.735 57.42 3.055 ;
      RECT 56.895 2.907 57.065 2.998 ;
      RECT 56.89 2.907 57.065 2.98 ;
      RECT 56.88 2.715 57.015 2.955 ;
      RECT 56.875 2.715 57.015 2.9 ;
      RECT 56.835 2.295 57.005 2.8 ;
      RECT 56.82 2.295 57.005 2.67 ;
      RECT 56.815 2.295 57.005 2.623 ;
      RECT 56.81 2.295 57.005 2.603 ;
      RECT 56.805 2.295 57.005 2.578 ;
      RECT 56.775 2.295 57.035 2.555 ;
      RECT 56.785 2.292 56.995 2.555 ;
      RECT 56.91 2.287 56.995 3.215 ;
      RECT 56.795 2.28 56.985 2.555 ;
      RECT 56.79 2.285 56.985 2.555 ;
      RECT 55.62 2.497 55.805 2.71 ;
      RECT 55.62 2.505 55.815 2.703 ;
      RECT 55.6 2.505 55.815 2.7 ;
      RECT 55.595 2.505 55.815 2.685 ;
      RECT 55.525 2.42 55.785 2.68 ;
      RECT 55.525 2.565 55.82 2.593 ;
      RECT 55.18 3.02 55.44 3.28 ;
      RECT 55.205 2.965 55.4 3.28 ;
      RECT 55.2 2.714 55.38 3.008 ;
      RECT 55.2 2.72 55.39 3.008 ;
      RECT 55.18 2.722 55.39 2.953 ;
      RECT 55.175 2.732 55.39 2.82 ;
      RECT 55.205 2.712 55.38 3.28 ;
      RECT 55.291 2.71 55.38 3.28 ;
      RECT 55.15 1.93 55.185 2.3 ;
      RECT 54.94 2.04 54.945 2.3 ;
      RECT 55.185 1.937 55.2 2.3 ;
      RECT 55.075 1.93 55.15 2.378 ;
      RECT 55.065 1.93 55.075 2.463 ;
      RECT 55.04 1.93 55.065 2.498 ;
      RECT 55 1.93 55.04 2.566 ;
      RECT 54.99 1.937 55 2.618 ;
      RECT 54.96 2.04 54.99 2.659 ;
      RECT 54.955 2.04 54.96 2.698 ;
      RECT 54.945 2.04 54.955 2.718 ;
      RECT 54.94 2.335 54.945 2.755 ;
      RECT 54.935 2.352 54.94 2.775 ;
      RECT 54.92 2.415 54.935 2.815 ;
      RECT 54.915 2.458 54.92 2.85 ;
      RECT 54.91 2.466 54.915 2.863 ;
      RECT 54.9 2.48 54.91 2.885 ;
      RECT 54.875 2.515 54.9 2.95 ;
      RECT 54.865 2.55 54.875 3.013 ;
      RECT 54.845 2.58 54.865 3.074 ;
      RECT 54.83 2.616 54.845 3.141 ;
      RECT 54.82 2.644 54.83 3.18 ;
      RECT 54.81 2.666 54.82 3.2 ;
      RECT 54.805 2.676 54.81 3.211 ;
      RECT 54.8 2.685 54.805 3.214 ;
      RECT 54.79 2.703 54.8 3.218 ;
      RECT 54.78 2.721 54.79 3.219 ;
      RECT 54.755 2.76 54.78 3.216 ;
      RECT 54.735 2.802 54.755 3.213 ;
      RECT 54.72 2.84 54.735 3.212 ;
      RECT 54.685 2.875 54.72 3.209 ;
      RECT 54.68 2.897 54.685 3.207 ;
      RECT 54.615 2.937 54.68 3.204 ;
      RECT 54.61 2.977 54.615 3.2 ;
      RECT 54.595 2.987 54.61 3.191 ;
      RECT 54.585 3.107 54.595 3.176 ;
      RECT 55.065 3.52 55.075 3.78 ;
      RECT 55.065 3.523 55.085 3.779 ;
      RECT 55.055 3.513 55.065 3.778 ;
      RECT 55.045 3.528 55.125 3.774 ;
      RECT 55.03 3.507 55.045 3.772 ;
      RECT 55.005 3.532 55.13 3.768 ;
      RECT 54.99 3.492 55.005 3.763 ;
      RECT 54.99 3.534 55.14 3.762 ;
      RECT 54.99 3.542 55.155 3.755 ;
      RECT 54.93 3.479 54.99 3.745 ;
      RECT 54.92 3.466 54.93 3.727 ;
      RECT 54.895 3.456 54.92 3.717 ;
      RECT 54.89 3.446 54.895 3.709 ;
      RECT 54.825 3.542 55.155 3.691 ;
      RECT 54.74 3.542 55.155 3.653 ;
      RECT 54.63 3.37 54.89 3.63 ;
      RECT 55.005 3.5 55.03 3.768 ;
      RECT 55.045 3.51 55.055 3.774 ;
      RECT 54.63 3.518 55.07 3.63 ;
      RECT 54.815 7.765 55.105 7.995 ;
      RECT 54.875 7.025 55.045 7.995 ;
      RECT 54.775 7.055 55.145 7.425 ;
      RECT 54.815 7.025 55.105 7.425 ;
      RECT 53.845 3.275 53.875 3.575 ;
      RECT 53.62 3.26 53.625 3.535 ;
      RECT 53.42 3.26 53.575 3.52 ;
      RECT 54.72 1.975 54.75 2.235 ;
      RECT 54.71 1.975 54.72 2.343 ;
      RECT 54.69 1.975 54.71 2.353 ;
      RECT 54.675 1.975 54.69 2.365 ;
      RECT 54.62 1.975 54.675 2.415 ;
      RECT 54.605 1.975 54.62 2.463 ;
      RECT 54.575 1.975 54.605 2.498 ;
      RECT 54.52 1.975 54.575 2.56 ;
      RECT 54.5 1.975 54.52 2.628 ;
      RECT 54.495 1.975 54.5 2.658 ;
      RECT 54.49 1.975 54.495 2.67 ;
      RECT 54.485 2.092 54.49 2.688 ;
      RECT 54.465 2.11 54.485 2.713 ;
      RECT 54.445 2.137 54.465 2.763 ;
      RECT 54.44 2.157 54.445 2.794 ;
      RECT 54.435 2.165 54.44 2.811 ;
      RECT 54.42 2.191 54.435 2.84 ;
      RECT 54.405 2.233 54.42 2.875 ;
      RECT 54.4 2.262 54.405 2.898 ;
      RECT 54.395 2.277 54.4 2.911 ;
      RECT 54.39 2.3 54.395 2.922 ;
      RECT 54.38 2.32 54.39 2.94 ;
      RECT 54.37 2.35 54.38 2.963 ;
      RECT 54.365 2.372 54.37 2.983 ;
      RECT 54.36 2.387 54.365 2.998 ;
      RECT 54.345 2.417 54.36 3.025 ;
      RECT 54.34 2.447 54.345 3.051 ;
      RECT 54.335 2.465 54.34 3.063 ;
      RECT 54.325 2.495 54.335 3.082 ;
      RECT 54.315 2.52 54.325 3.107 ;
      RECT 54.31 2.54 54.315 3.126 ;
      RECT 54.305 2.557 54.31 3.139 ;
      RECT 54.295 2.583 54.305 3.158 ;
      RECT 54.285 2.621 54.295 3.185 ;
      RECT 54.28 2.647 54.285 3.205 ;
      RECT 54.275 2.657 54.28 3.215 ;
      RECT 54.27 2.67 54.275 3.23 ;
      RECT 54.265 2.685 54.27 3.24 ;
      RECT 54.26 2.707 54.265 3.255 ;
      RECT 54.255 2.725 54.26 3.266 ;
      RECT 54.25 2.735 54.255 3.277 ;
      RECT 54.245 2.743 54.25 3.289 ;
      RECT 54.24 2.751 54.245 3.3 ;
      RECT 54.235 2.777 54.24 3.313 ;
      RECT 54.225 2.805 54.235 3.326 ;
      RECT 54.22 2.835 54.225 3.335 ;
      RECT 54.215 2.85 54.22 3.342 ;
      RECT 54.2 2.875 54.215 3.349 ;
      RECT 54.195 2.897 54.2 3.355 ;
      RECT 54.19 2.922 54.195 3.358 ;
      RECT 54.181 2.95 54.19 3.362 ;
      RECT 54.175 2.967 54.181 3.367 ;
      RECT 54.17 2.985 54.175 3.371 ;
      RECT 54.165 2.997 54.17 3.374 ;
      RECT 54.16 3.018 54.165 3.378 ;
      RECT 54.155 3.036 54.16 3.381 ;
      RECT 54.15 3.05 54.155 3.384 ;
      RECT 54.145 3.067 54.15 3.387 ;
      RECT 54.14 3.08 54.145 3.39 ;
      RECT 54.115 3.117 54.14 3.398 ;
      RECT 54.11 3.162 54.115 3.407 ;
      RECT 54.105 3.19 54.11 3.41 ;
      RECT 54.095 3.21 54.105 3.414 ;
      RECT 54.09 3.23 54.095 3.419 ;
      RECT 54.085 3.245 54.09 3.422 ;
      RECT 54.065 3.255 54.085 3.429 ;
      RECT 54 3.262 54.065 3.455 ;
      RECT 53.965 3.265 54 3.483 ;
      RECT 53.95 3.268 53.965 3.498 ;
      RECT 53.94 3.269 53.95 3.513 ;
      RECT 53.93 3.27 53.94 3.53 ;
      RECT 53.925 3.27 53.93 3.545 ;
      RECT 53.92 3.27 53.925 3.553 ;
      RECT 53.905 3.271 53.92 3.568 ;
      RECT 53.875 3.273 53.905 3.575 ;
      RECT 53.765 3.28 53.845 3.575 ;
      RECT 53.72 3.285 53.765 3.575 ;
      RECT 53.71 3.286 53.72 3.565 ;
      RECT 53.7 3.287 53.71 3.558 ;
      RECT 53.68 3.289 53.7 3.553 ;
      RECT 53.67 3.26 53.68 3.548 ;
      RECT 53.625 3.26 53.67 3.54 ;
      RECT 53.595 3.26 53.62 3.53 ;
      RECT 53.575 3.26 53.595 3.523 ;
      RECT 53.855 2.06 54.115 2.32 ;
      RECT 53.735 2.075 53.745 2.24 ;
      RECT 53.72 2.075 53.725 2.235 ;
      RECT 51.085 1.915 51.27 2.205 ;
      RECT 52.9 2.04 52.915 2.195 ;
      RECT 51.05 1.915 51.075 2.175 ;
      RECT 53.465 1.965 53.47 2.107 ;
      RECT 53.38 1.96 53.405 2.1 ;
      RECT 53.78 2.077 53.855 2.27 ;
      RECT 53.765 2.075 53.78 2.253 ;
      RECT 53.745 2.075 53.765 2.245 ;
      RECT 53.725 2.075 53.735 2.238 ;
      RECT 53.68 2.07 53.72 2.228 ;
      RECT 53.64 2.045 53.68 2.213 ;
      RECT 53.625 2.02 53.64 2.203 ;
      RECT 53.62 2.014 53.625 2.201 ;
      RECT 53.585 2.006 53.62 2.184 ;
      RECT 53.58 1.999 53.585 2.172 ;
      RECT 53.56 1.994 53.58 2.16 ;
      RECT 53.55 1.988 53.56 2.145 ;
      RECT 53.53 1.983 53.55 2.13 ;
      RECT 53.52 1.978 53.53 2.123 ;
      RECT 53.515 1.976 53.52 2.118 ;
      RECT 53.51 1.975 53.515 2.115 ;
      RECT 53.47 1.97 53.51 2.111 ;
      RECT 53.45 1.964 53.465 2.106 ;
      RECT 53.415 1.961 53.45 2.103 ;
      RECT 53.405 1.96 53.415 2.101 ;
      RECT 53.345 1.96 53.38 2.098 ;
      RECT 53.3 1.96 53.345 2.098 ;
      RECT 53.25 1.96 53.3 2.101 ;
      RECT 53.235 1.962 53.25 2.103 ;
      RECT 53.22 1.965 53.235 2.104 ;
      RECT 53.21 1.97 53.22 2.105 ;
      RECT 53.18 1.975 53.21 2.11 ;
      RECT 53.17 1.981 53.18 2.118 ;
      RECT 53.16 1.983 53.17 2.122 ;
      RECT 53.15 1.987 53.16 2.126 ;
      RECT 53.125 1.993 53.15 2.134 ;
      RECT 53.115 1.998 53.125 2.142 ;
      RECT 53.1 2.002 53.115 2.146 ;
      RECT 53.065 2.008 53.1 2.154 ;
      RECT 53.045 2.013 53.065 2.164 ;
      RECT 53.015 2.02 53.045 2.173 ;
      RECT 52.97 2.029 53.015 2.187 ;
      RECT 52.965 2.034 52.97 2.198 ;
      RECT 52.945 2.037 52.965 2.199 ;
      RECT 52.915 2.04 52.945 2.197 ;
      RECT 52.88 2.04 52.9 2.193 ;
      RECT 52.81 2.04 52.88 2.184 ;
      RECT 52.795 2.037 52.81 2.176 ;
      RECT 52.755 2.03 52.795 2.171 ;
      RECT 52.73 2.02 52.755 2.164 ;
      RECT 52.725 2.014 52.73 2.161 ;
      RECT 52.685 2.008 52.725 2.158 ;
      RECT 52.67 2.001 52.685 2.153 ;
      RECT 52.65 1.997 52.67 2.148 ;
      RECT 52.635 1.992 52.65 2.144 ;
      RECT 52.62 1.987 52.635 2.142 ;
      RECT 52.605 1.983 52.62 2.141 ;
      RECT 52.59 1.981 52.605 2.137 ;
      RECT 52.58 1.979 52.59 2.132 ;
      RECT 52.565 1.976 52.58 2.128 ;
      RECT 52.555 1.974 52.565 2.123 ;
      RECT 52.535 1.971 52.555 2.119 ;
      RECT 52.49 1.97 52.535 2.117 ;
      RECT 52.43 1.972 52.49 2.118 ;
      RECT 52.41 1.974 52.43 2.12 ;
      RECT 52.38 1.977 52.41 2.121 ;
      RECT 52.33 1.982 52.38 2.123 ;
      RECT 52.325 1.985 52.33 2.125 ;
      RECT 52.315 1.987 52.325 2.128 ;
      RECT 52.31 1.989 52.315 2.131 ;
      RECT 52.26 1.992 52.31 2.138 ;
      RECT 52.24 1.996 52.26 2.15 ;
      RECT 52.23 1.999 52.24 2.156 ;
      RECT 52.22 2 52.23 2.159 ;
      RECT 52.181 2.003 52.22 2.161 ;
      RECT 52.095 2.01 52.181 2.164 ;
      RECT 52.021 2.02 52.095 2.168 ;
      RECT 51.935 2.031 52.021 2.173 ;
      RECT 51.92 2.038 51.935 2.175 ;
      RECT 51.865 2.042 51.92 2.176 ;
      RECT 51.851 2.045 51.865 2.178 ;
      RECT 51.765 2.045 51.851 2.18 ;
      RECT 51.725 2.042 51.765 2.183 ;
      RECT 51.701 2.038 51.725 2.185 ;
      RECT 51.615 2.028 51.701 2.188 ;
      RECT 51.585 2.017 51.615 2.189 ;
      RECT 51.566 2.013 51.585 2.188 ;
      RECT 51.48 2.006 51.566 2.185 ;
      RECT 51.42 1.995 51.48 2.182 ;
      RECT 51.4 1.987 51.42 2.18 ;
      RECT 51.365 1.982 51.4 2.179 ;
      RECT 51.34 1.977 51.365 2.178 ;
      RECT 51.31 1.972 51.34 2.177 ;
      RECT 51.285 1.915 51.31 2.176 ;
      RECT 51.27 1.915 51.285 2.2 ;
      RECT 51.075 1.915 51.085 2.2 ;
      RECT 52.85 2.935 52.855 3.075 ;
      RECT 52.51 2.935 52.545 3.073 ;
      RECT 52.085 2.92 52.1 3.065 ;
      RECT 53.915 2.7 54.005 2.96 ;
      RECT 53.745 2.565 53.845 2.96 ;
      RECT 50.78 2.54 50.86 2.75 ;
      RECT 53.87 2.677 53.915 2.96 ;
      RECT 53.86 2.647 53.87 2.96 ;
      RECT 53.845 2.57 53.86 2.96 ;
      RECT 53.66 2.565 53.745 2.925 ;
      RECT 53.655 2.567 53.66 2.92 ;
      RECT 53.65 2.572 53.655 2.92 ;
      RECT 53.615 2.672 53.65 2.92 ;
      RECT 53.605 2.7 53.615 2.92 ;
      RECT 53.595 2.715 53.605 2.92 ;
      RECT 53.585 2.727 53.595 2.92 ;
      RECT 53.58 2.737 53.585 2.92 ;
      RECT 53.565 2.747 53.58 2.922 ;
      RECT 53.56 2.762 53.565 2.924 ;
      RECT 53.545 2.775 53.56 2.926 ;
      RECT 53.54 2.79 53.545 2.929 ;
      RECT 53.52 2.8 53.54 2.933 ;
      RECT 53.505 2.81 53.52 2.936 ;
      RECT 53.47 2.817 53.505 2.941 ;
      RECT 53.426 2.824 53.47 2.949 ;
      RECT 53.34 2.836 53.426 2.962 ;
      RECT 53.315 2.847 53.34 2.973 ;
      RECT 53.285 2.852 53.315 2.978 ;
      RECT 53.25 2.857 53.285 2.986 ;
      RECT 53.22 2.862 53.25 2.993 ;
      RECT 53.195 2.867 53.22 2.998 ;
      RECT 53.13 2.874 53.195 3.007 ;
      RECT 53.06 2.887 53.13 3.023 ;
      RECT 53.03 2.897 53.06 3.035 ;
      RECT 53.005 2.902 53.03 3.042 ;
      RECT 52.95 2.909 53.005 3.05 ;
      RECT 52.945 2.916 52.95 3.055 ;
      RECT 52.94 2.918 52.945 3.056 ;
      RECT 52.925 2.92 52.94 3.058 ;
      RECT 52.92 2.92 52.925 3.061 ;
      RECT 52.855 2.927 52.92 3.068 ;
      RECT 52.82 2.937 52.85 3.078 ;
      RECT 52.803 2.94 52.82 3.08 ;
      RECT 52.717 2.939 52.803 3.079 ;
      RECT 52.631 2.937 52.717 3.076 ;
      RECT 52.545 2.936 52.631 3.074 ;
      RECT 52.444 2.934 52.51 3.073 ;
      RECT 52.358 2.931 52.444 3.071 ;
      RECT 52.272 2.927 52.358 3.069 ;
      RECT 52.186 2.924 52.272 3.068 ;
      RECT 52.1 2.921 52.186 3.066 ;
      RECT 52 2.92 52.085 3.063 ;
      RECT 51.95 2.918 52 3.061 ;
      RECT 51.93 2.915 51.95 3.059 ;
      RECT 51.91 2.913 51.93 3.056 ;
      RECT 51.885 2.909 51.91 3.053 ;
      RECT 51.84 2.903 51.885 3.048 ;
      RECT 51.8 2.897 51.84 3.04 ;
      RECT 51.775 2.892 51.8 3.033 ;
      RECT 51.72 2.885 51.775 3.025 ;
      RECT 51.696 2.878 51.72 3.018 ;
      RECT 51.61 2.869 51.696 3.008 ;
      RECT 51.58 2.861 51.61 2.998 ;
      RECT 51.55 2.857 51.58 2.993 ;
      RECT 51.545 2.854 51.55 2.99 ;
      RECT 51.54 2.853 51.545 2.99 ;
      RECT 51.465 2.846 51.54 2.983 ;
      RECT 51.426 2.837 51.465 2.972 ;
      RECT 51.34 2.827 51.426 2.96 ;
      RECT 51.3 2.817 51.34 2.948 ;
      RECT 51.261 2.812 51.3 2.941 ;
      RECT 51.175 2.802 51.261 2.93 ;
      RECT 51.135 2.79 51.175 2.919 ;
      RECT 51.1 2.775 51.135 2.912 ;
      RECT 51.09 2.765 51.1 2.909 ;
      RECT 51.07 2.75 51.09 2.907 ;
      RECT 51.04 2.72 51.07 2.903 ;
      RECT 51.03 2.7 51.04 2.898 ;
      RECT 51.025 2.692 51.03 2.895 ;
      RECT 51.02 2.685 51.025 2.893 ;
      RECT 51.005 2.672 51.02 2.886 ;
      RECT 51 2.662 51.005 2.878 ;
      RECT 50.995 2.655 51 2.873 ;
      RECT 50.99 2.65 50.995 2.869 ;
      RECT 50.975 2.637 50.99 2.861 ;
      RECT 50.97 2.547 50.975 2.85 ;
      RECT 50.965 2.542 50.97 2.843 ;
      RECT 50.89 2.54 50.965 2.803 ;
      RECT 50.86 2.54 50.89 2.758 ;
      RECT 50.765 2.545 50.78 2.745 ;
      RECT 53.25 2.25 53.51 2.51 ;
      RECT 53.235 2.238 53.415 2.475 ;
      RECT 53.23 2.239 53.415 2.473 ;
      RECT 53.215 2.243 53.425 2.463 ;
      RECT 53.21 2.248 53.43 2.433 ;
      RECT 53.215 2.245 53.43 2.463 ;
      RECT 53.23 2.24 53.425 2.473 ;
      RECT 53.25 2.237 53.415 2.51 ;
      RECT 53.25 2.236 53.405 2.51 ;
      RECT 53.275 2.235 53.405 2.51 ;
      RECT 52.835 2.48 53.095 2.74 ;
      RECT 52.71 2.525 53.095 2.735 ;
      RECT 52.7 2.53 53.095 2.73 ;
      RECT 52.715 3.47 52.73 3.78 ;
      RECT 51.31 3.24 51.32 3.37 ;
      RECT 51.09 3.235 51.195 3.37 ;
      RECT 51.005 3.24 51.055 3.37 ;
      RECT 49.555 1.975 49.56 3.08 ;
      RECT 52.81 3.562 52.815 3.698 ;
      RECT 52.805 3.557 52.81 3.758 ;
      RECT 52.8 3.555 52.805 3.771 ;
      RECT 52.785 3.552 52.8 3.773 ;
      RECT 52.78 3.547 52.785 3.775 ;
      RECT 52.775 3.543 52.78 3.778 ;
      RECT 52.76 3.538 52.775 3.78 ;
      RECT 52.73 3.53 52.76 3.78 ;
      RECT 52.691 3.47 52.715 3.78 ;
      RECT 52.605 3.47 52.691 3.777 ;
      RECT 52.575 3.47 52.605 3.77 ;
      RECT 52.55 3.47 52.575 3.763 ;
      RECT 52.525 3.47 52.55 3.755 ;
      RECT 52.51 3.47 52.525 3.748 ;
      RECT 52.485 3.47 52.51 3.74 ;
      RECT 52.47 3.47 52.485 3.733 ;
      RECT 52.43 3.48 52.47 3.722 ;
      RECT 52.42 3.475 52.43 3.712 ;
      RECT 52.416 3.474 52.42 3.709 ;
      RECT 52.33 3.466 52.416 3.692 ;
      RECT 52.297 3.455 52.33 3.669 ;
      RECT 52.211 3.444 52.297 3.647 ;
      RECT 52.125 3.428 52.211 3.616 ;
      RECT 52.055 3.413 52.125 3.588 ;
      RECT 52.045 3.406 52.055 3.575 ;
      RECT 52.015 3.403 52.045 3.565 ;
      RECT 51.99 3.399 52.015 3.558 ;
      RECT 51.975 3.396 51.99 3.553 ;
      RECT 51.97 3.395 51.975 3.548 ;
      RECT 51.94 3.39 51.97 3.541 ;
      RECT 51.935 3.385 51.94 3.536 ;
      RECT 51.92 3.382 51.935 3.531 ;
      RECT 51.915 3.377 51.92 3.526 ;
      RECT 51.895 3.372 51.915 3.523 ;
      RECT 51.88 3.367 51.895 3.515 ;
      RECT 51.865 3.361 51.88 3.51 ;
      RECT 51.835 3.352 51.865 3.503 ;
      RECT 51.83 3.345 51.835 3.495 ;
      RECT 51.825 3.343 51.83 3.493 ;
      RECT 51.82 3.342 51.825 3.49 ;
      RECT 51.78 3.335 51.82 3.483 ;
      RECT 51.766 3.325 51.78 3.473 ;
      RECT 51.715 3.314 51.766 3.461 ;
      RECT 51.69 3.3 51.715 3.447 ;
      RECT 51.665 3.289 51.69 3.439 ;
      RECT 51.645 3.278 51.665 3.433 ;
      RECT 51.635 3.272 51.645 3.428 ;
      RECT 51.63 3.27 51.635 3.424 ;
      RECT 51.61 3.265 51.63 3.419 ;
      RECT 51.58 3.255 51.61 3.409 ;
      RECT 51.575 3.247 51.58 3.402 ;
      RECT 51.56 3.245 51.575 3.398 ;
      RECT 51.54 3.245 51.56 3.393 ;
      RECT 51.535 3.244 51.54 3.391 ;
      RECT 51.53 3.244 51.535 3.388 ;
      RECT 51.49 3.243 51.53 3.383 ;
      RECT 51.465 3.242 51.49 3.378 ;
      RECT 51.405 3.241 51.465 3.375 ;
      RECT 51.32 3.24 51.405 3.373 ;
      RECT 51.281 3.239 51.31 3.37 ;
      RECT 51.195 3.237 51.281 3.37 ;
      RECT 51.055 3.237 51.09 3.37 ;
      RECT 50.965 3.241 51.005 3.373 ;
      RECT 50.95 3.244 50.965 3.38 ;
      RECT 50.94 3.245 50.95 3.387 ;
      RECT 50.915 3.248 50.94 3.392 ;
      RECT 50.91 3.25 50.915 3.395 ;
      RECT 50.86 3.252 50.91 3.396 ;
      RECT 50.821 3.256 50.86 3.398 ;
      RECT 50.735 3.258 50.821 3.401 ;
      RECT 50.717 3.26 50.735 3.403 ;
      RECT 50.631 3.263 50.717 3.405 ;
      RECT 50.545 3.267 50.631 3.408 ;
      RECT 50.508 3.271 50.545 3.411 ;
      RECT 50.422 3.274 50.508 3.414 ;
      RECT 50.336 3.278 50.422 3.417 ;
      RECT 50.25 3.283 50.336 3.421 ;
      RECT 50.23 3.285 50.25 3.424 ;
      RECT 50.21 3.284 50.23 3.425 ;
      RECT 50.161 3.281 50.21 3.426 ;
      RECT 50.075 3.276 50.161 3.429 ;
      RECT 50.025 3.271 50.075 3.431 ;
      RECT 50.001 3.269 50.025 3.432 ;
      RECT 49.915 3.264 50.001 3.434 ;
      RECT 49.89 3.26 49.915 3.433 ;
      RECT 49.88 3.257 49.89 3.431 ;
      RECT 49.87 3.25 49.88 3.428 ;
      RECT 49.865 3.23 49.87 3.423 ;
      RECT 49.855 3.2 49.865 3.418 ;
      RECT 49.84 3.07 49.855 3.409 ;
      RECT 49.835 3.062 49.84 3.402 ;
      RECT 49.815 3.055 49.835 3.394 ;
      RECT 49.81 3.037 49.815 3.386 ;
      RECT 49.8 3.017 49.81 3.381 ;
      RECT 49.795 2.99 49.8 3.377 ;
      RECT 49.79 2.967 49.795 3.374 ;
      RECT 49.77 2.925 49.79 3.366 ;
      RECT 49.735 2.84 49.77 3.35 ;
      RECT 49.73 2.772 49.735 3.338 ;
      RECT 49.715 2.742 49.73 3.332 ;
      RECT 49.71 1.987 49.715 2.233 ;
      RECT 49.7 2.712 49.715 3.323 ;
      RECT 49.705 1.982 49.71 2.265 ;
      RECT 49.7 1.977 49.705 2.308 ;
      RECT 49.695 1.975 49.7 2.343 ;
      RECT 49.68 2.675 49.7 3.313 ;
      RECT 49.69 1.975 49.695 2.38 ;
      RECT 49.675 1.975 49.69 2.478 ;
      RECT 49.675 2.648 49.68 3.306 ;
      RECT 49.67 1.975 49.675 2.553 ;
      RECT 49.67 2.636 49.675 3.303 ;
      RECT 49.665 1.975 49.67 2.585 ;
      RECT 49.665 2.615 49.67 3.3 ;
      RECT 49.66 1.975 49.665 3.297 ;
      RECT 49.625 1.975 49.66 3.283 ;
      RECT 49.61 1.975 49.625 3.265 ;
      RECT 49.59 1.975 49.61 3.255 ;
      RECT 49.565 1.975 49.59 3.238 ;
      RECT 49.56 1.975 49.565 3.188 ;
      RECT 49.55 1.975 49.555 3.018 ;
      RECT 49.545 1.975 49.55 2.925 ;
      RECT 49.54 1.975 49.545 2.838 ;
      RECT 49.535 1.975 49.54 2.77 ;
      RECT 49.53 1.975 49.535 2.713 ;
      RECT 49.52 1.975 49.53 2.608 ;
      RECT 49.515 1.975 49.52 2.48 ;
      RECT 49.51 1.975 49.515 2.398 ;
      RECT 49.505 1.977 49.51 2.315 ;
      RECT 49.5 1.982 49.505 2.248 ;
      RECT 49.495 1.987 49.5 2.175 ;
      RECT 52.31 2.305 52.57 2.565 ;
      RECT 52.33 2.272 52.54 2.565 ;
      RECT 52.33 2.27 52.53 2.565 ;
      RECT 52.34 2.257 52.53 2.565 ;
      RECT 52.34 2.255 52.455 2.565 ;
      RECT 51.815 2.38 51.99 2.66 ;
      RECT 51.81 2.38 51.99 2.658 ;
      RECT 51.81 2.38 52.005 2.655 ;
      RECT 51.8 2.38 52.005 2.653 ;
      RECT 51.745 2.38 52.005 2.64 ;
      RECT 51.745 2.455 52.01 2.618 ;
      RECT 51.29 2.392 51.31 2.635 ;
      RECT 51.29 2.392 51.35 2.634 ;
      RECT 51.285 2.394 51.35 2.633 ;
      RECT 51.285 2.394 51.436 2.632 ;
      RECT 51.285 2.394 51.505 2.631 ;
      RECT 51.285 2.394 51.525 2.623 ;
      RECT 51.265 2.397 51.525 2.621 ;
      RECT 51.25 2.407 51.525 2.606 ;
      RECT 51.25 2.407 51.54 2.605 ;
      RECT 51.245 2.416 51.54 2.597 ;
      RECT 51.245 2.416 51.545 2.593 ;
      RECT 51.35 2.33 51.61 2.59 ;
      RECT 51.24 2.418 51.61 2.475 ;
      RECT 51.31 2.385 51.61 2.59 ;
      RECT 51.275 3.578 51.28 3.785 ;
      RECT 51.225 3.572 51.275 3.784 ;
      RECT 51.192 3.586 51.285 3.783 ;
      RECT 51.106 3.586 51.285 3.782 ;
      RECT 51.02 3.586 51.285 3.781 ;
      RECT 51.02 3.685 51.29 3.778 ;
      RECT 51.015 3.685 51.29 3.773 ;
      RECT 51.01 3.685 51.29 3.755 ;
      RECT 51.005 3.685 51.29 3.738 ;
      RECT 50.965 3.47 51.225 3.73 ;
      RECT 50.425 2.62 50.511 3.034 ;
      RECT 50.425 2.62 50.55 3.031 ;
      RECT 50.425 2.62 50.57 3.021 ;
      RECT 50.38 2.62 50.57 3.018 ;
      RECT 50.38 2.772 50.58 3.008 ;
      RECT 50.38 2.793 50.585 3.002 ;
      RECT 50.38 2.811 50.59 2.998 ;
      RECT 50.38 2.831 50.6 2.993 ;
      RECT 50.355 2.831 50.6 2.99 ;
      RECT 50.345 2.831 50.6 2.968 ;
      RECT 50.345 2.847 50.605 2.938 ;
      RECT 50.31 2.62 50.57 2.925 ;
      RECT 50.31 2.859 50.61 2.88 ;
      RECT 47.97 7.77 48.26 8 ;
      RECT 48.03 6.29 48.2 8 ;
      RECT 47.98 6.655 48.33 7.005 ;
      RECT 47.97 6.29 48.26 6.52 ;
      RECT 47.565 2.395 47.67 2.965 ;
      RECT 47.565 2.73 47.89 2.96 ;
      RECT 47.565 2.76 48.06 2.93 ;
      RECT 47.565 2.395 47.755 2.96 ;
      RECT 46.98 2.36 47.27 2.59 ;
      RECT 46.98 2.395 47.755 2.565 ;
      RECT 47.04 0.88 47.21 2.59 ;
      RECT 46.98 0.88 47.27 1.11 ;
      RECT 46.98 7.77 47.27 8 ;
      RECT 47.04 6.29 47.21 8 ;
      RECT 46.98 6.29 47.27 6.52 ;
      RECT 46.98 6.325 47.835 6.485 ;
      RECT 47.665 5.92 47.835 6.485 ;
      RECT 46.98 6.32 47.375 6.485 ;
      RECT 47.6 5.92 47.89 6.15 ;
      RECT 47.6 5.95 48.06 6.12 ;
      RECT 46.61 2.73 46.9 2.96 ;
      RECT 46.61 2.76 47.07 2.93 ;
      RECT 46.675 1.655 46.84 2.96 ;
      RECT 45.19 1.625 45.48 1.855 ;
      RECT 45.19 1.655 46.84 1.825 ;
      RECT 45.25 0.885 45.42 1.855 ;
      RECT 45.19 0.885 45.48 1.115 ;
      RECT 45.19 7.765 45.48 7.995 ;
      RECT 45.25 7.025 45.42 7.995 ;
      RECT 45.25 7.12 46.84 7.29 ;
      RECT 46.67 5.92 46.84 7.29 ;
      RECT 45.19 7.025 45.48 7.255 ;
      RECT 46.61 5.92 46.9 6.15 ;
      RECT 46.61 5.95 47.07 6.12 ;
      RECT 43.24 2.705 43.58 3.055 ;
      RECT 43.33 2.025 43.5 3.055 ;
      RECT 45.62 1.965 45.97 2.315 ;
      RECT 43.33 2.025 45.97 2.195 ;
      RECT 45.645 6.655 45.97 6.98 ;
      RECT 40.185 6.615 40.535 6.965 ;
      RECT 45.62 6.655 45.97 6.885 ;
      RECT 39.985 6.655 40.535 6.885 ;
      RECT 39.815 6.685 45.97 6.855 ;
      RECT 44.845 2.365 45.165 2.685 ;
      RECT 44.815 2.365 45.165 2.595 ;
      RECT 44.645 2.395 45.165 2.565 ;
      RECT 44.845 6.255 45.165 6.545 ;
      RECT 44.815 6.285 45.165 6.515 ;
      RECT 44.645 6.315 45.165 6.485 ;
      RECT 40.535 2.985 40.685 3.26 ;
      RECT 41.075 2.065 41.08 2.285 ;
      RECT 42.225 2.265 42.24 2.463 ;
      RECT 42.19 2.257 42.225 2.47 ;
      RECT 42.16 2.25 42.19 2.47 ;
      RECT 42.105 2.215 42.16 2.47 ;
      RECT 42.04 2.152 42.105 2.47 ;
      RECT 42.035 2.117 42.04 2.468 ;
      RECT 42.03 2.112 42.035 2.46 ;
      RECT 42.025 2.107 42.03 2.446 ;
      RECT 42.02 2.104 42.025 2.439 ;
      RECT 41.975 2.094 42.02 2.39 ;
      RECT 41.955 2.081 41.975 2.325 ;
      RECT 41.95 2.076 41.955 2.298 ;
      RECT 41.945 2.075 41.95 2.291 ;
      RECT 41.94 2.074 41.945 2.284 ;
      RECT 41.855 2.059 41.94 2.23 ;
      RECT 41.825 2.04 41.855 2.18 ;
      RECT 41.745 2.023 41.825 2.165 ;
      RECT 41.71 2.01 41.745 2.15 ;
      RECT 41.702 2.01 41.71 2.145 ;
      RECT 41.616 2.011 41.702 2.145 ;
      RECT 41.53 2.013 41.616 2.145 ;
      RECT 41.505 2.014 41.53 2.149 ;
      RECT 41.43 2.02 41.505 2.164 ;
      RECT 41.347 2.032 41.43 2.188 ;
      RECT 41.261 2.045 41.347 2.214 ;
      RECT 41.175 2.058 41.261 2.24 ;
      RECT 41.14 2.067 41.175 2.259 ;
      RECT 41.09 2.067 41.14 2.272 ;
      RECT 41.08 2.065 41.09 2.283 ;
      RECT 41.065 2.062 41.075 2.285 ;
      RECT 41.05 2.054 41.065 2.293 ;
      RECT 41.035 2.046 41.05 2.313 ;
      RECT 41.03 2.041 41.035 2.37 ;
      RECT 41.015 2.036 41.03 2.443 ;
      RECT 41.01 2.031 41.015 2.485 ;
      RECT 41.005 2.029 41.01 2.513 ;
      RECT 41 2.027 41.005 2.535 ;
      RECT 40.99 2.023 41 2.578 ;
      RECT 40.985 2.02 40.99 2.603 ;
      RECT 40.98 2.018 40.985 2.623 ;
      RECT 40.975 2.016 40.98 2.647 ;
      RECT 40.97 2.012 40.975 2.67 ;
      RECT 40.965 2.008 40.97 2.693 ;
      RECT 40.93 1.998 40.965 2.8 ;
      RECT 40.925 1.988 40.93 2.898 ;
      RECT 40.92 1.986 40.925 2.925 ;
      RECT 40.915 1.985 40.92 2.945 ;
      RECT 40.91 1.977 40.915 2.965 ;
      RECT 40.905 1.972 40.91 3 ;
      RECT 40.9 1.97 40.905 3.018 ;
      RECT 40.895 1.97 40.9 3.043 ;
      RECT 40.89 1.97 40.895 3.065 ;
      RECT 40.855 1.97 40.89 3.108 ;
      RECT 40.83 1.97 40.855 3.137 ;
      RECT 40.82 1.97 40.83 2.323 ;
      RECT 40.823 2.38 40.83 3.147 ;
      RECT 40.82 2.437 40.823 3.15 ;
      RECT 40.815 1.97 40.82 2.295 ;
      RECT 40.815 2.487 40.82 3.153 ;
      RECT 40.805 1.97 40.815 2.285 ;
      RECT 40.81 2.54 40.815 3.156 ;
      RECT 40.805 2.625 40.81 3.16 ;
      RECT 40.795 1.97 40.805 2.273 ;
      RECT 40.8 2.672 40.805 3.164 ;
      RECT 40.795 2.747 40.8 3.168 ;
      RECT 40.76 1.97 40.795 2.248 ;
      RECT 40.785 2.83 40.795 3.173 ;
      RECT 40.775 2.897 40.785 3.18 ;
      RECT 40.77 2.925 40.775 3.185 ;
      RECT 40.76 2.938 40.77 3.191 ;
      RECT 40.715 1.97 40.76 2.205 ;
      RECT 40.755 2.943 40.76 3.198 ;
      RECT 40.715 2.96 40.755 3.26 ;
      RECT 40.71 1.972 40.715 2.178 ;
      RECT 40.685 2.98 40.715 3.26 ;
      RECT 40.705 1.977 40.71 2.15 ;
      RECT 40.495 2.989 40.535 3.26 ;
      RECT 40.47 2.997 40.495 3.23 ;
      RECT 40.425 3.005 40.47 3.23 ;
      RECT 40.41 3.01 40.425 3.225 ;
      RECT 40.4 3.01 40.41 3.219 ;
      RECT 40.39 3.017 40.4 3.216 ;
      RECT 40.385 3.055 40.39 3.205 ;
      RECT 40.38 3.117 40.385 3.183 ;
      RECT 41.65 2.992 41.835 3.215 ;
      RECT 41.65 3.007 41.84 3.211 ;
      RECT 41.64 2.28 41.725 3.21 ;
      RECT 41.64 3.007 41.845 3.204 ;
      RECT 41.635 3.015 41.845 3.203 ;
      RECT 41.84 2.735 42.16 3.055 ;
      RECT 41.635 2.907 41.805 2.998 ;
      RECT 41.63 2.907 41.805 2.98 ;
      RECT 41.62 2.715 41.755 2.955 ;
      RECT 41.615 2.715 41.755 2.9 ;
      RECT 41.575 2.295 41.745 2.8 ;
      RECT 41.56 2.295 41.745 2.67 ;
      RECT 41.555 2.295 41.745 2.623 ;
      RECT 41.55 2.295 41.745 2.603 ;
      RECT 41.545 2.295 41.745 2.578 ;
      RECT 41.515 2.295 41.775 2.555 ;
      RECT 41.525 2.292 41.735 2.555 ;
      RECT 41.65 2.287 41.735 3.215 ;
      RECT 41.535 2.28 41.725 2.555 ;
      RECT 41.53 2.285 41.725 2.555 ;
      RECT 40.36 2.497 40.545 2.71 ;
      RECT 40.36 2.505 40.555 2.703 ;
      RECT 40.34 2.505 40.555 2.7 ;
      RECT 40.335 2.505 40.555 2.685 ;
      RECT 40.265 2.42 40.525 2.68 ;
      RECT 40.265 2.565 40.56 2.593 ;
      RECT 39.92 3.02 40.18 3.28 ;
      RECT 39.945 2.965 40.14 3.28 ;
      RECT 39.94 2.714 40.12 3.008 ;
      RECT 39.94 2.72 40.13 3.008 ;
      RECT 39.92 2.722 40.13 2.953 ;
      RECT 39.915 2.732 40.13 2.82 ;
      RECT 39.945 2.712 40.12 3.28 ;
      RECT 40.031 2.71 40.12 3.28 ;
      RECT 39.89 1.93 39.925 2.3 ;
      RECT 39.68 2.04 39.685 2.3 ;
      RECT 39.925 1.937 39.94 2.3 ;
      RECT 39.815 1.93 39.89 2.378 ;
      RECT 39.805 1.93 39.815 2.463 ;
      RECT 39.78 1.93 39.805 2.498 ;
      RECT 39.74 1.93 39.78 2.566 ;
      RECT 39.73 1.937 39.74 2.618 ;
      RECT 39.7 2.04 39.73 2.659 ;
      RECT 39.695 2.04 39.7 2.698 ;
      RECT 39.685 2.04 39.695 2.718 ;
      RECT 39.68 2.335 39.685 2.755 ;
      RECT 39.675 2.352 39.68 2.775 ;
      RECT 39.66 2.415 39.675 2.815 ;
      RECT 39.655 2.458 39.66 2.85 ;
      RECT 39.65 2.466 39.655 2.863 ;
      RECT 39.64 2.48 39.65 2.885 ;
      RECT 39.615 2.515 39.64 2.95 ;
      RECT 39.605 2.55 39.615 3.013 ;
      RECT 39.585 2.58 39.605 3.074 ;
      RECT 39.57 2.616 39.585 3.141 ;
      RECT 39.56 2.644 39.57 3.18 ;
      RECT 39.55 2.666 39.56 3.2 ;
      RECT 39.545 2.676 39.55 3.211 ;
      RECT 39.54 2.685 39.545 3.214 ;
      RECT 39.53 2.703 39.54 3.218 ;
      RECT 39.52 2.721 39.53 3.219 ;
      RECT 39.495 2.76 39.52 3.216 ;
      RECT 39.475 2.802 39.495 3.213 ;
      RECT 39.46 2.84 39.475 3.212 ;
      RECT 39.425 2.875 39.46 3.209 ;
      RECT 39.42 2.897 39.425 3.207 ;
      RECT 39.355 2.937 39.42 3.204 ;
      RECT 39.35 2.977 39.355 3.2 ;
      RECT 39.335 2.987 39.35 3.191 ;
      RECT 39.325 3.107 39.335 3.176 ;
      RECT 39.805 3.52 39.815 3.78 ;
      RECT 39.805 3.523 39.825 3.779 ;
      RECT 39.795 3.513 39.805 3.778 ;
      RECT 39.785 3.528 39.865 3.774 ;
      RECT 39.77 3.507 39.785 3.772 ;
      RECT 39.745 3.532 39.87 3.768 ;
      RECT 39.73 3.492 39.745 3.763 ;
      RECT 39.73 3.534 39.88 3.762 ;
      RECT 39.73 3.542 39.895 3.755 ;
      RECT 39.67 3.479 39.73 3.745 ;
      RECT 39.66 3.466 39.67 3.727 ;
      RECT 39.635 3.456 39.66 3.717 ;
      RECT 39.63 3.446 39.635 3.709 ;
      RECT 39.565 3.542 39.895 3.691 ;
      RECT 39.48 3.542 39.895 3.653 ;
      RECT 39.37 3.37 39.63 3.63 ;
      RECT 39.745 3.5 39.77 3.768 ;
      RECT 39.785 3.51 39.795 3.774 ;
      RECT 39.37 3.518 39.81 3.63 ;
      RECT 39.555 7.765 39.845 7.995 ;
      RECT 39.615 7.025 39.785 7.995 ;
      RECT 39.515 7.055 39.885 7.425 ;
      RECT 39.555 7.025 39.845 7.425 ;
      RECT 38.585 3.275 38.615 3.575 ;
      RECT 38.36 3.26 38.365 3.535 ;
      RECT 38.16 3.26 38.315 3.52 ;
      RECT 39.46 1.975 39.49 2.235 ;
      RECT 39.45 1.975 39.46 2.343 ;
      RECT 39.43 1.975 39.45 2.353 ;
      RECT 39.415 1.975 39.43 2.365 ;
      RECT 39.36 1.975 39.415 2.415 ;
      RECT 39.345 1.975 39.36 2.463 ;
      RECT 39.315 1.975 39.345 2.498 ;
      RECT 39.26 1.975 39.315 2.56 ;
      RECT 39.24 1.975 39.26 2.628 ;
      RECT 39.235 1.975 39.24 2.658 ;
      RECT 39.23 1.975 39.235 2.67 ;
      RECT 39.225 2.092 39.23 2.688 ;
      RECT 39.205 2.11 39.225 2.713 ;
      RECT 39.185 2.137 39.205 2.763 ;
      RECT 39.18 2.157 39.185 2.794 ;
      RECT 39.175 2.165 39.18 2.811 ;
      RECT 39.16 2.191 39.175 2.84 ;
      RECT 39.145 2.233 39.16 2.875 ;
      RECT 39.14 2.262 39.145 2.898 ;
      RECT 39.135 2.277 39.14 2.911 ;
      RECT 39.13 2.3 39.135 2.922 ;
      RECT 39.12 2.32 39.13 2.94 ;
      RECT 39.11 2.35 39.12 2.963 ;
      RECT 39.105 2.372 39.11 2.983 ;
      RECT 39.1 2.387 39.105 2.998 ;
      RECT 39.085 2.417 39.1 3.025 ;
      RECT 39.08 2.447 39.085 3.051 ;
      RECT 39.075 2.465 39.08 3.063 ;
      RECT 39.065 2.495 39.075 3.082 ;
      RECT 39.055 2.52 39.065 3.107 ;
      RECT 39.05 2.54 39.055 3.126 ;
      RECT 39.045 2.557 39.05 3.139 ;
      RECT 39.035 2.583 39.045 3.158 ;
      RECT 39.025 2.621 39.035 3.185 ;
      RECT 39.02 2.647 39.025 3.205 ;
      RECT 39.015 2.657 39.02 3.215 ;
      RECT 39.01 2.67 39.015 3.23 ;
      RECT 39.005 2.685 39.01 3.24 ;
      RECT 39 2.707 39.005 3.255 ;
      RECT 38.995 2.725 39 3.266 ;
      RECT 38.99 2.735 38.995 3.277 ;
      RECT 38.985 2.743 38.99 3.289 ;
      RECT 38.98 2.751 38.985 3.3 ;
      RECT 38.975 2.777 38.98 3.313 ;
      RECT 38.965 2.805 38.975 3.326 ;
      RECT 38.96 2.835 38.965 3.335 ;
      RECT 38.955 2.85 38.96 3.342 ;
      RECT 38.94 2.875 38.955 3.349 ;
      RECT 38.935 2.897 38.94 3.355 ;
      RECT 38.93 2.922 38.935 3.358 ;
      RECT 38.921 2.95 38.93 3.362 ;
      RECT 38.915 2.967 38.921 3.367 ;
      RECT 38.91 2.985 38.915 3.371 ;
      RECT 38.905 2.997 38.91 3.374 ;
      RECT 38.9 3.018 38.905 3.378 ;
      RECT 38.895 3.036 38.9 3.381 ;
      RECT 38.89 3.05 38.895 3.384 ;
      RECT 38.885 3.067 38.89 3.387 ;
      RECT 38.88 3.08 38.885 3.39 ;
      RECT 38.855 3.117 38.88 3.398 ;
      RECT 38.85 3.162 38.855 3.407 ;
      RECT 38.845 3.19 38.85 3.41 ;
      RECT 38.835 3.21 38.845 3.414 ;
      RECT 38.83 3.23 38.835 3.419 ;
      RECT 38.825 3.245 38.83 3.422 ;
      RECT 38.805 3.255 38.825 3.429 ;
      RECT 38.74 3.262 38.805 3.455 ;
      RECT 38.705 3.265 38.74 3.483 ;
      RECT 38.69 3.268 38.705 3.498 ;
      RECT 38.68 3.269 38.69 3.513 ;
      RECT 38.67 3.27 38.68 3.53 ;
      RECT 38.665 3.27 38.67 3.545 ;
      RECT 38.66 3.27 38.665 3.553 ;
      RECT 38.645 3.271 38.66 3.568 ;
      RECT 38.615 3.273 38.645 3.575 ;
      RECT 38.505 3.28 38.585 3.575 ;
      RECT 38.46 3.285 38.505 3.575 ;
      RECT 38.45 3.286 38.46 3.565 ;
      RECT 38.44 3.287 38.45 3.558 ;
      RECT 38.42 3.289 38.44 3.553 ;
      RECT 38.41 3.26 38.42 3.548 ;
      RECT 38.365 3.26 38.41 3.54 ;
      RECT 38.335 3.26 38.36 3.53 ;
      RECT 38.315 3.26 38.335 3.523 ;
      RECT 38.595 2.06 38.855 2.32 ;
      RECT 38.475 2.075 38.485 2.24 ;
      RECT 38.46 2.075 38.465 2.235 ;
      RECT 35.825 1.915 36.01 2.205 ;
      RECT 37.64 2.04 37.655 2.195 ;
      RECT 35.79 1.915 35.815 2.175 ;
      RECT 38.205 1.965 38.21 2.107 ;
      RECT 38.12 1.96 38.145 2.1 ;
      RECT 38.52 2.077 38.595 2.27 ;
      RECT 38.505 2.075 38.52 2.253 ;
      RECT 38.485 2.075 38.505 2.245 ;
      RECT 38.465 2.075 38.475 2.238 ;
      RECT 38.42 2.07 38.46 2.228 ;
      RECT 38.38 2.045 38.42 2.213 ;
      RECT 38.365 2.02 38.38 2.203 ;
      RECT 38.36 2.014 38.365 2.201 ;
      RECT 38.325 2.006 38.36 2.184 ;
      RECT 38.32 1.999 38.325 2.172 ;
      RECT 38.3 1.994 38.32 2.16 ;
      RECT 38.29 1.988 38.3 2.145 ;
      RECT 38.27 1.983 38.29 2.13 ;
      RECT 38.26 1.978 38.27 2.123 ;
      RECT 38.255 1.976 38.26 2.118 ;
      RECT 38.25 1.975 38.255 2.115 ;
      RECT 38.21 1.97 38.25 2.111 ;
      RECT 38.19 1.964 38.205 2.106 ;
      RECT 38.155 1.961 38.19 2.103 ;
      RECT 38.145 1.96 38.155 2.101 ;
      RECT 38.085 1.96 38.12 2.098 ;
      RECT 38.04 1.96 38.085 2.098 ;
      RECT 37.99 1.96 38.04 2.101 ;
      RECT 37.975 1.962 37.99 2.103 ;
      RECT 37.96 1.965 37.975 2.104 ;
      RECT 37.95 1.97 37.96 2.105 ;
      RECT 37.92 1.975 37.95 2.11 ;
      RECT 37.91 1.981 37.92 2.118 ;
      RECT 37.9 1.983 37.91 2.122 ;
      RECT 37.89 1.987 37.9 2.126 ;
      RECT 37.865 1.993 37.89 2.134 ;
      RECT 37.855 1.998 37.865 2.142 ;
      RECT 37.84 2.002 37.855 2.146 ;
      RECT 37.805 2.008 37.84 2.154 ;
      RECT 37.785 2.013 37.805 2.164 ;
      RECT 37.755 2.02 37.785 2.173 ;
      RECT 37.71 2.029 37.755 2.187 ;
      RECT 37.705 2.034 37.71 2.198 ;
      RECT 37.685 2.037 37.705 2.199 ;
      RECT 37.655 2.04 37.685 2.197 ;
      RECT 37.62 2.04 37.64 2.193 ;
      RECT 37.55 2.04 37.62 2.184 ;
      RECT 37.535 2.037 37.55 2.176 ;
      RECT 37.495 2.03 37.535 2.171 ;
      RECT 37.47 2.02 37.495 2.164 ;
      RECT 37.465 2.014 37.47 2.161 ;
      RECT 37.425 2.008 37.465 2.158 ;
      RECT 37.41 2.001 37.425 2.153 ;
      RECT 37.39 1.997 37.41 2.148 ;
      RECT 37.375 1.992 37.39 2.144 ;
      RECT 37.36 1.987 37.375 2.142 ;
      RECT 37.345 1.983 37.36 2.141 ;
      RECT 37.33 1.981 37.345 2.137 ;
      RECT 37.32 1.979 37.33 2.132 ;
      RECT 37.305 1.976 37.32 2.128 ;
      RECT 37.295 1.974 37.305 2.123 ;
      RECT 37.275 1.971 37.295 2.119 ;
      RECT 37.23 1.97 37.275 2.117 ;
      RECT 37.17 1.972 37.23 2.118 ;
      RECT 37.15 1.974 37.17 2.12 ;
      RECT 37.12 1.977 37.15 2.121 ;
      RECT 37.07 1.982 37.12 2.123 ;
      RECT 37.065 1.985 37.07 2.125 ;
      RECT 37.055 1.987 37.065 2.128 ;
      RECT 37.05 1.989 37.055 2.131 ;
      RECT 37 1.992 37.05 2.138 ;
      RECT 36.98 1.996 37 2.15 ;
      RECT 36.97 1.999 36.98 2.156 ;
      RECT 36.96 2 36.97 2.159 ;
      RECT 36.921 2.003 36.96 2.161 ;
      RECT 36.835 2.01 36.921 2.164 ;
      RECT 36.761 2.02 36.835 2.168 ;
      RECT 36.675 2.031 36.761 2.173 ;
      RECT 36.66 2.038 36.675 2.175 ;
      RECT 36.605 2.042 36.66 2.176 ;
      RECT 36.591 2.045 36.605 2.178 ;
      RECT 36.505 2.045 36.591 2.18 ;
      RECT 36.465 2.042 36.505 2.183 ;
      RECT 36.441 2.038 36.465 2.185 ;
      RECT 36.355 2.028 36.441 2.188 ;
      RECT 36.325 2.017 36.355 2.189 ;
      RECT 36.306 2.013 36.325 2.188 ;
      RECT 36.22 2.006 36.306 2.185 ;
      RECT 36.16 1.995 36.22 2.182 ;
      RECT 36.14 1.987 36.16 2.18 ;
      RECT 36.105 1.982 36.14 2.179 ;
      RECT 36.08 1.977 36.105 2.178 ;
      RECT 36.05 1.972 36.08 2.177 ;
      RECT 36.025 1.915 36.05 2.176 ;
      RECT 36.01 1.915 36.025 2.2 ;
      RECT 35.815 1.915 35.825 2.2 ;
      RECT 37.59 2.935 37.595 3.075 ;
      RECT 37.25 2.935 37.285 3.073 ;
      RECT 36.825 2.92 36.84 3.065 ;
      RECT 38.655 2.7 38.745 2.96 ;
      RECT 38.485 2.565 38.585 2.96 ;
      RECT 35.52 2.54 35.6 2.75 ;
      RECT 38.61 2.677 38.655 2.96 ;
      RECT 38.6 2.647 38.61 2.96 ;
      RECT 38.585 2.57 38.6 2.96 ;
      RECT 38.4 2.565 38.485 2.925 ;
      RECT 38.395 2.567 38.4 2.92 ;
      RECT 38.39 2.572 38.395 2.92 ;
      RECT 38.355 2.672 38.39 2.92 ;
      RECT 38.345 2.7 38.355 2.92 ;
      RECT 38.335 2.715 38.345 2.92 ;
      RECT 38.325 2.727 38.335 2.92 ;
      RECT 38.32 2.737 38.325 2.92 ;
      RECT 38.305 2.747 38.32 2.922 ;
      RECT 38.3 2.762 38.305 2.924 ;
      RECT 38.285 2.775 38.3 2.926 ;
      RECT 38.28 2.79 38.285 2.929 ;
      RECT 38.26 2.8 38.28 2.933 ;
      RECT 38.245 2.81 38.26 2.936 ;
      RECT 38.21 2.817 38.245 2.941 ;
      RECT 38.166 2.824 38.21 2.949 ;
      RECT 38.08 2.836 38.166 2.962 ;
      RECT 38.055 2.847 38.08 2.973 ;
      RECT 38.025 2.852 38.055 2.978 ;
      RECT 37.99 2.857 38.025 2.986 ;
      RECT 37.96 2.862 37.99 2.993 ;
      RECT 37.935 2.867 37.96 2.998 ;
      RECT 37.87 2.874 37.935 3.007 ;
      RECT 37.8 2.887 37.87 3.023 ;
      RECT 37.77 2.897 37.8 3.035 ;
      RECT 37.745 2.902 37.77 3.042 ;
      RECT 37.69 2.909 37.745 3.05 ;
      RECT 37.685 2.916 37.69 3.055 ;
      RECT 37.68 2.918 37.685 3.056 ;
      RECT 37.665 2.92 37.68 3.058 ;
      RECT 37.66 2.92 37.665 3.061 ;
      RECT 37.595 2.927 37.66 3.068 ;
      RECT 37.56 2.937 37.59 3.078 ;
      RECT 37.543 2.94 37.56 3.08 ;
      RECT 37.457 2.939 37.543 3.079 ;
      RECT 37.371 2.937 37.457 3.076 ;
      RECT 37.285 2.936 37.371 3.074 ;
      RECT 37.184 2.934 37.25 3.073 ;
      RECT 37.098 2.931 37.184 3.071 ;
      RECT 37.012 2.927 37.098 3.069 ;
      RECT 36.926 2.924 37.012 3.068 ;
      RECT 36.84 2.921 36.926 3.066 ;
      RECT 36.74 2.92 36.825 3.063 ;
      RECT 36.69 2.918 36.74 3.061 ;
      RECT 36.67 2.915 36.69 3.059 ;
      RECT 36.65 2.913 36.67 3.056 ;
      RECT 36.625 2.909 36.65 3.053 ;
      RECT 36.58 2.903 36.625 3.048 ;
      RECT 36.54 2.897 36.58 3.04 ;
      RECT 36.515 2.892 36.54 3.033 ;
      RECT 36.46 2.885 36.515 3.025 ;
      RECT 36.436 2.878 36.46 3.018 ;
      RECT 36.35 2.869 36.436 3.008 ;
      RECT 36.32 2.861 36.35 2.998 ;
      RECT 36.29 2.857 36.32 2.993 ;
      RECT 36.285 2.854 36.29 2.99 ;
      RECT 36.28 2.853 36.285 2.99 ;
      RECT 36.205 2.846 36.28 2.983 ;
      RECT 36.166 2.837 36.205 2.972 ;
      RECT 36.08 2.827 36.166 2.96 ;
      RECT 36.04 2.817 36.08 2.948 ;
      RECT 36.001 2.812 36.04 2.941 ;
      RECT 35.915 2.802 36.001 2.93 ;
      RECT 35.875 2.79 35.915 2.919 ;
      RECT 35.84 2.775 35.875 2.912 ;
      RECT 35.83 2.765 35.84 2.909 ;
      RECT 35.81 2.75 35.83 2.907 ;
      RECT 35.78 2.72 35.81 2.903 ;
      RECT 35.77 2.7 35.78 2.898 ;
      RECT 35.765 2.692 35.77 2.895 ;
      RECT 35.76 2.685 35.765 2.893 ;
      RECT 35.745 2.672 35.76 2.886 ;
      RECT 35.74 2.662 35.745 2.878 ;
      RECT 35.735 2.655 35.74 2.873 ;
      RECT 35.73 2.65 35.735 2.869 ;
      RECT 35.715 2.637 35.73 2.861 ;
      RECT 35.71 2.547 35.715 2.85 ;
      RECT 35.705 2.542 35.71 2.843 ;
      RECT 35.63 2.54 35.705 2.803 ;
      RECT 35.6 2.54 35.63 2.758 ;
      RECT 35.505 2.545 35.52 2.745 ;
      RECT 37.99 2.25 38.25 2.51 ;
      RECT 37.975 2.238 38.155 2.475 ;
      RECT 37.97 2.239 38.155 2.473 ;
      RECT 37.955 2.243 38.165 2.463 ;
      RECT 37.95 2.248 38.17 2.433 ;
      RECT 37.955 2.245 38.17 2.463 ;
      RECT 37.97 2.24 38.165 2.473 ;
      RECT 37.99 2.237 38.155 2.51 ;
      RECT 37.99 2.236 38.145 2.51 ;
      RECT 38.015 2.235 38.145 2.51 ;
      RECT 37.575 2.48 37.835 2.74 ;
      RECT 37.45 2.525 37.835 2.735 ;
      RECT 37.44 2.53 37.835 2.73 ;
      RECT 37.455 3.47 37.47 3.78 ;
      RECT 36.05 3.24 36.06 3.37 ;
      RECT 35.83 3.235 35.935 3.37 ;
      RECT 35.745 3.24 35.795 3.37 ;
      RECT 34.295 1.975 34.3 3.08 ;
      RECT 37.55 3.562 37.555 3.698 ;
      RECT 37.545 3.557 37.55 3.758 ;
      RECT 37.54 3.555 37.545 3.771 ;
      RECT 37.525 3.552 37.54 3.773 ;
      RECT 37.52 3.547 37.525 3.775 ;
      RECT 37.515 3.543 37.52 3.778 ;
      RECT 37.5 3.538 37.515 3.78 ;
      RECT 37.47 3.53 37.5 3.78 ;
      RECT 37.431 3.47 37.455 3.78 ;
      RECT 37.345 3.47 37.431 3.777 ;
      RECT 37.315 3.47 37.345 3.77 ;
      RECT 37.29 3.47 37.315 3.763 ;
      RECT 37.265 3.47 37.29 3.755 ;
      RECT 37.25 3.47 37.265 3.748 ;
      RECT 37.225 3.47 37.25 3.74 ;
      RECT 37.21 3.47 37.225 3.733 ;
      RECT 37.17 3.48 37.21 3.722 ;
      RECT 37.16 3.475 37.17 3.712 ;
      RECT 37.156 3.474 37.16 3.709 ;
      RECT 37.07 3.466 37.156 3.692 ;
      RECT 37.037 3.455 37.07 3.669 ;
      RECT 36.951 3.444 37.037 3.647 ;
      RECT 36.865 3.428 36.951 3.616 ;
      RECT 36.795 3.413 36.865 3.588 ;
      RECT 36.785 3.406 36.795 3.575 ;
      RECT 36.755 3.403 36.785 3.565 ;
      RECT 36.73 3.399 36.755 3.558 ;
      RECT 36.715 3.396 36.73 3.553 ;
      RECT 36.71 3.395 36.715 3.548 ;
      RECT 36.68 3.39 36.71 3.541 ;
      RECT 36.675 3.385 36.68 3.536 ;
      RECT 36.66 3.382 36.675 3.531 ;
      RECT 36.655 3.377 36.66 3.526 ;
      RECT 36.635 3.372 36.655 3.523 ;
      RECT 36.62 3.367 36.635 3.515 ;
      RECT 36.605 3.361 36.62 3.51 ;
      RECT 36.575 3.352 36.605 3.503 ;
      RECT 36.57 3.345 36.575 3.495 ;
      RECT 36.565 3.343 36.57 3.493 ;
      RECT 36.56 3.342 36.565 3.49 ;
      RECT 36.52 3.335 36.56 3.483 ;
      RECT 36.506 3.325 36.52 3.473 ;
      RECT 36.455 3.314 36.506 3.461 ;
      RECT 36.43 3.3 36.455 3.447 ;
      RECT 36.405 3.289 36.43 3.439 ;
      RECT 36.385 3.278 36.405 3.433 ;
      RECT 36.375 3.272 36.385 3.428 ;
      RECT 36.37 3.27 36.375 3.424 ;
      RECT 36.35 3.265 36.37 3.419 ;
      RECT 36.32 3.255 36.35 3.409 ;
      RECT 36.315 3.247 36.32 3.402 ;
      RECT 36.3 3.245 36.315 3.398 ;
      RECT 36.28 3.245 36.3 3.393 ;
      RECT 36.275 3.244 36.28 3.391 ;
      RECT 36.27 3.244 36.275 3.388 ;
      RECT 36.23 3.243 36.27 3.383 ;
      RECT 36.205 3.242 36.23 3.378 ;
      RECT 36.145 3.241 36.205 3.375 ;
      RECT 36.06 3.24 36.145 3.373 ;
      RECT 36.021 3.239 36.05 3.37 ;
      RECT 35.935 3.237 36.021 3.37 ;
      RECT 35.795 3.237 35.83 3.37 ;
      RECT 35.705 3.241 35.745 3.373 ;
      RECT 35.69 3.244 35.705 3.38 ;
      RECT 35.68 3.245 35.69 3.387 ;
      RECT 35.655 3.248 35.68 3.392 ;
      RECT 35.65 3.25 35.655 3.395 ;
      RECT 35.6 3.252 35.65 3.396 ;
      RECT 35.561 3.256 35.6 3.398 ;
      RECT 35.475 3.258 35.561 3.401 ;
      RECT 35.457 3.26 35.475 3.403 ;
      RECT 35.371 3.263 35.457 3.405 ;
      RECT 35.285 3.267 35.371 3.408 ;
      RECT 35.248 3.271 35.285 3.411 ;
      RECT 35.162 3.274 35.248 3.414 ;
      RECT 35.076 3.278 35.162 3.417 ;
      RECT 34.99 3.283 35.076 3.421 ;
      RECT 34.97 3.285 34.99 3.424 ;
      RECT 34.95 3.284 34.97 3.425 ;
      RECT 34.901 3.281 34.95 3.426 ;
      RECT 34.815 3.276 34.901 3.429 ;
      RECT 34.765 3.271 34.815 3.431 ;
      RECT 34.741 3.269 34.765 3.432 ;
      RECT 34.655 3.264 34.741 3.434 ;
      RECT 34.63 3.26 34.655 3.433 ;
      RECT 34.62 3.257 34.63 3.431 ;
      RECT 34.61 3.25 34.62 3.428 ;
      RECT 34.605 3.23 34.61 3.423 ;
      RECT 34.595 3.2 34.605 3.418 ;
      RECT 34.58 3.07 34.595 3.409 ;
      RECT 34.575 3.062 34.58 3.402 ;
      RECT 34.555 3.055 34.575 3.394 ;
      RECT 34.55 3.037 34.555 3.386 ;
      RECT 34.54 3.017 34.55 3.381 ;
      RECT 34.535 2.99 34.54 3.377 ;
      RECT 34.53 2.967 34.535 3.374 ;
      RECT 34.51 2.925 34.53 3.366 ;
      RECT 34.475 2.84 34.51 3.35 ;
      RECT 34.47 2.772 34.475 3.338 ;
      RECT 34.455 2.742 34.47 3.332 ;
      RECT 34.45 1.987 34.455 2.233 ;
      RECT 34.44 2.712 34.455 3.323 ;
      RECT 34.445 1.982 34.45 2.265 ;
      RECT 34.44 1.977 34.445 2.308 ;
      RECT 34.435 1.975 34.44 2.343 ;
      RECT 34.42 2.675 34.44 3.313 ;
      RECT 34.43 1.975 34.435 2.38 ;
      RECT 34.415 1.975 34.43 2.478 ;
      RECT 34.415 2.648 34.42 3.306 ;
      RECT 34.41 1.975 34.415 2.553 ;
      RECT 34.41 2.636 34.415 3.303 ;
      RECT 34.405 1.975 34.41 2.585 ;
      RECT 34.405 2.615 34.41 3.3 ;
      RECT 34.4 1.975 34.405 3.297 ;
      RECT 34.365 1.975 34.4 3.283 ;
      RECT 34.35 1.975 34.365 3.265 ;
      RECT 34.33 1.975 34.35 3.255 ;
      RECT 34.305 1.975 34.33 3.238 ;
      RECT 34.3 1.975 34.305 3.188 ;
      RECT 34.29 1.975 34.295 3.018 ;
      RECT 34.285 1.975 34.29 2.925 ;
      RECT 34.28 1.975 34.285 2.838 ;
      RECT 34.275 1.975 34.28 2.77 ;
      RECT 34.27 1.975 34.275 2.713 ;
      RECT 34.26 1.975 34.27 2.608 ;
      RECT 34.255 1.975 34.26 2.48 ;
      RECT 34.25 1.975 34.255 2.398 ;
      RECT 34.245 1.977 34.25 2.315 ;
      RECT 34.24 1.982 34.245 2.248 ;
      RECT 34.235 1.987 34.24 2.175 ;
      RECT 37.05 2.305 37.31 2.565 ;
      RECT 37.07 2.272 37.28 2.565 ;
      RECT 37.07 2.27 37.27 2.565 ;
      RECT 37.08 2.257 37.27 2.565 ;
      RECT 37.08 2.255 37.195 2.565 ;
      RECT 36.555 2.38 36.73 2.66 ;
      RECT 36.55 2.38 36.73 2.658 ;
      RECT 36.55 2.38 36.745 2.655 ;
      RECT 36.54 2.38 36.745 2.653 ;
      RECT 36.485 2.38 36.745 2.64 ;
      RECT 36.485 2.455 36.75 2.618 ;
      RECT 36.03 2.392 36.05 2.635 ;
      RECT 36.03 2.392 36.09 2.634 ;
      RECT 36.025 2.394 36.09 2.633 ;
      RECT 36.025 2.394 36.176 2.632 ;
      RECT 36.025 2.394 36.245 2.631 ;
      RECT 36.025 2.394 36.265 2.623 ;
      RECT 36.005 2.397 36.265 2.621 ;
      RECT 35.99 2.407 36.265 2.606 ;
      RECT 35.99 2.407 36.28 2.605 ;
      RECT 35.985 2.416 36.28 2.597 ;
      RECT 35.985 2.416 36.285 2.593 ;
      RECT 36.09 2.33 36.35 2.59 ;
      RECT 35.98 2.418 36.35 2.475 ;
      RECT 36.05 2.385 36.35 2.59 ;
      RECT 36.015 3.578 36.02 3.785 ;
      RECT 35.965 3.572 36.015 3.784 ;
      RECT 35.932 3.586 36.025 3.783 ;
      RECT 35.846 3.586 36.025 3.782 ;
      RECT 35.76 3.586 36.025 3.781 ;
      RECT 35.76 3.685 36.03 3.778 ;
      RECT 35.755 3.685 36.03 3.773 ;
      RECT 35.75 3.685 36.03 3.755 ;
      RECT 35.745 3.685 36.03 3.738 ;
      RECT 35.705 3.47 35.965 3.73 ;
      RECT 35.165 2.62 35.251 3.034 ;
      RECT 35.165 2.62 35.29 3.031 ;
      RECT 35.165 2.62 35.31 3.021 ;
      RECT 35.12 2.62 35.31 3.018 ;
      RECT 35.12 2.772 35.32 3.008 ;
      RECT 35.12 2.793 35.325 3.002 ;
      RECT 35.12 2.811 35.33 2.998 ;
      RECT 35.12 2.831 35.34 2.993 ;
      RECT 35.095 2.831 35.34 2.99 ;
      RECT 35.085 2.831 35.34 2.968 ;
      RECT 35.085 2.847 35.345 2.938 ;
      RECT 35.05 2.62 35.31 2.925 ;
      RECT 35.05 2.859 35.35 2.88 ;
      RECT 32.71 7.77 33 8 ;
      RECT 32.77 6.29 32.94 8 ;
      RECT 32.76 6.66 33.115 7.015 ;
      RECT 32.71 6.29 33 6.52 ;
      RECT 32.305 2.395 32.41 2.965 ;
      RECT 32.305 2.73 32.63 2.96 ;
      RECT 32.305 2.76 32.8 2.93 ;
      RECT 32.305 2.395 32.495 2.96 ;
      RECT 31.72 2.36 32.01 2.59 ;
      RECT 31.72 2.395 32.495 2.565 ;
      RECT 31.78 0.88 31.95 2.59 ;
      RECT 31.72 0.88 32.01 1.11 ;
      RECT 31.72 7.77 32.01 8 ;
      RECT 31.78 6.29 31.95 8 ;
      RECT 31.72 6.29 32.01 6.52 ;
      RECT 31.72 6.325 32.575 6.485 ;
      RECT 32.405 5.92 32.575 6.485 ;
      RECT 31.72 6.32 32.115 6.485 ;
      RECT 32.34 5.92 32.63 6.15 ;
      RECT 32.34 5.95 32.8 6.12 ;
      RECT 31.35 2.73 31.64 2.96 ;
      RECT 31.35 2.76 31.81 2.93 ;
      RECT 31.415 1.655 31.58 2.96 ;
      RECT 29.93 1.625 30.22 1.855 ;
      RECT 29.93 1.655 31.58 1.825 ;
      RECT 29.99 0.885 30.16 1.855 ;
      RECT 29.93 0.885 30.22 1.115 ;
      RECT 29.93 7.765 30.22 7.995 ;
      RECT 29.99 7.025 30.16 7.995 ;
      RECT 29.99 7.12 31.58 7.29 ;
      RECT 31.41 5.92 31.58 7.29 ;
      RECT 29.93 7.025 30.22 7.255 ;
      RECT 31.35 5.92 31.64 6.15 ;
      RECT 31.35 5.95 31.81 6.12 ;
      RECT 27.98 2.705 28.32 3.055 ;
      RECT 28.07 2.025 28.24 3.055 ;
      RECT 30.36 1.965 30.71 2.315 ;
      RECT 28.07 2.025 30.71 2.195 ;
      RECT 30.385 6.655 30.71 6.98 ;
      RECT 24.925 6.61 25.275 6.96 ;
      RECT 30.36 6.655 30.71 6.885 ;
      RECT 24.725 6.655 25.275 6.885 ;
      RECT 24.555 6.685 30.71 6.855 ;
      RECT 29.585 2.365 29.905 2.685 ;
      RECT 29.555 2.365 29.905 2.595 ;
      RECT 29.385 2.395 29.905 2.565 ;
      RECT 29.585 6.255 29.905 6.545 ;
      RECT 29.555 6.285 29.905 6.515 ;
      RECT 29.385 6.315 29.905 6.485 ;
      RECT 25.275 2.985 25.425 3.26 ;
      RECT 25.815 2.065 25.82 2.285 ;
      RECT 26.965 2.265 26.98 2.463 ;
      RECT 26.93 2.257 26.965 2.47 ;
      RECT 26.9 2.25 26.93 2.47 ;
      RECT 26.845 2.215 26.9 2.47 ;
      RECT 26.78 2.152 26.845 2.47 ;
      RECT 26.775 2.117 26.78 2.468 ;
      RECT 26.77 2.112 26.775 2.46 ;
      RECT 26.765 2.107 26.77 2.446 ;
      RECT 26.76 2.104 26.765 2.439 ;
      RECT 26.715 2.094 26.76 2.39 ;
      RECT 26.695 2.081 26.715 2.325 ;
      RECT 26.69 2.076 26.695 2.298 ;
      RECT 26.685 2.075 26.69 2.291 ;
      RECT 26.68 2.074 26.685 2.284 ;
      RECT 26.595 2.059 26.68 2.23 ;
      RECT 26.565 2.04 26.595 2.18 ;
      RECT 26.485 2.023 26.565 2.165 ;
      RECT 26.45 2.01 26.485 2.15 ;
      RECT 26.442 2.01 26.45 2.145 ;
      RECT 26.356 2.011 26.442 2.145 ;
      RECT 26.27 2.013 26.356 2.145 ;
      RECT 26.245 2.014 26.27 2.149 ;
      RECT 26.17 2.02 26.245 2.164 ;
      RECT 26.087 2.032 26.17 2.188 ;
      RECT 26.001 2.045 26.087 2.214 ;
      RECT 25.915 2.058 26.001 2.24 ;
      RECT 25.88 2.067 25.915 2.259 ;
      RECT 25.83 2.067 25.88 2.272 ;
      RECT 25.82 2.065 25.83 2.283 ;
      RECT 25.805 2.062 25.815 2.285 ;
      RECT 25.79 2.054 25.805 2.293 ;
      RECT 25.775 2.046 25.79 2.313 ;
      RECT 25.77 2.041 25.775 2.37 ;
      RECT 25.755 2.036 25.77 2.443 ;
      RECT 25.75 2.031 25.755 2.485 ;
      RECT 25.745 2.029 25.75 2.513 ;
      RECT 25.74 2.027 25.745 2.535 ;
      RECT 25.73 2.023 25.74 2.578 ;
      RECT 25.725 2.02 25.73 2.603 ;
      RECT 25.72 2.018 25.725 2.623 ;
      RECT 25.715 2.016 25.72 2.647 ;
      RECT 25.71 2.012 25.715 2.67 ;
      RECT 25.705 2.008 25.71 2.693 ;
      RECT 25.67 1.998 25.705 2.8 ;
      RECT 25.665 1.988 25.67 2.898 ;
      RECT 25.66 1.986 25.665 2.925 ;
      RECT 25.655 1.985 25.66 2.945 ;
      RECT 25.65 1.977 25.655 2.965 ;
      RECT 25.645 1.972 25.65 3 ;
      RECT 25.64 1.97 25.645 3.018 ;
      RECT 25.635 1.97 25.64 3.043 ;
      RECT 25.63 1.97 25.635 3.065 ;
      RECT 25.595 1.97 25.63 3.108 ;
      RECT 25.57 1.97 25.595 3.137 ;
      RECT 25.56 1.97 25.57 2.323 ;
      RECT 25.563 2.38 25.57 3.147 ;
      RECT 25.56 2.437 25.563 3.15 ;
      RECT 25.555 1.97 25.56 2.295 ;
      RECT 25.555 2.487 25.56 3.153 ;
      RECT 25.545 1.97 25.555 2.285 ;
      RECT 25.55 2.54 25.555 3.156 ;
      RECT 25.545 2.625 25.55 3.16 ;
      RECT 25.535 1.97 25.545 2.273 ;
      RECT 25.54 2.672 25.545 3.164 ;
      RECT 25.535 2.747 25.54 3.168 ;
      RECT 25.5 1.97 25.535 2.248 ;
      RECT 25.525 2.83 25.535 3.173 ;
      RECT 25.515 2.897 25.525 3.18 ;
      RECT 25.51 2.925 25.515 3.185 ;
      RECT 25.5 2.938 25.51 3.191 ;
      RECT 25.455 1.97 25.5 2.205 ;
      RECT 25.495 2.943 25.5 3.198 ;
      RECT 25.455 2.96 25.495 3.26 ;
      RECT 25.45 1.972 25.455 2.178 ;
      RECT 25.425 2.98 25.455 3.26 ;
      RECT 25.445 1.977 25.45 2.15 ;
      RECT 25.235 2.989 25.275 3.26 ;
      RECT 25.21 2.997 25.235 3.23 ;
      RECT 25.165 3.005 25.21 3.23 ;
      RECT 25.15 3.01 25.165 3.225 ;
      RECT 25.14 3.01 25.15 3.219 ;
      RECT 25.13 3.017 25.14 3.216 ;
      RECT 25.125 3.055 25.13 3.205 ;
      RECT 25.12 3.117 25.125 3.183 ;
      RECT 26.39 2.992 26.575 3.215 ;
      RECT 26.39 3.007 26.58 3.211 ;
      RECT 26.38 2.28 26.465 3.21 ;
      RECT 26.38 3.007 26.585 3.204 ;
      RECT 26.375 3.015 26.585 3.203 ;
      RECT 26.58 2.735 26.9 3.055 ;
      RECT 26.375 2.907 26.545 2.998 ;
      RECT 26.37 2.907 26.545 2.98 ;
      RECT 26.36 2.715 26.495 2.955 ;
      RECT 26.355 2.715 26.495 2.9 ;
      RECT 26.315 2.295 26.485 2.8 ;
      RECT 26.3 2.295 26.485 2.67 ;
      RECT 26.295 2.295 26.485 2.623 ;
      RECT 26.29 2.295 26.485 2.603 ;
      RECT 26.285 2.295 26.485 2.578 ;
      RECT 26.255 2.295 26.515 2.555 ;
      RECT 26.265 2.292 26.475 2.555 ;
      RECT 26.39 2.287 26.475 3.215 ;
      RECT 26.275 2.28 26.465 2.555 ;
      RECT 26.27 2.285 26.465 2.555 ;
      RECT 25.1 2.497 25.285 2.71 ;
      RECT 25.1 2.505 25.295 2.703 ;
      RECT 25.08 2.505 25.295 2.7 ;
      RECT 25.075 2.505 25.295 2.685 ;
      RECT 25.005 2.42 25.265 2.68 ;
      RECT 25.005 2.565 25.3 2.593 ;
      RECT 24.66 3.02 24.92 3.28 ;
      RECT 24.685 2.965 24.88 3.28 ;
      RECT 24.68 2.714 24.86 3.008 ;
      RECT 24.68 2.72 24.87 3.008 ;
      RECT 24.66 2.722 24.87 2.953 ;
      RECT 24.655 2.732 24.87 2.82 ;
      RECT 24.685 2.712 24.86 3.28 ;
      RECT 24.771 2.71 24.86 3.28 ;
      RECT 24.63 1.93 24.665 2.3 ;
      RECT 24.42 2.04 24.425 2.3 ;
      RECT 24.665 1.937 24.68 2.3 ;
      RECT 24.555 1.93 24.63 2.378 ;
      RECT 24.545 1.93 24.555 2.463 ;
      RECT 24.52 1.93 24.545 2.498 ;
      RECT 24.48 1.93 24.52 2.566 ;
      RECT 24.47 1.937 24.48 2.618 ;
      RECT 24.44 2.04 24.47 2.659 ;
      RECT 24.435 2.04 24.44 2.698 ;
      RECT 24.425 2.04 24.435 2.718 ;
      RECT 24.42 2.335 24.425 2.755 ;
      RECT 24.415 2.352 24.42 2.775 ;
      RECT 24.4 2.415 24.415 2.815 ;
      RECT 24.395 2.458 24.4 2.85 ;
      RECT 24.39 2.466 24.395 2.863 ;
      RECT 24.38 2.48 24.39 2.885 ;
      RECT 24.355 2.515 24.38 2.95 ;
      RECT 24.345 2.55 24.355 3.013 ;
      RECT 24.325 2.58 24.345 3.074 ;
      RECT 24.31 2.616 24.325 3.141 ;
      RECT 24.3 2.644 24.31 3.18 ;
      RECT 24.29 2.666 24.3 3.2 ;
      RECT 24.285 2.676 24.29 3.211 ;
      RECT 24.28 2.685 24.285 3.214 ;
      RECT 24.27 2.703 24.28 3.218 ;
      RECT 24.26 2.721 24.27 3.219 ;
      RECT 24.235 2.76 24.26 3.216 ;
      RECT 24.215 2.802 24.235 3.213 ;
      RECT 24.2 2.84 24.215 3.212 ;
      RECT 24.165 2.875 24.2 3.209 ;
      RECT 24.16 2.897 24.165 3.207 ;
      RECT 24.095 2.937 24.16 3.204 ;
      RECT 24.09 2.977 24.095 3.2 ;
      RECT 24.075 2.987 24.09 3.191 ;
      RECT 24.065 3.107 24.075 3.176 ;
      RECT 24.545 3.52 24.555 3.78 ;
      RECT 24.545 3.523 24.565 3.779 ;
      RECT 24.535 3.513 24.545 3.778 ;
      RECT 24.525 3.528 24.605 3.774 ;
      RECT 24.51 3.507 24.525 3.772 ;
      RECT 24.485 3.532 24.61 3.768 ;
      RECT 24.47 3.492 24.485 3.763 ;
      RECT 24.47 3.534 24.62 3.762 ;
      RECT 24.47 3.542 24.635 3.755 ;
      RECT 24.41 3.479 24.47 3.745 ;
      RECT 24.4 3.466 24.41 3.727 ;
      RECT 24.375 3.456 24.4 3.717 ;
      RECT 24.37 3.446 24.375 3.709 ;
      RECT 24.305 3.542 24.635 3.691 ;
      RECT 24.22 3.542 24.635 3.653 ;
      RECT 24.11 3.37 24.37 3.63 ;
      RECT 24.485 3.5 24.51 3.768 ;
      RECT 24.525 3.51 24.535 3.774 ;
      RECT 24.11 3.518 24.55 3.63 ;
      RECT 24.295 7.765 24.585 7.995 ;
      RECT 24.355 7.025 24.525 7.995 ;
      RECT 24.255 7.055 24.625 7.425 ;
      RECT 24.295 7.025 24.585 7.425 ;
      RECT 23.325 3.275 23.355 3.575 ;
      RECT 23.1 3.26 23.105 3.535 ;
      RECT 22.9 3.26 23.055 3.52 ;
      RECT 24.2 1.975 24.23 2.235 ;
      RECT 24.19 1.975 24.2 2.343 ;
      RECT 24.17 1.975 24.19 2.353 ;
      RECT 24.155 1.975 24.17 2.365 ;
      RECT 24.1 1.975 24.155 2.415 ;
      RECT 24.085 1.975 24.1 2.463 ;
      RECT 24.055 1.975 24.085 2.498 ;
      RECT 24 1.975 24.055 2.56 ;
      RECT 23.98 1.975 24 2.628 ;
      RECT 23.975 1.975 23.98 2.658 ;
      RECT 23.97 1.975 23.975 2.67 ;
      RECT 23.965 2.092 23.97 2.688 ;
      RECT 23.945 2.11 23.965 2.713 ;
      RECT 23.925 2.137 23.945 2.763 ;
      RECT 23.92 2.157 23.925 2.794 ;
      RECT 23.915 2.165 23.92 2.811 ;
      RECT 23.9 2.191 23.915 2.84 ;
      RECT 23.885 2.233 23.9 2.875 ;
      RECT 23.88 2.262 23.885 2.898 ;
      RECT 23.875 2.277 23.88 2.911 ;
      RECT 23.87 2.3 23.875 2.922 ;
      RECT 23.86 2.32 23.87 2.94 ;
      RECT 23.85 2.35 23.86 2.963 ;
      RECT 23.845 2.372 23.85 2.983 ;
      RECT 23.84 2.387 23.845 2.998 ;
      RECT 23.825 2.417 23.84 3.025 ;
      RECT 23.82 2.447 23.825 3.051 ;
      RECT 23.815 2.465 23.82 3.063 ;
      RECT 23.805 2.495 23.815 3.082 ;
      RECT 23.795 2.52 23.805 3.107 ;
      RECT 23.79 2.54 23.795 3.126 ;
      RECT 23.785 2.557 23.79 3.139 ;
      RECT 23.775 2.583 23.785 3.158 ;
      RECT 23.765 2.621 23.775 3.185 ;
      RECT 23.76 2.647 23.765 3.205 ;
      RECT 23.755 2.657 23.76 3.215 ;
      RECT 23.75 2.67 23.755 3.23 ;
      RECT 23.745 2.685 23.75 3.24 ;
      RECT 23.74 2.707 23.745 3.255 ;
      RECT 23.735 2.725 23.74 3.266 ;
      RECT 23.73 2.735 23.735 3.277 ;
      RECT 23.725 2.743 23.73 3.289 ;
      RECT 23.72 2.751 23.725 3.3 ;
      RECT 23.715 2.777 23.72 3.313 ;
      RECT 23.705 2.805 23.715 3.326 ;
      RECT 23.7 2.835 23.705 3.335 ;
      RECT 23.695 2.85 23.7 3.342 ;
      RECT 23.68 2.875 23.695 3.349 ;
      RECT 23.675 2.897 23.68 3.355 ;
      RECT 23.67 2.922 23.675 3.358 ;
      RECT 23.661 2.95 23.67 3.362 ;
      RECT 23.655 2.967 23.661 3.367 ;
      RECT 23.65 2.985 23.655 3.371 ;
      RECT 23.645 2.997 23.65 3.374 ;
      RECT 23.64 3.018 23.645 3.378 ;
      RECT 23.635 3.036 23.64 3.381 ;
      RECT 23.63 3.05 23.635 3.384 ;
      RECT 23.625 3.067 23.63 3.387 ;
      RECT 23.62 3.08 23.625 3.39 ;
      RECT 23.595 3.117 23.62 3.398 ;
      RECT 23.59 3.162 23.595 3.407 ;
      RECT 23.585 3.19 23.59 3.41 ;
      RECT 23.575 3.21 23.585 3.414 ;
      RECT 23.57 3.23 23.575 3.419 ;
      RECT 23.565 3.245 23.57 3.422 ;
      RECT 23.545 3.255 23.565 3.429 ;
      RECT 23.48 3.262 23.545 3.455 ;
      RECT 23.445 3.265 23.48 3.483 ;
      RECT 23.43 3.268 23.445 3.498 ;
      RECT 23.42 3.269 23.43 3.513 ;
      RECT 23.41 3.27 23.42 3.53 ;
      RECT 23.405 3.27 23.41 3.545 ;
      RECT 23.4 3.27 23.405 3.553 ;
      RECT 23.385 3.271 23.4 3.568 ;
      RECT 23.355 3.273 23.385 3.575 ;
      RECT 23.245 3.28 23.325 3.575 ;
      RECT 23.2 3.285 23.245 3.575 ;
      RECT 23.19 3.286 23.2 3.565 ;
      RECT 23.18 3.287 23.19 3.558 ;
      RECT 23.16 3.289 23.18 3.553 ;
      RECT 23.15 3.26 23.16 3.548 ;
      RECT 23.105 3.26 23.15 3.54 ;
      RECT 23.075 3.26 23.1 3.53 ;
      RECT 23.055 3.26 23.075 3.523 ;
      RECT 23.335 2.06 23.595 2.32 ;
      RECT 23.215 2.075 23.225 2.24 ;
      RECT 23.2 2.075 23.205 2.235 ;
      RECT 20.565 1.915 20.75 2.205 ;
      RECT 22.38 2.04 22.395 2.195 ;
      RECT 20.53 1.915 20.555 2.175 ;
      RECT 22.945 1.965 22.95 2.107 ;
      RECT 22.86 1.96 22.885 2.1 ;
      RECT 23.26 2.077 23.335 2.27 ;
      RECT 23.245 2.075 23.26 2.253 ;
      RECT 23.225 2.075 23.245 2.245 ;
      RECT 23.205 2.075 23.215 2.238 ;
      RECT 23.16 2.07 23.2 2.228 ;
      RECT 23.12 2.045 23.16 2.213 ;
      RECT 23.105 2.02 23.12 2.203 ;
      RECT 23.1 2.014 23.105 2.201 ;
      RECT 23.065 2.006 23.1 2.184 ;
      RECT 23.06 1.999 23.065 2.172 ;
      RECT 23.04 1.994 23.06 2.16 ;
      RECT 23.03 1.988 23.04 2.145 ;
      RECT 23.01 1.983 23.03 2.13 ;
      RECT 23 1.978 23.01 2.123 ;
      RECT 22.995 1.976 23 2.118 ;
      RECT 22.99 1.975 22.995 2.115 ;
      RECT 22.95 1.97 22.99 2.111 ;
      RECT 22.93 1.964 22.945 2.106 ;
      RECT 22.895 1.961 22.93 2.103 ;
      RECT 22.885 1.96 22.895 2.101 ;
      RECT 22.825 1.96 22.86 2.098 ;
      RECT 22.78 1.96 22.825 2.098 ;
      RECT 22.73 1.96 22.78 2.101 ;
      RECT 22.715 1.962 22.73 2.103 ;
      RECT 22.7 1.965 22.715 2.104 ;
      RECT 22.69 1.97 22.7 2.105 ;
      RECT 22.66 1.975 22.69 2.11 ;
      RECT 22.65 1.981 22.66 2.118 ;
      RECT 22.64 1.983 22.65 2.122 ;
      RECT 22.63 1.987 22.64 2.126 ;
      RECT 22.605 1.993 22.63 2.134 ;
      RECT 22.595 1.998 22.605 2.142 ;
      RECT 22.58 2.002 22.595 2.146 ;
      RECT 22.545 2.008 22.58 2.154 ;
      RECT 22.525 2.013 22.545 2.164 ;
      RECT 22.495 2.02 22.525 2.173 ;
      RECT 22.45 2.029 22.495 2.187 ;
      RECT 22.445 2.034 22.45 2.198 ;
      RECT 22.425 2.037 22.445 2.199 ;
      RECT 22.395 2.04 22.425 2.197 ;
      RECT 22.36 2.04 22.38 2.193 ;
      RECT 22.29 2.04 22.36 2.184 ;
      RECT 22.275 2.037 22.29 2.176 ;
      RECT 22.235 2.03 22.275 2.171 ;
      RECT 22.21 2.02 22.235 2.164 ;
      RECT 22.205 2.014 22.21 2.161 ;
      RECT 22.165 2.008 22.205 2.158 ;
      RECT 22.15 2.001 22.165 2.153 ;
      RECT 22.13 1.997 22.15 2.148 ;
      RECT 22.115 1.992 22.13 2.144 ;
      RECT 22.1 1.987 22.115 2.142 ;
      RECT 22.085 1.983 22.1 2.141 ;
      RECT 22.07 1.981 22.085 2.137 ;
      RECT 22.06 1.979 22.07 2.132 ;
      RECT 22.045 1.976 22.06 2.128 ;
      RECT 22.035 1.974 22.045 2.123 ;
      RECT 22.015 1.971 22.035 2.119 ;
      RECT 21.97 1.97 22.015 2.117 ;
      RECT 21.91 1.972 21.97 2.118 ;
      RECT 21.89 1.974 21.91 2.12 ;
      RECT 21.86 1.977 21.89 2.121 ;
      RECT 21.81 1.982 21.86 2.123 ;
      RECT 21.805 1.985 21.81 2.125 ;
      RECT 21.795 1.987 21.805 2.128 ;
      RECT 21.79 1.989 21.795 2.131 ;
      RECT 21.74 1.992 21.79 2.138 ;
      RECT 21.72 1.996 21.74 2.15 ;
      RECT 21.71 1.999 21.72 2.156 ;
      RECT 21.7 2 21.71 2.159 ;
      RECT 21.661 2.003 21.7 2.161 ;
      RECT 21.575 2.01 21.661 2.164 ;
      RECT 21.501 2.02 21.575 2.168 ;
      RECT 21.415 2.031 21.501 2.173 ;
      RECT 21.4 2.038 21.415 2.175 ;
      RECT 21.345 2.042 21.4 2.176 ;
      RECT 21.331 2.045 21.345 2.178 ;
      RECT 21.245 2.045 21.331 2.18 ;
      RECT 21.205 2.042 21.245 2.183 ;
      RECT 21.181 2.038 21.205 2.185 ;
      RECT 21.095 2.028 21.181 2.188 ;
      RECT 21.065 2.017 21.095 2.189 ;
      RECT 21.046 2.013 21.065 2.188 ;
      RECT 20.96 2.006 21.046 2.185 ;
      RECT 20.9 1.995 20.96 2.182 ;
      RECT 20.88 1.987 20.9 2.18 ;
      RECT 20.845 1.982 20.88 2.179 ;
      RECT 20.82 1.977 20.845 2.178 ;
      RECT 20.79 1.972 20.82 2.177 ;
      RECT 20.765 1.915 20.79 2.176 ;
      RECT 20.75 1.915 20.765 2.2 ;
      RECT 20.555 1.915 20.565 2.2 ;
      RECT 22.33 2.935 22.335 3.075 ;
      RECT 21.99 2.935 22.025 3.073 ;
      RECT 21.565 2.92 21.58 3.065 ;
      RECT 23.395 2.7 23.485 2.96 ;
      RECT 23.225 2.565 23.325 2.96 ;
      RECT 20.26 2.54 20.34 2.75 ;
      RECT 23.35 2.677 23.395 2.96 ;
      RECT 23.34 2.647 23.35 2.96 ;
      RECT 23.325 2.57 23.34 2.96 ;
      RECT 23.14 2.565 23.225 2.925 ;
      RECT 23.135 2.567 23.14 2.92 ;
      RECT 23.13 2.572 23.135 2.92 ;
      RECT 23.095 2.672 23.13 2.92 ;
      RECT 23.085 2.7 23.095 2.92 ;
      RECT 23.075 2.715 23.085 2.92 ;
      RECT 23.065 2.727 23.075 2.92 ;
      RECT 23.06 2.737 23.065 2.92 ;
      RECT 23.045 2.747 23.06 2.922 ;
      RECT 23.04 2.762 23.045 2.924 ;
      RECT 23.025 2.775 23.04 2.926 ;
      RECT 23.02 2.79 23.025 2.929 ;
      RECT 23 2.8 23.02 2.933 ;
      RECT 22.985 2.81 23 2.936 ;
      RECT 22.95 2.817 22.985 2.941 ;
      RECT 22.906 2.824 22.95 2.949 ;
      RECT 22.82 2.836 22.906 2.962 ;
      RECT 22.795 2.847 22.82 2.973 ;
      RECT 22.765 2.852 22.795 2.978 ;
      RECT 22.73 2.857 22.765 2.986 ;
      RECT 22.7 2.862 22.73 2.993 ;
      RECT 22.675 2.867 22.7 2.998 ;
      RECT 22.61 2.874 22.675 3.007 ;
      RECT 22.54 2.887 22.61 3.023 ;
      RECT 22.51 2.897 22.54 3.035 ;
      RECT 22.485 2.902 22.51 3.042 ;
      RECT 22.43 2.909 22.485 3.05 ;
      RECT 22.425 2.916 22.43 3.055 ;
      RECT 22.42 2.918 22.425 3.056 ;
      RECT 22.405 2.92 22.42 3.058 ;
      RECT 22.4 2.92 22.405 3.061 ;
      RECT 22.335 2.927 22.4 3.068 ;
      RECT 22.3 2.937 22.33 3.078 ;
      RECT 22.283 2.94 22.3 3.08 ;
      RECT 22.197 2.939 22.283 3.079 ;
      RECT 22.111 2.937 22.197 3.076 ;
      RECT 22.025 2.936 22.111 3.074 ;
      RECT 21.924 2.934 21.99 3.073 ;
      RECT 21.838 2.931 21.924 3.071 ;
      RECT 21.752 2.927 21.838 3.069 ;
      RECT 21.666 2.924 21.752 3.068 ;
      RECT 21.58 2.921 21.666 3.066 ;
      RECT 21.48 2.92 21.565 3.063 ;
      RECT 21.43 2.918 21.48 3.061 ;
      RECT 21.41 2.915 21.43 3.059 ;
      RECT 21.39 2.913 21.41 3.056 ;
      RECT 21.365 2.909 21.39 3.053 ;
      RECT 21.32 2.903 21.365 3.048 ;
      RECT 21.28 2.897 21.32 3.04 ;
      RECT 21.255 2.892 21.28 3.033 ;
      RECT 21.2 2.885 21.255 3.025 ;
      RECT 21.176 2.878 21.2 3.018 ;
      RECT 21.09 2.869 21.176 3.008 ;
      RECT 21.06 2.861 21.09 2.998 ;
      RECT 21.03 2.857 21.06 2.993 ;
      RECT 21.025 2.854 21.03 2.99 ;
      RECT 21.02 2.853 21.025 2.99 ;
      RECT 20.945 2.846 21.02 2.983 ;
      RECT 20.906 2.837 20.945 2.972 ;
      RECT 20.82 2.827 20.906 2.96 ;
      RECT 20.78 2.817 20.82 2.948 ;
      RECT 20.741 2.812 20.78 2.941 ;
      RECT 20.655 2.802 20.741 2.93 ;
      RECT 20.615 2.79 20.655 2.919 ;
      RECT 20.58 2.775 20.615 2.912 ;
      RECT 20.57 2.765 20.58 2.909 ;
      RECT 20.55 2.75 20.57 2.907 ;
      RECT 20.52 2.72 20.55 2.903 ;
      RECT 20.51 2.7 20.52 2.898 ;
      RECT 20.505 2.692 20.51 2.895 ;
      RECT 20.5 2.685 20.505 2.893 ;
      RECT 20.485 2.672 20.5 2.886 ;
      RECT 20.48 2.662 20.485 2.878 ;
      RECT 20.475 2.655 20.48 2.873 ;
      RECT 20.47 2.65 20.475 2.869 ;
      RECT 20.455 2.637 20.47 2.861 ;
      RECT 20.45 2.547 20.455 2.85 ;
      RECT 20.445 2.542 20.45 2.843 ;
      RECT 20.37 2.54 20.445 2.803 ;
      RECT 20.34 2.54 20.37 2.758 ;
      RECT 20.245 2.545 20.26 2.745 ;
      RECT 22.73 2.25 22.99 2.51 ;
      RECT 22.715 2.238 22.895 2.475 ;
      RECT 22.71 2.239 22.895 2.473 ;
      RECT 22.695 2.243 22.905 2.463 ;
      RECT 22.69 2.248 22.91 2.433 ;
      RECT 22.695 2.245 22.91 2.463 ;
      RECT 22.71 2.24 22.905 2.473 ;
      RECT 22.73 2.237 22.895 2.51 ;
      RECT 22.73 2.236 22.885 2.51 ;
      RECT 22.755 2.235 22.885 2.51 ;
      RECT 22.315 2.48 22.575 2.74 ;
      RECT 22.19 2.525 22.575 2.735 ;
      RECT 22.18 2.53 22.575 2.73 ;
      RECT 22.195 3.47 22.21 3.78 ;
      RECT 20.79 3.24 20.8 3.37 ;
      RECT 20.57 3.235 20.675 3.37 ;
      RECT 20.485 3.24 20.535 3.37 ;
      RECT 19.035 1.975 19.04 3.08 ;
      RECT 22.29 3.562 22.295 3.698 ;
      RECT 22.285 3.557 22.29 3.758 ;
      RECT 22.28 3.555 22.285 3.771 ;
      RECT 22.265 3.552 22.28 3.773 ;
      RECT 22.26 3.547 22.265 3.775 ;
      RECT 22.255 3.543 22.26 3.778 ;
      RECT 22.24 3.538 22.255 3.78 ;
      RECT 22.21 3.53 22.24 3.78 ;
      RECT 22.171 3.47 22.195 3.78 ;
      RECT 22.085 3.47 22.171 3.777 ;
      RECT 22.055 3.47 22.085 3.77 ;
      RECT 22.03 3.47 22.055 3.763 ;
      RECT 22.005 3.47 22.03 3.755 ;
      RECT 21.99 3.47 22.005 3.748 ;
      RECT 21.965 3.47 21.99 3.74 ;
      RECT 21.95 3.47 21.965 3.733 ;
      RECT 21.91 3.48 21.95 3.722 ;
      RECT 21.9 3.475 21.91 3.712 ;
      RECT 21.896 3.474 21.9 3.709 ;
      RECT 21.81 3.466 21.896 3.692 ;
      RECT 21.777 3.455 21.81 3.669 ;
      RECT 21.691 3.444 21.777 3.647 ;
      RECT 21.605 3.428 21.691 3.616 ;
      RECT 21.535 3.413 21.605 3.588 ;
      RECT 21.525 3.406 21.535 3.575 ;
      RECT 21.495 3.403 21.525 3.565 ;
      RECT 21.47 3.399 21.495 3.558 ;
      RECT 21.455 3.396 21.47 3.553 ;
      RECT 21.45 3.395 21.455 3.548 ;
      RECT 21.42 3.39 21.45 3.541 ;
      RECT 21.415 3.385 21.42 3.536 ;
      RECT 21.4 3.382 21.415 3.531 ;
      RECT 21.395 3.377 21.4 3.526 ;
      RECT 21.375 3.372 21.395 3.523 ;
      RECT 21.36 3.367 21.375 3.515 ;
      RECT 21.345 3.361 21.36 3.51 ;
      RECT 21.315 3.352 21.345 3.503 ;
      RECT 21.31 3.345 21.315 3.495 ;
      RECT 21.305 3.343 21.31 3.493 ;
      RECT 21.3 3.342 21.305 3.49 ;
      RECT 21.26 3.335 21.3 3.483 ;
      RECT 21.246 3.325 21.26 3.473 ;
      RECT 21.195 3.314 21.246 3.461 ;
      RECT 21.17 3.3 21.195 3.447 ;
      RECT 21.145 3.289 21.17 3.439 ;
      RECT 21.125 3.278 21.145 3.433 ;
      RECT 21.115 3.272 21.125 3.428 ;
      RECT 21.11 3.27 21.115 3.424 ;
      RECT 21.09 3.265 21.11 3.419 ;
      RECT 21.06 3.255 21.09 3.409 ;
      RECT 21.055 3.247 21.06 3.402 ;
      RECT 21.04 3.245 21.055 3.398 ;
      RECT 21.02 3.245 21.04 3.393 ;
      RECT 21.015 3.244 21.02 3.391 ;
      RECT 21.01 3.244 21.015 3.388 ;
      RECT 20.97 3.243 21.01 3.383 ;
      RECT 20.945 3.242 20.97 3.378 ;
      RECT 20.885 3.241 20.945 3.375 ;
      RECT 20.8 3.24 20.885 3.373 ;
      RECT 20.761 3.239 20.79 3.37 ;
      RECT 20.675 3.237 20.761 3.37 ;
      RECT 20.535 3.237 20.57 3.37 ;
      RECT 20.445 3.241 20.485 3.373 ;
      RECT 20.43 3.244 20.445 3.38 ;
      RECT 20.42 3.245 20.43 3.387 ;
      RECT 20.395 3.248 20.42 3.392 ;
      RECT 20.39 3.25 20.395 3.395 ;
      RECT 20.34 3.252 20.39 3.396 ;
      RECT 20.301 3.256 20.34 3.398 ;
      RECT 20.215 3.258 20.301 3.401 ;
      RECT 20.197 3.26 20.215 3.403 ;
      RECT 20.111 3.263 20.197 3.405 ;
      RECT 20.025 3.267 20.111 3.408 ;
      RECT 19.988 3.271 20.025 3.411 ;
      RECT 19.902 3.274 19.988 3.414 ;
      RECT 19.816 3.278 19.902 3.417 ;
      RECT 19.73 3.283 19.816 3.421 ;
      RECT 19.71 3.285 19.73 3.424 ;
      RECT 19.69 3.284 19.71 3.425 ;
      RECT 19.641 3.281 19.69 3.426 ;
      RECT 19.555 3.276 19.641 3.429 ;
      RECT 19.505 3.271 19.555 3.431 ;
      RECT 19.481 3.269 19.505 3.432 ;
      RECT 19.395 3.264 19.481 3.434 ;
      RECT 19.37 3.26 19.395 3.433 ;
      RECT 19.36 3.257 19.37 3.431 ;
      RECT 19.35 3.25 19.36 3.428 ;
      RECT 19.345 3.23 19.35 3.423 ;
      RECT 19.335 3.2 19.345 3.418 ;
      RECT 19.32 3.07 19.335 3.409 ;
      RECT 19.315 3.062 19.32 3.402 ;
      RECT 19.295 3.055 19.315 3.394 ;
      RECT 19.29 3.037 19.295 3.386 ;
      RECT 19.28 3.017 19.29 3.381 ;
      RECT 19.275 2.99 19.28 3.377 ;
      RECT 19.27 2.967 19.275 3.374 ;
      RECT 19.25 2.925 19.27 3.366 ;
      RECT 19.215 2.84 19.25 3.35 ;
      RECT 19.21 2.772 19.215 3.338 ;
      RECT 19.195 2.742 19.21 3.332 ;
      RECT 19.19 1.987 19.195 2.233 ;
      RECT 19.18 2.712 19.195 3.323 ;
      RECT 19.185 1.982 19.19 2.265 ;
      RECT 19.18 1.977 19.185 2.308 ;
      RECT 19.175 1.975 19.18 2.343 ;
      RECT 19.16 2.675 19.18 3.313 ;
      RECT 19.17 1.975 19.175 2.38 ;
      RECT 19.155 1.975 19.17 2.478 ;
      RECT 19.155 2.648 19.16 3.306 ;
      RECT 19.15 1.975 19.155 2.553 ;
      RECT 19.15 2.636 19.155 3.303 ;
      RECT 19.145 1.975 19.15 2.585 ;
      RECT 19.145 2.615 19.15 3.3 ;
      RECT 19.14 1.975 19.145 3.297 ;
      RECT 19.105 1.975 19.14 3.283 ;
      RECT 19.09 1.975 19.105 3.265 ;
      RECT 19.07 1.975 19.09 3.255 ;
      RECT 19.045 1.975 19.07 3.238 ;
      RECT 19.04 1.975 19.045 3.188 ;
      RECT 19.03 1.975 19.035 3.018 ;
      RECT 19.025 1.975 19.03 2.925 ;
      RECT 19.02 1.975 19.025 2.838 ;
      RECT 19.015 1.975 19.02 2.77 ;
      RECT 19.01 1.975 19.015 2.713 ;
      RECT 19 1.975 19.01 2.608 ;
      RECT 18.995 1.975 19 2.48 ;
      RECT 18.99 1.975 18.995 2.398 ;
      RECT 18.985 1.977 18.99 2.315 ;
      RECT 18.98 1.982 18.985 2.248 ;
      RECT 18.975 1.987 18.98 2.175 ;
      RECT 21.79 2.305 22.05 2.565 ;
      RECT 21.81 2.272 22.02 2.565 ;
      RECT 21.81 2.27 22.01 2.565 ;
      RECT 21.82 2.257 22.01 2.565 ;
      RECT 21.82 2.255 21.935 2.565 ;
      RECT 21.295 2.38 21.47 2.66 ;
      RECT 21.29 2.38 21.47 2.658 ;
      RECT 21.29 2.38 21.485 2.655 ;
      RECT 21.28 2.38 21.485 2.653 ;
      RECT 21.225 2.38 21.485 2.64 ;
      RECT 21.225 2.455 21.49 2.618 ;
      RECT 20.77 2.392 20.79 2.635 ;
      RECT 20.77 2.392 20.83 2.634 ;
      RECT 20.765 2.394 20.83 2.633 ;
      RECT 20.765 2.394 20.916 2.632 ;
      RECT 20.765 2.394 20.985 2.631 ;
      RECT 20.765 2.394 21.005 2.623 ;
      RECT 20.745 2.397 21.005 2.621 ;
      RECT 20.73 2.407 21.005 2.606 ;
      RECT 20.73 2.407 21.02 2.605 ;
      RECT 20.725 2.416 21.02 2.597 ;
      RECT 20.725 2.416 21.025 2.593 ;
      RECT 20.83 2.33 21.09 2.59 ;
      RECT 20.72 2.418 21.09 2.475 ;
      RECT 20.79 2.385 21.09 2.59 ;
      RECT 20.755 3.578 20.76 3.785 ;
      RECT 20.705 3.572 20.755 3.784 ;
      RECT 20.672 3.586 20.765 3.783 ;
      RECT 20.586 3.586 20.765 3.782 ;
      RECT 20.5 3.586 20.765 3.781 ;
      RECT 20.5 3.685 20.77 3.778 ;
      RECT 20.495 3.685 20.77 3.773 ;
      RECT 20.49 3.685 20.77 3.755 ;
      RECT 20.485 3.685 20.77 3.738 ;
      RECT 20.445 3.47 20.705 3.73 ;
      RECT 19.905 2.62 19.991 3.034 ;
      RECT 19.905 2.62 20.03 3.031 ;
      RECT 19.905 2.62 20.05 3.021 ;
      RECT 19.86 2.62 20.05 3.018 ;
      RECT 19.86 2.772 20.06 3.008 ;
      RECT 19.86 2.793 20.065 3.002 ;
      RECT 19.86 2.811 20.07 2.998 ;
      RECT 19.86 2.831 20.08 2.993 ;
      RECT 19.835 2.831 20.08 2.99 ;
      RECT 19.825 2.831 20.08 2.968 ;
      RECT 19.825 2.847 20.085 2.938 ;
      RECT 19.79 2.62 20.05 2.925 ;
      RECT 19.79 2.859 20.09 2.88 ;
      RECT 17.45 7.77 17.74 8 ;
      RECT 17.51 6.29 17.68 8 ;
      RECT 17.505 6.655 17.855 7.005 ;
      RECT 17.45 6.29 17.74 6.52 ;
      RECT 17.045 2.395 17.15 2.965 ;
      RECT 17.045 2.73 17.37 2.96 ;
      RECT 17.045 2.76 17.54 2.93 ;
      RECT 17.045 2.395 17.235 2.96 ;
      RECT 16.46 2.36 16.75 2.59 ;
      RECT 16.46 2.395 17.235 2.565 ;
      RECT 16.52 0.88 16.69 2.59 ;
      RECT 16.46 0.88 16.75 1.11 ;
      RECT 16.46 7.77 16.75 8 ;
      RECT 16.52 6.29 16.69 8 ;
      RECT 16.46 6.29 16.75 6.52 ;
      RECT 16.46 6.325 17.315 6.485 ;
      RECT 17.145 5.92 17.315 6.485 ;
      RECT 16.46 6.32 16.855 6.485 ;
      RECT 17.08 5.92 17.37 6.15 ;
      RECT 17.08 5.95 17.54 6.12 ;
      RECT 16.09 2.73 16.38 2.96 ;
      RECT 16.09 2.76 16.55 2.93 ;
      RECT 16.155 1.655 16.32 2.96 ;
      RECT 14.67 1.625 14.96 1.855 ;
      RECT 14.67 1.655 16.32 1.825 ;
      RECT 14.73 0.885 14.9 1.855 ;
      RECT 14.67 0.885 14.96 1.115 ;
      RECT 14.67 7.765 14.96 7.995 ;
      RECT 14.73 7.025 14.9 7.995 ;
      RECT 14.73 7.12 16.32 7.29 ;
      RECT 16.15 5.92 16.32 7.29 ;
      RECT 14.67 7.025 14.96 7.255 ;
      RECT 16.09 5.92 16.38 6.15 ;
      RECT 16.09 5.95 16.55 6.12 ;
      RECT 12.72 2.705 13.06 3.055 ;
      RECT 12.81 2.025 12.98 3.055 ;
      RECT 15.1 1.965 15.45 2.315 ;
      RECT 12.81 2.025 15.45 2.195 ;
      RECT 15.125 6.655 15.45 6.98 ;
      RECT 9.665 6.605 10.015 6.955 ;
      RECT 15.1 6.655 15.45 6.885 ;
      RECT 9.465 6.655 10.015 6.885 ;
      RECT 9.295 6.685 15.45 6.855 ;
      RECT 14.325 2.365 14.645 2.685 ;
      RECT 14.295 2.365 14.645 2.595 ;
      RECT 14.125 2.395 14.645 2.565 ;
      RECT 14.325 6.255 14.645 6.545 ;
      RECT 14.295 6.285 14.645 6.515 ;
      RECT 14.125 6.315 14.645 6.485 ;
      RECT 10.015 2.985 10.165 3.26 ;
      RECT 10.555 2.065 10.56 2.285 ;
      RECT 11.705 2.265 11.72 2.463 ;
      RECT 11.67 2.257 11.705 2.47 ;
      RECT 11.64 2.25 11.67 2.47 ;
      RECT 11.585 2.215 11.64 2.47 ;
      RECT 11.52 2.152 11.585 2.47 ;
      RECT 11.515 2.117 11.52 2.468 ;
      RECT 11.51 2.112 11.515 2.46 ;
      RECT 11.505 2.107 11.51 2.446 ;
      RECT 11.5 2.104 11.505 2.439 ;
      RECT 11.455 2.094 11.5 2.39 ;
      RECT 11.435 2.081 11.455 2.325 ;
      RECT 11.43 2.076 11.435 2.298 ;
      RECT 11.425 2.075 11.43 2.291 ;
      RECT 11.42 2.074 11.425 2.284 ;
      RECT 11.335 2.059 11.42 2.23 ;
      RECT 11.305 2.04 11.335 2.18 ;
      RECT 11.225 2.023 11.305 2.165 ;
      RECT 11.19 2.01 11.225 2.15 ;
      RECT 11.182 2.01 11.19 2.145 ;
      RECT 11.096 2.011 11.182 2.145 ;
      RECT 11.01 2.013 11.096 2.145 ;
      RECT 10.985 2.014 11.01 2.149 ;
      RECT 10.91 2.02 10.985 2.164 ;
      RECT 10.827 2.032 10.91 2.188 ;
      RECT 10.741 2.045 10.827 2.214 ;
      RECT 10.655 2.058 10.741 2.24 ;
      RECT 10.62 2.067 10.655 2.259 ;
      RECT 10.57 2.067 10.62 2.272 ;
      RECT 10.56 2.065 10.57 2.283 ;
      RECT 10.545 2.062 10.555 2.285 ;
      RECT 10.53 2.054 10.545 2.293 ;
      RECT 10.515 2.046 10.53 2.313 ;
      RECT 10.51 2.041 10.515 2.37 ;
      RECT 10.495 2.036 10.51 2.443 ;
      RECT 10.49 2.031 10.495 2.485 ;
      RECT 10.485 2.029 10.49 2.513 ;
      RECT 10.48 2.027 10.485 2.535 ;
      RECT 10.47 2.023 10.48 2.578 ;
      RECT 10.465 2.02 10.47 2.603 ;
      RECT 10.46 2.018 10.465 2.623 ;
      RECT 10.455 2.016 10.46 2.647 ;
      RECT 10.45 2.012 10.455 2.67 ;
      RECT 10.445 2.008 10.45 2.693 ;
      RECT 10.41 1.998 10.445 2.8 ;
      RECT 10.405 1.988 10.41 2.898 ;
      RECT 10.4 1.986 10.405 2.925 ;
      RECT 10.395 1.985 10.4 2.945 ;
      RECT 10.39 1.977 10.395 2.965 ;
      RECT 10.385 1.972 10.39 3 ;
      RECT 10.38 1.97 10.385 3.018 ;
      RECT 10.375 1.97 10.38 3.043 ;
      RECT 10.37 1.97 10.375 3.065 ;
      RECT 10.335 1.97 10.37 3.108 ;
      RECT 10.31 1.97 10.335 3.137 ;
      RECT 10.3 1.97 10.31 2.323 ;
      RECT 10.303 2.38 10.31 3.147 ;
      RECT 10.3 2.437 10.303 3.15 ;
      RECT 10.295 1.97 10.3 2.295 ;
      RECT 10.295 2.487 10.3 3.153 ;
      RECT 10.285 1.97 10.295 2.285 ;
      RECT 10.29 2.54 10.295 3.156 ;
      RECT 10.285 2.625 10.29 3.16 ;
      RECT 10.275 1.97 10.285 2.273 ;
      RECT 10.28 2.672 10.285 3.164 ;
      RECT 10.275 2.747 10.28 3.168 ;
      RECT 10.24 1.97 10.275 2.248 ;
      RECT 10.265 2.83 10.275 3.173 ;
      RECT 10.255 2.897 10.265 3.18 ;
      RECT 10.25 2.925 10.255 3.185 ;
      RECT 10.24 2.938 10.25 3.191 ;
      RECT 10.195 1.97 10.24 2.205 ;
      RECT 10.235 2.943 10.24 3.198 ;
      RECT 10.195 2.96 10.235 3.26 ;
      RECT 10.19 1.972 10.195 2.178 ;
      RECT 10.165 2.98 10.195 3.26 ;
      RECT 10.185 1.977 10.19 2.15 ;
      RECT 9.975 2.989 10.015 3.26 ;
      RECT 9.95 2.997 9.975 3.23 ;
      RECT 9.905 3.005 9.95 3.23 ;
      RECT 9.89 3.01 9.905 3.225 ;
      RECT 9.88 3.01 9.89 3.219 ;
      RECT 9.87 3.017 9.88 3.216 ;
      RECT 9.865 3.055 9.87 3.205 ;
      RECT 9.86 3.117 9.865 3.183 ;
      RECT 11.13 2.992 11.315 3.215 ;
      RECT 11.13 3.007 11.32 3.211 ;
      RECT 11.12 2.28 11.205 3.21 ;
      RECT 11.12 3.007 11.325 3.204 ;
      RECT 11.115 3.015 11.325 3.203 ;
      RECT 11.32 2.735 11.64 3.055 ;
      RECT 11.115 2.907 11.285 2.998 ;
      RECT 11.11 2.907 11.285 2.98 ;
      RECT 11.1 2.715 11.235 2.955 ;
      RECT 11.095 2.715 11.235 2.9 ;
      RECT 11.055 2.295 11.225 2.8 ;
      RECT 11.04 2.295 11.225 2.67 ;
      RECT 11.035 2.295 11.225 2.623 ;
      RECT 11.03 2.295 11.225 2.603 ;
      RECT 11.025 2.295 11.225 2.578 ;
      RECT 10.995 2.295 11.255 2.555 ;
      RECT 11.005 2.292 11.215 2.555 ;
      RECT 11.13 2.287 11.215 3.215 ;
      RECT 11.015 2.28 11.205 2.555 ;
      RECT 11.01 2.285 11.205 2.555 ;
      RECT 9.84 2.497 10.025 2.71 ;
      RECT 9.84 2.505 10.035 2.703 ;
      RECT 9.82 2.505 10.035 2.7 ;
      RECT 9.815 2.505 10.035 2.685 ;
      RECT 9.745 2.42 10.005 2.68 ;
      RECT 9.745 2.565 10.04 2.593 ;
      RECT 9.4 3.02 9.66 3.28 ;
      RECT 9.425 2.965 9.62 3.28 ;
      RECT 9.42 2.714 9.6 3.008 ;
      RECT 9.42 2.72 9.61 3.008 ;
      RECT 9.4 2.722 9.61 2.953 ;
      RECT 9.395 2.732 9.61 2.82 ;
      RECT 9.425 2.712 9.6 3.28 ;
      RECT 9.511 2.71 9.6 3.28 ;
      RECT 9.37 1.93 9.405 2.3 ;
      RECT 9.16 2.04 9.165 2.3 ;
      RECT 9.405 1.937 9.42 2.3 ;
      RECT 9.295 1.93 9.37 2.378 ;
      RECT 9.285 1.93 9.295 2.463 ;
      RECT 9.26 1.93 9.285 2.498 ;
      RECT 9.22 1.93 9.26 2.566 ;
      RECT 9.21 1.937 9.22 2.618 ;
      RECT 9.18 2.04 9.21 2.659 ;
      RECT 9.175 2.04 9.18 2.698 ;
      RECT 9.165 2.04 9.175 2.718 ;
      RECT 9.16 2.335 9.165 2.755 ;
      RECT 9.155 2.352 9.16 2.775 ;
      RECT 9.14 2.415 9.155 2.815 ;
      RECT 9.135 2.458 9.14 2.85 ;
      RECT 9.13 2.466 9.135 2.863 ;
      RECT 9.12 2.48 9.13 2.885 ;
      RECT 9.095 2.515 9.12 2.95 ;
      RECT 9.085 2.55 9.095 3.013 ;
      RECT 9.065 2.58 9.085 3.074 ;
      RECT 9.05 2.616 9.065 3.141 ;
      RECT 9.04 2.644 9.05 3.18 ;
      RECT 9.03 2.666 9.04 3.2 ;
      RECT 9.025 2.676 9.03 3.211 ;
      RECT 9.02 2.685 9.025 3.214 ;
      RECT 9.01 2.703 9.02 3.218 ;
      RECT 9 2.721 9.01 3.219 ;
      RECT 8.975 2.76 9 3.216 ;
      RECT 8.955 2.802 8.975 3.213 ;
      RECT 8.94 2.84 8.955 3.212 ;
      RECT 8.905 2.875 8.94 3.209 ;
      RECT 8.9 2.897 8.905 3.207 ;
      RECT 8.835 2.937 8.9 3.204 ;
      RECT 8.83 2.977 8.835 3.2 ;
      RECT 8.815 2.987 8.83 3.191 ;
      RECT 8.805 3.107 8.815 3.176 ;
      RECT 9.285 3.52 9.295 3.78 ;
      RECT 9.285 3.523 9.305 3.779 ;
      RECT 9.275 3.513 9.285 3.778 ;
      RECT 9.265 3.528 9.345 3.774 ;
      RECT 9.25 3.507 9.265 3.772 ;
      RECT 9.225 3.532 9.35 3.768 ;
      RECT 9.21 3.492 9.225 3.763 ;
      RECT 9.21 3.534 9.36 3.762 ;
      RECT 9.21 3.542 9.375 3.755 ;
      RECT 9.15 3.479 9.21 3.745 ;
      RECT 9.14 3.466 9.15 3.727 ;
      RECT 9.115 3.456 9.14 3.717 ;
      RECT 9.11 3.446 9.115 3.709 ;
      RECT 9.045 3.542 9.375 3.691 ;
      RECT 8.96 3.542 9.375 3.653 ;
      RECT 8.85 3.37 9.11 3.63 ;
      RECT 9.225 3.5 9.25 3.768 ;
      RECT 9.265 3.51 9.275 3.774 ;
      RECT 8.85 3.518 9.29 3.63 ;
      RECT 9.035 7.765 9.325 7.995 ;
      RECT 9.095 7.025 9.265 7.995 ;
      RECT 8.995 7.055 9.365 7.425 ;
      RECT 9.035 7.025 9.325 7.425 ;
      RECT 8.065 3.275 8.095 3.575 ;
      RECT 7.84 3.26 7.845 3.535 ;
      RECT 7.64 3.26 7.795 3.52 ;
      RECT 8.94 1.975 8.97 2.235 ;
      RECT 8.93 1.975 8.94 2.343 ;
      RECT 8.91 1.975 8.93 2.353 ;
      RECT 8.895 1.975 8.91 2.365 ;
      RECT 8.84 1.975 8.895 2.415 ;
      RECT 8.825 1.975 8.84 2.463 ;
      RECT 8.795 1.975 8.825 2.498 ;
      RECT 8.74 1.975 8.795 2.56 ;
      RECT 8.72 1.975 8.74 2.628 ;
      RECT 8.715 1.975 8.72 2.658 ;
      RECT 8.71 1.975 8.715 2.67 ;
      RECT 8.705 2.092 8.71 2.688 ;
      RECT 8.685 2.11 8.705 2.713 ;
      RECT 8.665 2.137 8.685 2.763 ;
      RECT 8.66 2.157 8.665 2.794 ;
      RECT 8.655 2.165 8.66 2.811 ;
      RECT 8.64 2.191 8.655 2.84 ;
      RECT 8.625 2.233 8.64 2.875 ;
      RECT 8.62 2.262 8.625 2.898 ;
      RECT 8.615 2.277 8.62 2.911 ;
      RECT 8.61 2.3 8.615 2.922 ;
      RECT 8.6 2.32 8.61 2.94 ;
      RECT 8.59 2.35 8.6 2.963 ;
      RECT 8.585 2.372 8.59 2.983 ;
      RECT 8.58 2.387 8.585 2.998 ;
      RECT 8.565 2.417 8.58 3.025 ;
      RECT 8.56 2.447 8.565 3.051 ;
      RECT 8.555 2.465 8.56 3.063 ;
      RECT 8.545 2.495 8.555 3.082 ;
      RECT 8.535 2.52 8.545 3.107 ;
      RECT 8.53 2.54 8.535 3.126 ;
      RECT 8.525 2.557 8.53 3.139 ;
      RECT 8.515 2.583 8.525 3.158 ;
      RECT 8.505 2.621 8.515 3.185 ;
      RECT 8.5 2.647 8.505 3.205 ;
      RECT 8.495 2.657 8.5 3.215 ;
      RECT 8.49 2.67 8.495 3.23 ;
      RECT 8.485 2.685 8.49 3.24 ;
      RECT 8.48 2.707 8.485 3.255 ;
      RECT 8.475 2.725 8.48 3.266 ;
      RECT 8.47 2.735 8.475 3.277 ;
      RECT 8.465 2.743 8.47 3.289 ;
      RECT 8.46 2.751 8.465 3.3 ;
      RECT 8.455 2.777 8.46 3.313 ;
      RECT 8.445 2.805 8.455 3.326 ;
      RECT 8.44 2.835 8.445 3.335 ;
      RECT 8.435 2.85 8.44 3.342 ;
      RECT 8.42 2.875 8.435 3.349 ;
      RECT 8.415 2.897 8.42 3.355 ;
      RECT 8.41 2.922 8.415 3.358 ;
      RECT 8.401 2.95 8.41 3.362 ;
      RECT 8.395 2.967 8.401 3.367 ;
      RECT 8.39 2.985 8.395 3.371 ;
      RECT 8.385 2.997 8.39 3.374 ;
      RECT 8.38 3.018 8.385 3.378 ;
      RECT 8.375 3.036 8.38 3.381 ;
      RECT 8.37 3.05 8.375 3.384 ;
      RECT 8.365 3.067 8.37 3.387 ;
      RECT 8.36 3.08 8.365 3.39 ;
      RECT 8.335 3.117 8.36 3.398 ;
      RECT 8.33 3.162 8.335 3.407 ;
      RECT 8.325 3.19 8.33 3.41 ;
      RECT 8.315 3.21 8.325 3.414 ;
      RECT 8.31 3.23 8.315 3.419 ;
      RECT 8.305 3.245 8.31 3.422 ;
      RECT 8.285 3.255 8.305 3.429 ;
      RECT 8.22 3.262 8.285 3.455 ;
      RECT 8.185 3.265 8.22 3.483 ;
      RECT 8.17 3.268 8.185 3.498 ;
      RECT 8.16 3.269 8.17 3.513 ;
      RECT 8.15 3.27 8.16 3.53 ;
      RECT 8.145 3.27 8.15 3.545 ;
      RECT 8.14 3.27 8.145 3.553 ;
      RECT 8.125 3.271 8.14 3.568 ;
      RECT 8.095 3.273 8.125 3.575 ;
      RECT 7.985 3.28 8.065 3.575 ;
      RECT 7.94 3.285 7.985 3.575 ;
      RECT 7.93 3.286 7.94 3.565 ;
      RECT 7.92 3.287 7.93 3.558 ;
      RECT 7.9 3.289 7.92 3.553 ;
      RECT 7.89 3.26 7.9 3.548 ;
      RECT 7.845 3.26 7.89 3.54 ;
      RECT 7.815 3.26 7.84 3.53 ;
      RECT 7.795 3.26 7.815 3.523 ;
      RECT 8.075 2.06 8.335 2.32 ;
      RECT 7.955 2.075 7.965 2.24 ;
      RECT 7.94 2.075 7.945 2.235 ;
      RECT 5.305 1.915 5.49 2.205 ;
      RECT 7.12 2.04 7.135 2.195 ;
      RECT 5.27 1.915 5.295 2.175 ;
      RECT 7.685 1.965 7.69 2.107 ;
      RECT 7.6 1.96 7.625 2.1 ;
      RECT 8 2.077 8.075 2.27 ;
      RECT 7.985 2.075 8 2.253 ;
      RECT 7.965 2.075 7.985 2.245 ;
      RECT 7.945 2.075 7.955 2.238 ;
      RECT 7.9 2.07 7.94 2.228 ;
      RECT 7.86 2.045 7.9 2.213 ;
      RECT 7.845 2.02 7.86 2.203 ;
      RECT 7.84 2.014 7.845 2.201 ;
      RECT 7.805 2.006 7.84 2.184 ;
      RECT 7.8 1.999 7.805 2.172 ;
      RECT 7.78 1.994 7.8 2.16 ;
      RECT 7.77 1.988 7.78 2.145 ;
      RECT 7.75 1.983 7.77 2.13 ;
      RECT 7.74 1.978 7.75 2.123 ;
      RECT 7.735 1.976 7.74 2.118 ;
      RECT 7.73 1.975 7.735 2.115 ;
      RECT 7.69 1.97 7.73 2.111 ;
      RECT 7.67 1.964 7.685 2.106 ;
      RECT 7.635 1.961 7.67 2.103 ;
      RECT 7.625 1.96 7.635 2.101 ;
      RECT 7.565 1.96 7.6 2.098 ;
      RECT 7.52 1.96 7.565 2.098 ;
      RECT 7.47 1.96 7.52 2.101 ;
      RECT 7.455 1.962 7.47 2.103 ;
      RECT 7.44 1.965 7.455 2.104 ;
      RECT 7.43 1.97 7.44 2.105 ;
      RECT 7.4 1.975 7.43 2.11 ;
      RECT 7.39 1.981 7.4 2.118 ;
      RECT 7.38 1.983 7.39 2.122 ;
      RECT 7.37 1.987 7.38 2.126 ;
      RECT 7.345 1.993 7.37 2.134 ;
      RECT 7.335 1.998 7.345 2.142 ;
      RECT 7.32 2.002 7.335 2.146 ;
      RECT 7.285 2.008 7.32 2.154 ;
      RECT 7.265 2.013 7.285 2.164 ;
      RECT 7.235 2.02 7.265 2.173 ;
      RECT 7.19 2.029 7.235 2.187 ;
      RECT 7.185 2.034 7.19 2.198 ;
      RECT 7.165 2.037 7.185 2.199 ;
      RECT 7.135 2.04 7.165 2.197 ;
      RECT 7.1 2.04 7.12 2.193 ;
      RECT 7.03 2.04 7.1 2.184 ;
      RECT 7.015 2.037 7.03 2.176 ;
      RECT 6.975 2.03 7.015 2.171 ;
      RECT 6.95 2.02 6.975 2.164 ;
      RECT 6.945 2.014 6.95 2.161 ;
      RECT 6.905 2.008 6.945 2.158 ;
      RECT 6.89 2.001 6.905 2.153 ;
      RECT 6.87 1.997 6.89 2.148 ;
      RECT 6.855 1.992 6.87 2.144 ;
      RECT 6.84 1.987 6.855 2.142 ;
      RECT 6.825 1.983 6.84 2.141 ;
      RECT 6.81 1.981 6.825 2.137 ;
      RECT 6.8 1.979 6.81 2.132 ;
      RECT 6.785 1.976 6.8 2.128 ;
      RECT 6.775 1.974 6.785 2.123 ;
      RECT 6.755 1.971 6.775 2.119 ;
      RECT 6.71 1.97 6.755 2.117 ;
      RECT 6.65 1.972 6.71 2.118 ;
      RECT 6.63 1.974 6.65 2.12 ;
      RECT 6.6 1.977 6.63 2.121 ;
      RECT 6.55 1.982 6.6 2.123 ;
      RECT 6.545 1.985 6.55 2.125 ;
      RECT 6.535 1.987 6.545 2.128 ;
      RECT 6.53 1.989 6.535 2.131 ;
      RECT 6.48 1.992 6.53 2.138 ;
      RECT 6.46 1.996 6.48 2.15 ;
      RECT 6.45 1.999 6.46 2.156 ;
      RECT 6.44 2 6.45 2.159 ;
      RECT 6.401 2.003 6.44 2.161 ;
      RECT 6.315 2.01 6.401 2.164 ;
      RECT 6.241 2.02 6.315 2.168 ;
      RECT 6.155 2.031 6.241 2.173 ;
      RECT 6.14 2.038 6.155 2.175 ;
      RECT 6.085 2.042 6.14 2.176 ;
      RECT 6.071 2.045 6.085 2.178 ;
      RECT 5.985 2.045 6.071 2.18 ;
      RECT 5.945 2.042 5.985 2.183 ;
      RECT 5.921 2.038 5.945 2.185 ;
      RECT 5.835 2.028 5.921 2.188 ;
      RECT 5.805 2.017 5.835 2.189 ;
      RECT 5.786 2.013 5.805 2.188 ;
      RECT 5.7 2.006 5.786 2.185 ;
      RECT 5.64 1.995 5.7 2.182 ;
      RECT 5.62 1.987 5.64 2.18 ;
      RECT 5.585 1.982 5.62 2.179 ;
      RECT 5.56 1.977 5.585 2.178 ;
      RECT 5.53 1.972 5.56 2.177 ;
      RECT 5.505 1.915 5.53 2.176 ;
      RECT 5.49 1.915 5.505 2.2 ;
      RECT 5.295 1.915 5.305 2.2 ;
      RECT 7.07 2.935 7.075 3.075 ;
      RECT 6.73 2.935 6.765 3.073 ;
      RECT 6.305 2.92 6.32 3.065 ;
      RECT 8.135 2.7 8.225 2.96 ;
      RECT 7.965 2.565 8.065 2.96 ;
      RECT 5 2.54 5.08 2.75 ;
      RECT 8.09 2.677 8.135 2.96 ;
      RECT 8.08 2.647 8.09 2.96 ;
      RECT 8.065 2.57 8.08 2.96 ;
      RECT 7.88 2.565 7.965 2.925 ;
      RECT 7.875 2.567 7.88 2.92 ;
      RECT 7.87 2.572 7.875 2.92 ;
      RECT 7.835 2.672 7.87 2.92 ;
      RECT 7.825 2.7 7.835 2.92 ;
      RECT 7.815 2.715 7.825 2.92 ;
      RECT 7.805 2.727 7.815 2.92 ;
      RECT 7.8 2.737 7.805 2.92 ;
      RECT 7.785 2.747 7.8 2.922 ;
      RECT 7.78 2.762 7.785 2.924 ;
      RECT 7.765 2.775 7.78 2.926 ;
      RECT 7.76 2.79 7.765 2.929 ;
      RECT 7.74 2.8 7.76 2.933 ;
      RECT 7.725 2.81 7.74 2.936 ;
      RECT 7.69 2.817 7.725 2.941 ;
      RECT 7.646 2.824 7.69 2.949 ;
      RECT 7.56 2.836 7.646 2.962 ;
      RECT 7.535 2.847 7.56 2.973 ;
      RECT 7.505 2.852 7.535 2.978 ;
      RECT 7.47 2.857 7.505 2.986 ;
      RECT 7.44 2.862 7.47 2.993 ;
      RECT 7.415 2.867 7.44 2.998 ;
      RECT 7.35 2.874 7.415 3.007 ;
      RECT 7.28 2.887 7.35 3.023 ;
      RECT 7.25 2.897 7.28 3.035 ;
      RECT 7.225 2.902 7.25 3.042 ;
      RECT 7.17 2.909 7.225 3.05 ;
      RECT 7.165 2.916 7.17 3.055 ;
      RECT 7.16 2.918 7.165 3.056 ;
      RECT 7.145 2.92 7.16 3.058 ;
      RECT 7.14 2.92 7.145 3.061 ;
      RECT 7.075 2.927 7.14 3.068 ;
      RECT 7.04 2.937 7.07 3.078 ;
      RECT 7.023 2.94 7.04 3.08 ;
      RECT 6.937 2.939 7.023 3.079 ;
      RECT 6.851 2.937 6.937 3.076 ;
      RECT 6.765 2.936 6.851 3.074 ;
      RECT 6.664 2.934 6.73 3.073 ;
      RECT 6.578 2.931 6.664 3.071 ;
      RECT 6.492 2.927 6.578 3.069 ;
      RECT 6.406 2.924 6.492 3.068 ;
      RECT 6.32 2.921 6.406 3.066 ;
      RECT 6.22 2.92 6.305 3.063 ;
      RECT 6.17 2.918 6.22 3.061 ;
      RECT 6.15 2.915 6.17 3.059 ;
      RECT 6.13 2.913 6.15 3.056 ;
      RECT 6.105 2.909 6.13 3.053 ;
      RECT 6.06 2.903 6.105 3.048 ;
      RECT 6.02 2.897 6.06 3.04 ;
      RECT 5.995 2.892 6.02 3.033 ;
      RECT 5.94 2.885 5.995 3.025 ;
      RECT 5.916 2.878 5.94 3.018 ;
      RECT 5.83 2.869 5.916 3.008 ;
      RECT 5.8 2.861 5.83 2.998 ;
      RECT 5.77 2.857 5.8 2.993 ;
      RECT 5.765 2.854 5.77 2.99 ;
      RECT 5.76 2.853 5.765 2.99 ;
      RECT 5.685 2.846 5.76 2.983 ;
      RECT 5.646 2.837 5.685 2.972 ;
      RECT 5.56 2.827 5.646 2.96 ;
      RECT 5.52 2.817 5.56 2.948 ;
      RECT 5.481 2.812 5.52 2.941 ;
      RECT 5.395 2.802 5.481 2.93 ;
      RECT 5.355 2.79 5.395 2.919 ;
      RECT 5.32 2.775 5.355 2.912 ;
      RECT 5.31 2.765 5.32 2.909 ;
      RECT 5.29 2.75 5.31 2.907 ;
      RECT 5.26 2.72 5.29 2.903 ;
      RECT 5.25 2.7 5.26 2.898 ;
      RECT 5.245 2.692 5.25 2.895 ;
      RECT 5.24 2.685 5.245 2.893 ;
      RECT 5.225 2.672 5.24 2.886 ;
      RECT 5.22 2.662 5.225 2.878 ;
      RECT 5.215 2.655 5.22 2.873 ;
      RECT 5.21 2.65 5.215 2.869 ;
      RECT 5.195 2.637 5.21 2.861 ;
      RECT 5.19 2.547 5.195 2.85 ;
      RECT 5.185 2.542 5.19 2.843 ;
      RECT 5.11 2.54 5.185 2.803 ;
      RECT 5.08 2.54 5.11 2.758 ;
      RECT 4.985 2.545 5 2.745 ;
      RECT 7.47 2.25 7.73 2.51 ;
      RECT 7.455 2.238 7.635 2.475 ;
      RECT 7.45 2.239 7.635 2.473 ;
      RECT 7.435 2.243 7.645 2.463 ;
      RECT 7.43 2.248 7.65 2.433 ;
      RECT 7.435 2.245 7.65 2.463 ;
      RECT 7.45 2.24 7.645 2.473 ;
      RECT 7.47 2.237 7.635 2.51 ;
      RECT 7.47 2.236 7.625 2.51 ;
      RECT 7.495 2.235 7.625 2.51 ;
      RECT 7.055 2.48 7.315 2.74 ;
      RECT 6.93 2.525 7.315 2.735 ;
      RECT 6.92 2.53 7.315 2.73 ;
      RECT 6.935 3.47 6.95 3.78 ;
      RECT 5.53 3.24 5.54 3.37 ;
      RECT 5.31 3.235 5.415 3.37 ;
      RECT 5.225 3.24 5.275 3.37 ;
      RECT 3.775 1.975 3.78 3.08 ;
      RECT 7.03 3.562 7.035 3.698 ;
      RECT 7.025 3.557 7.03 3.758 ;
      RECT 7.02 3.555 7.025 3.771 ;
      RECT 7.005 3.552 7.02 3.773 ;
      RECT 7 3.547 7.005 3.775 ;
      RECT 6.995 3.543 7 3.778 ;
      RECT 6.98 3.538 6.995 3.78 ;
      RECT 6.95 3.53 6.98 3.78 ;
      RECT 6.911 3.47 6.935 3.78 ;
      RECT 6.825 3.47 6.911 3.777 ;
      RECT 6.795 3.47 6.825 3.77 ;
      RECT 6.77 3.47 6.795 3.763 ;
      RECT 6.745 3.47 6.77 3.755 ;
      RECT 6.73 3.47 6.745 3.748 ;
      RECT 6.705 3.47 6.73 3.74 ;
      RECT 6.69 3.47 6.705 3.733 ;
      RECT 6.65 3.48 6.69 3.722 ;
      RECT 6.64 3.475 6.65 3.712 ;
      RECT 6.636 3.474 6.64 3.709 ;
      RECT 6.55 3.466 6.636 3.692 ;
      RECT 6.517 3.455 6.55 3.669 ;
      RECT 6.431 3.444 6.517 3.647 ;
      RECT 6.345 3.428 6.431 3.616 ;
      RECT 6.275 3.413 6.345 3.588 ;
      RECT 6.265 3.406 6.275 3.575 ;
      RECT 6.235 3.403 6.265 3.565 ;
      RECT 6.21 3.399 6.235 3.558 ;
      RECT 6.195 3.396 6.21 3.553 ;
      RECT 6.19 3.395 6.195 3.548 ;
      RECT 6.16 3.39 6.19 3.541 ;
      RECT 6.155 3.385 6.16 3.536 ;
      RECT 6.14 3.382 6.155 3.531 ;
      RECT 6.135 3.377 6.14 3.526 ;
      RECT 6.115 3.372 6.135 3.523 ;
      RECT 6.1 3.367 6.115 3.515 ;
      RECT 6.085 3.361 6.1 3.51 ;
      RECT 6.055 3.352 6.085 3.503 ;
      RECT 6.05 3.345 6.055 3.495 ;
      RECT 6.045 3.343 6.05 3.493 ;
      RECT 6.04 3.342 6.045 3.49 ;
      RECT 6 3.335 6.04 3.483 ;
      RECT 5.986 3.325 6 3.473 ;
      RECT 5.935 3.314 5.986 3.461 ;
      RECT 5.91 3.3 5.935 3.447 ;
      RECT 5.885 3.289 5.91 3.439 ;
      RECT 5.865 3.278 5.885 3.433 ;
      RECT 5.855 3.272 5.865 3.428 ;
      RECT 5.85 3.27 5.855 3.424 ;
      RECT 5.83 3.265 5.85 3.419 ;
      RECT 5.8 3.255 5.83 3.409 ;
      RECT 5.795 3.247 5.8 3.402 ;
      RECT 5.78 3.245 5.795 3.398 ;
      RECT 5.76 3.245 5.78 3.393 ;
      RECT 5.755 3.244 5.76 3.391 ;
      RECT 5.75 3.244 5.755 3.388 ;
      RECT 5.71 3.243 5.75 3.383 ;
      RECT 5.685 3.242 5.71 3.378 ;
      RECT 5.625 3.241 5.685 3.375 ;
      RECT 5.54 3.24 5.625 3.373 ;
      RECT 5.501 3.239 5.53 3.37 ;
      RECT 5.415 3.237 5.501 3.37 ;
      RECT 5.275 3.237 5.31 3.37 ;
      RECT 5.185 3.241 5.225 3.373 ;
      RECT 5.17 3.244 5.185 3.38 ;
      RECT 5.16 3.245 5.17 3.387 ;
      RECT 5.135 3.248 5.16 3.392 ;
      RECT 5.13 3.25 5.135 3.395 ;
      RECT 5.08 3.252 5.13 3.396 ;
      RECT 5.041 3.256 5.08 3.398 ;
      RECT 4.955 3.258 5.041 3.401 ;
      RECT 4.937 3.26 4.955 3.403 ;
      RECT 4.851 3.263 4.937 3.405 ;
      RECT 4.765 3.267 4.851 3.408 ;
      RECT 4.728 3.271 4.765 3.411 ;
      RECT 4.642 3.274 4.728 3.414 ;
      RECT 4.556 3.278 4.642 3.417 ;
      RECT 4.47 3.283 4.556 3.421 ;
      RECT 4.45 3.285 4.47 3.424 ;
      RECT 4.43 3.284 4.45 3.425 ;
      RECT 4.381 3.281 4.43 3.426 ;
      RECT 4.295 3.276 4.381 3.429 ;
      RECT 4.245 3.271 4.295 3.431 ;
      RECT 4.221 3.269 4.245 3.432 ;
      RECT 4.135 3.264 4.221 3.434 ;
      RECT 4.11 3.26 4.135 3.433 ;
      RECT 4.1 3.257 4.11 3.431 ;
      RECT 4.09 3.25 4.1 3.428 ;
      RECT 4.085 3.23 4.09 3.423 ;
      RECT 4.075 3.2 4.085 3.418 ;
      RECT 4.06 3.07 4.075 3.409 ;
      RECT 4.055 3.062 4.06 3.402 ;
      RECT 4.035 3.055 4.055 3.394 ;
      RECT 4.03 3.037 4.035 3.386 ;
      RECT 4.02 3.017 4.03 3.381 ;
      RECT 4.015 2.99 4.02 3.377 ;
      RECT 4.01 2.967 4.015 3.374 ;
      RECT 3.99 2.925 4.01 3.366 ;
      RECT 3.955 2.84 3.99 3.35 ;
      RECT 3.95 2.772 3.955 3.338 ;
      RECT 3.935 2.742 3.95 3.332 ;
      RECT 3.93 1.987 3.935 2.233 ;
      RECT 3.92 2.712 3.935 3.323 ;
      RECT 3.925 1.982 3.93 2.265 ;
      RECT 3.92 1.977 3.925 2.308 ;
      RECT 3.915 1.975 3.92 2.343 ;
      RECT 3.9 2.675 3.92 3.313 ;
      RECT 3.91 1.975 3.915 2.38 ;
      RECT 3.895 1.975 3.91 2.478 ;
      RECT 3.895 2.648 3.9 3.306 ;
      RECT 3.89 1.975 3.895 2.553 ;
      RECT 3.89 2.636 3.895 3.303 ;
      RECT 3.885 1.975 3.89 2.585 ;
      RECT 3.885 2.615 3.89 3.3 ;
      RECT 3.88 1.975 3.885 3.297 ;
      RECT 3.845 1.975 3.88 3.283 ;
      RECT 3.83 1.975 3.845 3.265 ;
      RECT 3.81 1.975 3.83 3.255 ;
      RECT 3.785 1.975 3.81 3.238 ;
      RECT 3.78 1.975 3.785 3.188 ;
      RECT 3.77 1.975 3.775 3.018 ;
      RECT 3.765 1.975 3.77 2.925 ;
      RECT 3.76 1.975 3.765 2.838 ;
      RECT 3.755 1.975 3.76 2.77 ;
      RECT 3.75 1.975 3.755 2.713 ;
      RECT 3.74 1.975 3.75 2.608 ;
      RECT 3.735 1.975 3.74 2.48 ;
      RECT 3.73 1.975 3.735 2.398 ;
      RECT 3.725 1.977 3.73 2.315 ;
      RECT 3.72 1.982 3.725 2.248 ;
      RECT 3.715 1.987 3.72 2.175 ;
      RECT 6.53 2.305 6.79 2.565 ;
      RECT 6.55 2.272 6.76 2.565 ;
      RECT 6.55 2.27 6.75 2.565 ;
      RECT 6.56 2.257 6.75 2.565 ;
      RECT 6.56 2.255 6.675 2.565 ;
      RECT 6.035 2.38 6.21 2.66 ;
      RECT 6.03 2.38 6.21 2.658 ;
      RECT 6.03 2.38 6.225 2.655 ;
      RECT 6.02 2.38 6.225 2.653 ;
      RECT 5.965 2.38 6.225 2.64 ;
      RECT 5.965 2.455 6.23 2.618 ;
      RECT 5.51 2.392 5.53 2.635 ;
      RECT 5.51 2.392 5.57 2.634 ;
      RECT 5.505 2.394 5.57 2.633 ;
      RECT 5.505 2.394 5.656 2.632 ;
      RECT 5.505 2.394 5.725 2.631 ;
      RECT 5.505 2.394 5.745 2.623 ;
      RECT 5.485 2.397 5.745 2.621 ;
      RECT 5.47 2.407 5.745 2.606 ;
      RECT 5.47 2.407 5.76 2.605 ;
      RECT 5.465 2.416 5.76 2.597 ;
      RECT 5.465 2.416 5.765 2.593 ;
      RECT 5.57 2.33 5.83 2.59 ;
      RECT 5.46 2.418 5.83 2.475 ;
      RECT 5.53 2.385 5.83 2.59 ;
      RECT 5.495 3.578 5.5 3.785 ;
      RECT 5.445 3.572 5.495 3.784 ;
      RECT 5.412 3.586 5.505 3.783 ;
      RECT 5.326 3.586 5.505 3.782 ;
      RECT 5.24 3.586 5.505 3.781 ;
      RECT 5.24 3.685 5.51 3.778 ;
      RECT 5.235 3.685 5.51 3.773 ;
      RECT 5.23 3.685 5.51 3.755 ;
      RECT 5.225 3.685 5.51 3.738 ;
      RECT 5.185 3.47 5.445 3.73 ;
      RECT 4.645 2.62 4.731 3.034 ;
      RECT 4.645 2.62 4.77 3.031 ;
      RECT 4.645 2.62 4.79 3.021 ;
      RECT 4.6 2.62 4.79 3.018 ;
      RECT 4.6 2.772 4.8 3.008 ;
      RECT 4.6 2.793 4.805 3.002 ;
      RECT 4.6 2.811 4.81 2.998 ;
      RECT 4.6 2.831 4.82 2.993 ;
      RECT 4.575 2.831 4.82 2.99 ;
      RECT 4.565 2.831 4.82 2.968 ;
      RECT 4.565 2.847 4.825 2.938 ;
      RECT 4.53 2.62 4.79 2.925 ;
      RECT 4.53 2.859 4.83 2.88 ;
      RECT 1.54 7.765 1.83 7.995 ;
      RECT 1.6 7.025 1.77 7.995 ;
      RECT 1.51 7.025 1.86 7.315 ;
      RECT 1.135 6.285 1.485 6.575 ;
      RECT 0.995 6.315 1.485 6.485 ;
      RECT 68.155 3.265 68.415 3.525 ;
      RECT 52.895 3.265 53.155 3.525 ;
      RECT 37.635 3.265 37.895 3.525 ;
      RECT 22.375 3.265 22.635 3.525 ;
      RECT 7.115 3.265 7.375 3.525 ;
    LAYER mcon ;
      RECT 78.55 6.32 78.72 6.49 ;
      RECT 78.555 6.315 78.725 6.485 ;
      RECT 63.29 6.32 63.46 6.49 ;
      RECT 63.295 6.315 63.465 6.485 ;
      RECT 48.03 6.32 48.2 6.49 ;
      RECT 48.035 6.315 48.205 6.485 ;
      RECT 32.77 6.32 32.94 6.49 ;
      RECT 32.775 6.315 32.945 6.485 ;
      RECT 17.51 6.32 17.68 6.49 ;
      RECT 17.515 6.315 17.685 6.485 ;
      RECT 78.55 7.8 78.72 7.97 ;
      RECT 78.2 0.1 78.37 0.27 ;
      RECT 78.2 8.61 78.37 8.78 ;
      RECT 78.18 2.76 78.35 2.93 ;
      RECT 78.18 5.95 78.35 6.12 ;
      RECT 77.56 0.91 77.73 1.08 ;
      RECT 77.56 2.39 77.73 2.56 ;
      RECT 77.56 6.32 77.73 6.49 ;
      RECT 77.56 7.8 77.73 7.97 ;
      RECT 77.21 0.1 77.38 0.27 ;
      RECT 77.21 8.61 77.38 8.78 ;
      RECT 77.19 2.76 77.36 2.93 ;
      RECT 77.19 5.95 77.36 6.12 ;
      RECT 76.51 0.105 76.68 0.275 ;
      RECT 76.51 8.605 76.68 8.775 ;
      RECT 76.2 2.025 76.37 2.195 ;
      RECT 76.2 6.685 76.37 6.855 ;
      RECT 75.83 0.105 76 0.275 ;
      RECT 75.83 8.605 76 8.775 ;
      RECT 75.77 0.915 75.94 1.085 ;
      RECT 75.77 1.655 75.94 1.825 ;
      RECT 75.77 7.055 75.94 7.225 ;
      RECT 75.77 7.795 75.94 7.965 ;
      RECT 75.395 2.395 75.565 2.565 ;
      RECT 75.395 6.315 75.565 6.485 ;
      RECT 75.15 0.105 75.32 0.275 ;
      RECT 75.15 8.605 75.32 8.775 ;
      RECT 74.47 0.105 74.64 0.275 ;
      RECT 74.47 8.605 74.64 8.775 ;
      RECT 73.01 1.415 73.18 1.585 ;
      RECT 72.57 2.28 72.74 2.45 ;
      RECT 72.55 1.415 72.72 1.585 ;
      RECT 72.175 3.025 72.345 3.195 ;
      RECT 72.09 1.415 72.26 1.585 ;
      RECT 72.065 2.3 72.235 2.47 ;
      RECT 71.63 1.415 71.8 1.585 ;
      RECT 71.245 1.99 71.415 2.16 ;
      RECT 71.17 1.415 71.34 1.585 ;
      RECT 70.93 3.03 71.1 3.2 ;
      RECT 70.885 2.52 71.055 2.69 ;
      RECT 70.875 8.605 71.045 8.775 ;
      RECT 70.71 1.415 70.88 1.585 ;
      RECT 70.565 6.685 70.735 6.855 ;
      RECT 70.46 2.73 70.63 2.9 ;
      RECT 70.27 1.95 70.44 2.12 ;
      RECT 70.25 1.415 70.42 1.585 ;
      RECT 70.22 3.56 70.39 3.73 ;
      RECT 70.195 8.605 70.365 8.775 ;
      RECT 70.135 7.055 70.305 7.225 ;
      RECT 70.135 7.795 70.305 7.965 ;
      RECT 69.885 3 70.055 3.17 ;
      RECT 69.79 1.415 69.96 1.585 ;
      RECT 69.79 2.16 69.96 2.33 ;
      RECT 69.76 6.315 69.93 6.485 ;
      RECT 69.515 8.605 69.685 8.775 ;
      RECT 69.33 1.415 69.5 1.585 ;
      RECT 68.99 3.385 69.16 3.555 ;
      RECT 68.93 2.585 69.1 2.755 ;
      RECT 68.87 1.415 69.04 1.585 ;
      RECT 68.835 8.605 69.005 8.775 ;
      RECT 68.49 2.255 68.66 2.425 ;
      RECT 68.41 1.415 68.58 1.585 ;
      RECT 68.225 3.305 68.395 3.475 ;
      RECT 67.98 2.545 68.15 2.715 ;
      RECT 67.95 1.415 68.12 1.585 ;
      RECT 67.885 3.575 68.055 3.745 ;
      RECT 67.61 2.27 67.78 2.44 ;
      RECT 67.49 1.415 67.66 1.585 ;
      RECT 67.08 2.47 67.25 2.64 ;
      RECT 67.03 1.415 67.2 1.585 ;
      RECT 66.57 1.415 66.74 1.585 ;
      RECT 66.56 2.415 66.73 2.585 ;
      RECT 66.355 2.015 66.525 2.185 ;
      RECT 66.355 3.595 66.525 3.765 ;
      RECT 66.11 1.415 66.28 1.585 ;
      RECT 66.045 2.56 66.215 2.73 ;
      RECT 65.65 1.415 65.82 1.585 ;
      RECT 65.635 2.785 65.805 2.955 ;
      RECT 65.19 1.415 65.36 1.585 ;
      RECT 64.925 3.085 65.095 3.255 ;
      RECT 64.78 1.995 64.95 2.165 ;
      RECT 64.73 1.415 64.9 1.585 ;
      RECT 63.29 7.8 63.46 7.97 ;
      RECT 62.94 0.1 63.11 0.27 ;
      RECT 62.94 8.61 63.11 8.78 ;
      RECT 62.92 2.76 63.09 2.93 ;
      RECT 62.92 5.95 63.09 6.12 ;
      RECT 62.3 0.91 62.47 1.08 ;
      RECT 62.3 2.39 62.47 2.56 ;
      RECT 62.3 6.32 62.47 6.49 ;
      RECT 62.3 7.8 62.47 7.97 ;
      RECT 61.95 0.1 62.12 0.27 ;
      RECT 61.95 8.61 62.12 8.78 ;
      RECT 61.93 2.76 62.1 2.93 ;
      RECT 61.93 5.95 62.1 6.12 ;
      RECT 61.25 0.105 61.42 0.275 ;
      RECT 61.25 8.605 61.42 8.775 ;
      RECT 60.94 2.025 61.11 2.195 ;
      RECT 60.94 6.685 61.11 6.855 ;
      RECT 60.57 0.105 60.74 0.275 ;
      RECT 60.57 8.605 60.74 8.775 ;
      RECT 60.51 0.915 60.68 1.085 ;
      RECT 60.51 1.655 60.68 1.825 ;
      RECT 60.51 7.055 60.68 7.225 ;
      RECT 60.51 7.795 60.68 7.965 ;
      RECT 60.135 2.395 60.305 2.565 ;
      RECT 60.135 6.315 60.305 6.485 ;
      RECT 59.89 0.105 60.06 0.275 ;
      RECT 59.89 8.605 60.06 8.775 ;
      RECT 59.21 0.105 59.38 0.275 ;
      RECT 59.21 8.605 59.38 8.775 ;
      RECT 57.75 1.415 57.92 1.585 ;
      RECT 57.31 2.28 57.48 2.45 ;
      RECT 57.29 1.415 57.46 1.585 ;
      RECT 56.915 3.025 57.085 3.195 ;
      RECT 56.83 1.415 57 1.585 ;
      RECT 56.805 2.3 56.975 2.47 ;
      RECT 56.37 1.415 56.54 1.585 ;
      RECT 55.985 1.99 56.155 2.16 ;
      RECT 55.91 1.415 56.08 1.585 ;
      RECT 55.67 3.03 55.84 3.2 ;
      RECT 55.625 2.52 55.795 2.69 ;
      RECT 55.615 8.605 55.785 8.775 ;
      RECT 55.45 1.415 55.62 1.585 ;
      RECT 55.305 6.685 55.475 6.855 ;
      RECT 55.2 2.73 55.37 2.9 ;
      RECT 55.01 1.95 55.18 2.12 ;
      RECT 54.99 1.415 55.16 1.585 ;
      RECT 54.96 3.56 55.13 3.73 ;
      RECT 54.935 8.605 55.105 8.775 ;
      RECT 54.875 7.055 55.045 7.225 ;
      RECT 54.875 7.795 55.045 7.965 ;
      RECT 54.625 3 54.795 3.17 ;
      RECT 54.53 1.415 54.7 1.585 ;
      RECT 54.53 2.16 54.7 2.33 ;
      RECT 54.5 6.315 54.67 6.485 ;
      RECT 54.255 8.605 54.425 8.775 ;
      RECT 54.07 1.415 54.24 1.585 ;
      RECT 53.73 3.385 53.9 3.555 ;
      RECT 53.67 2.585 53.84 2.755 ;
      RECT 53.61 1.415 53.78 1.585 ;
      RECT 53.575 8.605 53.745 8.775 ;
      RECT 53.23 2.255 53.4 2.425 ;
      RECT 53.15 1.415 53.32 1.585 ;
      RECT 52.965 3.305 53.135 3.475 ;
      RECT 52.72 2.545 52.89 2.715 ;
      RECT 52.69 1.415 52.86 1.585 ;
      RECT 52.625 3.575 52.795 3.745 ;
      RECT 52.35 2.27 52.52 2.44 ;
      RECT 52.23 1.415 52.4 1.585 ;
      RECT 51.82 2.47 51.99 2.64 ;
      RECT 51.77 1.415 51.94 1.585 ;
      RECT 51.31 1.415 51.48 1.585 ;
      RECT 51.3 2.415 51.47 2.585 ;
      RECT 51.095 2.015 51.265 2.185 ;
      RECT 51.095 3.595 51.265 3.765 ;
      RECT 50.85 1.415 51.02 1.585 ;
      RECT 50.785 2.56 50.955 2.73 ;
      RECT 50.39 1.415 50.56 1.585 ;
      RECT 50.375 2.785 50.545 2.955 ;
      RECT 49.93 1.415 50.1 1.585 ;
      RECT 49.665 3.085 49.835 3.255 ;
      RECT 49.52 1.995 49.69 2.165 ;
      RECT 49.47 1.415 49.64 1.585 ;
      RECT 48.03 7.8 48.2 7.97 ;
      RECT 47.68 0.1 47.85 0.27 ;
      RECT 47.68 8.61 47.85 8.78 ;
      RECT 47.66 2.76 47.83 2.93 ;
      RECT 47.66 5.95 47.83 6.12 ;
      RECT 47.04 0.91 47.21 1.08 ;
      RECT 47.04 2.39 47.21 2.56 ;
      RECT 47.04 6.32 47.21 6.49 ;
      RECT 47.04 7.8 47.21 7.97 ;
      RECT 46.69 0.1 46.86 0.27 ;
      RECT 46.69 8.61 46.86 8.78 ;
      RECT 46.67 2.76 46.84 2.93 ;
      RECT 46.67 5.95 46.84 6.12 ;
      RECT 45.99 0.105 46.16 0.275 ;
      RECT 45.99 8.605 46.16 8.775 ;
      RECT 45.68 2.025 45.85 2.195 ;
      RECT 45.68 6.685 45.85 6.855 ;
      RECT 45.31 0.105 45.48 0.275 ;
      RECT 45.31 8.605 45.48 8.775 ;
      RECT 45.25 0.915 45.42 1.085 ;
      RECT 45.25 1.655 45.42 1.825 ;
      RECT 45.25 7.055 45.42 7.225 ;
      RECT 45.25 7.795 45.42 7.965 ;
      RECT 44.875 2.395 45.045 2.565 ;
      RECT 44.875 6.315 45.045 6.485 ;
      RECT 44.63 0.105 44.8 0.275 ;
      RECT 44.63 8.605 44.8 8.775 ;
      RECT 43.95 0.105 44.12 0.275 ;
      RECT 43.95 8.605 44.12 8.775 ;
      RECT 42.49 1.415 42.66 1.585 ;
      RECT 42.05 2.28 42.22 2.45 ;
      RECT 42.03 1.415 42.2 1.585 ;
      RECT 41.655 3.025 41.825 3.195 ;
      RECT 41.57 1.415 41.74 1.585 ;
      RECT 41.545 2.3 41.715 2.47 ;
      RECT 41.11 1.415 41.28 1.585 ;
      RECT 40.725 1.99 40.895 2.16 ;
      RECT 40.65 1.415 40.82 1.585 ;
      RECT 40.41 3.03 40.58 3.2 ;
      RECT 40.365 2.52 40.535 2.69 ;
      RECT 40.355 8.605 40.525 8.775 ;
      RECT 40.19 1.415 40.36 1.585 ;
      RECT 40.045 6.685 40.215 6.855 ;
      RECT 39.94 2.73 40.11 2.9 ;
      RECT 39.75 1.95 39.92 2.12 ;
      RECT 39.73 1.415 39.9 1.585 ;
      RECT 39.7 3.56 39.87 3.73 ;
      RECT 39.675 8.605 39.845 8.775 ;
      RECT 39.615 7.055 39.785 7.225 ;
      RECT 39.615 7.795 39.785 7.965 ;
      RECT 39.365 3 39.535 3.17 ;
      RECT 39.27 1.415 39.44 1.585 ;
      RECT 39.27 2.16 39.44 2.33 ;
      RECT 39.24 6.315 39.41 6.485 ;
      RECT 38.995 8.605 39.165 8.775 ;
      RECT 38.81 1.415 38.98 1.585 ;
      RECT 38.47 3.385 38.64 3.555 ;
      RECT 38.41 2.585 38.58 2.755 ;
      RECT 38.35 1.415 38.52 1.585 ;
      RECT 38.315 8.605 38.485 8.775 ;
      RECT 37.97 2.255 38.14 2.425 ;
      RECT 37.89 1.415 38.06 1.585 ;
      RECT 37.705 3.305 37.875 3.475 ;
      RECT 37.46 2.545 37.63 2.715 ;
      RECT 37.43 1.415 37.6 1.585 ;
      RECT 37.365 3.575 37.535 3.745 ;
      RECT 37.09 2.27 37.26 2.44 ;
      RECT 36.97 1.415 37.14 1.585 ;
      RECT 36.56 2.47 36.73 2.64 ;
      RECT 36.51 1.415 36.68 1.585 ;
      RECT 36.05 1.415 36.22 1.585 ;
      RECT 36.04 2.415 36.21 2.585 ;
      RECT 35.835 2.015 36.005 2.185 ;
      RECT 35.835 3.595 36.005 3.765 ;
      RECT 35.59 1.415 35.76 1.585 ;
      RECT 35.525 2.56 35.695 2.73 ;
      RECT 35.13 1.415 35.3 1.585 ;
      RECT 35.115 2.785 35.285 2.955 ;
      RECT 34.67 1.415 34.84 1.585 ;
      RECT 34.405 3.085 34.575 3.255 ;
      RECT 34.26 1.995 34.43 2.165 ;
      RECT 34.21 1.415 34.38 1.585 ;
      RECT 32.77 7.8 32.94 7.97 ;
      RECT 32.42 0.1 32.59 0.27 ;
      RECT 32.42 8.61 32.59 8.78 ;
      RECT 32.4 2.76 32.57 2.93 ;
      RECT 32.4 5.95 32.57 6.12 ;
      RECT 31.78 0.91 31.95 1.08 ;
      RECT 31.78 2.39 31.95 2.56 ;
      RECT 31.78 6.32 31.95 6.49 ;
      RECT 31.78 7.8 31.95 7.97 ;
      RECT 31.43 0.1 31.6 0.27 ;
      RECT 31.43 8.61 31.6 8.78 ;
      RECT 31.41 2.76 31.58 2.93 ;
      RECT 31.41 5.95 31.58 6.12 ;
      RECT 30.73 0.105 30.9 0.275 ;
      RECT 30.73 8.605 30.9 8.775 ;
      RECT 30.42 2.025 30.59 2.195 ;
      RECT 30.42 6.685 30.59 6.855 ;
      RECT 30.05 0.105 30.22 0.275 ;
      RECT 30.05 8.605 30.22 8.775 ;
      RECT 29.99 0.915 30.16 1.085 ;
      RECT 29.99 1.655 30.16 1.825 ;
      RECT 29.99 7.055 30.16 7.225 ;
      RECT 29.99 7.795 30.16 7.965 ;
      RECT 29.615 2.395 29.785 2.565 ;
      RECT 29.615 6.315 29.785 6.485 ;
      RECT 29.37 0.105 29.54 0.275 ;
      RECT 29.37 8.605 29.54 8.775 ;
      RECT 28.69 0.105 28.86 0.275 ;
      RECT 28.69 8.605 28.86 8.775 ;
      RECT 27.23 1.415 27.4 1.585 ;
      RECT 26.79 2.28 26.96 2.45 ;
      RECT 26.77 1.415 26.94 1.585 ;
      RECT 26.395 3.025 26.565 3.195 ;
      RECT 26.31 1.415 26.48 1.585 ;
      RECT 26.285 2.3 26.455 2.47 ;
      RECT 25.85 1.415 26.02 1.585 ;
      RECT 25.465 1.99 25.635 2.16 ;
      RECT 25.39 1.415 25.56 1.585 ;
      RECT 25.15 3.03 25.32 3.2 ;
      RECT 25.105 2.52 25.275 2.69 ;
      RECT 25.095 8.605 25.265 8.775 ;
      RECT 24.93 1.415 25.1 1.585 ;
      RECT 24.785 6.685 24.955 6.855 ;
      RECT 24.68 2.73 24.85 2.9 ;
      RECT 24.49 1.95 24.66 2.12 ;
      RECT 24.47 1.415 24.64 1.585 ;
      RECT 24.44 3.56 24.61 3.73 ;
      RECT 24.415 8.605 24.585 8.775 ;
      RECT 24.355 7.055 24.525 7.225 ;
      RECT 24.355 7.795 24.525 7.965 ;
      RECT 24.105 3 24.275 3.17 ;
      RECT 24.01 1.415 24.18 1.585 ;
      RECT 24.01 2.16 24.18 2.33 ;
      RECT 23.98 6.315 24.15 6.485 ;
      RECT 23.735 8.605 23.905 8.775 ;
      RECT 23.55 1.415 23.72 1.585 ;
      RECT 23.21 3.385 23.38 3.555 ;
      RECT 23.15 2.585 23.32 2.755 ;
      RECT 23.09 1.415 23.26 1.585 ;
      RECT 23.055 8.605 23.225 8.775 ;
      RECT 22.71 2.255 22.88 2.425 ;
      RECT 22.63 1.415 22.8 1.585 ;
      RECT 22.445 3.305 22.615 3.475 ;
      RECT 22.2 2.545 22.37 2.715 ;
      RECT 22.17 1.415 22.34 1.585 ;
      RECT 22.105 3.575 22.275 3.745 ;
      RECT 21.83 2.27 22 2.44 ;
      RECT 21.71 1.415 21.88 1.585 ;
      RECT 21.3 2.47 21.47 2.64 ;
      RECT 21.25 1.415 21.42 1.585 ;
      RECT 20.79 1.415 20.96 1.585 ;
      RECT 20.78 2.415 20.95 2.585 ;
      RECT 20.575 2.015 20.745 2.185 ;
      RECT 20.575 3.595 20.745 3.765 ;
      RECT 20.33 1.415 20.5 1.585 ;
      RECT 20.265 2.56 20.435 2.73 ;
      RECT 19.87 1.415 20.04 1.585 ;
      RECT 19.855 2.785 20.025 2.955 ;
      RECT 19.41 1.415 19.58 1.585 ;
      RECT 19.145 3.085 19.315 3.255 ;
      RECT 19 1.995 19.17 2.165 ;
      RECT 18.95 1.415 19.12 1.585 ;
      RECT 17.51 7.8 17.68 7.97 ;
      RECT 17.16 0.1 17.33 0.27 ;
      RECT 17.16 8.61 17.33 8.78 ;
      RECT 17.14 2.76 17.31 2.93 ;
      RECT 17.14 5.95 17.31 6.12 ;
      RECT 16.52 0.91 16.69 1.08 ;
      RECT 16.52 2.39 16.69 2.56 ;
      RECT 16.52 6.32 16.69 6.49 ;
      RECT 16.52 7.8 16.69 7.97 ;
      RECT 16.17 0.1 16.34 0.27 ;
      RECT 16.17 8.61 16.34 8.78 ;
      RECT 16.15 2.76 16.32 2.93 ;
      RECT 16.15 5.95 16.32 6.12 ;
      RECT 15.47 0.105 15.64 0.275 ;
      RECT 15.47 8.605 15.64 8.775 ;
      RECT 15.16 2.025 15.33 2.195 ;
      RECT 15.16 6.685 15.33 6.855 ;
      RECT 14.79 0.105 14.96 0.275 ;
      RECT 14.79 8.605 14.96 8.775 ;
      RECT 14.73 0.915 14.9 1.085 ;
      RECT 14.73 1.655 14.9 1.825 ;
      RECT 14.73 7.055 14.9 7.225 ;
      RECT 14.73 7.795 14.9 7.965 ;
      RECT 14.355 2.395 14.525 2.565 ;
      RECT 14.355 6.315 14.525 6.485 ;
      RECT 14.11 0.105 14.28 0.275 ;
      RECT 14.11 8.605 14.28 8.775 ;
      RECT 13.43 0.105 13.6 0.275 ;
      RECT 13.43 8.605 13.6 8.775 ;
      RECT 11.97 1.415 12.14 1.585 ;
      RECT 11.53 2.28 11.7 2.45 ;
      RECT 11.51 1.415 11.68 1.585 ;
      RECT 11.135 3.025 11.305 3.195 ;
      RECT 11.05 1.415 11.22 1.585 ;
      RECT 11.025 2.3 11.195 2.47 ;
      RECT 10.59 1.415 10.76 1.585 ;
      RECT 10.205 1.99 10.375 2.16 ;
      RECT 10.13 1.415 10.3 1.585 ;
      RECT 9.89 3.03 10.06 3.2 ;
      RECT 9.845 2.52 10.015 2.69 ;
      RECT 9.835 8.605 10.005 8.775 ;
      RECT 9.67 1.415 9.84 1.585 ;
      RECT 9.525 6.685 9.695 6.855 ;
      RECT 9.42 2.73 9.59 2.9 ;
      RECT 9.23 1.95 9.4 2.12 ;
      RECT 9.21 1.415 9.38 1.585 ;
      RECT 9.18 3.56 9.35 3.73 ;
      RECT 9.155 8.605 9.325 8.775 ;
      RECT 9.095 7.055 9.265 7.225 ;
      RECT 9.095 7.795 9.265 7.965 ;
      RECT 8.845 3 9.015 3.17 ;
      RECT 8.75 1.415 8.92 1.585 ;
      RECT 8.75 2.16 8.92 2.33 ;
      RECT 8.72 6.315 8.89 6.485 ;
      RECT 8.475 8.605 8.645 8.775 ;
      RECT 8.29 1.415 8.46 1.585 ;
      RECT 7.95 3.385 8.12 3.555 ;
      RECT 7.89 2.585 8.06 2.755 ;
      RECT 7.83 1.415 8 1.585 ;
      RECT 7.795 8.605 7.965 8.775 ;
      RECT 7.45 2.255 7.62 2.425 ;
      RECT 7.37 1.415 7.54 1.585 ;
      RECT 7.185 3.305 7.355 3.475 ;
      RECT 6.94 2.545 7.11 2.715 ;
      RECT 6.91 1.415 7.08 1.585 ;
      RECT 6.845 3.575 7.015 3.745 ;
      RECT 6.57 2.27 6.74 2.44 ;
      RECT 6.45 1.415 6.62 1.585 ;
      RECT 6.04 2.47 6.21 2.64 ;
      RECT 5.99 1.415 6.16 1.585 ;
      RECT 5.53 1.415 5.7 1.585 ;
      RECT 5.52 2.415 5.69 2.585 ;
      RECT 5.315 2.015 5.485 2.185 ;
      RECT 5.315 3.595 5.485 3.765 ;
      RECT 5.07 1.415 5.24 1.585 ;
      RECT 5.005 2.56 5.175 2.73 ;
      RECT 4.61 1.415 4.78 1.585 ;
      RECT 4.595 2.785 4.765 2.955 ;
      RECT 4.15 1.415 4.32 1.585 ;
      RECT 3.885 3.085 4.055 3.255 ;
      RECT 3.74 1.995 3.91 2.165 ;
      RECT 3.69 1.415 3.86 1.585 ;
      RECT 2.34 8.605 2.51 8.775 ;
      RECT 1.66 8.605 1.83 8.775 ;
      RECT 1.6 7.055 1.77 7.225 ;
      RECT 1.6 7.795 1.77 7.965 ;
      RECT 1.225 6.315 1.395 6.485 ;
      RECT 0.98 8.605 1.15 8.775 ;
      RECT 0.3 8.605 0.47 8.775 ;
    LAYER li1 ;
      RECT 72.555 0 72.725 2.085 ;
      RECT 71.615 0 71.785 2.085 ;
      RECT 70.655 0 70.825 2.085 ;
      RECT 68.735 0 68.905 2.085 ;
      RECT 67.775 0 67.945 2.085 ;
      RECT 65.855 0 66.025 2.085 ;
      RECT 57.295 0 57.465 2.085 ;
      RECT 56.355 0 56.525 2.085 ;
      RECT 55.395 0 55.565 2.085 ;
      RECT 53.475 0 53.645 2.085 ;
      RECT 52.515 0 52.685 2.085 ;
      RECT 50.595 0 50.765 2.085 ;
      RECT 42.035 0 42.205 2.085 ;
      RECT 41.095 0 41.265 2.085 ;
      RECT 40.135 0 40.305 2.085 ;
      RECT 38.215 0 38.385 2.085 ;
      RECT 37.255 0 37.425 2.085 ;
      RECT 35.335 0 35.505 2.085 ;
      RECT 26.775 0 26.945 2.085 ;
      RECT 25.835 0 26.005 2.085 ;
      RECT 24.875 0 25.045 2.085 ;
      RECT 22.955 0 23.125 2.085 ;
      RECT 21.995 0 22.165 2.085 ;
      RECT 20.075 0 20.245 2.085 ;
      RECT 11.515 0 11.685 2.085 ;
      RECT 10.575 0 10.745 2.085 ;
      RECT 9.615 0 9.785 2.085 ;
      RECT 7.695 0 7.865 2.085 ;
      RECT 6.735 0 6.905 2.085 ;
      RECT 4.815 0 4.985 2.085 ;
      RECT 69.61 0 69.805 1.595 ;
      RECT 65.855 0 66.13 1.595 ;
      RECT 54.35 0 54.545 1.595 ;
      RECT 50.595 0 50.87 1.595 ;
      RECT 39.09 0 39.285 1.595 ;
      RECT 35.335 0 35.61 1.595 ;
      RECT 23.83 0 24.025 1.595 ;
      RECT 20.075 0 20.35 1.595 ;
      RECT 8.57 0 8.765 1.595 ;
      RECT 4.815 0 5.09 1.595 ;
      RECT 64.585 0 73.325 1.585 ;
      RECT 49.325 0 58.065 1.585 ;
      RECT 34.065 0 42.805 1.585 ;
      RECT 18.805 0 27.545 1.585 ;
      RECT 3.545 0 12.285 1.585 ;
      RECT 74.39 0 74.56 0.935 ;
      RECT 59.13 0 59.3 0.935 ;
      RECT 43.87 0 44.04 0.935 ;
      RECT 28.61 0 28.78 0.935 ;
      RECT 13.35 0 13.52 0.935 ;
      RECT 78.12 0 78.29 0.93 ;
      RECT 77.13 0 77.3 0.93 ;
      RECT 62.86 0 63.03 0.93 ;
      RECT 61.87 0 62.04 0.93 ;
      RECT 47.6 0 47.77 0.93 ;
      RECT 46.61 0 46.78 0.93 ;
      RECT 32.34 0 32.51 0.93 ;
      RECT 31.35 0 31.52 0.93 ;
      RECT 17.08 0 17.25 0.93 ;
      RECT 16.09 0 16.26 0.93 ;
      RECT 78.915 0 79.095 0.305 ;
      RECT 63.655 0 76.965 0.305 ;
      RECT 48.395 0 61.705 0.305 ;
      RECT 33.135 0 46.445 0.305 ;
      RECT 17.875 0 31.185 0.305 ;
      RECT 0 0 15.925 0.305 ;
      RECT 0 0 79.095 0.3 ;
      RECT 0 8.58 79.095 8.88 ;
      RECT 78.915 8.575 79.095 8.88 ;
      RECT 78.12 7.95 78.29 8.88 ;
      RECT 77.13 7.95 77.3 8.88 ;
      RECT 63.655 8.575 76.965 8.88 ;
      RECT 62.86 7.95 63.03 8.88 ;
      RECT 61.87 7.95 62.04 8.88 ;
      RECT 48.395 8.575 61.705 8.88 ;
      RECT 47.6 7.95 47.77 8.88 ;
      RECT 46.61 7.95 46.78 8.88 ;
      RECT 33.135 8.575 46.445 8.88 ;
      RECT 32.34 7.95 32.51 8.88 ;
      RECT 31.35 7.95 31.52 8.88 ;
      RECT 17.875 8.575 31.185 8.88 ;
      RECT 17.08 7.95 17.25 8.88 ;
      RECT 16.09 7.95 16.26 8.88 ;
      RECT 0 8.575 15.925 8.88 ;
      RECT 74.39 7.945 74.56 8.88 ;
      RECT 68.755 7.945 68.925 8.88 ;
      RECT 59.13 7.945 59.3 8.88 ;
      RECT 53.495 7.945 53.665 8.88 ;
      RECT 43.87 7.945 44.04 8.88 ;
      RECT 38.235 7.945 38.405 8.88 ;
      RECT 28.61 7.945 28.78 8.88 ;
      RECT 22.975 7.945 23.145 8.88 ;
      RECT 13.35 7.945 13.52 8.88 ;
      RECT 7.715 7.945 7.885 8.88 ;
      RECT 0.005 8.565 0.81 8.88 ;
      RECT 0.22 8.545 0.47 8.88 ;
      RECT 0.22 7.945 0.39 8.88 ;
      RECT 78.55 5.02 78.72 6.49 ;
      RECT 78.55 6.315 78.725 6.485 ;
      RECT 78.18 1.74 78.35 2.93 ;
      RECT 78.18 1.74 78.65 1.91 ;
      RECT 78.18 6.97 78.65 7.14 ;
      RECT 78.18 5.95 78.35 7.14 ;
      RECT 77.19 1.74 77.36 2.93 ;
      RECT 77.19 1.74 77.66 1.91 ;
      RECT 77.19 6.97 77.66 7.14 ;
      RECT 77.19 5.95 77.36 7.14 ;
      RECT 75.34 2.635 75.51 3.865 ;
      RECT 75.395 0.855 75.565 2.805 ;
      RECT 75.34 0.575 75.51 1.025 ;
      RECT 75.34 7.855 75.51 8.305 ;
      RECT 75.395 6.075 75.565 8.025 ;
      RECT 75.34 5.015 75.51 6.245 ;
      RECT 74.82 0.575 74.99 3.865 ;
      RECT 74.82 2.075 75.225 2.405 ;
      RECT 74.82 1.235 75.225 1.565 ;
      RECT 74.82 5.015 74.99 8.305 ;
      RECT 74.82 7.315 75.225 7.645 ;
      RECT 74.82 6.475 75.225 6.805 ;
      RECT 72.745 3.126 72.75 3.298 ;
      RECT 72.74 3.119 72.745 3.388 ;
      RECT 72.735 3.113 72.74 3.407 ;
      RECT 72.715 3.107 72.735 3.417 ;
      RECT 72.7 3.102 72.715 3.425 ;
      RECT 72.663 3.096 72.7 3.423 ;
      RECT 72.577 3.082 72.663 3.419 ;
      RECT 72.491 3.064 72.577 3.414 ;
      RECT 72.405 3.045 72.491 3.408 ;
      RECT 72.375 3.033 72.405 3.404 ;
      RECT 72.355 3.027 72.375 3.403 ;
      RECT 72.29 3.025 72.355 3.401 ;
      RECT 72.275 3.025 72.29 3.393 ;
      RECT 72.26 3.025 72.275 3.38 ;
      RECT 72.255 3.025 72.26 3.37 ;
      RECT 72.24 3.025 72.255 3.348 ;
      RECT 72.225 3.025 72.24 3.315 ;
      RECT 72.22 3.025 72.225 3.293 ;
      RECT 72.21 3.025 72.22 3.275 ;
      RECT 72.195 3.025 72.21 3.253 ;
      RECT 72.175 3.025 72.195 3.215 ;
      RECT 72.525 2.31 72.56 2.749 ;
      RECT 72.525 2.31 72.565 2.748 ;
      RECT 72.47 2.37 72.565 2.747 ;
      RECT 72.335 2.542 72.565 2.746 ;
      RECT 72.445 2.42 72.565 2.746 ;
      RECT 72.335 2.542 72.59 2.736 ;
      RECT 72.39 2.487 72.67 2.653 ;
      RECT 72.565 2.281 72.57 2.744 ;
      RECT 72.42 2.457 72.71 2.53 ;
      RECT 72.435 2.44 72.565 2.746 ;
      RECT 72.57 2.28 72.74 2.468 ;
      RECT 72.56 2.283 72.74 2.468 ;
      RECT 72.065 2.16 72.235 2.47 ;
      RECT 72.065 2.16 72.24 2.443 ;
      RECT 72.065 2.16 72.245 2.42 ;
      RECT 72.065 2.16 72.255 2.37 ;
      RECT 72.06 2.265 72.255 2.34 ;
      RECT 72.095 1.835 72.265 2.313 ;
      RECT 72.095 1.835 72.28 2.234 ;
      RECT 72.085 2.045 72.28 2.234 ;
      RECT 72.095 1.845 72.29 2.149 ;
      RECT 72.025 2.587 72.03 2.79 ;
      RECT 72.015 2.575 72.025 2.9 ;
      RECT 71.99 2.575 72.015 2.94 ;
      RECT 71.91 2.575 71.99 3.025 ;
      RECT 71.9 2.575 71.91 3.095 ;
      RECT 71.875 2.575 71.9 3.118 ;
      RECT 71.855 2.575 71.875 3.153 ;
      RECT 71.81 2.585 71.855 3.196 ;
      RECT 71.8 2.597 71.81 3.233 ;
      RECT 71.78 2.611 71.8 3.253 ;
      RECT 71.77 2.629 71.78 3.269 ;
      RECT 71.755 2.655 71.77 3.279 ;
      RECT 71.74 2.696 71.755 3.293 ;
      RECT 71.73 2.731 71.74 3.303 ;
      RECT 71.725 2.747 71.73 3.308 ;
      RECT 71.715 2.762 71.725 3.313 ;
      RECT 71.695 2.805 71.715 3.323 ;
      RECT 71.675 2.842 71.695 3.336 ;
      RECT 71.64 2.865 71.675 3.354 ;
      RECT 71.63 2.879 71.64 3.37 ;
      RECT 71.61 2.889 71.63 3.38 ;
      RECT 71.605 2.898 71.61 3.388 ;
      RECT 71.595 2.905 71.605 3.395 ;
      RECT 71.585 2.912 71.595 3.403 ;
      RECT 71.57 2.922 71.585 3.411 ;
      RECT 71.56 2.936 71.57 3.421 ;
      RECT 71.55 2.948 71.56 3.433 ;
      RECT 71.535 2.97 71.55 3.446 ;
      RECT 71.525 2.992 71.535 3.457 ;
      RECT 71.515 3.012 71.525 3.466 ;
      RECT 71.51 3.027 71.515 3.473 ;
      RECT 71.48 3.06 71.51 3.487 ;
      RECT 71.47 3.095 71.48 3.502 ;
      RECT 71.465 3.102 71.47 3.508 ;
      RECT 71.445 3.117 71.465 3.515 ;
      RECT 71.44 3.132 71.445 3.523 ;
      RECT 71.435 3.141 71.44 3.528 ;
      RECT 71.42 3.147 71.435 3.535 ;
      RECT 71.415 3.153 71.42 3.543 ;
      RECT 71.41 3.157 71.415 3.55 ;
      RECT 71.405 3.161 71.41 3.56 ;
      RECT 71.395 3.166 71.405 3.57 ;
      RECT 71.375 3.177 71.395 3.598 ;
      RECT 71.36 3.189 71.375 3.625 ;
      RECT 71.34 3.202 71.36 3.65 ;
      RECT 71.32 3.217 71.34 3.674 ;
      RECT 71.305 3.232 71.32 3.689 ;
      RECT 71.3 3.243 71.305 3.698 ;
      RECT 71.235 3.288 71.3 3.708 ;
      RECT 71.2 3.347 71.235 3.721 ;
      RECT 71.195 3.37 71.2 3.727 ;
      RECT 71.19 3.377 71.195 3.729 ;
      RECT 71.175 3.387 71.19 3.732 ;
      RECT 71.145 3.412 71.175 3.736 ;
      RECT 71.14 3.43 71.145 3.74 ;
      RECT 71.135 3.437 71.14 3.741 ;
      RECT 71.115 3.445 71.135 3.745 ;
      RECT 71.105 3.452 71.115 3.749 ;
      RECT 71.061 3.463 71.105 3.756 ;
      RECT 70.975 3.491 71.061 3.772 ;
      RECT 70.915 3.515 70.975 3.79 ;
      RECT 70.87 3.525 70.915 3.804 ;
      RECT 70.811 3.533 70.87 3.818 ;
      RECT 70.725 3.54 70.811 3.837 ;
      RECT 70.7 3.545 70.725 3.852 ;
      RECT 70.62 3.548 70.7 3.855 ;
      RECT 70.54 3.552 70.62 3.842 ;
      RECT 70.531 3.555 70.54 3.827 ;
      RECT 70.445 3.555 70.531 3.812 ;
      RECT 70.385 3.557 70.445 3.789 ;
      RECT 70.381 3.56 70.385 3.779 ;
      RECT 70.295 3.56 70.381 3.764 ;
      RECT 70.22 3.56 70.295 3.74 ;
      RECT 71.535 2.569 71.545 2.745 ;
      RECT 71.49 2.536 71.535 2.745 ;
      RECT 71.445 2.487 71.49 2.745 ;
      RECT 71.415 2.457 71.445 2.746 ;
      RECT 71.41 2.44 71.415 2.747 ;
      RECT 71.385 2.42 71.41 2.748 ;
      RECT 71.37 2.395 71.385 2.749 ;
      RECT 71.365 2.382 71.37 2.75 ;
      RECT 71.36 2.376 71.365 2.748 ;
      RECT 71.355 2.368 71.36 2.742 ;
      RECT 71.33 2.36 71.355 2.722 ;
      RECT 71.31 2.349 71.33 2.693 ;
      RECT 71.28 2.334 71.31 2.664 ;
      RECT 71.26 2.32 71.28 2.636 ;
      RECT 71.25 2.314 71.26 2.615 ;
      RECT 71.245 2.311 71.25 2.598 ;
      RECT 71.24 2.308 71.245 2.583 ;
      RECT 71.225 2.303 71.24 2.548 ;
      RECT 71.22 2.299 71.225 2.515 ;
      RECT 71.2 2.294 71.22 2.491 ;
      RECT 71.17 2.286 71.2 2.456 ;
      RECT 71.155 2.28 71.17 2.433 ;
      RECT 71.115 2.273 71.155 2.418 ;
      RECT 71.09 2.265 71.115 2.398 ;
      RECT 71.07 2.26 71.09 2.388 ;
      RECT 71.035 2.254 71.07 2.383 ;
      RECT 70.99 2.245 71.035 2.382 ;
      RECT 70.96 2.241 70.99 2.384 ;
      RECT 70.875 2.249 70.96 2.388 ;
      RECT 70.805 2.26 70.875 2.41 ;
      RECT 70.792 2.266 70.805 2.433 ;
      RECT 70.706 2.273 70.792 2.455 ;
      RECT 70.62 2.285 70.706 2.492 ;
      RECT 70.62 2.662 70.63 2.9 ;
      RECT 70.615 2.291 70.62 2.515 ;
      RECT 70.61 2.547 70.62 2.9 ;
      RECT 70.61 2.292 70.615 2.52 ;
      RECT 70.605 2.293 70.61 2.9 ;
      RECT 70.581 2.295 70.605 2.901 ;
      RECT 70.495 2.303 70.581 2.903 ;
      RECT 70.475 2.317 70.495 2.906 ;
      RECT 70.47 2.345 70.475 2.907 ;
      RECT 70.465 2.357 70.47 2.908 ;
      RECT 70.46 2.372 70.465 2.909 ;
      RECT 70.45 2.402 70.46 2.91 ;
      RECT 70.445 2.44 70.45 2.908 ;
      RECT 70.44 2.46 70.445 2.903 ;
      RECT 70.425 2.495 70.44 2.888 ;
      RECT 70.415 2.547 70.425 2.868 ;
      RECT 70.41 2.577 70.415 2.856 ;
      RECT 70.395 2.59 70.41 2.839 ;
      RECT 70.37 2.594 70.395 2.806 ;
      RECT 70.355 2.592 70.37 2.783 ;
      RECT 70.34 2.591 70.355 2.78 ;
      RECT 70.28 2.589 70.34 2.778 ;
      RECT 70.27 2.587 70.28 2.773 ;
      RECT 70.23 2.586 70.27 2.77 ;
      RECT 70.16 2.583 70.23 2.768 ;
      RECT 70.105 2.581 70.16 2.763 ;
      RECT 70.035 2.575 70.105 2.758 ;
      RECT 70.026 2.575 70.035 2.755 ;
      RECT 69.94 2.575 70.026 2.75 ;
      RECT 69.935 2.575 69.94 2.745 ;
      RECT 71.24 1.81 71.415 2.16 ;
      RECT 71.24 1.825 71.425 2.158 ;
      RECT 71.215 1.775 71.36 2.155 ;
      RECT 71.195 1.776 71.36 2.148 ;
      RECT 71.185 1.777 71.37 2.143 ;
      RECT 71.155 1.778 71.37 2.13 ;
      RECT 71.105 1.779 71.37 2.106 ;
      RECT 71.1 1.781 71.37 2.091 ;
      RECT 71.1 1.847 71.43 2.085 ;
      RECT 71.08 1.788 71.385 2.065 ;
      RECT 71.07 1.797 71.395 1.92 ;
      RECT 71.08 1.792 71.395 2.065 ;
      RECT 71.1 1.782 71.385 2.091 ;
      RECT 70.685 3.107 70.855 3.395 ;
      RECT 70.68 3.125 70.865 3.39 ;
      RECT 70.645 3.133 70.93 3.31 ;
      RECT 70.645 3.133 71.016 3.3 ;
      RECT 70.645 3.133 71.07 3.246 ;
      RECT 70.93 3.03 71.1 3.214 ;
      RECT 70.645 3.185 71.105 3.202 ;
      RECT 70.63 3.155 71.1 3.198 ;
      RECT 70.89 3.037 70.93 3.349 ;
      RECT 70.77 3.074 71.1 3.214 ;
      RECT 70.865 3.049 70.89 3.375 ;
      RECT 70.855 3.056 71.1 3.214 ;
      RECT 70.986 2.52 71.055 2.779 ;
      RECT 70.986 2.575 71.06 2.778 ;
      RECT 70.9 2.575 71.06 2.777 ;
      RECT 70.895 2.575 71.065 2.77 ;
      RECT 70.885 2.52 71.055 2.765 ;
      RECT 70.265 1.819 70.44 2.12 ;
      RECT 70.25 1.807 70.265 2.105 ;
      RECT 70.22 1.806 70.25 2.058 ;
      RECT 70.22 1.824 70.445 2.053 ;
      RECT 70.205 1.808 70.265 2.018 ;
      RECT 70.2 1.83 70.455 1.918 ;
      RECT 70.2 1.813 70.351 1.918 ;
      RECT 70.2 1.815 70.355 1.918 ;
      RECT 70.205 1.811 70.351 2.018 ;
      RECT 70.31 3.047 70.315 3.395 ;
      RECT 70.3 3.037 70.31 3.401 ;
      RECT 70.265 3.027 70.3 3.403 ;
      RECT 70.227 3.022 70.265 3.407 ;
      RECT 70.141 3.015 70.227 3.414 ;
      RECT 70.055 3.005 70.141 3.424 ;
      RECT 70.01 3 70.055 3.432 ;
      RECT 70.006 3 70.01 3.436 ;
      RECT 69.92 3 70.006 3.443 ;
      RECT 69.905 3 69.92 3.443 ;
      RECT 69.895 2.998 69.905 3.415 ;
      RECT 69.885 2.994 69.895 3.358 ;
      RECT 69.865 2.988 69.885 3.29 ;
      RECT 69.86 2.984 69.865 3.238 ;
      RECT 69.85 2.983 69.86 3.205 ;
      RECT 69.8 2.981 69.85 3.19 ;
      RECT 69.775 2.979 69.8 3.185 ;
      RECT 69.732 2.977 69.775 3.181 ;
      RECT 69.646 2.973 69.732 3.169 ;
      RECT 69.56 2.968 69.646 3.153 ;
      RECT 69.53 2.965 69.56 3.14 ;
      RECT 69.505 2.964 69.53 3.128 ;
      RECT 69.5 2.964 69.505 3.118 ;
      RECT 69.46 2.963 69.5 3.11 ;
      RECT 69.445 2.962 69.46 3.103 ;
      RECT 69.395 2.961 69.445 3.095 ;
      RECT 69.393 2.96 69.395 3.09 ;
      RECT 69.307 2.958 69.393 3.09 ;
      RECT 69.221 2.953 69.307 3.09 ;
      RECT 69.135 2.949 69.221 3.09 ;
      RECT 69.086 2.945 69.135 3.088 ;
      RECT 69 2.942 69.086 3.083 ;
      RECT 68.977 2.939 69 3.079 ;
      RECT 68.891 2.936 68.977 3.074 ;
      RECT 68.805 2.932 68.891 3.065 ;
      RECT 68.78 2.925 68.805 3.06 ;
      RECT 68.72 2.89 68.78 3.057 ;
      RECT 68.7 2.815 68.72 3.054 ;
      RECT 68.695 2.757 68.7 3.053 ;
      RECT 68.67 2.697 68.695 3.052 ;
      RECT 68.595 2.575 68.67 3.048 ;
      RECT 68.585 2.575 68.595 3.04 ;
      RECT 68.57 2.575 68.585 3.03 ;
      RECT 68.555 2.575 68.57 3 ;
      RECT 68.54 2.575 68.555 2.945 ;
      RECT 68.525 2.575 68.54 2.883 ;
      RECT 68.5 2.575 68.525 2.808 ;
      RECT 68.495 2.575 68.5 2.758 ;
      RECT 69.84 2.12 69.86 2.429 ;
      RECT 69.826 2.122 69.875 2.426 ;
      RECT 69.826 2.127 69.895 2.417 ;
      RECT 69.74 2.125 69.875 2.411 ;
      RECT 69.74 2.133 69.93 2.394 ;
      RECT 69.705 2.135 69.93 2.393 ;
      RECT 69.675 2.143 69.93 2.384 ;
      RECT 69.665 2.148 69.95 2.37 ;
      RECT 69.705 2.138 69.95 2.37 ;
      RECT 69.705 2.141 69.96 2.358 ;
      RECT 69.675 2.143 69.97 2.345 ;
      RECT 69.675 2.147 69.98 2.288 ;
      RECT 69.665 2.152 69.985 2.203 ;
      RECT 69.826 2.12 69.86 2.426 ;
      RECT 69.705 7.855 69.875 8.305 ;
      RECT 69.76 6.075 69.93 8.025 ;
      RECT 69.705 5.015 69.875 6.245 ;
      RECT 69.265 2.223 69.27 2.435 ;
      RECT 69.14 2.22 69.155 2.435 ;
      RECT 68.605 2.25 68.675 2.435 ;
      RECT 68.49 2.25 68.525 2.43 ;
      RECT 69.611 2.552 69.63 2.746 ;
      RECT 69.525 2.507 69.611 2.747 ;
      RECT 69.515 2.46 69.525 2.749 ;
      RECT 69.51 2.44 69.515 2.75 ;
      RECT 69.49 2.405 69.51 2.751 ;
      RECT 69.475 2.355 69.49 2.752 ;
      RECT 69.455 2.292 69.475 2.753 ;
      RECT 69.445 2.255 69.455 2.754 ;
      RECT 69.43 2.244 69.445 2.755 ;
      RECT 69.425 2.236 69.43 2.753 ;
      RECT 69.415 2.235 69.425 2.745 ;
      RECT 69.385 2.232 69.415 2.724 ;
      RECT 69.31 2.227 69.385 2.669 ;
      RECT 69.295 2.223 69.31 2.615 ;
      RECT 69.285 2.223 69.295 2.51 ;
      RECT 69.27 2.223 69.285 2.443 ;
      RECT 69.255 2.223 69.265 2.433 ;
      RECT 69.2 2.222 69.255 2.43 ;
      RECT 69.155 2.22 69.2 2.433 ;
      RECT 69.127 2.22 69.14 2.436 ;
      RECT 69.041 2.224 69.127 2.438 ;
      RECT 68.955 2.23 69.041 2.443 ;
      RECT 68.935 2.234 68.955 2.445 ;
      RECT 68.933 2.235 68.935 2.444 ;
      RECT 68.847 2.237 68.933 2.443 ;
      RECT 68.761 2.242 68.847 2.44 ;
      RECT 68.675 2.247 68.761 2.437 ;
      RECT 68.525 2.25 68.605 2.433 ;
      RECT 69.185 5.015 69.355 8.305 ;
      RECT 69.185 7.315 69.59 7.645 ;
      RECT 69.185 6.475 69.59 6.805 ;
      RECT 69.301 3.225 69.35 3.559 ;
      RECT 69.301 3.225 69.355 3.558 ;
      RECT 69.215 3.225 69.355 3.557 ;
      RECT 68.99 3.333 69.36 3.555 ;
      RECT 69.215 3.225 69.385 3.548 ;
      RECT 69.185 3.237 69.39 3.539 ;
      RECT 69.17 3.255 69.395 3.536 ;
      RECT 68.985 3.339 69.395 3.463 ;
      RECT 68.98 3.346 69.395 3.423 ;
      RECT 68.995 3.312 69.395 3.536 ;
      RECT 69.156 3.258 69.36 3.555 ;
      RECT 69.07 3.278 69.395 3.536 ;
      RECT 69.17 3.252 69.39 3.539 ;
      RECT 68.94 2.576 69.13 2.77 ;
      RECT 68.935 2.578 69.13 2.769 ;
      RECT 68.93 2.582 69.145 2.766 ;
      RECT 68.945 2.575 69.145 2.766 ;
      RECT 68.93 2.685 69.15 2.761 ;
      RECT 68.225 3.185 68.316 3.483 ;
      RECT 68.22 3.187 68.395 3.478 ;
      RECT 68.225 3.185 68.395 3.478 ;
      RECT 68.22 3.191 68.415 3.476 ;
      RECT 68.22 3.246 68.455 3.475 ;
      RECT 68.22 3.281 68.47 3.469 ;
      RECT 68.22 3.315 68.48 3.459 ;
      RECT 68.21 3.195 68.415 3.31 ;
      RECT 68.21 3.215 68.43 3.31 ;
      RECT 68.21 3.198 68.42 3.31 ;
      RECT 68.435 1.966 68.44 2.028 ;
      RECT 68.43 1.888 68.435 2.051 ;
      RECT 68.425 1.845 68.43 2.062 ;
      RECT 68.42 1.835 68.425 2.074 ;
      RECT 68.415 1.835 68.42 2.083 ;
      RECT 68.39 1.835 68.415 2.115 ;
      RECT 68.385 1.835 68.39 2.148 ;
      RECT 68.37 1.835 68.385 2.173 ;
      RECT 68.36 1.835 68.37 2.2 ;
      RECT 68.355 1.835 68.36 2.213 ;
      RECT 68.35 1.835 68.355 2.228 ;
      RECT 68.34 1.835 68.35 2.243 ;
      RECT 68.335 1.835 68.34 2.263 ;
      RECT 68.31 1.835 68.335 2.298 ;
      RECT 68.265 1.835 68.31 2.343 ;
      RECT 68.255 1.835 68.265 2.356 ;
      RECT 68.17 1.92 68.255 2.363 ;
      RECT 68.135 2.042 68.17 2.372 ;
      RECT 68.13 2.082 68.135 2.376 ;
      RECT 68.11 2.105 68.13 2.378 ;
      RECT 68.105 2.135 68.11 2.381 ;
      RECT 68.095 2.147 68.105 2.382 ;
      RECT 68.05 2.17 68.095 2.387 ;
      RECT 68.01 2.2 68.05 2.395 ;
      RECT 67.975 2.212 68.01 2.401 ;
      RECT 67.97 2.217 67.975 2.405 ;
      RECT 67.9 2.227 67.97 2.412 ;
      RECT 67.86 2.237 67.9 2.422 ;
      RECT 67.84 2.242 67.86 2.428 ;
      RECT 67.83 2.246 67.84 2.433 ;
      RECT 67.825 2.249 67.83 2.436 ;
      RECT 67.815 2.25 67.825 2.437 ;
      RECT 67.79 2.252 67.815 2.441 ;
      RECT 67.78 2.257 67.79 2.444 ;
      RECT 67.735 2.265 67.78 2.445 ;
      RECT 67.61 2.27 67.735 2.445 ;
      RECT 68.165 2.567 68.185 2.749 ;
      RECT 68.116 2.552 68.165 2.748 ;
      RECT 68.03 2.567 68.185 2.746 ;
      RECT 68.015 2.567 68.185 2.745 ;
      RECT 67.98 2.545 68.15 2.73 ;
      RECT 68.05 3.565 68.065 3.774 ;
      RECT 68.05 3.573 68.07 3.773 ;
      RECT 67.995 3.573 68.07 3.772 ;
      RECT 67.975 3.577 68.075 3.77 ;
      RECT 67.955 3.527 67.995 3.769 ;
      RECT 67.9 3.585 68.08 3.767 ;
      RECT 67.865 3.542 67.995 3.765 ;
      RECT 67.861 3.545 68.05 3.764 ;
      RECT 67.775 3.553 68.05 3.762 ;
      RECT 67.775 3.597 68.085 3.755 ;
      RECT 67.765 3.69 68.085 3.753 ;
      RECT 67.775 3.609 68.09 3.738 ;
      RECT 67.775 3.63 68.105 3.708 ;
      RECT 67.775 3.657 68.11 3.678 ;
      RECT 67.9 3.535 67.995 3.767 ;
      RECT 67.53 2.58 67.535 3.118 ;
      RECT 67.335 2.91 67.34 3.105 ;
      RECT 65.635 2.575 65.65 2.955 ;
      RECT 67.7 2.575 67.705 2.745 ;
      RECT 67.695 2.575 67.7 2.755 ;
      RECT 67.69 2.575 67.695 2.768 ;
      RECT 67.665 2.575 67.69 2.81 ;
      RECT 67.64 2.575 67.665 2.883 ;
      RECT 67.625 2.575 67.64 2.935 ;
      RECT 67.62 2.575 67.625 2.965 ;
      RECT 67.595 2.575 67.62 3.005 ;
      RECT 67.58 2.575 67.595 3.06 ;
      RECT 67.575 2.575 67.58 3.093 ;
      RECT 67.55 2.575 67.575 3.113 ;
      RECT 67.535 2.575 67.55 3.119 ;
      RECT 67.465 2.61 67.53 3.115 ;
      RECT 67.415 2.665 67.465 3.11 ;
      RECT 67.405 2.697 67.415 3.108 ;
      RECT 67.4 2.722 67.405 3.108 ;
      RECT 67.38 2.795 67.4 3.108 ;
      RECT 67.37 2.875 67.38 3.107 ;
      RECT 67.355 2.905 67.37 3.107 ;
      RECT 67.34 2.91 67.355 3.106 ;
      RECT 67.28 2.912 67.335 3.103 ;
      RECT 67.25 2.917 67.28 3.099 ;
      RECT 67.248 2.92 67.25 3.098 ;
      RECT 67.162 2.922 67.248 3.095 ;
      RECT 67.076 2.928 67.162 3.089 ;
      RECT 66.99 2.933 67.076 3.083 ;
      RECT 66.917 2.938 66.99 3.084 ;
      RECT 66.831 2.944 66.917 3.092 ;
      RECT 66.745 2.95 66.831 3.101 ;
      RECT 66.725 2.954 66.745 3.106 ;
      RECT 66.678 2.956 66.725 3.109 ;
      RECT 66.592 2.961 66.678 3.115 ;
      RECT 66.506 2.966 66.592 3.124 ;
      RECT 66.42 2.972 66.506 3.132 ;
      RECT 66.335 2.97 66.42 3.141 ;
      RECT 66.331 2.965 66.335 3.145 ;
      RECT 66.245 2.96 66.331 3.137 ;
      RECT 66.181 2.951 66.245 3.125 ;
      RECT 66.095 2.942 66.181 3.112 ;
      RECT 66.071 2.935 66.095 3.103 ;
      RECT 65.985 2.929 66.071 3.09 ;
      RECT 65.945 2.922 65.985 3.076 ;
      RECT 65.94 2.912 65.945 3.072 ;
      RECT 65.93 2.9 65.94 3.071 ;
      RECT 65.91 2.87 65.93 3.068 ;
      RECT 65.855 2.79 65.91 3.062 ;
      RECT 65.835 2.709 65.855 3.057 ;
      RECT 65.815 2.667 65.835 3.053 ;
      RECT 65.79 2.62 65.815 3.047 ;
      RECT 65.785 2.595 65.79 3.044 ;
      RECT 65.75 2.575 65.785 3.039 ;
      RECT 65.741 2.575 65.75 3.032 ;
      RECT 65.655 2.575 65.741 3.002 ;
      RECT 65.65 2.575 65.655 2.965 ;
      RECT 65.615 2.575 65.635 2.887 ;
      RECT 65.61 2.617 65.615 2.852 ;
      RECT 65.605 2.692 65.61 2.808 ;
      RECT 67.055 2.497 67.23 2.745 ;
      RECT 67.055 2.497 67.235 2.743 ;
      RECT 67.05 2.529 67.235 2.703 ;
      RECT 67.08 2.47 67.25 2.69 ;
      RECT 67.045 2.547 67.25 2.623 ;
      RECT 66.355 2.01 66.525 2.185 ;
      RECT 66.355 2.01 66.697 2.177 ;
      RECT 66.355 2.01 66.78 2.171 ;
      RECT 66.355 2.01 66.815 2.167 ;
      RECT 66.355 2.01 66.835 2.166 ;
      RECT 66.355 2.01 66.921 2.162 ;
      RECT 66.815 1.835 66.985 2.157 ;
      RECT 66.39 1.942 67.015 2.155 ;
      RECT 66.38 1.997 67.02 2.153 ;
      RECT 66.355 2.033 67.03 2.148 ;
      RECT 66.355 2.06 67.035 2.078 ;
      RECT 66.42 1.885 66.995 2.155 ;
      RECT 66.611 1.87 66.995 2.155 ;
      RECT 66.445 1.873 66.995 2.155 ;
      RECT 66.525 1.871 66.611 2.182 ;
      RECT 66.611 1.868 66.99 2.155 ;
      RECT 66.795 1.845 66.99 2.155 ;
      RECT 66.697 1.866 66.99 2.155 ;
      RECT 66.78 1.86 66.795 2.168 ;
      RECT 66.93 3.225 66.935 3.425 ;
      RECT 66.395 3.29 66.44 3.425 ;
      RECT 66.965 3.225 66.985 3.398 ;
      RECT 66.935 3.225 66.965 3.413 ;
      RECT 66.87 3.225 66.93 3.45 ;
      RECT 66.855 3.225 66.87 3.48 ;
      RECT 66.84 3.225 66.855 3.493 ;
      RECT 66.82 3.225 66.84 3.508 ;
      RECT 66.815 3.225 66.82 3.517 ;
      RECT 66.805 3.229 66.815 3.522 ;
      RECT 66.79 3.239 66.805 3.533 ;
      RECT 66.765 3.255 66.79 3.543 ;
      RECT 66.755 3.269 66.765 3.545 ;
      RECT 66.735 3.281 66.755 3.542 ;
      RECT 66.705 3.302 66.735 3.536 ;
      RECT 66.695 3.314 66.705 3.531 ;
      RECT 66.685 3.312 66.695 3.528 ;
      RECT 66.67 3.311 66.685 3.523 ;
      RECT 66.665 3.31 66.67 3.518 ;
      RECT 66.63 3.308 66.665 3.508 ;
      RECT 66.61 3.305 66.63 3.49 ;
      RECT 66.6 3.303 66.61 3.485 ;
      RECT 66.59 3.302 66.6 3.48 ;
      RECT 66.555 3.3 66.59 3.468 ;
      RECT 66.5 3.296 66.555 3.448 ;
      RECT 66.49 3.294 66.5 3.433 ;
      RECT 66.485 3.294 66.49 3.428 ;
      RECT 66.44 3.292 66.485 3.425 ;
      RECT 66.345 3.29 66.395 3.429 ;
      RECT 66.335 3.291 66.345 3.434 ;
      RECT 66.275 3.298 66.335 3.448 ;
      RECT 66.25 3.306 66.275 3.468 ;
      RECT 66.24 3.31 66.25 3.48 ;
      RECT 66.235 3.311 66.24 3.485 ;
      RECT 66.22 3.313 66.235 3.488 ;
      RECT 66.205 3.315 66.22 3.493 ;
      RECT 66.2 3.315 66.205 3.496 ;
      RECT 66.155 3.32 66.2 3.507 ;
      RECT 66.15 3.324 66.155 3.519 ;
      RECT 66.125 3.32 66.15 3.523 ;
      RECT 66.115 3.316 66.125 3.527 ;
      RECT 66.105 3.315 66.115 3.531 ;
      RECT 66.09 3.305 66.105 3.537 ;
      RECT 66.085 3.293 66.09 3.541 ;
      RECT 66.08 3.29 66.085 3.542 ;
      RECT 66.075 3.287 66.08 3.544 ;
      RECT 66.06 3.275 66.075 3.543 ;
      RECT 66.045 3.257 66.06 3.54 ;
      RECT 66.025 3.236 66.045 3.533 ;
      RECT 65.96 3.225 66.025 3.505 ;
      RECT 65.956 3.225 65.96 3.484 ;
      RECT 65.87 3.225 65.956 3.454 ;
      RECT 65.855 3.225 65.87 3.41 ;
      RECT 66.43 2.325 66.435 2.56 ;
      RECT 65.56 2.241 65.565 2.445 ;
      RECT 66.14 2.27 66.145 2.425 ;
      RECT 66.06 2.25 66.065 2.425 ;
      RECT 66.73 2.392 66.745 2.745 ;
      RECT 66.656 2.377 66.73 2.745 ;
      RECT 66.57 2.36 66.656 2.745 ;
      RECT 66.56 2.35 66.57 2.743 ;
      RECT 66.555 2.348 66.56 2.738 ;
      RECT 66.54 2.346 66.555 2.724 ;
      RECT 66.47 2.338 66.54 2.664 ;
      RECT 66.45 2.329 66.47 2.598 ;
      RECT 66.445 2.326 66.45 2.578 ;
      RECT 66.435 2.325 66.445 2.568 ;
      RECT 66.425 2.325 66.43 2.552 ;
      RECT 66.415 2.324 66.425 2.542 ;
      RECT 66.405 2.322 66.415 2.53 ;
      RECT 66.39 2.319 66.405 2.51 ;
      RECT 66.38 2.317 66.39 2.495 ;
      RECT 66.36 2.314 66.38 2.483 ;
      RECT 66.355 2.312 66.36 2.473 ;
      RECT 66.33 2.31 66.355 2.46 ;
      RECT 66.3 2.305 66.33 2.445 ;
      RECT 66.22 2.296 66.3 2.436 ;
      RECT 66.175 2.285 66.22 2.429 ;
      RECT 66.155 2.276 66.175 2.426 ;
      RECT 66.145 2.271 66.155 2.425 ;
      RECT 66.1 2.265 66.14 2.425 ;
      RECT 66.085 2.257 66.1 2.425 ;
      RECT 66.065 2.252 66.085 2.425 ;
      RECT 66.045 2.249 66.06 2.425 ;
      RECT 65.962 2.248 66.045 2.424 ;
      RECT 65.876 2.247 65.962 2.42 ;
      RECT 65.79 2.245 65.876 2.417 ;
      RECT 65.737 2.244 65.79 2.419 ;
      RECT 65.651 2.243 65.737 2.428 ;
      RECT 65.565 2.242 65.651 2.44 ;
      RECT 65.545 2.241 65.56 2.448 ;
      RECT 65.465 2.24 65.545 2.46 ;
      RECT 65.44 2.24 65.465 2.473 ;
      RECT 65.415 2.24 65.44 2.488 ;
      RECT 65.41 2.24 65.415 2.51 ;
      RECT 65.405 2.24 65.41 2.528 ;
      RECT 65.4 2.24 65.405 2.545 ;
      RECT 65.395 2.24 65.4 2.558 ;
      RECT 65.39 2.24 65.395 2.568 ;
      RECT 65.35 2.24 65.39 2.653 ;
      RECT 65.335 2.24 65.35 2.738 ;
      RECT 65.325 2.241 65.335 2.75 ;
      RECT 65.29 2.246 65.325 2.755 ;
      RECT 65.25 2.255 65.29 2.755 ;
      RECT 65.235 2.265 65.25 2.755 ;
      RECT 65.23 2.275 65.235 2.755 ;
      RECT 65.21 2.302 65.23 2.755 ;
      RECT 65.16 2.385 65.21 2.755 ;
      RECT 65.155 2.447 65.16 2.755 ;
      RECT 65.145 2.46 65.155 2.755 ;
      RECT 65.135 2.482 65.145 2.755 ;
      RECT 65.125 2.507 65.135 2.75 ;
      RECT 65.12 2.545 65.125 2.743 ;
      RECT 65.11 2.655 65.12 2.738 ;
      RECT 66.505 3.576 66.52 3.835 ;
      RECT 66.505 3.591 66.525 3.834 ;
      RECT 66.421 3.591 66.525 3.832 ;
      RECT 66.421 3.605 66.53 3.831 ;
      RECT 66.335 3.647 66.535 3.828 ;
      RECT 66.33 3.59 66.52 3.823 ;
      RECT 66.33 3.661 66.54 3.82 ;
      RECT 66.325 3.692 66.54 3.818 ;
      RECT 66.33 3.689 66.555 3.808 ;
      RECT 66.325 3.735 66.57 3.793 ;
      RECT 66.325 3.763 66.575 3.778 ;
      RECT 66.335 3.565 66.505 3.828 ;
      RECT 66.095 2.575 66.265 2.745 ;
      RECT 66.06 2.575 66.265 2.74 ;
      RECT 66.05 2.575 66.265 2.733 ;
      RECT 66.045 2.56 66.215 2.73 ;
      RECT 64.875 3.097 65.14 3.54 ;
      RECT 64.87 3.068 65.085 3.538 ;
      RECT 64.865 3.222 65.145 3.533 ;
      RECT 64.87 3.117 65.145 3.533 ;
      RECT 64.87 3.128 65.155 3.52 ;
      RECT 64.87 3.075 65.115 3.538 ;
      RECT 64.875 3.062 65.085 3.54 ;
      RECT 64.875 3.06 65.035 3.54 ;
      RECT 64.976 3.052 65.035 3.54 ;
      RECT 64.89 3.053 65.035 3.54 ;
      RECT 64.976 3.051 65.025 3.54 ;
      RECT 64.78 1.866 64.955 2.165 ;
      RECT 64.83 1.828 64.955 2.165 ;
      RECT 64.815 1.83 65.041 2.157 ;
      RECT 64.815 1.833 65.08 2.144 ;
      RECT 64.815 1.834 65.09 2.13 ;
      RECT 64.77 1.885 65.09 2.12 ;
      RECT 64.815 1.835 65.095 2.115 ;
      RECT 64.77 2.045 65.1 2.105 ;
      RECT 64.755 1.905 65.095 2.045 ;
      RECT 64.75 1.921 65.095 1.985 ;
      RECT 64.795 1.845 65.095 2.115 ;
      RECT 64.83 1.826 64.916 2.165 ;
      RECT 63.29 5.02 63.46 6.49 ;
      RECT 63.29 6.315 63.465 6.485 ;
      RECT 62.92 1.74 63.09 2.93 ;
      RECT 62.92 1.74 63.39 1.91 ;
      RECT 62.92 6.97 63.39 7.14 ;
      RECT 62.92 5.95 63.09 7.14 ;
      RECT 61.93 1.74 62.1 2.93 ;
      RECT 61.93 1.74 62.4 1.91 ;
      RECT 61.93 6.97 62.4 7.14 ;
      RECT 61.93 5.95 62.1 7.14 ;
      RECT 60.08 2.635 60.25 3.865 ;
      RECT 60.135 0.855 60.305 2.805 ;
      RECT 60.08 0.575 60.25 1.025 ;
      RECT 60.08 7.855 60.25 8.305 ;
      RECT 60.135 6.075 60.305 8.025 ;
      RECT 60.08 5.015 60.25 6.245 ;
      RECT 59.56 0.575 59.73 3.865 ;
      RECT 59.56 2.075 59.965 2.405 ;
      RECT 59.56 1.235 59.965 1.565 ;
      RECT 59.56 5.015 59.73 8.305 ;
      RECT 59.56 7.315 59.965 7.645 ;
      RECT 59.56 6.475 59.965 6.805 ;
      RECT 57.485 3.126 57.49 3.298 ;
      RECT 57.48 3.119 57.485 3.388 ;
      RECT 57.475 3.113 57.48 3.407 ;
      RECT 57.455 3.107 57.475 3.417 ;
      RECT 57.44 3.102 57.455 3.425 ;
      RECT 57.403 3.096 57.44 3.423 ;
      RECT 57.317 3.082 57.403 3.419 ;
      RECT 57.231 3.064 57.317 3.414 ;
      RECT 57.145 3.045 57.231 3.408 ;
      RECT 57.115 3.033 57.145 3.404 ;
      RECT 57.095 3.027 57.115 3.403 ;
      RECT 57.03 3.025 57.095 3.401 ;
      RECT 57.015 3.025 57.03 3.393 ;
      RECT 57 3.025 57.015 3.38 ;
      RECT 56.995 3.025 57 3.37 ;
      RECT 56.98 3.025 56.995 3.348 ;
      RECT 56.965 3.025 56.98 3.315 ;
      RECT 56.96 3.025 56.965 3.293 ;
      RECT 56.95 3.025 56.96 3.275 ;
      RECT 56.935 3.025 56.95 3.253 ;
      RECT 56.915 3.025 56.935 3.215 ;
      RECT 57.265 2.31 57.3 2.749 ;
      RECT 57.265 2.31 57.305 2.748 ;
      RECT 57.21 2.37 57.305 2.747 ;
      RECT 57.075 2.542 57.305 2.746 ;
      RECT 57.185 2.42 57.305 2.746 ;
      RECT 57.075 2.542 57.33 2.736 ;
      RECT 57.13 2.487 57.41 2.653 ;
      RECT 57.305 2.281 57.31 2.744 ;
      RECT 57.16 2.457 57.45 2.53 ;
      RECT 57.175 2.44 57.305 2.746 ;
      RECT 57.31 2.28 57.48 2.468 ;
      RECT 57.3 2.283 57.48 2.468 ;
      RECT 56.805 2.16 56.975 2.47 ;
      RECT 56.805 2.16 56.98 2.443 ;
      RECT 56.805 2.16 56.985 2.42 ;
      RECT 56.805 2.16 56.995 2.37 ;
      RECT 56.8 2.265 56.995 2.34 ;
      RECT 56.835 1.835 57.005 2.313 ;
      RECT 56.835 1.835 57.02 2.234 ;
      RECT 56.825 2.045 57.02 2.234 ;
      RECT 56.835 1.845 57.03 2.149 ;
      RECT 56.765 2.587 56.77 2.79 ;
      RECT 56.755 2.575 56.765 2.9 ;
      RECT 56.73 2.575 56.755 2.94 ;
      RECT 56.65 2.575 56.73 3.025 ;
      RECT 56.64 2.575 56.65 3.095 ;
      RECT 56.615 2.575 56.64 3.118 ;
      RECT 56.595 2.575 56.615 3.153 ;
      RECT 56.55 2.585 56.595 3.196 ;
      RECT 56.54 2.597 56.55 3.233 ;
      RECT 56.52 2.611 56.54 3.253 ;
      RECT 56.51 2.629 56.52 3.269 ;
      RECT 56.495 2.655 56.51 3.279 ;
      RECT 56.48 2.696 56.495 3.293 ;
      RECT 56.47 2.731 56.48 3.303 ;
      RECT 56.465 2.747 56.47 3.308 ;
      RECT 56.455 2.762 56.465 3.313 ;
      RECT 56.435 2.805 56.455 3.323 ;
      RECT 56.415 2.842 56.435 3.336 ;
      RECT 56.38 2.865 56.415 3.354 ;
      RECT 56.37 2.879 56.38 3.37 ;
      RECT 56.35 2.889 56.37 3.38 ;
      RECT 56.345 2.898 56.35 3.388 ;
      RECT 56.335 2.905 56.345 3.395 ;
      RECT 56.325 2.912 56.335 3.403 ;
      RECT 56.31 2.922 56.325 3.411 ;
      RECT 56.3 2.936 56.31 3.421 ;
      RECT 56.29 2.948 56.3 3.433 ;
      RECT 56.275 2.97 56.29 3.446 ;
      RECT 56.265 2.992 56.275 3.457 ;
      RECT 56.255 3.012 56.265 3.466 ;
      RECT 56.25 3.027 56.255 3.473 ;
      RECT 56.22 3.06 56.25 3.487 ;
      RECT 56.21 3.095 56.22 3.502 ;
      RECT 56.205 3.102 56.21 3.508 ;
      RECT 56.185 3.117 56.205 3.515 ;
      RECT 56.18 3.132 56.185 3.523 ;
      RECT 56.175 3.141 56.18 3.528 ;
      RECT 56.16 3.147 56.175 3.535 ;
      RECT 56.155 3.153 56.16 3.543 ;
      RECT 56.15 3.157 56.155 3.55 ;
      RECT 56.145 3.161 56.15 3.56 ;
      RECT 56.135 3.166 56.145 3.57 ;
      RECT 56.115 3.177 56.135 3.598 ;
      RECT 56.1 3.189 56.115 3.625 ;
      RECT 56.08 3.202 56.1 3.65 ;
      RECT 56.06 3.217 56.08 3.674 ;
      RECT 56.045 3.232 56.06 3.689 ;
      RECT 56.04 3.243 56.045 3.698 ;
      RECT 55.975 3.288 56.04 3.708 ;
      RECT 55.94 3.347 55.975 3.721 ;
      RECT 55.935 3.37 55.94 3.727 ;
      RECT 55.93 3.377 55.935 3.729 ;
      RECT 55.915 3.387 55.93 3.732 ;
      RECT 55.885 3.412 55.915 3.736 ;
      RECT 55.88 3.43 55.885 3.74 ;
      RECT 55.875 3.437 55.88 3.741 ;
      RECT 55.855 3.445 55.875 3.745 ;
      RECT 55.845 3.452 55.855 3.749 ;
      RECT 55.801 3.463 55.845 3.756 ;
      RECT 55.715 3.491 55.801 3.772 ;
      RECT 55.655 3.515 55.715 3.79 ;
      RECT 55.61 3.525 55.655 3.804 ;
      RECT 55.551 3.533 55.61 3.818 ;
      RECT 55.465 3.54 55.551 3.837 ;
      RECT 55.44 3.545 55.465 3.852 ;
      RECT 55.36 3.548 55.44 3.855 ;
      RECT 55.28 3.552 55.36 3.842 ;
      RECT 55.271 3.555 55.28 3.827 ;
      RECT 55.185 3.555 55.271 3.812 ;
      RECT 55.125 3.557 55.185 3.789 ;
      RECT 55.121 3.56 55.125 3.779 ;
      RECT 55.035 3.56 55.121 3.764 ;
      RECT 54.96 3.56 55.035 3.74 ;
      RECT 56.275 2.569 56.285 2.745 ;
      RECT 56.23 2.536 56.275 2.745 ;
      RECT 56.185 2.487 56.23 2.745 ;
      RECT 56.155 2.457 56.185 2.746 ;
      RECT 56.15 2.44 56.155 2.747 ;
      RECT 56.125 2.42 56.15 2.748 ;
      RECT 56.11 2.395 56.125 2.749 ;
      RECT 56.105 2.382 56.11 2.75 ;
      RECT 56.1 2.376 56.105 2.748 ;
      RECT 56.095 2.368 56.1 2.742 ;
      RECT 56.07 2.36 56.095 2.722 ;
      RECT 56.05 2.349 56.07 2.693 ;
      RECT 56.02 2.334 56.05 2.664 ;
      RECT 56 2.32 56.02 2.636 ;
      RECT 55.99 2.314 56 2.615 ;
      RECT 55.985 2.311 55.99 2.598 ;
      RECT 55.98 2.308 55.985 2.583 ;
      RECT 55.965 2.303 55.98 2.548 ;
      RECT 55.96 2.299 55.965 2.515 ;
      RECT 55.94 2.294 55.96 2.491 ;
      RECT 55.91 2.286 55.94 2.456 ;
      RECT 55.895 2.28 55.91 2.433 ;
      RECT 55.855 2.273 55.895 2.418 ;
      RECT 55.83 2.265 55.855 2.398 ;
      RECT 55.81 2.26 55.83 2.388 ;
      RECT 55.775 2.254 55.81 2.383 ;
      RECT 55.73 2.245 55.775 2.382 ;
      RECT 55.7 2.241 55.73 2.384 ;
      RECT 55.615 2.249 55.7 2.388 ;
      RECT 55.545 2.26 55.615 2.41 ;
      RECT 55.532 2.266 55.545 2.433 ;
      RECT 55.446 2.273 55.532 2.455 ;
      RECT 55.36 2.285 55.446 2.492 ;
      RECT 55.36 2.662 55.37 2.9 ;
      RECT 55.355 2.291 55.36 2.515 ;
      RECT 55.35 2.547 55.36 2.9 ;
      RECT 55.35 2.292 55.355 2.52 ;
      RECT 55.345 2.293 55.35 2.9 ;
      RECT 55.321 2.295 55.345 2.901 ;
      RECT 55.235 2.303 55.321 2.903 ;
      RECT 55.215 2.317 55.235 2.906 ;
      RECT 55.21 2.345 55.215 2.907 ;
      RECT 55.205 2.357 55.21 2.908 ;
      RECT 55.2 2.372 55.205 2.909 ;
      RECT 55.19 2.402 55.2 2.91 ;
      RECT 55.185 2.44 55.19 2.908 ;
      RECT 55.18 2.46 55.185 2.903 ;
      RECT 55.165 2.495 55.18 2.888 ;
      RECT 55.155 2.547 55.165 2.868 ;
      RECT 55.15 2.577 55.155 2.856 ;
      RECT 55.135 2.59 55.15 2.839 ;
      RECT 55.11 2.594 55.135 2.806 ;
      RECT 55.095 2.592 55.11 2.783 ;
      RECT 55.08 2.591 55.095 2.78 ;
      RECT 55.02 2.589 55.08 2.778 ;
      RECT 55.01 2.587 55.02 2.773 ;
      RECT 54.97 2.586 55.01 2.77 ;
      RECT 54.9 2.583 54.97 2.768 ;
      RECT 54.845 2.581 54.9 2.763 ;
      RECT 54.775 2.575 54.845 2.758 ;
      RECT 54.766 2.575 54.775 2.755 ;
      RECT 54.68 2.575 54.766 2.75 ;
      RECT 54.675 2.575 54.68 2.745 ;
      RECT 55.98 1.81 56.155 2.16 ;
      RECT 55.98 1.825 56.165 2.158 ;
      RECT 55.955 1.775 56.1 2.155 ;
      RECT 55.935 1.776 56.1 2.148 ;
      RECT 55.925 1.777 56.11 2.143 ;
      RECT 55.895 1.778 56.11 2.13 ;
      RECT 55.845 1.779 56.11 2.106 ;
      RECT 55.84 1.781 56.11 2.091 ;
      RECT 55.84 1.847 56.17 2.085 ;
      RECT 55.82 1.788 56.125 2.065 ;
      RECT 55.81 1.797 56.135 1.92 ;
      RECT 55.82 1.792 56.135 2.065 ;
      RECT 55.84 1.782 56.125 2.091 ;
      RECT 55.425 3.107 55.595 3.395 ;
      RECT 55.42 3.125 55.605 3.39 ;
      RECT 55.385 3.133 55.67 3.31 ;
      RECT 55.385 3.133 55.756 3.3 ;
      RECT 55.385 3.133 55.81 3.246 ;
      RECT 55.67 3.03 55.84 3.214 ;
      RECT 55.385 3.185 55.845 3.202 ;
      RECT 55.37 3.155 55.84 3.198 ;
      RECT 55.63 3.037 55.67 3.349 ;
      RECT 55.51 3.074 55.84 3.214 ;
      RECT 55.605 3.049 55.63 3.375 ;
      RECT 55.595 3.056 55.84 3.214 ;
      RECT 55.726 2.52 55.795 2.779 ;
      RECT 55.726 2.575 55.8 2.778 ;
      RECT 55.64 2.575 55.8 2.777 ;
      RECT 55.635 2.575 55.805 2.77 ;
      RECT 55.625 2.52 55.795 2.765 ;
      RECT 55.005 1.819 55.18 2.12 ;
      RECT 54.99 1.807 55.005 2.105 ;
      RECT 54.96 1.806 54.99 2.058 ;
      RECT 54.96 1.824 55.185 2.053 ;
      RECT 54.945 1.808 55.005 2.018 ;
      RECT 54.94 1.83 55.195 1.918 ;
      RECT 54.94 1.813 55.091 1.918 ;
      RECT 54.94 1.815 55.095 1.918 ;
      RECT 54.945 1.811 55.091 2.018 ;
      RECT 55.05 3.047 55.055 3.395 ;
      RECT 55.04 3.037 55.05 3.401 ;
      RECT 55.005 3.027 55.04 3.403 ;
      RECT 54.967 3.022 55.005 3.407 ;
      RECT 54.881 3.015 54.967 3.414 ;
      RECT 54.795 3.005 54.881 3.424 ;
      RECT 54.75 3 54.795 3.432 ;
      RECT 54.746 3 54.75 3.436 ;
      RECT 54.66 3 54.746 3.443 ;
      RECT 54.645 3 54.66 3.443 ;
      RECT 54.635 2.998 54.645 3.415 ;
      RECT 54.625 2.994 54.635 3.358 ;
      RECT 54.605 2.988 54.625 3.29 ;
      RECT 54.6 2.984 54.605 3.238 ;
      RECT 54.59 2.983 54.6 3.205 ;
      RECT 54.54 2.981 54.59 3.19 ;
      RECT 54.515 2.979 54.54 3.185 ;
      RECT 54.472 2.977 54.515 3.181 ;
      RECT 54.386 2.973 54.472 3.169 ;
      RECT 54.3 2.968 54.386 3.153 ;
      RECT 54.27 2.965 54.3 3.14 ;
      RECT 54.245 2.964 54.27 3.128 ;
      RECT 54.24 2.964 54.245 3.118 ;
      RECT 54.2 2.963 54.24 3.11 ;
      RECT 54.185 2.962 54.2 3.103 ;
      RECT 54.135 2.961 54.185 3.095 ;
      RECT 54.133 2.96 54.135 3.09 ;
      RECT 54.047 2.958 54.133 3.09 ;
      RECT 53.961 2.953 54.047 3.09 ;
      RECT 53.875 2.949 53.961 3.09 ;
      RECT 53.826 2.945 53.875 3.088 ;
      RECT 53.74 2.942 53.826 3.083 ;
      RECT 53.717 2.939 53.74 3.079 ;
      RECT 53.631 2.936 53.717 3.074 ;
      RECT 53.545 2.932 53.631 3.065 ;
      RECT 53.52 2.925 53.545 3.06 ;
      RECT 53.46 2.89 53.52 3.057 ;
      RECT 53.44 2.815 53.46 3.054 ;
      RECT 53.435 2.757 53.44 3.053 ;
      RECT 53.41 2.697 53.435 3.052 ;
      RECT 53.335 2.575 53.41 3.048 ;
      RECT 53.325 2.575 53.335 3.04 ;
      RECT 53.31 2.575 53.325 3.03 ;
      RECT 53.295 2.575 53.31 3 ;
      RECT 53.28 2.575 53.295 2.945 ;
      RECT 53.265 2.575 53.28 2.883 ;
      RECT 53.24 2.575 53.265 2.808 ;
      RECT 53.235 2.575 53.24 2.758 ;
      RECT 54.58 2.12 54.6 2.429 ;
      RECT 54.566 2.122 54.615 2.426 ;
      RECT 54.566 2.127 54.635 2.417 ;
      RECT 54.48 2.125 54.615 2.411 ;
      RECT 54.48 2.133 54.67 2.394 ;
      RECT 54.445 2.135 54.67 2.393 ;
      RECT 54.415 2.143 54.67 2.384 ;
      RECT 54.405 2.148 54.69 2.37 ;
      RECT 54.445 2.138 54.69 2.37 ;
      RECT 54.445 2.141 54.7 2.358 ;
      RECT 54.415 2.143 54.71 2.345 ;
      RECT 54.415 2.147 54.72 2.288 ;
      RECT 54.405 2.152 54.725 2.203 ;
      RECT 54.566 2.12 54.6 2.426 ;
      RECT 54.445 7.855 54.615 8.305 ;
      RECT 54.5 6.075 54.67 8.025 ;
      RECT 54.445 5.015 54.615 6.245 ;
      RECT 54.005 2.223 54.01 2.435 ;
      RECT 53.88 2.22 53.895 2.435 ;
      RECT 53.345 2.25 53.415 2.435 ;
      RECT 53.23 2.25 53.265 2.43 ;
      RECT 54.351 2.552 54.37 2.746 ;
      RECT 54.265 2.507 54.351 2.747 ;
      RECT 54.255 2.46 54.265 2.749 ;
      RECT 54.25 2.44 54.255 2.75 ;
      RECT 54.23 2.405 54.25 2.751 ;
      RECT 54.215 2.355 54.23 2.752 ;
      RECT 54.195 2.292 54.215 2.753 ;
      RECT 54.185 2.255 54.195 2.754 ;
      RECT 54.17 2.244 54.185 2.755 ;
      RECT 54.165 2.236 54.17 2.753 ;
      RECT 54.155 2.235 54.165 2.745 ;
      RECT 54.125 2.232 54.155 2.724 ;
      RECT 54.05 2.227 54.125 2.669 ;
      RECT 54.035 2.223 54.05 2.615 ;
      RECT 54.025 2.223 54.035 2.51 ;
      RECT 54.01 2.223 54.025 2.443 ;
      RECT 53.995 2.223 54.005 2.433 ;
      RECT 53.94 2.222 53.995 2.43 ;
      RECT 53.895 2.22 53.94 2.433 ;
      RECT 53.867 2.22 53.88 2.436 ;
      RECT 53.781 2.224 53.867 2.438 ;
      RECT 53.695 2.23 53.781 2.443 ;
      RECT 53.675 2.234 53.695 2.445 ;
      RECT 53.673 2.235 53.675 2.444 ;
      RECT 53.587 2.237 53.673 2.443 ;
      RECT 53.501 2.242 53.587 2.44 ;
      RECT 53.415 2.247 53.501 2.437 ;
      RECT 53.265 2.25 53.345 2.433 ;
      RECT 53.925 5.015 54.095 8.305 ;
      RECT 53.925 7.315 54.33 7.645 ;
      RECT 53.925 6.475 54.33 6.805 ;
      RECT 54.041 3.225 54.09 3.559 ;
      RECT 54.041 3.225 54.095 3.558 ;
      RECT 53.955 3.225 54.095 3.557 ;
      RECT 53.73 3.333 54.1 3.555 ;
      RECT 53.955 3.225 54.125 3.548 ;
      RECT 53.925 3.237 54.13 3.539 ;
      RECT 53.91 3.255 54.135 3.536 ;
      RECT 53.725 3.339 54.135 3.463 ;
      RECT 53.72 3.346 54.135 3.423 ;
      RECT 53.735 3.312 54.135 3.536 ;
      RECT 53.896 3.258 54.1 3.555 ;
      RECT 53.81 3.278 54.135 3.536 ;
      RECT 53.91 3.252 54.13 3.539 ;
      RECT 53.68 2.576 53.87 2.77 ;
      RECT 53.675 2.578 53.87 2.769 ;
      RECT 53.67 2.582 53.885 2.766 ;
      RECT 53.685 2.575 53.885 2.766 ;
      RECT 53.67 2.685 53.89 2.761 ;
      RECT 52.965 3.185 53.056 3.483 ;
      RECT 52.96 3.187 53.135 3.478 ;
      RECT 52.965 3.185 53.135 3.478 ;
      RECT 52.96 3.191 53.155 3.476 ;
      RECT 52.96 3.246 53.195 3.475 ;
      RECT 52.96 3.281 53.21 3.469 ;
      RECT 52.96 3.315 53.22 3.459 ;
      RECT 52.95 3.195 53.155 3.31 ;
      RECT 52.95 3.215 53.17 3.31 ;
      RECT 52.95 3.198 53.16 3.31 ;
      RECT 53.175 1.966 53.18 2.028 ;
      RECT 53.17 1.888 53.175 2.051 ;
      RECT 53.165 1.845 53.17 2.062 ;
      RECT 53.16 1.835 53.165 2.074 ;
      RECT 53.155 1.835 53.16 2.083 ;
      RECT 53.13 1.835 53.155 2.115 ;
      RECT 53.125 1.835 53.13 2.148 ;
      RECT 53.11 1.835 53.125 2.173 ;
      RECT 53.1 1.835 53.11 2.2 ;
      RECT 53.095 1.835 53.1 2.213 ;
      RECT 53.09 1.835 53.095 2.228 ;
      RECT 53.08 1.835 53.09 2.243 ;
      RECT 53.075 1.835 53.08 2.263 ;
      RECT 53.05 1.835 53.075 2.298 ;
      RECT 53.005 1.835 53.05 2.343 ;
      RECT 52.995 1.835 53.005 2.356 ;
      RECT 52.91 1.92 52.995 2.363 ;
      RECT 52.875 2.042 52.91 2.372 ;
      RECT 52.87 2.082 52.875 2.376 ;
      RECT 52.85 2.105 52.87 2.378 ;
      RECT 52.845 2.135 52.85 2.381 ;
      RECT 52.835 2.147 52.845 2.382 ;
      RECT 52.79 2.17 52.835 2.387 ;
      RECT 52.75 2.2 52.79 2.395 ;
      RECT 52.715 2.212 52.75 2.401 ;
      RECT 52.71 2.217 52.715 2.405 ;
      RECT 52.64 2.227 52.71 2.412 ;
      RECT 52.6 2.237 52.64 2.422 ;
      RECT 52.58 2.242 52.6 2.428 ;
      RECT 52.57 2.246 52.58 2.433 ;
      RECT 52.565 2.249 52.57 2.436 ;
      RECT 52.555 2.25 52.565 2.437 ;
      RECT 52.53 2.252 52.555 2.441 ;
      RECT 52.52 2.257 52.53 2.444 ;
      RECT 52.475 2.265 52.52 2.445 ;
      RECT 52.35 2.27 52.475 2.445 ;
      RECT 52.905 2.567 52.925 2.749 ;
      RECT 52.856 2.552 52.905 2.748 ;
      RECT 52.77 2.567 52.925 2.746 ;
      RECT 52.755 2.567 52.925 2.745 ;
      RECT 52.72 2.545 52.89 2.73 ;
      RECT 52.79 3.565 52.805 3.774 ;
      RECT 52.79 3.573 52.81 3.773 ;
      RECT 52.735 3.573 52.81 3.772 ;
      RECT 52.715 3.577 52.815 3.77 ;
      RECT 52.695 3.527 52.735 3.769 ;
      RECT 52.64 3.585 52.82 3.767 ;
      RECT 52.605 3.542 52.735 3.765 ;
      RECT 52.601 3.545 52.79 3.764 ;
      RECT 52.515 3.553 52.79 3.762 ;
      RECT 52.515 3.597 52.825 3.755 ;
      RECT 52.505 3.69 52.825 3.753 ;
      RECT 52.515 3.609 52.83 3.738 ;
      RECT 52.515 3.63 52.845 3.708 ;
      RECT 52.515 3.657 52.85 3.678 ;
      RECT 52.64 3.535 52.735 3.767 ;
      RECT 52.27 2.58 52.275 3.118 ;
      RECT 52.075 2.91 52.08 3.105 ;
      RECT 50.375 2.575 50.39 2.955 ;
      RECT 52.44 2.575 52.445 2.745 ;
      RECT 52.435 2.575 52.44 2.755 ;
      RECT 52.43 2.575 52.435 2.768 ;
      RECT 52.405 2.575 52.43 2.81 ;
      RECT 52.38 2.575 52.405 2.883 ;
      RECT 52.365 2.575 52.38 2.935 ;
      RECT 52.36 2.575 52.365 2.965 ;
      RECT 52.335 2.575 52.36 3.005 ;
      RECT 52.32 2.575 52.335 3.06 ;
      RECT 52.315 2.575 52.32 3.093 ;
      RECT 52.29 2.575 52.315 3.113 ;
      RECT 52.275 2.575 52.29 3.119 ;
      RECT 52.205 2.61 52.27 3.115 ;
      RECT 52.155 2.665 52.205 3.11 ;
      RECT 52.145 2.697 52.155 3.108 ;
      RECT 52.14 2.722 52.145 3.108 ;
      RECT 52.12 2.795 52.14 3.108 ;
      RECT 52.11 2.875 52.12 3.107 ;
      RECT 52.095 2.905 52.11 3.107 ;
      RECT 52.08 2.91 52.095 3.106 ;
      RECT 52.02 2.912 52.075 3.103 ;
      RECT 51.99 2.917 52.02 3.099 ;
      RECT 51.988 2.92 51.99 3.098 ;
      RECT 51.902 2.922 51.988 3.095 ;
      RECT 51.816 2.928 51.902 3.089 ;
      RECT 51.73 2.933 51.816 3.083 ;
      RECT 51.657 2.938 51.73 3.084 ;
      RECT 51.571 2.944 51.657 3.092 ;
      RECT 51.485 2.95 51.571 3.101 ;
      RECT 51.465 2.954 51.485 3.106 ;
      RECT 51.418 2.956 51.465 3.109 ;
      RECT 51.332 2.961 51.418 3.115 ;
      RECT 51.246 2.966 51.332 3.124 ;
      RECT 51.16 2.972 51.246 3.132 ;
      RECT 51.075 2.97 51.16 3.141 ;
      RECT 51.071 2.965 51.075 3.145 ;
      RECT 50.985 2.96 51.071 3.137 ;
      RECT 50.921 2.951 50.985 3.125 ;
      RECT 50.835 2.942 50.921 3.112 ;
      RECT 50.811 2.935 50.835 3.103 ;
      RECT 50.725 2.929 50.811 3.09 ;
      RECT 50.685 2.922 50.725 3.076 ;
      RECT 50.68 2.912 50.685 3.072 ;
      RECT 50.67 2.9 50.68 3.071 ;
      RECT 50.65 2.87 50.67 3.068 ;
      RECT 50.595 2.79 50.65 3.062 ;
      RECT 50.575 2.709 50.595 3.057 ;
      RECT 50.555 2.667 50.575 3.053 ;
      RECT 50.53 2.62 50.555 3.047 ;
      RECT 50.525 2.595 50.53 3.044 ;
      RECT 50.49 2.575 50.525 3.039 ;
      RECT 50.481 2.575 50.49 3.032 ;
      RECT 50.395 2.575 50.481 3.002 ;
      RECT 50.39 2.575 50.395 2.965 ;
      RECT 50.355 2.575 50.375 2.887 ;
      RECT 50.35 2.617 50.355 2.852 ;
      RECT 50.345 2.692 50.35 2.808 ;
      RECT 51.795 2.497 51.97 2.745 ;
      RECT 51.795 2.497 51.975 2.743 ;
      RECT 51.79 2.529 51.975 2.703 ;
      RECT 51.82 2.47 51.99 2.69 ;
      RECT 51.785 2.547 51.99 2.623 ;
      RECT 51.095 2.01 51.265 2.185 ;
      RECT 51.095 2.01 51.437 2.177 ;
      RECT 51.095 2.01 51.52 2.171 ;
      RECT 51.095 2.01 51.555 2.167 ;
      RECT 51.095 2.01 51.575 2.166 ;
      RECT 51.095 2.01 51.661 2.162 ;
      RECT 51.555 1.835 51.725 2.157 ;
      RECT 51.13 1.942 51.755 2.155 ;
      RECT 51.12 1.997 51.76 2.153 ;
      RECT 51.095 2.033 51.77 2.148 ;
      RECT 51.095 2.06 51.775 2.078 ;
      RECT 51.16 1.885 51.735 2.155 ;
      RECT 51.351 1.87 51.735 2.155 ;
      RECT 51.185 1.873 51.735 2.155 ;
      RECT 51.265 1.871 51.351 2.182 ;
      RECT 51.351 1.868 51.73 2.155 ;
      RECT 51.535 1.845 51.73 2.155 ;
      RECT 51.437 1.866 51.73 2.155 ;
      RECT 51.52 1.86 51.535 2.168 ;
      RECT 51.67 3.225 51.675 3.425 ;
      RECT 51.135 3.29 51.18 3.425 ;
      RECT 51.705 3.225 51.725 3.398 ;
      RECT 51.675 3.225 51.705 3.413 ;
      RECT 51.61 3.225 51.67 3.45 ;
      RECT 51.595 3.225 51.61 3.48 ;
      RECT 51.58 3.225 51.595 3.493 ;
      RECT 51.56 3.225 51.58 3.508 ;
      RECT 51.555 3.225 51.56 3.517 ;
      RECT 51.545 3.229 51.555 3.522 ;
      RECT 51.53 3.239 51.545 3.533 ;
      RECT 51.505 3.255 51.53 3.543 ;
      RECT 51.495 3.269 51.505 3.545 ;
      RECT 51.475 3.281 51.495 3.542 ;
      RECT 51.445 3.302 51.475 3.536 ;
      RECT 51.435 3.314 51.445 3.531 ;
      RECT 51.425 3.312 51.435 3.528 ;
      RECT 51.41 3.311 51.425 3.523 ;
      RECT 51.405 3.31 51.41 3.518 ;
      RECT 51.37 3.308 51.405 3.508 ;
      RECT 51.35 3.305 51.37 3.49 ;
      RECT 51.34 3.303 51.35 3.485 ;
      RECT 51.33 3.302 51.34 3.48 ;
      RECT 51.295 3.3 51.33 3.468 ;
      RECT 51.24 3.296 51.295 3.448 ;
      RECT 51.23 3.294 51.24 3.433 ;
      RECT 51.225 3.294 51.23 3.428 ;
      RECT 51.18 3.292 51.225 3.425 ;
      RECT 51.085 3.29 51.135 3.429 ;
      RECT 51.075 3.291 51.085 3.434 ;
      RECT 51.015 3.298 51.075 3.448 ;
      RECT 50.99 3.306 51.015 3.468 ;
      RECT 50.98 3.31 50.99 3.48 ;
      RECT 50.975 3.311 50.98 3.485 ;
      RECT 50.96 3.313 50.975 3.488 ;
      RECT 50.945 3.315 50.96 3.493 ;
      RECT 50.94 3.315 50.945 3.496 ;
      RECT 50.895 3.32 50.94 3.507 ;
      RECT 50.89 3.324 50.895 3.519 ;
      RECT 50.865 3.32 50.89 3.523 ;
      RECT 50.855 3.316 50.865 3.527 ;
      RECT 50.845 3.315 50.855 3.531 ;
      RECT 50.83 3.305 50.845 3.537 ;
      RECT 50.825 3.293 50.83 3.541 ;
      RECT 50.82 3.29 50.825 3.542 ;
      RECT 50.815 3.287 50.82 3.544 ;
      RECT 50.8 3.275 50.815 3.543 ;
      RECT 50.785 3.257 50.8 3.54 ;
      RECT 50.765 3.236 50.785 3.533 ;
      RECT 50.7 3.225 50.765 3.505 ;
      RECT 50.696 3.225 50.7 3.484 ;
      RECT 50.61 3.225 50.696 3.454 ;
      RECT 50.595 3.225 50.61 3.41 ;
      RECT 51.17 2.325 51.175 2.56 ;
      RECT 50.3 2.241 50.305 2.445 ;
      RECT 50.88 2.27 50.885 2.425 ;
      RECT 50.8 2.25 50.805 2.425 ;
      RECT 51.47 2.392 51.485 2.745 ;
      RECT 51.396 2.377 51.47 2.745 ;
      RECT 51.31 2.36 51.396 2.745 ;
      RECT 51.3 2.35 51.31 2.743 ;
      RECT 51.295 2.348 51.3 2.738 ;
      RECT 51.28 2.346 51.295 2.724 ;
      RECT 51.21 2.338 51.28 2.664 ;
      RECT 51.19 2.329 51.21 2.598 ;
      RECT 51.185 2.326 51.19 2.578 ;
      RECT 51.175 2.325 51.185 2.568 ;
      RECT 51.165 2.325 51.17 2.552 ;
      RECT 51.155 2.324 51.165 2.542 ;
      RECT 51.145 2.322 51.155 2.53 ;
      RECT 51.13 2.319 51.145 2.51 ;
      RECT 51.12 2.317 51.13 2.495 ;
      RECT 51.1 2.314 51.12 2.483 ;
      RECT 51.095 2.312 51.1 2.473 ;
      RECT 51.07 2.31 51.095 2.46 ;
      RECT 51.04 2.305 51.07 2.445 ;
      RECT 50.96 2.296 51.04 2.436 ;
      RECT 50.915 2.285 50.96 2.429 ;
      RECT 50.895 2.276 50.915 2.426 ;
      RECT 50.885 2.271 50.895 2.425 ;
      RECT 50.84 2.265 50.88 2.425 ;
      RECT 50.825 2.257 50.84 2.425 ;
      RECT 50.805 2.252 50.825 2.425 ;
      RECT 50.785 2.249 50.8 2.425 ;
      RECT 50.702 2.248 50.785 2.424 ;
      RECT 50.616 2.247 50.702 2.42 ;
      RECT 50.53 2.245 50.616 2.417 ;
      RECT 50.477 2.244 50.53 2.419 ;
      RECT 50.391 2.243 50.477 2.428 ;
      RECT 50.305 2.242 50.391 2.44 ;
      RECT 50.285 2.241 50.3 2.448 ;
      RECT 50.205 2.24 50.285 2.46 ;
      RECT 50.18 2.24 50.205 2.473 ;
      RECT 50.155 2.24 50.18 2.488 ;
      RECT 50.15 2.24 50.155 2.51 ;
      RECT 50.145 2.24 50.15 2.528 ;
      RECT 50.14 2.24 50.145 2.545 ;
      RECT 50.135 2.24 50.14 2.558 ;
      RECT 50.13 2.24 50.135 2.568 ;
      RECT 50.09 2.24 50.13 2.653 ;
      RECT 50.075 2.24 50.09 2.738 ;
      RECT 50.065 2.241 50.075 2.75 ;
      RECT 50.03 2.246 50.065 2.755 ;
      RECT 49.99 2.255 50.03 2.755 ;
      RECT 49.975 2.265 49.99 2.755 ;
      RECT 49.97 2.275 49.975 2.755 ;
      RECT 49.95 2.302 49.97 2.755 ;
      RECT 49.9 2.385 49.95 2.755 ;
      RECT 49.895 2.447 49.9 2.755 ;
      RECT 49.885 2.46 49.895 2.755 ;
      RECT 49.875 2.482 49.885 2.755 ;
      RECT 49.865 2.507 49.875 2.75 ;
      RECT 49.86 2.545 49.865 2.743 ;
      RECT 49.85 2.655 49.86 2.738 ;
      RECT 51.245 3.576 51.26 3.835 ;
      RECT 51.245 3.591 51.265 3.834 ;
      RECT 51.161 3.591 51.265 3.832 ;
      RECT 51.161 3.605 51.27 3.831 ;
      RECT 51.075 3.647 51.275 3.828 ;
      RECT 51.07 3.59 51.26 3.823 ;
      RECT 51.07 3.661 51.28 3.82 ;
      RECT 51.065 3.692 51.28 3.818 ;
      RECT 51.07 3.689 51.295 3.808 ;
      RECT 51.065 3.735 51.31 3.793 ;
      RECT 51.065 3.763 51.315 3.778 ;
      RECT 51.075 3.565 51.245 3.828 ;
      RECT 50.835 2.575 51.005 2.745 ;
      RECT 50.8 2.575 51.005 2.74 ;
      RECT 50.79 2.575 51.005 2.733 ;
      RECT 50.785 2.56 50.955 2.73 ;
      RECT 49.615 3.097 49.88 3.54 ;
      RECT 49.61 3.068 49.825 3.538 ;
      RECT 49.605 3.222 49.885 3.533 ;
      RECT 49.61 3.117 49.885 3.533 ;
      RECT 49.61 3.128 49.895 3.52 ;
      RECT 49.61 3.075 49.855 3.538 ;
      RECT 49.615 3.062 49.825 3.54 ;
      RECT 49.615 3.06 49.775 3.54 ;
      RECT 49.716 3.052 49.775 3.54 ;
      RECT 49.63 3.053 49.775 3.54 ;
      RECT 49.716 3.051 49.765 3.54 ;
      RECT 49.52 1.866 49.695 2.165 ;
      RECT 49.57 1.828 49.695 2.165 ;
      RECT 49.555 1.83 49.781 2.157 ;
      RECT 49.555 1.833 49.82 2.144 ;
      RECT 49.555 1.834 49.83 2.13 ;
      RECT 49.51 1.885 49.83 2.12 ;
      RECT 49.555 1.835 49.835 2.115 ;
      RECT 49.51 2.045 49.84 2.105 ;
      RECT 49.495 1.905 49.835 2.045 ;
      RECT 49.49 1.921 49.835 1.985 ;
      RECT 49.535 1.845 49.835 2.115 ;
      RECT 49.57 1.826 49.656 2.165 ;
      RECT 48.03 5.02 48.2 6.49 ;
      RECT 48.03 6.315 48.205 6.485 ;
      RECT 47.66 1.74 47.83 2.93 ;
      RECT 47.66 1.74 48.13 1.91 ;
      RECT 47.66 6.97 48.13 7.14 ;
      RECT 47.66 5.95 47.83 7.14 ;
      RECT 46.67 1.74 46.84 2.93 ;
      RECT 46.67 1.74 47.14 1.91 ;
      RECT 46.67 6.97 47.14 7.14 ;
      RECT 46.67 5.95 46.84 7.14 ;
      RECT 44.82 2.635 44.99 3.865 ;
      RECT 44.875 0.855 45.045 2.805 ;
      RECT 44.82 0.575 44.99 1.025 ;
      RECT 44.82 7.855 44.99 8.305 ;
      RECT 44.875 6.075 45.045 8.025 ;
      RECT 44.82 5.015 44.99 6.245 ;
      RECT 44.3 0.575 44.47 3.865 ;
      RECT 44.3 2.075 44.705 2.405 ;
      RECT 44.3 1.235 44.705 1.565 ;
      RECT 44.3 5.015 44.47 8.305 ;
      RECT 44.3 7.315 44.705 7.645 ;
      RECT 44.3 6.475 44.705 6.805 ;
      RECT 42.225 3.126 42.23 3.298 ;
      RECT 42.22 3.119 42.225 3.388 ;
      RECT 42.215 3.113 42.22 3.407 ;
      RECT 42.195 3.107 42.215 3.417 ;
      RECT 42.18 3.102 42.195 3.425 ;
      RECT 42.143 3.096 42.18 3.423 ;
      RECT 42.057 3.082 42.143 3.419 ;
      RECT 41.971 3.064 42.057 3.414 ;
      RECT 41.885 3.045 41.971 3.408 ;
      RECT 41.855 3.033 41.885 3.404 ;
      RECT 41.835 3.027 41.855 3.403 ;
      RECT 41.77 3.025 41.835 3.401 ;
      RECT 41.755 3.025 41.77 3.393 ;
      RECT 41.74 3.025 41.755 3.38 ;
      RECT 41.735 3.025 41.74 3.37 ;
      RECT 41.72 3.025 41.735 3.348 ;
      RECT 41.705 3.025 41.72 3.315 ;
      RECT 41.7 3.025 41.705 3.293 ;
      RECT 41.69 3.025 41.7 3.275 ;
      RECT 41.675 3.025 41.69 3.253 ;
      RECT 41.655 3.025 41.675 3.215 ;
      RECT 42.005 2.31 42.04 2.749 ;
      RECT 42.005 2.31 42.045 2.748 ;
      RECT 41.95 2.37 42.045 2.747 ;
      RECT 41.815 2.542 42.045 2.746 ;
      RECT 41.925 2.42 42.045 2.746 ;
      RECT 41.815 2.542 42.07 2.736 ;
      RECT 41.87 2.487 42.15 2.653 ;
      RECT 42.045 2.281 42.05 2.744 ;
      RECT 41.9 2.457 42.19 2.53 ;
      RECT 41.915 2.44 42.045 2.746 ;
      RECT 42.05 2.28 42.22 2.468 ;
      RECT 42.04 2.283 42.22 2.468 ;
      RECT 41.545 2.16 41.715 2.47 ;
      RECT 41.545 2.16 41.72 2.443 ;
      RECT 41.545 2.16 41.725 2.42 ;
      RECT 41.545 2.16 41.735 2.37 ;
      RECT 41.54 2.265 41.735 2.34 ;
      RECT 41.575 1.835 41.745 2.313 ;
      RECT 41.575 1.835 41.76 2.234 ;
      RECT 41.565 2.045 41.76 2.234 ;
      RECT 41.575 1.845 41.77 2.149 ;
      RECT 41.505 2.587 41.51 2.79 ;
      RECT 41.495 2.575 41.505 2.9 ;
      RECT 41.47 2.575 41.495 2.94 ;
      RECT 41.39 2.575 41.47 3.025 ;
      RECT 41.38 2.575 41.39 3.095 ;
      RECT 41.355 2.575 41.38 3.118 ;
      RECT 41.335 2.575 41.355 3.153 ;
      RECT 41.29 2.585 41.335 3.196 ;
      RECT 41.28 2.597 41.29 3.233 ;
      RECT 41.26 2.611 41.28 3.253 ;
      RECT 41.25 2.629 41.26 3.269 ;
      RECT 41.235 2.655 41.25 3.279 ;
      RECT 41.22 2.696 41.235 3.293 ;
      RECT 41.21 2.731 41.22 3.303 ;
      RECT 41.205 2.747 41.21 3.308 ;
      RECT 41.195 2.762 41.205 3.313 ;
      RECT 41.175 2.805 41.195 3.323 ;
      RECT 41.155 2.842 41.175 3.336 ;
      RECT 41.12 2.865 41.155 3.354 ;
      RECT 41.11 2.879 41.12 3.37 ;
      RECT 41.09 2.889 41.11 3.38 ;
      RECT 41.085 2.898 41.09 3.388 ;
      RECT 41.075 2.905 41.085 3.395 ;
      RECT 41.065 2.912 41.075 3.403 ;
      RECT 41.05 2.922 41.065 3.411 ;
      RECT 41.04 2.936 41.05 3.421 ;
      RECT 41.03 2.948 41.04 3.433 ;
      RECT 41.015 2.97 41.03 3.446 ;
      RECT 41.005 2.992 41.015 3.457 ;
      RECT 40.995 3.012 41.005 3.466 ;
      RECT 40.99 3.027 40.995 3.473 ;
      RECT 40.96 3.06 40.99 3.487 ;
      RECT 40.95 3.095 40.96 3.502 ;
      RECT 40.945 3.102 40.95 3.508 ;
      RECT 40.925 3.117 40.945 3.515 ;
      RECT 40.92 3.132 40.925 3.523 ;
      RECT 40.915 3.141 40.92 3.528 ;
      RECT 40.9 3.147 40.915 3.535 ;
      RECT 40.895 3.153 40.9 3.543 ;
      RECT 40.89 3.157 40.895 3.55 ;
      RECT 40.885 3.161 40.89 3.56 ;
      RECT 40.875 3.166 40.885 3.57 ;
      RECT 40.855 3.177 40.875 3.598 ;
      RECT 40.84 3.189 40.855 3.625 ;
      RECT 40.82 3.202 40.84 3.65 ;
      RECT 40.8 3.217 40.82 3.674 ;
      RECT 40.785 3.232 40.8 3.689 ;
      RECT 40.78 3.243 40.785 3.698 ;
      RECT 40.715 3.288 40.78 3.708 ;
      RECT 40.68 3.347 40.715 3.721 ;
      RECT 40.675 3.37 40.68 3.727 ;
      RECT 40.67 3.377 40.675 3.729 ;
      RECT 40.655 3.387 40.67 3.732 ;
      RECT 40.625 3.412 40.655 3.736 ;
      RECT 40.62 3.43 40.625 3.74 ;
      RECT 40.615 3.437 40.62 3.741 ;
      RECT 40.595 3.445 40.615 3.745 ;
      RECT 40.585 3.452 40.595 3.749 ;
      RECT 40.541 3.463 40.585 3.756 ;
      RECT 40.455 3.491 40.541 3.772 ;
      RECT 40.395 3.515 40.455 3.79 ;
      RECT 40.35 3.525 40.395 3.804 ;
      RECT 40.291 3.533 40.35 3.818 ;
      RECT 40.205 3.54 40.291 3.837 ;
      RECT 40.18 3.545 40.205 3.852 ;
      RECT 40.1 3.548 40.18 3.855 ;
      RECT 40.02 3.552 40.1 3.842 ;
      RECT 40.011 3.555 40.02 3.827 ;
      RECT 39.925 3.555 40.011 3.812 ;
      RECT 39.865 3.557 39.925 3.789 ;
      RECT 39.861 3.56 39.865 3.779 ;
      RECT 39.775 3.56 39.861 3.764 ;
      RECT 39.7 3.56 39.775 3.74 ;
      RECT 41.015 2.569 41.025 2.745 ;
      RECT 40.97 2.536 41.015 2.745 ;
      RECT 40.925 2.487 40.97 2.745 ;
      RECT 40.895 2.457 40.925 2.746 ;
      RECT 40.89 2.44 40.895 2.747 ;
      RECT 40.865 2.42 40.89 2.748 ;
      RECT 40.85 2.395 40.865 2.749 ;
      RECT 40.845 2.382 40.85 2.75 ;
      RECT 40.84 2.376 40.845 2.748 ;
      RECT 40.835 2.368 40.84 2.742 ;
      RECT 40.81 2.36 40.835 2.722 ;
      RECT 40.79 2.349 40.81 2.693 ;
      RECT 40.76 2.334 40.79 2.664 ;
      RECT 40.74 2.32 40.76 2.636 ;
      RECT 40.73 2.314 40.74 2.615 ;
      RECT 40.725 2.311 40.73 2.598 ;
      RECT 40.72 2.308 40.725 2.583 ;
      RECT 40.705 2.303 40.72 2.548 ;
      RECT 40.7 2.299 40.705 2.515 ;
      RECT 40.68 2.294 40.7 2.491 ;
      RECT 40.65 2.286 40.68 2.456 ;
      RECT 40.635 2.28 40.65 2.433 ;
      RECT 40.595 2.273 40.635 2.418 ;
      RECT 40.57 2.265 40.595 2.398 ;
      RECT 40.55 2.26 40.57 2.388 ;
      RECT 40.515 2.254 40.55 2.383 ;
      RECT 40.47 2.245 40.515 2.382 ;
      RECT 40.44 2.241 40.47 2.384 ;
      RECT 40.355 2.249 40.44 2.388 ;
      RECT 40.285 2.26 40.355 2.41 ;
      RECT 40.272 2.266 40.285 2.433 ;
      RECT 40.186 2.273 40.272 2.455 ;
      RECT 40.1 2.285 40.186 2.492 ;
      RECT 40.1 2.662 40.11 2.9 ;
      RECT 40.095 2.291 40.1 2.515 ;
      RECT 40.09 2.547 40.1 2.9 ;
      RECT 40.09 2.292 40.095 2.52 ;
      RECT 40.085 2.293 40.09 2.9 ;
      RECT 40.061 2.295 40.085 2.901 ;
      RECT 39.975 2.303 40.061 2.903 ;
      RECT 39.955 2.317 39.975 2.906 ;
      RECT 39.95 2.345 39.955 2.907 ;
      RECT 39.945 2.357 39.95 2.908 ;
      RECT 39.94 2.372 39.945 2.909 ;
      RECT 39.93 2.402 39.94 2.91 ;
      RECT 39.925 2.44 39.93 2.908 ;
      RECT 39.92 2.46 39.925 2.903 ;
      RECT 39.905 2.495 39.92 2.888 ;
      RECT 39.895 2.547 39.905 2.868 ;
      RECT 39.89 2.577 39.895 2.856 ;
      RECT 39.875 2.59 39.89 2.839 ;
      RECT 39.85 2.594 39.875 2.806 ;
      RECT 39.835 2.592 39.85 2.783 ;
      RECT 39.82 2.591 39.835 2.78 ;
      RECT 39.76 2.589 39.82 2.778 ;
      RECT 39.75 2.587 39.76 2.773 ;
      RECT 39.71 2.586 39.75 2.77 ;
      RECT 39.64 2.583 39.71 2.768 ;
      RECT 39.585 2.581 39.64 2.763 ;
      RECT 39.515 2.575 39.585 2.758 ;
      RECT 39.506 2.575 39.515 2.755 ;
      RECT 39.42 2.575 39.506 2.75 ;
      RECT 39.415 2.575 39.42 2.745 ;
      RECT 40.72 1.81 40.895 2.16 ;
      RECT 40.72 1.825 40.905 2.158 ;
      RECT 40.695 1.775 40.84 2.155 ;
      RECT 40.675 1.776 40.84 2.148 ;
      RECT 40.665 1.777 40.85 2.143 ;
      RECT 40.635 1.778 40.85 2.13 ;
      RECT 40.585 1.779 40.85 2.106 ;
      RECT 40.58 1.781 40.85 2.091 ;
      RECT 40.58 1.847 40.91 2.085 ;
      RECT 40.56 1.788 40.865 2.065 ;
      RECT 40.55 1.797 40.875 1.92 ;
      RECT 40.56 1.792 40.875 2.065 ;
      RECT 40.58 1.782 40.865 2.091 ;
      RECT 40.165 3.107 40.335 3.395 ;
      RECT 40.16 3.125 40.345 3.39 ;
      RECT 40.125 3.133 40.41 3.31 ;
      RECT 40.125 3.133 40.496 3.3 ;
      RECT 40.125 3.133 40.55 3.246 ;
      RECT 40.41 3.03 40.58 3.214 ;
      RECT 40.125 3.185 40.585 3.202 ;
      RECT 40.11 3.155 40.58 3.198 ;
      RECT 40.37 3.037 40.41 3.349 ;
      RECT 40.25 3.074 40.58 3.214 ;
      RECT 40.345 3.049 40.37 3.375 ;
      RECT 40.335 3.056 40.58 3.214 ;
      RECT 40.466 2.52 40.535 2.779 ;
      RECT 40.466 2.575 40.54 2.778 ;
      RECT 40.38 2.575 40.54 2.777 ;
      RECT 40.375 2.575 40.545 2.77 ;
      RECT 40.365 2.52 40.535 2.765 ;
      RECT 39.745 1.819 39.92 2.12 ;
      RECT 39.73 1.807 39.745 2.105 ;
      RECT 39.7 1.806 39.73 2.058 ;
      RECT 39.7 1.824 39.925 2.053 ;
      RECT 39.685 1.808 39.745 2.018 ;
      RECT 39.68 1.83 39.935 1.918 ;
      RECT 39.68 1.813 39.831 1.918 ;
      RECT 39.68 1.815 39.835 1.918 ;
      RECT 39.685 1.811 39.831 2.018 ;
      RECT 39.79 3.047 39.795 3.395 ;
      RECT 39.78 3.037 39.79 3.401 ;
      RECT 39.745 3.027 39.78 3.403 ;
      RECT 39.707 3.022 39.745 3.407 ;
      RECT 39.621 3.015 39.707 3.414 ;
      RECT 39.535 3.005 39.621 3.424 ;
      RECT 39.49 3 39.535 3.432 ;
      RECT 39.486 3 39.49 3.436 ;
      RECT 39.4 3 39.486 3.443 ;
      RECT 39.385 3 39.4 3.443 ;
      RECT 39.375 2.998 39.385 3.415 ;
      RECT 39.365 2.994 39.375 3.358 ;
      RECT 39.345 2.988 39.365 3.29 ;
      RECT 39.34 2.984 39.345 3.238 ;
      RECT 39.33 2.983 39.34 3.205 ;
      RECT 39.28 2.981 39.33 3.19 ;
      RECT 39.255 2.979 39.28 3.185 ;
      RECT 39.212 2.977 39.255 3.181 ;
      RECT 39.126 2.973 39.212 3.169 ;
      RECT 39.04 2.968 39.126 3.153 ;
      RECT 39.01 2.965 39.04 3.14 ;
      RECT 38.985 2.964 39.01 3.128 ;
      RECT 38.98 2.964 38.985 3.118 ;
      RECT 38.94 2.963 38.98 3.11 ;
      RECT 38.925 2.962 38.94 3.103 ;
      RECT 38.875 2.961 38.925 3.095 ;
      RECT 38.873 2.96 38.875 3.09 ;
      RECT 38.787 2.958 38.873 3.09 ;
      RECT 38.701 2.953 38.787 3.09 ;
      RECT 38.615 2.949 38.701 3.09 ;
      RECT 38.566 2.945 38.615 3.088 ;
      RECT 38.48 2.942 38.566 3.083 ;
      RECT 38.457 2.939 38.48 3.079 ;
      RECT 38.371 2.936 38.457 3.074 ;
      RECT 38.285 2.932 38.371 3.065 ;
      RECT 38.26 2.925 38.285 3.06 ;
      RECT 38.2 2.89 38.26 3.057 ;
      RECT 38.18 2.815 38.2 3.054 ;
      RECT 38.175 2.757 38.18 3.053 ;
      RECT 38.15 2.697 38.175 3.052 ;
      RECT 38.075 2.575 38.15 3.048 ;
      RECT 38.065 2.575 38.075 3.04 ;
      RECT 38.05 2.575 38.065 3.03 ;
      RECT 38.035 2.575 38.05 3 ;
      RECT 38.02 2.575 38.035 2.945 ;
      RECT 38.005 2.575 38.02 2.883 ;
      RECT 37.98 2.575 38.005 2.808 ;
      RECT 37.975 2.575 37.98 2.758 ;
      RECT 39.32 2.12 39.34 2.429 ;
      RECT 39.306 2.122 39.355 2.426 ;
      RECT 39.306 2.127 39.375 2.417 ;
      RECT 39.22 2.125 39.355 2.411 ;
      RECT 39.22 2.133 39.41 2.394 ;
      RECT 39.185 2.135 39.41 2.393 ;
      RECT 39.155 2.143 39.41 2.384 ;
      RECT 39.145 2.148 39.43 2.37 ;
      RECT 39.185 2.138 39.43 2.37 ;
      RECT 39.185 2.141 39.44 2.358 ;
      RECT 39.155 2.143 39.45 2.345 ;
      RECT 39.155 2.147 39.46 2.288 ;
      RECT 39.145 2.152 39.465 2.203 ;
      RECT 39.306 2.12 39.34 2.426 ;
      RECT 39.185 7.855 39.355 8.305 ;
      RECT 39.24 6.075 39.41 8.025 ;
      RECT 39.185 5.015 39.355 6.245 ;
      RECT 38.745 2.223 38.75 2.435 ;
      RECT 38.62 2.22 38.635 2.435 ;
      RECT 38.085 2.25 38.155 2.435 ;
      RECT 37.97 2.25 38.005 2.43 ;
      RECT 39.091 2.552 39.11 2.746 ;
      RECT 39.005 2.507 39.091 2.747 ;
      RECT 38.995 2.46 39.005 2.749 ;
      RECT 38.99 2.44 38.995 2.75 ;
      RECT 38.97 2.405 38.99 2.751 ;
      RECT 38.955 2.355 38.97 2.752 ;
      RECT 38.935 2.292 38.955 2.753 ;
      RECT 38.925 2.255 38.935 2.754 ;
      RECT 38.91 2.244 38.925 2.755 ;
      RECT 38.905 2.236 38.91 2.753 ;
      RECT 38.895 2.235 38.905 2.745 ;
      RECT 38.865 2.232 38.895 2.724 ;
      RECT 38.79 2.227 38.865 2.669 ;
      RECT 38.775 2.223 38.79 2.615 ;
      RECT 38.765 2.223 38.775 2.51 ;
      RECT 38.75 2.223 38.765 2.443 ;
      RECT 38.735 2.223 38.745 2.433 ;
      RECT 38.68 2.222 38.735 2.43 ;
      RECT 38.635 2.22 38.68 2.433 ;
      RECT 38.607 2.22 38.62 2.436 ;
      RECT 38.521 2.224 38.607 2.438 ;
      RECT 38.435 2.23 38.521 2.443 ;
      RECT 38.415 2.234 38.435 2.445 ;
      RECT 38.413 2.235 38.415 2.444 ;
      RECT 38.327 2.237 38.413 2.443 ;
      RECT 38.241 2.242 38.327 2.44 ;
      RECT 38.155 2.247 38.241 2.437 ;
      RECT 38.005 2.25 38.085 2.433 ;
      RECT 38.665 5.015 38.835 8.305 ;
      RECT 38.665 7.315 39.07 7.645 ;
      RECT 38.665 6.475 39.07 6.805 ;
      RECT 38.781 3.225 38.83 3.559 ;
      RECT 38.781 3.225 38.835 3.558 ;
      RECT 38.695 3.225 38.835 3.557 ;
      RECT 38.47 3.333 38.84 3.555 ;
      RECT 38.695 3.225 38.865 3.548 ;
      RECT 38.665 3.237 38.87 3.539 ;
      RECT 38.65 3.255 38.875 3.536 ;
      RECT 38.465 3.339 38.875 3.463 ;
      RECT 38.46 3.346 38.875 3.423 ;
      RECT 38.475 3.312 38.875 3.536 ;
      RECT 38.636 3.258 38.84 3.555 ;
      RECT 38.55 3.278 38.875 3.536 ;
      RECT 38.65 3.252 38.87 3.539 ;
      RECT 38.42 2.576 38.61 2.77 ;
      RECT 38.415 2.578 38.61 2.769 ;
      RECT 38.41 2.582 38.625 2.766 ;
      RECT 38.425 2.575 38.625 2.766 ;
      RECT 38.41 2.685 38.63 2.761 ;
      RECT 37.705 3.185 37.796 3.483 ;
      RECT 37.7 3.187 37.875 3.478 ;
      RECT 37.705 3.185 37.875 3.478 ;
      RECT 37.7 3.191 37.895 3.476 ;
      RECT 37.7 3.246 37.935 3.475 ;
      RECT 37.7 3.281 37.95 3.469 ;
      RECT 37.7 3.315 37.96 3.459 ;
      RECT 37.69 3.195 37.895 3.31 ;
      RECT 37.69 3.215 37.91 3.31 ;
      RECT 37.69 3.198 37.9 3.31 ;
      RECT 37.915 1.966 37.92 2.028 ;
      RECT 37.91 1.888 37.915 2.051 ;
      RECT 37.905 1.845 37.91 2.062 ;
      RECT 37.9 1.835 37.905 2.074 ;
      RECT 37.895 1.835 37.9 2.083 ;
      RECT 37.87 1.835 37.895 2.115 ;
      RECT 37.865 1.835 37.87 2.148 ;
      RECT 37.85 1.835 37.865 2.173 ;
      RECT 37.84 1.835 37.85 2.2 ;
      RECT 37.835 1.835 37.84 2.213 ;
      RECT 37.83 1.835 37.835 2.228 ;
      RECT 37.82 1.835 37.83 2.243 ;
      RECT 37.815 1.835 37.82 2.263 ;
      RECT 37.79 1.835 37.815 2.298 ;
      RECT 37.745 1.835 37.79 2.343 ;
      RECT 37.735 1.835 37.745 2.356 ;
      RECT 37.65 1.92 37.735 2.363 ;
      RECT 37.615 2.042 37.65 2.372 ;
      RECT 37.61 2.082 37.615 2.376 ;
      RECT 37.59 2.105 37.61 2.378 ;
      RECT 37.585 2.135 37.59 2.381 ;
      RECT 37.575 2.147 37.585 2.382 ;
      RECT 37.53 2.17 37.575 2.387 ;
      RECT 37.49 2.2 37.53 2.395 ;
      RECT 37.455 2.212 37.49 2.401 ;
      RECT 37.45 2.217 37.455 2.405 ;
      RECT 37.38 2.227 37.45 2.412 ;
      RECT 37.34 2.237 37.38 2.422 ;
      RECT 37.32 2.242 37.34 2.428 ;
      RECT 37.31 2.246 37.32 2.433 ;
      RECT 37.305 2.249 37.31 2.436 ;
      RECT 37.295 2.25 37.305 2.437 ;
      RECT 37.27 2.252 37.295 2.441 ;
      RECT 37.26 2.257 37.27 2.444 ;
      RECT 37.215 2.265 37.26 2.445 ;
      RECT 37.09 2.27 37.215 2.445 ;
      RECT 37.645 2.567 37.665 2.749 ;
      RECT 37.596 2.552 37.645 2.748 ;
      RECT 37.51 2.567 37.665 2.746 ;
      RECT 37.495 2.567 37.665 2.745 ;
      RECT 37.46 2.545 37.63 2.73 ;
      RECT 37.53 3.565 37.545 3.774 ;
      RECT 37.53 3.573 37.55 3.773 ;
      RECT 37.475 3.573 37.55 3.772 ;
      RECT 37.455 3.577 37.555 3.77 ;
      RECT 37.435 3.527 37.475 3.769 ;
      RECT 37.38 3.585 37.56 3.767 ;
      RECT 37.345 3.542 37.475 3.765 ;
      RECT 37.341 3.545 37.53 3.764 ;
      RECT 37.255 3.553 37.53 3.762 ;
      RECT 37.255 3.597 37.565 3.755 ;
      RECT 37.245 3.69 37.565 3.753 ;
      RECT 37.255 3.609 37.57 3.738 ;
      RECT 37.255 3.63 37.585 3.708 ;
      RECT 37.255 3.657 37.59 3.678 ;
      RECT 37.38 3.535 37.475 3.767 ;
      RECT 37.01 2.58 37.015 3.118 ;
      RECT 36.815 2.91 36.82 3.105 ;
      RECT 35.115 2.575 35.13 2.955 ;
      RECT 37.18 2.575 37.185 2.745 ;
      RECT 37.175 2.575 37.18 2.755 ;
      RECT 37.17 2.575 37.175 2.768 ;
      RECT 37.145 2.575 37.17 2.81 ;
      RECT 37.12 2.575 37.145 2.883 ;
      RECT 37.105 2.575 37.12 2.935 ;
      RECT 37.1 2.575 37.105 2.965 ;
      RECT 37.075 2.575 37.1 3.005 ;
      RECT 37.06 2.575 37.075 3.06 ;
      RECT 37.055 2.575 37.06 3.093 ;
      RECT 37.03 2.575 37.055 3.113 ;
      RECT 37.015 2.575 37.03 3.119 ;
      RECT 36.945 2.61 37.01 3.115 ;
      RECT 36.895 2.665 36.945 3.11 ;
      RECT 36.885 2.697 36.895 3.108 ;
      RECT 36.88 2.722 36.885 3.108 ;
      RECT 36.86 2.795 36.88 3.108 ;
      RECT 36.85 2.875 36.86 3.107 ;
      RECT 36.835 2.905 36.85 3.107 ;
      RECT 36.82 2.91 36.835 3.106 ;
      RECT 36.76 2.912 36.815 3.103 ;
      RECT 36.73 2.917 36.76 3.099 ;
      RECT 36.728 2.92 36.73 3.098 ;
      RECT 36.642 2.922 36.728 3.095 ;
      RECT 36.556 2.928 36.642 3.089 ;
      RECT 36.47 2.933 36.556 3.083 ;
      RECT 36.397 2.938 36.47 3.084 ;
      RECT 36.311 2.944 36.397 3.092 ;
      RECT 36.225 2.95 36.311 3.101 ;
      RECT 36.205 2.954 36.225 3.106 ;
      RECT 36.158 2.956 36.205 3.109 ;
      RECT 36.072 2.961 36.158 3.115 ;
      RECT 35.986 2.966 36.072 3.124 ;
      RECT 35.9 2.972 35.986 3.132 ;
      RECT 35.815 2.97 35.9 3.141 ;
      RECT 35.811 2.965 35.815 3.145 ;
      RECT 35.725 2.96 35.811 3.137 ;
      RECT 35.661 2.951 35.725 3.125 ;
      RECT 35.575 2.942 35.661 3.112 ;
      RECT 35.551 2.935 35.575 3.103 ;
      RECT 35.465 2.929 35.551 3.09 ;
      RECT 35.425 2.922 35.465 3.076 ;
      RECT 35.42 2.912 35.425 3.072 ;
      RECT 35.41 2.9 35.42 3.071 ;
      RECT 35.39 2.87 35.41 3.068 ;
      RECT 35.335 2.79 35.39 3.062 ;
      RECT 35.315 2.709 35.335 3.057 ;
      RECT 35.295 2.667 35.315 3.053 ;
      RECT 35.27 2.62 35.295 3.047 ;
      RECT 35.265 2.595 35.27 3.044 ;
      RECT 35.23 2.575 35.265 3.039 ;
      RECT 35.221 2.575 35.23 3.032 ;
      RECT 35.135 2.575 35.221 3.002 ;
      RECT 35.13 2.575 35.135 2.965 ;
      RECT 35.095 2.575 35.115 2.887 ;
      RECT 35.09 2.617 35.095 2.852 ;
      RECT 35.085 2.692 35.09 2.808 ;
      RECT 36.535 2.497 36.71 2.745 ;
      RECT 36.535 2.497 36.715 2.743 ;
      RECT 36.53 2.529 36.715 2.703 ;
      RECT 36.56 2.47 36.73 2.69 ;
      RECT 36.525 2.547 36.73 2.623 ;
      RECT 35.835 2.01 36.005 2.185 ;
      RECT 35.835 2.01 36.177 2.177 ;
      RECT 35.835 2.01 36.26 2.171 ;
      RECT 35.835 2.01 36.295 2.167 ;
      RECT 35.835 2.01 36.315 2.166 ;
      RECT 35.835 2.01 36.401 2.162 ;
      RECT 36.295 1.835 36.465 2.157 ;
      RECT 35.87 1.942 36.495 2.155 ;
      RECT 35.86 1.997 36.5 2.153 ;
      RECT 35.835 2.033 36.51 2.148 ;
      RECT 35.835 2.06 36.515 2.078 ;
      RECT 35.9 1.885 36.475 2.155 ;
      RECT 36.091 1.87 36.475 2.155 ;
      RECT 35.925 1.873 36.475 2.155 ;
      RECT 36.005 1.871 36.091 2.182 ;
      RECT 36.091 1.868 36.47 2.155 ;
      RECT 36.275 1.845 36.47 2.155 ;
      RECT 36.177 1.866 36.47 2.155 ;
      RECT 36.26 1.86 36.275 2.168 ;
      RECT 36.41 3.225 36.415 3.425 ;
      RECT 35.875 3.29 35.92 3.425 ;
      RECT 36.445 3.225 36.465 3.398 ;
      RECT 36.415 3.225 36.445 3.413 ;
      RECT 36.35 3.225 36.41 3.45 ;
      RECT 36.335 3.225 36.35 3.48 ;
      RECT 36.32 3.225 36.335 3.493 ;
      RECT 36.3 3.225 36.32 3.508 ;
      RECT 36.295 3.225 36.3 3.517 ;
      RECT 36.285 3.229 36.295 3.522 ;
      RECT 36.27 3.239 36.285 3.533 ;
      RECT 36.245 3.255 36.27 3.543 ;
      RECT 36.235 3.269 36.245 3.545 ;
      RECT 36.215 3.281 36.235 3.542 ;
      RECT 36.185 3.302 36.215 3.536 ;
      RECT 36.175 3.314 36.185 3.531 ;
      RECT 36.165 3.312 36.175 3.528 ;
      RECT 36.15 3.311 36.165 3.523 ;
      RECT 36.145 3.31 36.15 3.518 ;
      RECT 36.11 3.308 36.145 3.508 ;
      RECT 36.09 3.305 36.11 3.49 ;
      RECT 36.08 3.303 36.09 3.485 ;
      RECT 36.07 3.302 36.08 3.48 ;
      RECT 36.035 3.3 36.07 3.468 ;
      RECT 35.98 3.296 36.035 3.448 ;
      RECT 35.97 3.294 35.98 3.433 ;
      RECT 35.965 3.294 35.97 3.428 ;
      RECT 35.92 3.292 35.965 3.425 ;
      RECT 35.825 3.29 35.875 3.429 ;
      RECT 35.815 3.291 35.825 3.434 ;
      RECT 35.755 3.298 35.815 3.448 ;
      RECT 35.73 3.306 35.755 3.468 ;
      RECT 35.72 3.31 35.73 3.48 ;
      RECT 35.715 3.311 35.72 3.485 ;
      RECT 35.7 3.313 35.715 3.488 ;
      RECT 35.685 3.315 35.7 3.493 ;
      RECT 35.68 3.315 35.685 3.496 ;
      RECT 35.635 3.32 35.68 3.507 ;
      RECT 35.63 3.324 35.635 3.519 ;
      RECT 35.605 3.32 35.63 3.523 ;
      RECT 35.595 3.316 35.605 3.527 ;
      RECT 35.585 3.315 35.595 3.531 ;
      RECT 35.57 3.305 35.585 3.537 ;
      RECT 35.565 3.293 35.57 3.541 ;
      RECT 35.56 3.29 35.565 3.542 ;
      RECT 35.555 3.287 35.56 3.544 ;
      RECT 35.54 3.275 35.555 3.543 ;
      RECT 35.525 3.257 35.54 3.54 ;
      RECT 35.505 3.236 35.525 3.533 ;
      RECT 35.44 3.225 35.505 3.505 ;
      RECT 35.436 3.225 35.44 3.484 ;
      RECT 35.35 3.225 35.436 3.454 ;
      RECT 35.335 3.225 35.35 3.41 ;
      RECT 35.91 2.325 35.915 2.56 ;
      RECT 35.04 2.241 35.045 2.445 ;
      RECT 35.62 2.27 35.625 2.425 ;
      RECT 35.54 2.25 35.545 2.425 ;
      RECT 36.21 2.392 36.225 2.745 ;
      RECT 36.136 2.377 36.21 2.745 ;
      RECT 36.05 2.36 36.136 2.745 ;
      RECT 36.04 2.35 36.05 2.743 ;
      RECT 36.035 2.348 36.04 2.738 ;
      RECT 36.02 2.346 36.035 2.724 ;
      RECT 35.95 2.338 36.02 2.664 ;
      RECT 35.93 2.329 35.95 2.598 ;
      RECT 35.925 2.326 35.93 2.578 ;
      RECT 35.915 2.325 35.925 2.568 ;
      RECT 35.905 2.325 35.91 2.552 ;
      RECT 35.895 2.324 35.905 2.542 ;
      RECT 35.885 2.322 35.895 2.53 ;
      RECT 35.87 2.319 35.885 2.51 ;
      RECT 35.86 2.317 35.87 2.495 ;
      RECT 35.84 2.314 35.86 2.483 ;
      RECT 35.835 2.312 35.84 2.473 ;
      RECT 35.81 2.31 35.835 2.46 ;
      RECT 35.78 2.305 35.81 2.445 ;
      RECT 35.7 2.296 35.78 2.436 ;
      RECT 35.655 2.285 35.7 2.429 ;
      RECT 35.635 2.276 35.655 2.426 ;
      RECT 35.625 2.271 35.635 2.425 ;
      RECT 35.58 2.265 35.62 2.425 ;
      RECT 35.565 2.257 35.58 2.425 ;
      RECT 35.545 2.252 35.565 2.425 ;
      RECT 35.525 2.249 35.54 2.425 ;
      RECT 35.442 2.248 35.525 2.424 ;
      RECT 35.356 2.247 35.442 2.42 ;
      RECT 35.27 2.245 35.356 2.417 ;
      RECT 35.217 2.244 35.27 2.419 ;
      RECT 35.131 2.243 35.217 2.428 ;
      RECT 35.045 2.242 35.131 2.44 ;
      RECT 35.025 2.241 35.04 2.448 ;
      RECT 34.945 2.24 35.025 2.46 ;
      RECT 34.92 2.24 34.945 2.473 ;
      RECT 34.895 2.24 34.92 2.488 ;
      RECT 34.89 2.24 34.895 2.51 ;
      RECT 34.885 2.24 34.89 2.528 ;
      RECT 34.88 2.24 34.885 2.545 ;
      RECT 34.875 2.24 34.88 2.558 ;
      RECT 34.87 2.24 34.875 2.568 ;
      RECT 34.83 2.24 34.87 2.653 ;
      RECT 34.815 2.24 34.83 2.738 ;
      RECT 34.805 2.241 34.815 2.75 ;
      RECT 34.77 2.246 34.805 2.755 ;
      RECT 34.73 2.255 34.77 2.755 ;
      RECT 34.715 2.265 34.73 2.755 ;
      RECT 34.71 2.275 34.715 2.755 ;
      RECT 34.69 2.302 34.71 2.755 ;
      RECT 34.64 2.385 34.69 2.755 ;
      RECT 34.635 2.447 34.64 2.755 ;
      RECT 34.625 2.46 34.635 2.755 ;
      RECT 34.615 2.482 34.625 2.755 ;
      RECT 34.605 2.507 34.615 2.75 ;
      RECT 34.6 2.545 34.605 2.743 ;
      RECT 34.59 2.655 34.6 2.738 ;
      RECT 35.985 3.576 36 3.835 ;
      RECT 35.985 3.591 36.005 3.834 ;
      RECT 35.901 3.591 36.005 3.832 ;
      RECT 35.901 3.605 36.01 3.831 ;
      RECT 35.815 3.647 36.015 3.828 ;
      RECT 35.81 3.59 36 3.823 ;
      RECT 35.81 3.661 36.02 3.82 ;
      RECT 35.805 3.692 36.02 3.818 ;
      RECT 35.81 3.689 36.035 3.808 ;
      RECT 35.805 3.735 36.05 3.793 ;
      RECT 35.805 3.763 36.055 3.778 ;
      RECT 35.815 3.565 35.985 3.828 ;
      RECT 35.575 2.575 35.745 2.745 ;
      RECT 35.54 2.575 35.745 2.74 ;
      RECT 35.53 2.575 35.745 2.733 ;
      RECT 35.525 2.56 35.695 2.73 ;
      RECT 34.355 3.097 34.62 3.54 ;
      RECT 34.35 3.068 34.565 3.538 ;
      RECT 34.345 3.222 34.625 3.533 ;
      RECT 34.35 3.117 34.625 3.533 ;
      RECT 34.35 3.128 34.635 3.52 ;
      RECT 34.35 3.075 34.595 3.538 ;
      RECT 34.355 3.062 34.565 3.54 ;
      RECT 34.355 3.06 34.515 3.54 ;
      RECT 34.456 3.052 34.515 3.54 ;
      RECT 34.37 3.053 34.515 3.54 ;
      RECT 34.456 3.051 34.505 3.54 ;
      RECT 34.26 1.866 34.435 2.165 ;
      RECT 34.31 1.828 34.435 2.165 ;
      RECT 34.295 1.83 34.521 2.157 ;
      RECT 34.295 1.833 34.56 2.144 ;
      RECT 34.295 1.834 34.57 2.13 ;
      RECT 34.25 1.885 34.57 2.12 ;
      RECT 34.295 1.835 34.575 2.115 ;
      RECT 34.25 2.045 34.58 2.105 ;
      RECT 34.235 1.905 34.575 2.045 ;
      RECT 34.23 1.921 34.575 1.985 ;
      RECT 34.275 1.845 34.575 2.115 ;
      RECT 34.31 1.826 34.396 2.165 ;
      RECT 32.77 5.02 32.94 6.49 ;
      RECT 32.77 6.315 32.945 6.485 ;
      RECT 32.4 1.74 32.57 2.93 ;
      RECT 32.4 1.74 32.87 1.91 ;
      RECT 32.4 6.97 32.87 7.14 ;
      RECT 32.4 5.95 32.57 7.14 ;
      RECT 31.41 1.74 31.58 2.93 ;
      RECT 31.41 1.74 31.88 1.91 ;
      RECT 31.41 6.97 31.88 7.14 ;
      RECT 31.41 5.95 31.58 7.14 ;
      RECT 29.56 2.635 29.73 3.865 ;
      RECT 29.615 0.855 29.785 2.805 ;
      RECT 29.56 0.575 29.73 1.025 ;
      RECT 29.56 7.855 29.73 8.305 ;
      RECT 29.615 6.075 29.785 8.025 ;
      RECT 29.56 5.015 29.73 6.245 ;
      RECT 29.04 0.575 29.21 3.865 ;
      RECT 29.04 2.075 29.445 2.405 ;
      RECT 29.04 1.235 29.445 1.565 ;
      RECT 29.04 5.015 29.21 8.305 ;
      RECT 29.04 7.315 29.445 7.645 ;
      RECT 29.04 6.475 29.445 6.805 ;
      RECT 26.965 3.126 26.97 3.298 ;
      RECT 26.96 3.119 26.965 3.388 ;
      RECT 26.955 3.113 26.96 3.407 ;
      RECT 26.935 3.107 26.955 3.417 ;
      RECT 26.92 3.102 26.935 3.425 ;
      RECT 26.883 3.096 26.92 3.423 ;
      RECT 26.797 3.082 26.883 3.419 ;
      RECT 26.711 3.064 26.797 3.414 ;
      RECT 26.625 3.045 26.711 3.408 ;
      RECT 26.595 3.033 26.625 3.404 ;
      RECT 26.575 3.027 26.595 3.403 ;
      RECT 26.51 3.025 26.575 3.401 ;
      RECT 26.495 3.025 26.51 3.393 ;
      RECT 26.48 3.025 26.495 3.38 ;
      RECT 26.475 3.025 26.48 3.37 ;
      RECT 26.46 3.025 26.475 3.348 ;
      RECT 26.445 3.025 26.46 3.315 ;
      RECT 26.44 3.025 26.445 3.293 ;
      RECT 26.43 3.025 26.44 3.275 ;
      RECT 26.415 3.025 26.43 3.253 ;
      RECT 26.395 3.025 26.415 3.215 ;
      RECT 26.745 2.31 26.78 2.749 ;
      RECT 26.745 2.31 26.785 2.748 ;
      RECT 26.69 2.37 26.785 2.747 ;
      RECT 26.555 2.542 26.785 2.746 ;
      RECT 26.665 2.42 26.785 2.746 ;
      RECT 26.555 2.542 26.81 2.736 ;
      RECT 26.61 2.487 26.89 2.653 ;
      RECT 26.785 2.281 26.79 2.744 ;
      RECT 26.64 2.457 26.93 2.53 ;
      RECT 26.655 2.44 26.785 2.746 ;
      RECT 26.79 2.28 26.96 2.468 ;
      RECT 26.78 2.283 26.96 2.468 ;
      RECT 26.285 2.16 26.455 2.47 ;
      RECT 26.285 2.16 26.46 2.443 ;
      RECT 26.285 2.16 26.465 2.42 ;
      RECT 26.285 2.16 26.475 2.37 ;
      RECT 26.28 2.265 26.475 2.34 ;
      RECT 26.315 1.835 26.485 2.313 ;
      RECT 26.315 1.835 26.5 2.234 ;
      RECT 26.305 2.045 26.5 2.234 ;
      RECT 26.315 1.845 26.51 2.149 ;
      RECT 26.245 2.587 26.25 2.79 ;
      RECT 26.235 2.575 26.245 2.9 ;
      RECT 26.21 2.575 26.235 2.94 ;
      RECT 26.13 2.575 26.21 3.025 ;
      RECT 26.12 2.575 26.13 3.095 ;
      RECT 26.095 2.575 26.12 3.118 ;
      RECT 26.075 2.575 26.095 3.153 ;
      RECT 26.03 2.585 26.075 3.196 ;
      RECT 26.02 2.597 26.03 3.233 ;
      RECT 26 2.611 26.02 3.253 ;
      RECT 25.99 2.629 26 3.269 ;
      RECT 25.975 2.655 25.99 3.279 ;
      RECT 25.96 2.696 25.975 3.293 ;
      RECT 25.95 2.731 25.96 3.303 ;
      RECT 25.945 2.747 25.95 3.308 ;
      RECT 25.935 2.762 25.945 3.313 ;
      RECT 25.915 2.805 25.935 3.323 ;
      RECT 25.895 2.842 25.915 3.336 ;
      RECT 25.86 2.865 25.895 3.354 ;
      RECT 25.85 2.879 25.86 3.37 ;
      RECT 25.83 2.889 25.85 3.38 ;
      RECT 25.825 2.898 25.83 3.388 ;
      RECT 25.815 2.905 25.825 3.395 ;
      RECT 25.805 2.912 25.815 3.403 ;
      RECT 25.79 2.922 25.805 3.411 ;
      RECT 25.78 2.936 25.79 3.421 ;
      RECT 25.77 2.948 25.78 3.433 ;
      RECT 25.755 2.97 25.77 3.446 ;
      RECT 25.745 2.992 25.755 3.457 ;
      RECT 25.735 3.012 25.745 3.466 ;
      RECT 25.73 3.027 25.735 3.473 ;
      RECT 25.7 3.06 25.73 3.487 ;
      RECT 25.69 3.095 25.7 3.502 ;
      RECT 25.685 3.102 25.69 3.508 ;
      RECT 25.665 3.117 25.685 3.515 ;
      RECT 25.66 3.132 25.665 3.523 ;
      RECT 25.655 3.141 25.66 3.528 ;
      RECT 25.64 3.147 25.655 3.535 ;
      RECT 25.635 3.153 25.64 3.543 ;
      RECT 25.63 3.157 25.635 3.55 ;
      RECT 25.625 3.161 25.63 3.56 ;
      RECT 25.615 3.166 25.625 3.57 ;
      RECT 25.595 3.177 25.615 3.598 ;
      RECT 25.58 3.189 25.595 3.625 ;
      RECT 25.56 3.202 25.58 3.65 ;
      RECT 25.54 3.217 25.56 3.674 ;
      RECT 25.525 3.232 25.54 3.689 ;
      RECT 25.52 3.243 25.525 3.698 ;
      RECT 25.455 3.288 25.52 3.708 ;
      RECT 25.42 3.347 25.455 3.721 ;
      RECT 25.415 3.37 25.42 3.727 ;
      RECT 25.41 3.377 25.415 3.729 ;
      RECT 25.395 3.387 25.41 3.732 ;
      RECT 25.365 3.412 25.395 3.736 ;
      RECT 25.36 3.43 25.365 3.74 ;
      RECT 25.355 3.437 25.36 3.741 ;
      RECT 25.335 3.445 25.355 3.745 ;
      RECT 25.325 3.452 25.335 3.749 ;
      RECT 25.281 3.463 25.325 3.756 ;
      RECT 25.195 3.491 25.281 3.772 ;
      RECT 25.135 3.515 25.195 3.79 ;
      RECT 25.09 3.525 25.135 3.804 ;
      RECT 25.031 3.533 25.09 3.818 ;
      RECT 24.945 3.54 25.031 3.837 ;
      RECT 24.92 3.545 24.945 3.852 ;
      RECT 24.84 3.548 24.92 3.855 ;
      RECT 24.76 3.552 24.84 3.842 ;
      RECT 24.751 3.555 24.76 3.827 ;
      RECT 24.665 3.555 24.751 3.812 ;
      RECT 24.605 3.557 24.665 3.789 ;
      RECT 24.601 3.56 24.605 3.779 ;
      RECT 24.515 3.56 24.601 3.764 ;
      RECT 24.44 3.56 24.515 3.74 ;
      RECT 25.755 2.569 25.765 2.745 ;
      RECT 25.71 2.536 25.755 2.745 ;
      RECT 25.665 2.487 25.71 2.745 ;
      RECT 25.635 2.457 25.665 2.746 ;
      RECT 25.63 2.44 25.635 2.747 ;
      RECT 25.605 2.42 25.63 2.748 ;
      RECT 25.59 2.395 25.605 2.749 ;
      RECT 25.585 2.382 25.59 2.75 ;
      RECT 25.58 2.376 25.585 2.748 ;
      RECT 25.575 2.368 25.58 2.742 ;
      RECT 25.55 2.36 25.575 2.722 ;
      RECT 25.53 2.349 25.55 2.693 ;
      RECT 25.5 2.334 25.53 2.664 ;
      RECT 25.48 2.32 25.5 2.636 ;
      RECT 25.47 2.314 25.48 2.615 ;
      RECT 25.465 2.311 25.47 2.598 ;
      RECT 25.46 2.308 25.465 2.583 ;
      RECT 25.445 2.303 25.46 2.548 ;
      RECT 25.44 2.299 25.445 2.515 ;
      RECT 25.42 2.294 25.44 2.491 ;
      RECT 25.39 2.286 25.42 2.456 ;
      RECT 25.375 2.28 25.39 2.433 ;
      RECT 25.335 2.273 25.375 2.418 ;
      RECT 25.31 2.265 25.335 2.398 ;
      RECT 25.29 2.26 25.31 2.388 ;
      RECT 25.255 2.254 25.29 2.383 ;
      RECT 25.21 2.245 25.255 2.382 ;
      RECT 25.18 2.241 25.21 2.384 ;
      RECT 25.095 2.249 25.18 2.388 ;
      RECT 25.025 2.26 25.095 2.41 ;
      RECT 25.012 2.266 25.025 2.433 ;
      RECT 24.926 2.273 25.012 2.455 ;
      RECT 24.84 2.285 24.926 2.492 ;
      RECT 24.84 2.662 24.85 2.9 ;
      RECT 24.835 2.291 24.84 2.515 ;
      RECT 24.83 2.547 24.84 2.9 ;
      RECT 24.83 2.292 24.835 2.52 ;
      RECT 24.825 2.293 24.83 2.9 ;
      RECT 24.801 2.295 24.825 2.901 ;
      RECT 24.715 2.303 24.801 2.903 ;
      RECT 24.695 2.317 24.715 2.906 ;
      RECT 24.69 2.345 24.695 2.907 ;
      RECT 24.685 2.357 24.69 2.908 ;
      RECT 24.68 2.372 24.685 2.909 ;
      RECT 24.67 2.402 24.68 2.91 ;
      RECT 24.665 2.44 24.67 2.908 ;
      RECT 24.66 2.46 24.665 2.903 ;
      RECT 24.645 2.495 24.66 2.888 ;
      RECT 24.635 2.547 24.645 2.868 ;
      RECT 24.63 2.577 24.635 2.856 ;
      RECT 24.615 2.59 24.63 2.839 ;
      RECT 24.59 2.594 24.615 2.806 ;
      RECT 24.575 2.592 24.59 2.783 ;
      RECT 24.56 2.591 24.575 2.78 ;
      RECT 24.5 2.589 24.56 2.778 ;
      RECT 24.49 2.587 24.5 2.773 ;
      RECT 24.45 2.586 24.49 2.77 ;
      RECT 24.38 2.583 24.45 2.768 ;
      RECT 24.325 2.581 24.38 2.763 ;
      RECT 24.255 2.575 24.325 2.758 ;
      RECT 24.246 2.575 24.255 2.755 ;
      RECT 24.16 2.575 24.246 2.75 ;
      RECT 24.155 2.575 24.16 2.745 ;
      RECT 25.46 1.81 25.635 2.16 ;
      RECT 25.46 1.825 25.645 2.158 ;
      RECT 25.435 1.775 25.58 2.155 ;
      RECT 25.415 1.776 25.58 2.148 ;
      RECT 25.405 1.777 25.59 2.143 ;
      RECT 25.375 1.778 25.59 2.13 ;
      RECT 25.325 1.779 25.59 2.106 ;
      RECT 25.32 1.781 25.59 2.091 ;
      RECT 25.32 1.847 25.65 2.085 ;
      RECT 25.3 1.788 25.605 2.065 ;
      RECT 25.29 1.797 25.615 1.92 ;
      RECT 25.3 1.792 25.615 2.065 ;
      RECT 25.32 1.782 25.605 2.091 ;
      RECT 24.905 3.107 25.075 3.395 ;
      RECT 24.9 3.125 25.085 3.39 ;
      RECT 24.865 3.133 25.15 3.31 ;
      RECT 24.865 3.133 25.236 3.3 ;
      RECT 24.865 3.133 25.29 3.246 ;
      RECT 25.15 3.03 25.32 3.214 ;
      RECT 24.865 3.185 25.325 3.202 ;
      RECT 24.85 3.155 25.32 3.198 ;
      RECT 25.11 3.037 25.15 3.349 ;
      RECT 24.99 3.074 25.32 3.214 ;
      RECT 25.085 3.049 25.11 3.375 ;
      RECT 25.075 3.056 25.32 3.214 ;
      RECT 25.206 2.52 25.275 2.779 ;
      RECT 25.206 2.575 25.28 2.778 ;
      RECT 25.12 2.575 25.28 2.777 ;
      RECT 25.115 2.575 25.285 2.77 ;
      RECT 25.105 2.52 25.275 2.765 ;
      RECT 24.485 1.819 24.66 2.12 ;
      RECT 24.47 1.807 24.485 2.105 ;
      RECT 24.44 1.806 24.47 2.058 ;
      RECT 24.44 1.824 24.665 2.053 ;
      RECT 24.425 1.808 24.485 2.018 ;
      RECT 24.42 1.83 24.675 1.918 ;
      RECT 24.42 1.813 24.571 1.918 ;
      RECT 24.42 1.815 24.575 1.918 ;
      RECT 24.425 1.811 24.571 2.018 ;
      RECT 24.53 3.047 24.535 3.395 ;
      RECT 24.52 3.037 24.53 3.401 ;
      RECT 24.485 3.027 24.52 3.403 ;
      RECT 24.447 3.022 24.485 3.407 ;
      RECT 24.361 3.015 24.447 3.414 ;
      RECT 24.275 3.005 24.361 3.424 ;
      RECT 24.23 3 24.275 3.432 ;
      RECT 24.226 3 24.23 3.436 ;
      RECT 24.14 3 24.226 3.443 ;
      RECT 24.125 3 24.14 3.443 ;
      RECT 24.115 2.998 24.125 3.415 ;
      RECT 24.105 2.994 24.115 3.358 ;
      RECT 24.085 2.988 24.105 3.29 ;
      RECT 24.08 2.984 24.085 3.238 ;
      RECT 24.07 2.983 24.08 3.205 ;
      RECT 24.02 2.981 24.07 3.19 ;
      RECT 23.995 2.979 24.02 3.185 ;
      RECT 23.952 2.977 23.995 3.181 ;
      RECT 23.866 2.973 23.952 3.169 ;
      RECT 23.78 2.968 23.866 3.153 ;
      RECT 23.75 2.965 23.78 3.14 ;
      RECT 23.725 2.964 23.75 3.128 ;
      RECT 23.72 2.964 23.725 3.118 ;
      RECT 23.68 2.963 23.72 3.11 ;
      RECT 23.665 2.962 23.68 3.103 ;
      RECT 23.615 2.961 23.665 3.095 ;
      RECT 23.613 2.96 23.615 3.09 ;
      RECT 23.527 2.958 23.613 3.09 ;
      RECT 23.441 2.953 23.527 3.09 ;
      RECT 23.355 2.949 23.441 3.09 ;
      RECT 23.306 2.945 23.355 3.088 ;
      RECT 23.22 2.942 23.306 3.083 ;
      RECT 23.197 2.939 23.22 3.079 ;
      RECT 23.111 2.936 23.197 3.074 ;
      RECT 23.025 2.932 23.111 3.065 ;
      RECT 23 2.925 23.025 3.06 ;
      RECT 22.94 2.89 23 3.057 ;
      RECT 22.92 2.815 22.94 3.054 ;
      RECT 22.915 2.757 22.92 3.053 ;
      RECT 22.89 2.697 22.915 3.052 ;
      RECT 22.815 2.575 22.89 3.048 ;
      RECT 22.805 2.575 22.815 3.04 ;
      RECT 22.79 2.575 22.805 3.03 ;
      RECT 22.775 2.575 22.79 3 ;
      RECT 22.76 2.575 22.775 2.945 ;
      RECT 22.745 2.575 22.76 2.883 ;
      RECT 22.72 2.575 22.745 2.808 ;
      RECT 22.715 2.575 22.72 2.758 ;
      RECT 24.06 2.12 24.08 2.429 ;
      RECT 24.046 2.122 24.095 2.426 ;
      RECT 24.046 2.127 24.115 2.417 ;
      RECT 23.96 2.125 24.095 2.411 ;
      RECT 23.96 2.133 24.15 2.394 ;
      RECT 23.925 2.135 24.15 2.393 ;
      RECT 23.895 2.143 24.15 2.384 ;
      RECT 23.885 2.148 24.17 2.37 ;
      RECT 23.925 2.138 24.17 2.37 ;
      RECT 23.925 2.141 24.18 2.358 ;
      RECT 23.895 2.143 24.19 2.345 ;
      RECT 23.895 2.147 24.2 2.288 ;
      RECT 23.885 2.152 24.205 2.203 ;
      RECT 24.046 2.12 24.08 2.426 ;
      RECT 23.925 7.855 24.095 8.305 ;
      RECT 23.98 6.075 24.15 8.025 ;
      RECT 23.925 5.015 24.095 6.245 ;
      RECT 23.485 2.223 23.49 2.435 ;
      RECT 23.36 2.22 23.375 2.435 ;
      RECT 22.825 2.25 22.895 2.435 ;
      RECT 22.71 2.25 22.745 2.43 ;
      RECT 23.831 2.552 23.85 2.746 ;
      RECT 23.745 2.507 23.831 2.747 ;
      RECT 23.735 2.46 23.745 2.749 ;
      RECT 23.73 2.44 23.735 2.75 ;
      RECT 23.71 2.405 23.73 2.751 ;
      RECT 23.695 2.355 23.71 2.752 ;
      RECT 23.675 2.292 23.695 2.753 ;
      RECT 23.665 2.255 23.675 2.754 ;
      RECT 23.65 2.244 23.665 2.755 ;
      RECT 23.645 2.236 23.65 2.753 ;
      RECT 23.635 2.235 23.645 2.745 ;
      RECT 23.605 2.232 23.635 2.724 ;
      RECT 23.53 2.227 23.605 2.669 ;
      RECT 23.515 2.223 23.53 2.615 ;
      RECT 23.505 2.223 23.515 2.51 ;
      RECT 23.49 2.223 23.505 2.443 ;
      RECT 23.475 2.223 23.485 2.433 ;
      RECT 23.42 2.222 23.475 2.43 ;
      RECT 23.375 2.22 23.42 2.433 ;
      RECT 23.347 2.22 23.36 2.436 ;
      RECT 23.261 2.224 23.347 2.438 ;
      RECT 23.175 2.23 23.261 2.443 ;
      RECT 23.155 2.234 23.175 2.445 ;
      RECT 23.153 2.235 23.155 2.444 ;
      RECT 23.067 2.237 23.153 2.443 ;
      RECT 22.981 2.242 23.067 2.44 ;
      RECT 22.895 2.247 22.981 2.437 ;
      RECT 22.745 2.25 22.825 2.433 ;
      RECT 23.405 5.015 23.575 8.305 ;
      RECT 23.405 7.315 23.81 7.645 ;
      RECT 23.405 6.475 23.81 6.805 ;
      RECT 23.521 3.225 23.57 3.559 ;
      RECT 23.521 3.225 23.575 3.558 ;
      RECT 23.435 3.225 23.575 3.557 ;
      RECT 23.21 3.333 23.58 3.555 ;
      RECT 23.435 3.225 23.605 3.548 ;
      RECT 23.405 3.237 23.61 3.539 ;
      RECT 23.39 3.255 23.615 3.536 ;
      RECT 23.205 3.339 23.615 3.463 ;
      RECT 23.2 3.346 23.615 3.423 ;
      RECT 23.215 3.312 23.615 3.536 ;
      RECT 23.376 3.258 23.58 3.555 ;
      RECT 23.29 3.278 23.615 3.536 ;
      RECT 23.39 3.252 23.61 3.539 ;
      RECT 23.16 2.576 23.35 2.77 ;
      RECT 23.155 2.578 23.35 2.769 ;
      RECT 23.15 2.582 23.365 2.766 ;
      RECT 23.165 2.575 23.365 2.766 ;
      RECT 23.15 2.685 23.37 2.761 ;
      RECT 22.445 3.185 22.536 3.483 ;
      RECT 22.44 3.187 22.615 3.478 ;
      RECT 22.445 3.185 22.615 3.478 ;
      RECT 22.44 3.191 22.635 3.476 ;
      RECT 22.44 3.246 22.675 3.475 ;
      RECT 22.44 3.281 22.69 3.469 ;
      RECT 22.44 3.315 22.7 3.459 ;
      RECT 22.43 3.195 22.635 3.31 ;
      RECT 22.43 3.215 22.65 3.31 ;
      RECT 22.43 3.198 22.64 3.31 ;
      RECT 22.655 1.966 22.66 2.028 ;
      RECT 22.65 1.888 22.655 2.051 ;
      RECT 22.645 1.845 22.65 2.062 ;
      RECT 22.64 1.835 22.645 2.074 ;
      RECT 22.635 1.835 22.64 2.083 ;
      RECT 22.61 1.835 22.635 2.115 ;
      RECT 22.605 1.835 22.61 2.148 ;
      RECT 22.59 1.835 22.605 2.173 ;
      RECT 22.58 1.835 22.59 2.2 ;
      RECT 22.575 1.835 22.58 2.213 ;
      RECT 22.57 1.835 22.575 2.228 ;
      RECT 22.56 1.835 22.57 2.243 ;
      RECT 22.555 1.835 22.56 2.263 ;
      RECT 22.53 1.835 22.555 2.298 ;
      RECT 22.485 1.835 22.53 2.343 ;
      RECT 22.475 1.835 22.485 2.356 ;
      RECT 22.39 1.92 22.475 2.363 ;
      RECT 22.355 2.042 22.39 2.372 ;
      RECT 22.35 2.082 22.355 2.376 ;
      RECT 22.33 2.105 22.35 2.378 ;
      RECT 22.325 2.135 22.33 2.381 ;
      RECT 22.315 2.147 22.325 2.382 ;
      RECT 22.27 2.17 22.315 2.387 ;
      RECT 22.23 2.2 22.27 2.395 ;
      RECT 22.195 2.212 22.23 2.401 ;
      RECT 22.19 2.217 22.195 2.405 ;
      RECT 22.12 2.227 22.19 2.412 ;
      RECT 22.08 2.237 22.12 2.422 ;
      RECT 22.06 2.242 22.08 2.428 ;
      RECT 22.05 2.246 22.06 2.433 ;
      RECT 22.045 2.249 22.05 2.436 ;
      RECT 22.035 2.25 22.045 2.437 ;
      RECT 22.01 2.252 22.035 2.441 ;
      RECT 22 2.257 22.01 2.444 ;
      RECT 21.955 2.265 22 2.445 ;
      RECT 21.83 2.27 21.955 2.445 ;
      RECT 22.385 2.567 22.405 2.749 ;
      RECT 22.336 2.552 22.385 2.748 ;
      RECT 22.25 2.567 22.405 2.746 ;
      RECT 22.235 2.567 22.405 2.745 ;
      RECT 22.2 2.545 22.37 2.73 ;
      RECT 22.27 3.565 22.285 3.774 ;
      RECT 22.27 3.573 22.29 3.773 ;
      RECT 22.215 3.573 22.29 3.772 ;
      RECT 22.195 3.577 22.295 3.77 ;
      RECT 22.175 3.527 22.215 3.769 ;
      RECT 22.12 3.585 22.3 3.767 ;
      RECT 22.085 3.542 22.215 3.765 ;
      RECT 22.081 3.545 22.27 3.764 ;
      RECT 21.995 3.553 22.27 3.762 ;
      RECT 21.995 3.597 22.305 3.755 ;
      RECT 21.985 3.69 22.305 3.753 ;
      RECT 21.995 3.609 22.31 3.738 ;
      RECT 21.995 3.63 22.325 3.708 ;
      RECT 21.995 3.657 22.33 3.678 ;
      RECT 22.12 3.535 22.215 3.767 ;
      RECT 21.75 2.58 21.755 3.118 ;
      RECT 21.555 2.91 21.56 3.105 ;
      RECT 19.855 2.575 19.87 2.955 ;
      RECT 21.92 2.575 21.925 2.745 ;
      RECT 21.915 2.575 21.92 2.755 ;
      RECT 21.91 2.575 21.915 2.768 ;
      RECT 21.885 2.575 21.91 2.81 ;
      RECT 21.86 2.575 21.885 2.883 ;
      RECT 21.845 2.575 21.86 2.935 ;
      RECT 21.84 2.575 21.845 2.965 ;
      RECT 21.815 2.575 21.84 3.005 ;
      RECT 21.8 2.575 21.815 3.06 ;
      RECT 21.795 2.575 21.8 3.093 ;
      RECT 21.77 2.575 21.795 3.113 ;
      RECT 21.755 2.575 21.77 3.119 ;
      RECT 21.685 2.61 21.75 3.115 ;
      RECT 21.635 2.665 21.685 3.11 ;
      RECT 21.625 2.697 21.635 3.108 ;
      RECT 21.62 2.722 21.625 3.108 ;
      RECT 21.6 2.795 21.62 3.108 ;
      RECT 21.59 2.875 21.6 3.107 ;
      RECT 21.575 2.905 21.59 3.107 ;
      RECT 21.56 2.91 21.575 3.106 ;
      RECT 21.5 2.912 21.555 3.103 ;
      RECT 21.47 2.917 21.5 3.099 ;
      RECT 21.468 2.92 21.47 3.098 ;
      RECT 21.382 2.922 21.468 3.095 ;
      RECT 21.296 2.928 21.382 3.089 ;
      RECT 21.21 2.933 21.296 3.083 ;
      RECT 21.137 2.938 21.21 3.084 ;
      RECT 21.051 2.944 21.137 3.092 ;
      RECT 20.965 2.95 21.051 3.101 ;
      RECT 20.945 2.954 20.965 3.106 ;
      RECT 20.898 2.956 20.945 3.109 ;
      RECT 20.812 2.961 20.898 3.115 ;
      RECT 20.726 2.966 20.812 3.124 ;
      RECT 20.64 2.972 20.726 3.132 ;
      RECT 20.555 2.97 20.64 3.141 ;
      RECT 20.551 2.965 20.555 3.145 ;
      RECT 20.465 2.96 20.551 3.137 ;
      RECT 20.401 2.951 20.465 3.125 ;
      RECT 20.315 2.942 20.401 3.112 ;
      RECT 20.291 2.935 20.315 3.103 ;
      RECT 20.205 2.929 20.291 3.09 ;
      RECT 20.165 2.922 20.205 3.076 ;
      RECT 20.16 2.912 20.165 3.072 ;
      RECT 20.15 2.9 20.16 3.071 ;
      RECT 20.13 2.87 20.15 3.068 ;
      RECT 20.075 2.79 20.13 3.062 ;
      RECT 20.055 2.709 20.075 3.057 ;
      RECT 20.035 2.667 20.055 3.053 ;
      RECT 20.01 2.62 20.035 3.047 ;
      RECT 20.005 2.595 20.01 3.044 ;
      RECT 19.97 2.575 20.005 3.039 ;
      RECT 19.961 2.575 19.97 3.032 ;
      RECT 19.875 2.575 19.961 3.002 ;
      RECT 19.87 2.575 19.875 2.965 ;
      RECT 19.835 2.575 19.855 2.887 ;
      RECT 19.83 2.617 19.835 2.852 ;
      RECT 19.825 2.692 19.83 2.808 ;
      RECT 21.275 2.497 21.45 2.745 ;
      RECT 21.275 2.497 21.455 2.743 ;
      RECT 21.27 2.529 21.455 2.703 ;
      RECT 21.3 2.47 21.47 2.69 ;
      RECT 21.265 2.547 21.47 2.623 ;
      RECT 20.575 2.01 20.745 2.185 ;
      RECT 20.575 2.01 20.917 2.177 ;
      RECT 20.575 2.01 21 2.171 ;
      RECT 20.575 2.01 21.035 2.167 ;
      RECT 20.575 2.01 21.055 2.166 ;
      RECT 20.575 2.01 21.141 2.162 ;
      RECT 21.035 1.835 21.205 2.157 ;
      RECT 20.61 1.942 21.235 2.155 ;
      RECT 20.6 1.997 21.24 2.153 ;
      RECT 20.575 2.033 21.25 2.148 ;
      RECT 20.575 2.06 21.255 2.078 ;
      RECT 20.64 1.885 21.215 2.155 ;
      RECT 20.831 1.87 21.215 2.155 ;
      RECT 20.665 1.873 21.215 2.155 ;
      RECT 20.745 1.871 20.831 2.182 ;
      RECT 20.831 1.868 21.21 2.155 ;
      RECT 21.015 1.845 21.21 2.155 ;
      RECT 20.917 1.866 21.21 2.155 ;
      RECT 21 1.86 21.015 2.168 ;
      RECT 21.15 3.225 21.155 3.425 ;
      RECT 20.615 3.29 20.66 3.425 ;
      RECT 21.185 3.225 21.205 3.398 ;
      RECT 21.155 3.225 21.185 3.413 ;
      RECT 21.09 3.225 21.15 3.45 ;
      RECT 21.075 3.225 21.09 3.48 ;
      RECT 21.06 3.225 21.075 3.493 ;
      RECT 21.04 3.225 21.06 3.508 ;
      RECT 21.035 3.225 21.04 3.517 ;
      RECT 21.025 3.229 21.035 3.522 ;
      RECT 21.01 3.239 21.025 3.533 ;
      RECT 20.985 3.255 21.01 3.543 ;
      RECT 20.975 3.269 20.985 3.545 ;
      RECT 20.955 3.281 20.975 3.542 ;
      RECT 20.925 3.302 20.955 3.536 ;
      RECT 20.915 3.314 20.925 3.531 ;
      RECT 20.905 3.312 20.915 3.528 ;
      RECT 20.89 3.311 20.905 3.523 ;
      RECT 20.885 3.31 20.89 3.518 ;
      RECT 20.85 3.308 20.885 3.508 ;
      RECT 20.83 3.305 20.85 3.49 ;
      RECT 20.82 3.303 20.83 3.485 ;
      RECT 20.81 3.302 20.82 3.48 ;
      RECT 20.775 3.3 20.81 3.468 ;
      RECT 20.72 3.296 20.775 3.448 ;
      RECT 20.71 3.294 20.72 3.433 ;
      RECT 20.705 3.294 20.71 3.428 ;
      RECT 20.66 3.292 20.705 3.425 ;
      RECT 20.565 3.29 20.615 3.429 ;
      RECT 20.555 3.291 20.565 3.434 ;
      RECT 20.495 3.298 20.555 3.448 ;
      RECT 20.47 3.306 20.495 3.468 ;
      RECT 20.46 3.31 20.47 3.48 ;
      RECT 20.455 3.311 20.46 3.485 ;
      RECT 20.44 3.313 20.455 3.488 ;
      RECT 20.425 3.315 20.44 3.493 ;
      RECT 20.42 3.315 20.425 3.496 ;
      RECT 20.375 3.32 20.42 3.507 ;
      RECT 20.37 3.324 20.375 3.519 ;
      RECT 20.345 3.32 20.37 3.523 ;
      RECT 20.335 3.316 20.345 3.527 ;
      RECT 20.325 3.315 20.335 3.531 ;
      RECT 20.31 3.305 20.325 3.537 ;
      RECT 20.305 3.293 20.31 3.541 ;
      RECT 20.3 3.29 20.305 3.542 ;
      RECT 20.295 3.287 20.3 3.544 ;
      RECT 20.28 3.275 20.295 3.543 ;
      RECT 20.265 3.257 20.28 3.54 ;
      RECT 20.245 3.236 20.265 3.533 ;
      RECT 20.18 3.225 20.245 3.505 ;
      RECT 20.176 3.225 20.18 3.484 ;
      RECT 20.09 3.225 20.176 3.454 ;
      RECT 20.075 3.225 20.09 3.41 ;
      RECT 20.65 2.325 20.655 2.56 ;
      RECT 19.78 2.241 19.785 2.445 ;
      RECT 20.36 2.27 20.365 2.425 ;
      RECT 20.28 2.25 20.285 2.425 ;
      RECT 20.95 2.392 20.965 2.745 ;
      RECT 20.876 2.377 20.95 2.745 ;
      RECT 20.79 2.36 20.876 2.745 ;
      RECT 20.78 2.35 20.79 2.743 ;
      RECT 20.775 2.348 20.78 2.738 ;
      RECT 20.76 2.346 20.775 2.724 ;
      RECT 20.69 2.338 20.76 2.664 ;
      RECT 20.67 2.329 20.69 2.598 ;
      RECT 20.665 2.326 20.67 2.578 ;
      RECT 20.655 2.325 20.665 2.568 ;
      RECT 20.645 2.325 20.65 2.552 ;
      RECT 20.635 2.324 20.645 2.542 ;
      RECT 20.625 2.322 20.635 2.53 ;
      RECT 20.61 2.319 20.625 2.51 ;
      RECT 20.6 2.317 20.61 2.495 ;
      RECT 20.58 2.314 20.6 2.483 ;
      RECT 20.575 2.312 20.58 2.473 ;
      RECT 20.55 2.31 20.575 2.46 ;
      RECT 20.52 2.305 20.55 2.445 ;
      RECT 20.44 2.296 20.52 2.436 ;
      RECT 20.395 2.285 20.44 2.429 ;
      RECT 20.375 2.276 20.395 2.426 ;
      RECT 20.365 2.271 20.375 2.425 ;
      RECT 20.32 2.265 20.36 2.425 ;
      RECT 20.305 2.257 20.32 2.425 ;
      RECT 20.285 2.252 20.305 2.425 ;
      RECT 20.265 2.249 20.28 2.425 ;
      RECT 20.182 2.248 20.265 2.424 ;
      RECT 20.096 2.247 20.182 2.42 ;
      RECT 20.01 2.245 20.096 2.417 ;
      RECT 19.957 2.244 20.01 2.419 ;
      RECT 19.871 2.243 19.957 2.428 ;
      RECT 19.785 2.242 19.871 2.44 ;
      RECT 19.765 2.241 19.78 2.448 ;
      RECT 19.685 2.24 19.765 2.46 ;
      RECT 19.66 2.24 19.685 2.473 ;
      RECT 19.635 2.24 19.66 2.488 ;
      RECT 19.63 2.24 19.635 2.51 ;
      RECT 19.625 2.24 19.63 2.528 ;
      RECT 19.62 2.24 19.625 2.545 ;
      RECT 19.615 2.24 19.62 2.558 ;
      RECT 19.61 2.24 19.615 2.568 ;
      RECT 19.57 2.24 19.61 2.653 ;
      RECT 19.555 2.24 19.57 2.738 ;
      RECT 19.545 2.241 19.555 2.75 ;
      RECT 19.51 2.246 19.545 2.755 ;
      RECT 19.47 2.255 19.51 2.755 ;
      RECT 19.455 2.265 19.47 2.755 ;
      RECT 19.45 2.275 19.455 2.755 ;
      RECT 19.43 2.302 19.45 2.755 ;
      RECT 19.38 2.385 19.43 2.755 ;
      RECT 19.375 2.447 19.38 2.755 ;
      RECT 19.365 2.46 19.375 2.755 ;
      RECT 19.355 2.482 19.365 2.755 ;
      RECT 19.345 2.507 19.355 2.75 ;
      RECT 19.34 2.545 19.345 2.743 ;
      RECT 19.33 2.655 19.34 2.738 ;
      RECT 20.725 3.576 20.74 3.835 ;
      RECT 20.725 3.591 20.745 3.834 ;
      RECT 20.641 3.591 20.745 3.832 ;
      RECT 20.641 3.605 20.75 3.831 ;
      RECT 20.555 3.647 20.755 3.828 ;
      RECT 20.55 3.59 20.74 3.823 ;
      RECT 20.55 3.661 20.76 3.82 ;
      RECT 20.545 3.692 20.76 3.818 ;
      RECT 20.55 3.689 20.775 3.808 ;
      RECT 20.545 3.735 20.79 3.793 ;
      RECT 20.545 3.763 20.795 3.778 ;
      RECT 20.555 3.565 20.725 3.828 ;
      RECT 20.315 2.575 20.485 2.745 ;
      RECT 20.28 2.575 20.485 2.74 ;
      RECT 20.27 2.575 20.485 2.733 ;
      RECT 20.265 2.56 20.435 2.73 ;
      RECT 19.095 3.097 19.36 3.54 ;
      RECT 19.09 3.068 19.305 3.538 ;
      RECT 19.085 3.222 19.365 3.533 ;
      RECT 19.09 3.117 19.365 3.533 ;
      RECT 19.09 3.128 19.375 3.52 ;
      RECT 19.09 3.075 19.335 3.538 ;
      RECT 19.095 3.062 19.305 3.54 ;
      RECT 19.095 3.06 19.255 3.54 ;
      RECT 19.196 3.052 19.255 3.54 ;
      RECT 19.11 3.053 19.255 3.54 ;
      RECT 19.196 3.051 19.245 3.54 ;
      RECT 19 1.866 19.175 2.165 ;
      RECT 19.05 1.828 19.175 2.165 ;
      RECT 19.035 1.83 19.261 2.157 ;
      RECT 19.035 1.833 19.3 2.144 ;
      RECT 19.035 1.834 19.31 2.13 ;
      RECT 18.99 1.885 19.31 2.12 ;
      RECT 19.035 1.835 19.315 2.115 ;
      RECT 18.99 2.045 19.32 2.105 ;
      RECT 18.975 1.905 19.315 2.045 ;
      RECT 18.97 1.921 19.315 1.985 ;
      RECT 19.015 1.845 19.315 2.115 ;
      RECT 19.05 1.826 19.136 2.165 ;
      RECT 17.51 5.02 17.68 6.49 ;
      RECT 17.51 6.315 17.685 6.485 ;
      RECT 17.14 1.74 17.31 2.93 ;
      RECT 17.14 1.74 17.61 1.91 ;
      RECT 17.14 6.97 17.61 7.14 ;
      RECT 17.14 5.95 17.31 7.14 ;
      RECT 16.15 1.74 16.32 2.93 ;
      RECT 16.15 1.74 16.62 1.91 ;
      RECT 16.15 6.97 16.62 7.14 ;
      RECT 16.15 5.95 16.32 7.14 ;
      RECT 14.3 2.635 14.47 3.865 ;
      RECT 14.355 0.855 14.525 2.805 ;
      RECT 14.3 0.575 14.47 1.025 ;
      RECT 14.3 7.855 14.47 8.305 ;
      RECT 14.355 6.075 14.525 8.025 ;
      RECT 14.3 5.015 14.47 6.245 ;
      RECT 13.78 0.575 13.95 3.865 ;
      RECT 13.78 2.075 14.185 2.405 ;
      RECT 13.78 1.235 14.185 1.565 ;
      RECT 13.78 5.015 13.95 8.305 ;
      RECT 13.78 7.315 14.185 7.645 ;
      RECT 13.78 6.475 14.185 6.805 ;
      RECT 11.705 3.126 11.71 3.298 ;
      RECT 11.7 3.119 11.705 3.388 ;
      RECT 11.695 3.113 11.7 3.407 ;
      RECT 11.675 3.107 11.695 3.417 ;
      RECT 11.66 3.102 11.675 3.425 ;
      RECT 11.623 3.096 11.66 3.423 ;
      RECT 11.537 3.082 11.623 3.419 ;
      RECT 11.451 3.064 11.537 3.414 ;
      RECT 11.365 3.045 11.451 3.408 ;
      RECT 11.335 3.033 11.365 3.404 ;
      RECT 11.315 3.027 11.335 3.403 ;
      RECT 11.25 3.025 11.315 3.401 ;
      RECT 11.235 3.025 11.25 3.393 ;
      RECT 11.22 3.025 11.235 3.38 ;
      RECT 11.215 3.025 11.22 3.37 ;
      RECT 11.2 3.025 11.215 3.348 ;
      RECT 11.185 3.025 11.2 3.315 ;
      RECT 11.18 3.025 11.185 3.293 ;
      RECT 11.17 3.025 11.18 3.275 ;
      RECT 11.155 3.025 11.17 3.253 ;
      RECT 11.135 3.025 11.155 3.215 ;
      RECT 11.485 2.31 11.52 2.749 ;
      RECT 11.485 2.31 11.525 2.748 ;
      RECT 11.43 2.37 11.525 2.747 ;
      RECT 11.295 2.542 11.525 2.746 ;
      RECT 11.405 2.42 11.525 2.746 ;
      RECT 11.295 2.542 11.55 2.736 ;
      RECT 11.35 2.487 11.63 2.653 ;
      RECT 11.525 2.281 11.53 2.744 ;
      RECT 11.38 2.457 11.67 2.53 ;
      RECT 11.395 2.44 11.525 2.746 ;
      RECT 11.53 2.28 11.7 2.468 ;
      RECT 11.52 2.283 11.7 2.468 ;
      RECT 11.025 2.16 11.195 2.47 ;
      RECT 11.025 2.16 11.2 2.443 ;
      RECT 11.025 2.16 11.205 2.42 ;
      RECT 11.025 2.16 11.215 2.37 ;
      RECT 11.02 2.265 11.215 2.34 ;
      RECT 11.055 1.835 11.225 2.313 ;
      RECT 11.055 1.835 11.24 2.234 ;
      RECT 11.045 2.045 11.24 2.234 ;
      RECT 11.055 1.845 11.25 2.149 ;
      RECT 10.985 2.587 10.99 2.79 ;
      RECT 10.975 2.575 10.985 2.9 ;
      RECT 10.95 2.575 10.975 2.94 ;
      RECT 10.87 2.575 10.95 3.025 ;
      RECT 10.86 2.575 10.87 3.095 ;
      RECT 10.835 2.575 10.86 3.118 ;
      RECT 10.815 2.575 10.835 3.153 ;
      RECT 10.77 2.585 10.815 3.196 ;
      RECT 10.76 2.597 10.77 3.233 ;
      RECT 10.74 2.611 10.76 3.253 ;
      RECT 10.73 2.629 10.74 3.269 ;
      RECT 10.715 2.655 10.73 3.279 ;
      RECT 10.7 2.696 10.715 3.293 ;
      RECT 10.69 2.731 10.7 3.303 ;
      RECT 10.685 2.747 10.69 3.308 ;
      RECT 10.675 2.762 10.685 3.313 ;
      RECT 10.655 2.805 10.675 3.323 ;
      RECT 10.635 2.842 10.655 3.336 ;
      RECT 10.6 2.865 10.635 3.354 ;
      RECT 10.59 2.879 10.6 3.37 ;
      RECT 10.57 2.889 10.59 3.38 ;
      RECT 10.565 2.898 10.57 3.388 ;
      RECT 10.555 2.905 10.565 3.395 ;
      RECT 10.545 2.912 10.555 3.403 ;
      RECT 10.53 2.922 10.545 3.411 ;
      RECT 10.52 2.936 10.53 3.421 ;
      RECT 10.51 2.948 10.52 3.433 ;
      RECT 10.495 2.97 10.51 3.446 ;
      RECT 10.485 2.992 10.495 3.457 ;
      RECT 10.475 3.012 10.485 3.466 ;
      RECT 10.47 3.027 10.475 3.473 ;
      RECT 10.44 3.06 10.47 3.487 ;
      RECT 10.43 3.095 10.44 3.502 ;
      RECT 10.425 3.102 10.43 3.508 ;
      RECT 10.405 3.117 10.425 3.515 ;
      RECT 10.4 3.132 10.405 3.523 ;
      RECT 10.395 3.141 10.4 3.528 ;
      RECT 10.38 3.147 10.395 3.535 ;
      RECT 10.375 3.153 10.38 3.543 ;
      RECT 10.37 3.157 10.375 3.55 ;
      RECT 10.365 3.161 10.37 3.56 ;
      RECT 10.355 3.166 10.365 3.57 ;
      RECT 10.335 3.177 10.355 3.598 ;
      RECT 10.32 3.189 10.335 3.625 ;
      RECT 10.3 3.202 10.32 3.65 ;
      RECT 10.28 3.217 10.3 3.674 ;
      RECT 10.265 3.232 10.28 3.689 ;
      RECT 10.26 3.243 10.265 3.698 ;
      RECT 10.195 3.288 10.26 3.708 ;
      RECT 10.16 3.347 10.195 3.721 ;
      RECT 10.155 3.37 10.16 3.727 ;
      RECT 10.15 3.377 10.155 3.729 ;
      RECT 10.135 3.387 10.15 3.732 ;
      RECT 10.105 3.412 10.135 3.736 ;
      RECT 10.1 3.43 10.105 3.74 ;
      RECT 10.095 3.437 10.1 3.741 ;
      RECT 10.075 3.445 10.095 3.745 ;
      RECT 10.065 3.452 10.075 3.749 ;
      RECT 10.021 3.463 10.065 3.756 ;
      RECT 9.935 3.491 10.021 3.772 ;
      RECT 9.875 3.515 9.935 3.79 ;
      RECT 9.83 3.525 9.875 3.804 ;
      RECT 9.771 3.533 9.83 3.818 ;
      RECT 9.685 3.54 9.771 3.837 ;
      RECT 9.66 3.545 9.685 3.852 ;
      RECT 9.58 3.548 9.66 3.855 ;
      RECT 9.5 3.552 9.58 3.842 ;
      RECT 9.491 3.555 9.5 3.827 ;
      RECT 9.405 3.555 9.491 3.812 ;
      RECT 9.345 3.557 9.405 3.789 ;
      RECT 9.341 3.56 9.345 3.779 ;
      RECT 9.255 3.56 9.341 3.764 ;
      RECT 9.18 3.56 9.255 3.74 ;
      RECT 10.495 2.569 10.505 2.745 ;
      RECT 10.45 2.536 10.495 2.745 ;
      RECT 10.405 2.487 10.45 2.745 ;
      RECT 10.375 2.457 10.405 2.746 ;
      RECT 10.37 2.44 10.375 2.747 ;
      RECT 10.345 2.42 10.37 2.748 ;
      RECT 10.33 2.395 10.345 2.749 ;
      RECT 10.325 2.382 10.33 2.75 ;
      RECT 10.32 2.376 10.325 2.748 ;
      RECT 10.315 2.368 10.32 2.742 ;
      RECT 10.29 2.36 10.315 2.722 ;
      RECT 10.27 2.349 10.29 2.693 ;
      RECT 10.24 2.334 10.27 2.664 ;
      RECT 10.22 2.32 10.24 2.636 ;
      RECT 10.21 2.314 10.22 2.615 ;
      RECT 10.205 2.311 10.21 2.598 ;
      RECT 10.2 2.308 10.205 2.583 ;
      RECT 10.185 2.303 10.2 2.548 ;
      RECT 10.18 2.299 10.185 2.515 ;
      RECT 10.16 2.294 10.18 2.491 ;
      RECT 10.13 2.286 10.16 2.456 ;
      RECT 10.115 2.28 10.13 2.433 ;
      RECT 10.075 2.273 10.115 2.418 ;
      RECT 10.05 2.265 10.075 2.398 ;
      RECT 10.03 2.26 10.05 2.388 ;
      RECT 9.995 2.254 10.03 2.383 ;
      RECT 9.95 2.245 9.995 2.382 ;
      RECT 9.92 2.241 9.95 2.384 ;
      RECT 9.835 2.249 9.92 2.388 ;
      RECT 9.765 2.26 9.835 2.41 ;
      RECT 9.752 2.266 9.765 2.433 ;
      RECT 9.666 2.273 9.752 2.455 ;
      RECT 9.58 2.285 9.666 2.492 ;
      RECT 9.58 2.662 9.59 2.9 ;
      RECT 9.575 2.291 9.58 2.515 ;
      RECT 9.57 2.547 9.58 2.9 ;
      RECT 9.57 2.292 9.575 2.52 ;
      RECT 9.565 2.293 9.57 2.9 ;
      RECT 9.541 2.295 9.565 2.901 ;
      RECT 9.455 2.303 9.541 2.903 ;
      RECT 9.435 2.317 9.455 2.906 ;
      RECT 9.43 2.345 9.435 2.907 ;
      RECT 9.425 2.357 9.43 2.908 ;
      RECT 9.42 2.372 9.425 2.909 ;
      RECT 9.41 2.402 9.42 2.91 ;
      RECT 9.405 2.44 9.41 2.908 ;
      RECT 9.4 2.46 9.405 2.903 ;
      RECT 9.385 2.495 9.4 2.888 ;
      RECT 9.375 2.547 9.385 2.868 ;
      RECT 9.37 2.577 9.375 2.856 ;
      RECT 9.355 2.59 9.37 2.839 ;
      RECT 9.33 2.594 9.355 2.806 ;
      RECT 9.315 2.592 9.33 2.783 ;
      RECT 9.3 2.591 9.315 2.78 ;
      RECT 9.24 2.589 9.3 2.778 ;
      RECT 9.23 2.587 9.24 2.773 ;
      RECT 9.19 2.586 9.23 2.77 ;
      RECT 9.12 2.583 9.19 2.768 ;
      RECT 9.065 2.581 9.12 2.763 ;
      RECT 8.995 2.575 9.065 2.758 ;
      RECT 8.986 2.575 8.995 2.755 ;
      RECT 8.9 2.575 8.986 2.75 ;
      RECT 8.895 2.575 8.9 2.745 ;
      RECT 10.2 1.81 10.375 2.16 ;
      RECT 10.2 1.825 10.385 2.158 ;
      RECT 10.175 1.775 10.32 2.155 ;
      RECT 10.155 1.776 10.32 2.148 ;
      RECT 10.145 1.777 10.33 2.143 ;
      RECT 10.115 1.778 10.33 2.13 ;
      RECT 10.065 1.779 10.33 2.106 ;
      RECT 10.06 1.781 10.33 2.091 ;
      RECT 10.06 1.847 10.39 2.085 ;
      RECT 10.04 1.788 10.345 2.065 ;
      RECT 10.03 1.797 10.355 1.92 ;
      RECT 10.04 1.792 10.355 2.065 ;
      RECT 10.06 1.782 10.345 2.091 ;
      RECT 9.645 3.107 9.815 3.395 ;
      RECT 9.64 3.125 9.825 3.39 ;
      RECT 9.605 3.133 9.89 3.31 ;
      RECT 9.605 3.133 9.976 3.3 ;
      RECT 9.605 3.133 10.03 3.246 ;
      RECT 9.89 3.03 10.06 3.214 ;
      RECT 9.605 3.185 10.065 3.202 ;
      RECT 9.59 3.155 10.06 3.198 ;
      RECT 9.85 3.037 9.89 3.349 ;
      RECT 9.73 3.074 10.06 3.214 ;
      RECT 9.825 3.049 9.85 3.375 ;
      RECT 9.815 3.056 10.06 3.214 ;
      RECT 9.946 2.52 10.015 2.779 ;
      RECT 9.946 2.575 10.02 2.778 ;
      RECT 9.86 2.575 10.02 2.777 ;
      RECT 9.855 2.575 10.025 2.77 ;
      RECT 9.845 2.52 10.015 2.765 ;
      RECT 9.225 1.819 9.4 2.12 ;
      RECT 9.21 1.807 9.225 2.105 ;
      RECT 9.18 1.806 9.21 2.058 ;
      RECT 9.18 1.824 9.405 2.053 ;
      RECT 9.165 1.808 9.225 2.018 ;
      RECT 9.16 1.83 9.415 1.918 ;
      RECT 9.16 1.813 9.311 1.918 ;
      RECT 9.16 1.815 9.315 1.918 ;
      RECT 9.165 1.811 9.311 2.018 ;
      RECT 9.27 3.047 9.275 3.395 ;
      RECT 9.26 3.037 9.27 3.401 ;
      RECT 9.225 3.027 9.26 3.403 ;
      RECT 9.187 3.022 9.225 3.407 ;
      RECT 9.101 3.015 9.187 3.414 ;
      RECT 9.015 3.005 9.101 3.424 ;
      RECT 8.97 3 9.015 3.432 ;
      RECT 8.966 3 8.97 3.436 ;
      RECT 8.88 3 8.966 3.443 ;
      RECT 8.865 3 8.88 3.443 ;
      RECT 8.855 2.998 8.865 3.415 ;
      RECT 8.845 2.994 8.855 3.358 ;
      RECT 8.825 2.988 8.845 3.29 ;
      RECT 8.82 2.984 8.825 3.238 ;
      RECT 8.81 2.983 8.82 3.205 ;
      RECT 8.76 2.981 8.81 3.19 ;
      RECT 8.735 2.979 8.76 3.185 ;
      RECT 8.692 2.977 8.735 3.181 ;
      RECT 8.606 2.973 8.692 3.169 ;
      RECT 8.52 2.968 8.606 3.153 ;
      RECT 8.49 2.965 8.52 3.14 ;
      RECT 8.465 2.964 8.49 3.128 ;
      RECT 8.46 2.964 8.465 3.118 ;
      RECT 8.42 2.963 8.46 3.11 ;
      RECT 8.405 2.962 8.42 3.103 ;
      RECT 8.355 2.961 8.405 3.095 ;
      RECT 8.353 2.96 8.355 3.09 ;
      RECT 8.267 2.958 8.353 3.09 ;
      RECT 8.181 2.953 8.267 3.09 ;
      RECT 8.095 2.949 8.181 3.09 ;
      RECT 8.046 2.945 8.095 3.088 ;
      RECT 7.96 2.942 8.046 3.083 ;
      RECT 7.937 2.939 7.96 3.079 ;
      RECT 7.851 2.936 7.937 3.074 ;
      RECT 7.765 2.932 7.851 3.065 ;
      RECT 7.74 2.925 7.765 3.06 ;
      RECT 7.68 2.89 7.74 3.057 ;
      RECT 7.66 2.815 7.68 3.054 ;
      RECT 7.655 2.757 7.66 3.053 ;
      RECT 7.63 2.697 7.655 3.052 ;
      RECT 7.555 2.575 7.63 3.048 ;
      RECT 7.545 2.575 7.555 3.04 ;
      RECT 7.53 2.575 7.545 3.03 ;
      RECT 7.515 2.575 7.53 3 ;
      RECT 7.5 2.575 7.515 2.945 ;
      RECT 7.485 2.575 7.5 2.883 ;
      RECT 7.46 2.575 7.485 2.808 ;
      RECT 7.455 2.575 7.46 2.758 ;
      RECT 8.8 2.12 8.82 2.429 ;
      RECT 8.786 2.122 8.835 2.426 ;
      RECT 8.786 2.127 8.855 2.417 ;
      RECT 8.7 2.125 8.835 2.411 ;
      RECT 8.7 2.133 8.89 2.394 ;
      RECT 8.665 2.135 8.89 2.393 ;
      RECT 8.635 2.143 8.89 2.384 ;
      RECT 8.625 2.148 8.91 2.37 ;
      RECT 8.665 2.138 8.91 2.37 ;
      RECT 8.665 2.141 8.92 2.358 ;
      RECT 8.635 2.143 8.93 2.345 ;
      RECT 8.635 2.147 8.94 2.288 ;
      RECT 8.625 2.152 8.945 2.203 ;
      RECT 8.786 2.12 8.82 2.426 ;
      RECT 8.665 7.855 8.835 8.305 ;
      RECT 8.72 6.075 8.89 8.025 ;
      RECT 8.665 5.015 8.835 6.245 ;
      RECT 8.225 2.223 8.23 2.435 ;
      RECT 8.1 2.22 8.115 2.435 ;
      RECT 7.565 2.25 7.635 2.435 ;
      RECT 7.45 2.25 7.485 2.43 ;
      RECT 8.571 2.552 8.59 2.746 ;
      RECT 8.485 2.507 8.571 2.747 ;
      RECT 8.475 2.46 8.485 2.749 ;
      RECT 8.47 2.44 8.475 2.75 ;
      RECT 8.45 2.405 8.47 2.751 ;
      RECT 8.435 2.355 8.45 2.752 ;
      RECT 8.415 2.292 8.435 2.753 ;
      RECT 8.405 2.255 8.415 2.754 ;
      RECT 8.39 2.244 8.405 2.755 ;
      RECT 8.385 2.236 8.39 2.753 ;
      RECT 8.375 2.235 8.385 2.745 ;
      RECT 8.345 2.232 8.375 2.724 ;
      RECT 8.27 2.227 8.345 2.669 ;
      RECT 8.255 2.223 8.27 2.615 ;
      RECT 8.245 2.223 8.255 2.51 ;
      RECT 8.23 2.223 8.245 2.443 ;
      RECT 8.215 2.223 8.225 2.433 ;
      RECT 8.16 2.222 8.215 2.43 ;
      RECT 8.115 2.22 8.16 2.433 ;
      RECT 8.087 2.22 8.1 2.436 ;
      RECT 8.001 2.224 8.087 2.438 ;
      RECT 7.915 2.23 8.001 2.443 ;
      RECT 7.895 2.234 7.915 2.445 ;
      RECT 7.893 2.235 7.895 2.444 ;
      RECT 7.807 2.237 7.893 2.443 ;
      RECT 7.721 2.242 7.807 2.44 ;
      RECT 7.635 2.247 7.721 2.437 ;
      RECT 7.485 2.25 7.565 2.433 ;
      RECT 8.145 5.015 8.315 8.305 ;
      RECT 8.145 7.315 8.55 7.645 ;
      RECT 8.145 6.475 8.55 6.805 ;
      RECT 8.261 3.225 8.31 3.559 ;
      RECT 8.261 3.225 8.315 3.558 ;
      RECT 8.175 3.225 8.315 3.557 ;
      RECT 7.95 3.333 8.32 3.555 ;
      RECT 8.175 3.225 8.345 3.548 ;
      RECT 8.145 3.237 8.35 3.539 ;
      RECT 8.13 3.255 8.355 3.536 ;
      RECT 7.945 3.339 8.355 3.463 ;
      RECT 7.94 3.346 8.355 3.423 ;
      RECT 7.955 3.312 8.355 3.536 ;
      RECT 8.116 3.258 8.32 3.555 ;
      RECT 8.03 3.278 8.355 3.536 ;
      RECT 8.13 3.252 8.35 3.539 ;
      RECT 7.9 2.576 8.09 2.77 ;
      RECT 7.895 2.578 8.09 2.769 ;
      RECT 7.89 2.582 8.105 2.766 ;
      RECT 7.905 2.575 8.105 2.766 ;
      RECT 7.89 2.685 8.11 2.761 ;
      RECT 7.185 3.185 7.276 3.483 ;
      RECT 7.18 3.187 7.355 3.478 ;
      RECT 7.185 3.185 7.355 3.478 ;
      RECT 7.18 3.191 7.375 3.476 ;
      RECT 7.18 3.246 7.415 3.475 ;
      RECT 7.18 3.281 7.43 3.469 ;
      RECT 7.18 3.315 7.44 3.459 ;
      RECT 7.17 3.195 7.375 3.31 ;
      RECT 7.17 3.215 7.39 3.31 ;
      RECT 7.17 3.198 7.38 3.31 ;
      RECT 7.395 1.966 7.4 2.028 ;
      RECT 7.39 1.888 7.395 2.051 ;
      RECT 7.385 1.845 7.39 2.062 ;
      RECT 7.38 1.835 7.385 2.074 ;
      RECT 7.375 1.835 7.38 2.083 ;
      RECT 7.35 1.835 7.375 2.115 ;
      RECT 7.345 1.835 7.35 2.148 ;
      RECT 7.33 1.835 7.345 2.173 ;
      RECT 7.32 1.835 7.33 2.2 ;
      RECT 7.315 1.835 7.32 2.213 ;
      RECT 7.31 1.835 7.315 2.228 ;
      RECT 7.3 1.835 7.31 2.243 ;
      RECT 7.295 1.835 7.3 2.263 ;
      RECT 7.27 1.835 7.295 2.298 ;
      RECT 7.225 1.835 7.27 2.343 ;
      RECT 7.215 1.835 7.225 2.356 ;
      RECT 7.13 1.92 7.215 2.363 ;
      RECT 7.095 2.042 7.13 2.372 ;
      RECT 7.09 2.082 7.095 2.376 ;
      RECT 7.07 2.105 7.09 2.378 ;
      RECT 7.065 2.135 7.07 2.381 ;
      RECT 7.055 2.147 7.065 2.382 ;
      RECT 7.01 2.17 7.055 2.387 ;
      RECT 6.97 2.2 7.01 2.395 ;
      RECT 6.935 2.212 6.97 2.401 ;
      RECT 6.93 2.217 6.935 2.405 ;
      RECT 6.86 2.227 6.93 2.412 ;
      RECT 6.82 2.237 6.86 2.422 ;
      RECT 6.8 2.242 6.82 2.428 ;
      RECT 6.79 2.246 6.8 2.433 ;
      RECT 6.785 2.249 6.79 2.436 ;
      RECT 6.775 2.25 6.785 2.437 ;
      RECT 6.75 2.252 6.775 2.441 ;
      RECT 6.74 2.257 6.75 2.444 ;
      RECT 6.695 2.265 6.74 2.445 ;
      RECT 6.57 2.27 6.695 2.445 ;
      RECT 7.125 2.567 7.145 2.749 ;
      RECT 7.076 2.552 7.125 2.748 ;
      RECT 6.99 2.567 7.145 2.746 ;
      RECT 6.975 2.567 7.145 2.745 ;
      RECT 6.94 2.545 7.11 2.73 ;
      RECT 7.01 3.565 7.025 3.774 ;
      RECT 7.01 3.573 7.03 3.773 ;
      RECT 6.955 3.573 7.03 3.772 ;
      RECT 6.935 3.577 7.035 3.77 ;
      RECT 6.915 3.527 6.955 3.769 ;
      RECT 6.86 3.585 7.04 3.767 ;
      RECT 6.825 3.542 6.955 3.765 ;
      RECT 6.821 3.545 7.01 3.764 ;
      RECT 6.735 3.553 7.01 3.762 ;
      RECT 6.735 3.597 7.045 3.755 ;
      RECT 6.725 3.69 7.045 3.753 ;
      RECT 6.735 3.609 7.05 3.738 ;
      RECT 6.735 3.63 7.065 3.708 ;
      RECT 6.735 3.657 7.07 3.678 ;
      RECT 6.86 3.535 6.955 3.767 ;
      RECT 6.49 2.58 6.495 3.118 ;
      RECT 6.295 2.91 6.3 3.105 ;
      RECT 4.595 2.575 4.61 2.955 ;
      RECT 6.66 2.575 6.665 2.745 ;
      RECT 6.655 2.575 6.66 2.755 ;
      RECT 6.65 2.575 6.655 2.768 ;
      RECT 6.625 2.575 6.65 2.81 ;
      RECT 6.6 2.575 6.625 2.883 ;
      RECT 6.585 2.575 6.6 2.935 ;
      RECT 6.58 2.575 6.585 2.965 ;
      RECT 6.555 2.575 6.58 3.005 ;
      RECT 6.54 2.575 6.555 3.06 ;
      RECT 6.535 2.575 6.54 3.093 ;
      RECT 6.51 2.575 6.535 3.113 ;
      RECT 6.495 2.575 6.51 3.119 ;
      RECT 6.425 2.61 6.49 3.115 ;
      RECT 6.375 2.665 6.425 3.11 ;
      RECT 6.365 2.697 6.375 3.108 ;
      RECT 6.36 2.722 6.365 3.108 ;
      RECT 6.34 2.795 6.36 3.108 ;
      RECT 6.33 2.875 6.34 3.107 ;
      RECT 6.315 2.905 6.33 3.107 ;
      RECT 6.3 2.91 6.315 3.106 ;
      RECT 6.24 2.912 6.295 3.103 ;
      RECT 6.21 2.917 6.24 3.099 ;
      RECT 6.208 2.92 6.21 3.098 ;
      RECT 6.122 2.922 6.208 3.095 ;
      RECT 6.036 2.928 6.122 3.089 ;
      RECT 5.95 2.933 6.036 3.083 ;
      RECT 5.877 2.938 5.95 3.084 ;
      RECT 5.791 2.944 5.877 3.092 ;
      RECT 5.705 2.95 5.791 3.101 ;
      RECT 5.685 2.954 5.705 3.106 ;
      RECT 5.638 2.956 5.685 3.109 ;
      RECT 5.552 2.961 5.638 3.115 ;
      RECT 5.466 2.966 5.552 3.124 ;
      RECT 5.38 2.972 5.466 3.132 ;
      RECT 5.295 2.97 5.38 3.141 ;
      RECT 5.291 2.965 5.295 3.145 ;
      RECT 5.205 2.96 5.291 3.137 ;
      RECT 5.141 2.951 5.205 3.125 ;
      RECT 5.055 2.942 5.141 3.112 ;
      RECT 5.031 2.935 5.055 3.103 ;
      RECT 4.945 2.929 5.031 3.09 ;
      RECT 4.905 2.922 4.945 3.076 ;
      RECT 4.9 2.912 4.905 3.072 ;
      RECT 4.89 2.9 4.9 3.071 ;
      RECT 4.87 2.87 4.89 3.068 ;
      RECT 4.815 2.79 4.87 3.062 ;
      RECT 4.795 2.709 4.815 3.057 ;
      RECT 4.775 2.667 4.795 3.053 ;
      RECT 4.75 2.62 4.775 3.047 ;
      RECT 4.745 2.595 4.75 3.044 ;
      RECT 4.71 2.575 4.745 3.039 ;
      RECT 4.701 2.575 4.71 3.032 ;
      RECT 4.615 2.575 4.701 3.002 ;
      RECT 4.61 2.575 4.615 2.965 ;
      RECT 4.575 2.575 4.595 2.887 ;
      RECT 4.57 2.617 4.575 2.852 ;
      RECT 4.565 2.692 4.57 2.808 ;
      RECT 6.015 2.497 6.19 2.745 ;
      RECT 6.015 2.497 6.195 2.743 ;
      RECT 6.01 2.529 6.195 2.703 ;
      RECT 6.04 2.47 6.21 2.69 ;
      RECT 6.005 2.547 6.21 2.623 ;
      RECT 5.315 2.01 5.485 2.185 ;
      RECT 5.315 2.01 5.657 2.177 ;
      RECT 5.315 2.01 5.74 2.171 ;
      RECT 5.315 2.01 5.775 2.167 ;
      RECT 5.315 2.01 5.795 2.166 ;
      RECT 5.315 2.01 5.881 2.162 ;
      RECT 5.775 1.835 5.945 2.157 ;
      RECT 5.35 1.942 5.975 2.155 ;
      RECT 5.34 1.997 5.98 2.153 ;
      RECT 5.315 2.033 5.99 2.148 ;
      RECT 5.315 2.06 5.995 2.078 ;
      RECT 5.38 1.885 5.955 2.155 ;
      RECT 5.571 1.87 5.955 2.155 ;
      RECT 5.405 1.873 5.955 2.155 ;
      RECT 5.485 1.871 5.571 2.182 ;
      RECT 5.571 1.868 5.95 2.155 ;
      RECT 5.755 1.845 5.95 2.155 ;
      RECT 5.657 1.866 5.95 2.155 ;
      RECT 5.74 1.86 5.755 2.168 ;
      RECT 5.89 3.225 5.895 3.425 ;
      RECT 5.355 3.29 5.4 3.425 ;
      RECT 5.925 3.225 5.945 3.398 ;
      RECT 5.895 3.225 5.925 3.413 ;
      RECT 5.83 3.225 5.89 3.45 ;
      RECT 5.815 3.225 5.83 3.48 ;
      RECT 5.8 3.225 5.815 3.493 ;
      RECT 5.78 3.225 5.8 3.508 ;
      RECT 5.775 3.225 5.78 3.517 ;
      RECT 5.765 3.229 5.775 3.522 ;
      RECT 5.75 3.239 5.765 3.533 ;
      RECT 5.725 3.255 5.75 3.543 ;
      RECT 5.715 3.269 5.725 3.545 ;
      RECT 5.695 3.281 5.715 3.542 ;
      RECT 5.665 3.302 5.695 3.536 ;
      RECT 5.655 3.314 5.665 3.531 ;
      RECT 5.645 3.312 5.655 3.528 ;
      RECT 5.63 3.311 5.645 3.523 ;
      RECT 5.625 3.31 5.63 3.518 ;
      RECT 5.59 3.308 5.625 3.508 ;
      RECT 5.57 3.305 5.59 3.49 ;
      RECT 5.56 3.303 5.57 3.485 ;
      RECT 5.55 3.302 5.56 3.48 ;
      RECT 5.515 3.3 5.55 3.468 ;
      RECT 5.46 3.296 5.515 3.448 ;
      RECT 5.45 3.294 5.46 3.433 ;
      RECT 5.445 3.294 5.45 3.428 ;
      RECT 5.4 3.292 5.445 3.425 ;
      RECT 5.305 3.29 5.355 3.429 ;
      RECT 5.295 3.291 5.305 3.434 ;
      RECT 5.235 3.298 5.295 3.448 ;
      RECT 5.21 3.306 5.235 3.468 ;
      RECT 5.2 3.31 5.21 3.48 ;
      RECT 5.195 3.311 5.2 3.485 ;
      RECT 5.18 3.313 5.195 3.488 ;
      RECT 5.165 3.315 5.18 3.493 ;
      RECT 5.16 3.315 5.165 3.496 ;
      RECT 5.115 3.32 5.16 3.507 ;
      RECT 5.11 3.324 5.115 3.519 ;
      RECT 5.085 3.32 5.11 3.523 ;
      RECT 5.075 3.316 5.085 3.527 ;
      RECT 5.065 3.315 5.075 3.531 ;
      RECT 5.05 3.305 5.065 3.537 ;
      RECT 5.045 3.293 5.05 3.541 ;
      RECT 5.04 3.29 5.045 3.542 ;
      RECT 5.035 3.287 5.04 3.544 ;
      RECT 5.02 3.275 5.035 3.543 ;
      RECT 5.005 3.257 5.02 3.54 ;
      RECT 4.985 3.236 5.005 3.533 ;
      RECT 4.92 3.225 4.985 3.505 ;
      RECT 4.916 3.225 4.92 3.484 ;
      RECT 4.83 3.225 4.916 3.454 ;
      RECT 4.815 3.225 4.83 3.41 ;
      RECT 5.39 2.325 5.395 2.56 ;
      RECT 4.52 2.241 4.525 2.445 ;
      RECT 5.1 2.27 5.105 2.425 ;
      RECT 5.02 2.25 5.025 2.425 ;
      RECT 5.69 2.392 5.705 2.745 ;
      RECT 5.616 2.377 5.69 2.745 ;
      RECT 5.53 2.36 5.616 2.745 ;
      RECT 5.52 2.35 5.53 2.743 ;
      RECT 5.515 2.348 5.52 2.738 ;
      RECT 5.5 2.346 5.515 2.724 ;
      RECT 5.43 2.338 5.5 2.664 ;
      RECT 5.41 2.329 5.43 2.598 ;
      RECT 5.405 2.326 5.41 2.578 ;
      RECT 5.395 2.325 5.405 2.568 ;
      RECT 5.385 2.325 5.39 2.552 ;
      RECT 5.375 2.324 5.385 2.542 ;
      RECT 5.365 2.322 5.375 2.53 ;
      RECT 5.35 2.319 5.365 2.51 ;
      RECT 5.34 2.317 5.35 2.495 ;
      RECT 5.32 2.314 5.34 2.483 ;
      RECT 5.315 2.312 5.32 2.473 ;
      RECT 5.29 2.31 5.315 2.46 ;
      RECT 5.26 2.305 5.29 2.445 ;
      RECT 5.18 2.296 5.26 2.436 ;
      RECT 5.135 2.285 5.18 2.429 ;
      RECT 5.115 2.276 5.135 2.426 ;
      RECT 5.105 2.271 5.115 2.425 ;
      RECT 5.06 2.265 5.1 2.425 ;
      RECT 5.045 2.257 5.06 2.425 ;
      RECT 5.025 2.252 5.045 2.425 ;
      RECT 5.005 2.249 5.02 2.425 ;
      RECT 4.922 2.248 5.005 2.424 ;
      RECT 4.836 2.247 4.922 2.42 ;
      RECT 4.75 2.245 4.836 2.417 ;
      RECT 4.697 2.244 4.75 2.419 ;
      RECT 4.611 2.243 4.697 2.428 ;
      RECT 4.525 2.242 4.611 2.44 ;
      RECT 4.505 2.241 4.52 2.448 ;
      RECT 4.425 2.24 4.505 2.46 ;
      RECT 4.4 2.24 4.425 2.473 ;
      RECT 4.375 2.24 4.4 2.488 ;
      RECT 4.37 2.24 4.375 2.51 ;
      RECT 4.365 2.24 4.37 2.528 ;
      RECT 4.36 2.24 4.365 2.545 ;
      RECT 4.355 2.24 4.36 2.558 ;
      RECT 4.35 2.24 4.355 2.568 ;
      RECT 4.31 2.24 4.35 2.653 ;
      RECT 4.295 2.24 4.31 2.738 ;
      RECT 4.285 2.241 4.295 2.75 ;
      RECT 4.25 2.246 4.285 2.755 ;
      RECT 4.21 2.255 4.25 2.755 ;
      RECT 4.195 2.265 4.21 2.755 ;
      RECT 4.19 2.275 4.195 2.755 ;
      RECT 4.17 2.302 4.19 2.755 ;
      RECT 4.12 2.385 4.17 2.755 ;
      RECT 4.115 2.447 4.12 2.755 ;
      RECT 4.105 2.46 4.115 2.755 ;
      RECT 4.095 2.482 4.105 2.755 ;
      RECT 4.085 2.507 4.095 2.75 ;
      RECT 4.08 2.545 4.085 2.743 ;
      RECT 4.07 2.655 4.08 2.738 ;
      RECT 5.465 3.576 5.48 3.835 ;
      RECT 5.465 3.591 5.485 3.834 ;
      RECT 5.381 3.591 5.485 3.832 ;
      RECT 5.381 3.605 5.49 3.831 ;
      RECT 5.295 3.647 5.495 3.828 ;
      RECT 5.29 3.59 5.48 3.823 ;
      RECT 5.29 3.661 5.5 3.82 ;
      RECT 5.285 3.692 5.5 3.818 ;
      RECT 5.29 3.689 5.515 3.808 ;
      RECT 5.285 3.735 5.53 3.793 ;
      RECT 5.285 3.763 5.535 3.778 ;
      RECT 5.295 3.565 5.465 3.828 ;
      RECT 5.055 2.575 5.225 2.745 ;
      RECT 5.02 2.575 5.225 2.74 ;
      RECT 5.01 2.575 5.225 2.733 ;
      RECT 5.005 2.56 5.175 2.73 ;
      RECT 3.835 3.097 4.1 3.54 ;
      RECT 3.83 3.068 4.045 3.538 ;
      RECT 3.825 3.222 4.105 3.533 ;
      RECT 3.83 3.117 4.105 3.533 ;
      RECT 3.83 3.128 4.115 3.52 ;
      RECT 3.83 3.075 4.075 3.538 ;
      RECT 3.835 3.062 4.045 3.54 ;
      RECT 3.835 3.06 3.995 3.54 ;
      RECT 3.936 3.052 3.995 3.54 ;
      RECT 3.85 3.053 3.995 3.54 ;
      RECT 3.936 3.051 3.985 3.54 ;
      RECT 3.74 1.866 3.915 2.165 ;
      RECT 3.79 1.828 3.915 2.165 ;
      RECT 3.775 1.83 4.001 2.157 ;
      RECT 3.775 1.833 4.04 2.144 ;
      RECT 3.775 1.834 4.05 2.13 ;
      RECT 3.73 1.885 4.05 2.12 ;
      RECT 3.775 1.835 4.055 2.115 ;
      RECT 3.73 2.045 4.06 2.105 ;
      RECT 3.715 1.905 4.055 2.045 ;
      RECT 3.71 1.921 4.055 1.985 ;
      RECT 3.755 1.845 4.055 2.115 ;
      RECT 3.79 1.826 3.876 2.165 ;
      RECT 1.17 7.855 1.34 8.305 ;
      RECT 1.225 6.075 1.395 8.025 ;
      RECT 1.17 5.015 1.34 6.245 ;
      RECT 0.65 5.015 0.82 8.305 ;
      RECT 0.65 7.315 1.055 7.645 ;
      RECT 0.65 6.475 1.055 6.805 ;
      RECT 78.55 7.8 78.72 8.31 ;
      RECT 77.56 0.57 77.73 1.08 ;
      RECT 77.56 2.39 77.73 3.86 ;
      RECT 77.56 5.02 77.73 6.49 ;
      RECT 77.56 7.8 77.73 8.31 ;
      RECT 76.2 0.575 76.37 3.865 ;
      RECT 76.2 5.015 76.37 8.305 ;
      RECT 75.77 0.575 75.94 1.085 ;
      RECT 75.77 1.655 75.94 3.865 ;
      RECT 75.77 5.015 75.94 7.225 ;
      RECT 75.77 7.795 75.94 8.305 ;
      RECT 70.565 5.015 70.735 8.305 ;
      RECT 70.135 5.015 70.305 7.225 ;
      RECT 70.135 7.795 70.305 8.305 ;
      RECT 63.29 7.8 63.46 8.31 ;
      RECT 62.3 0.57 62.47 1.08 ;
      RECT 62.3 2.39 62.47 3.86 ;
      RECT 62.3 5.02 62.47 6.49 ;
      RECT 62.3 7.8 62.47 8.31 ;
      RECT 60.94 0.575 61.11 3.865 ;
      RECT 60.94 5.015 61.11 8.305 ;
      RECT 60.51 0.575 60.68 1.085 ;
      RECT 60.51 1.655 60.68 3.865 ;
      RECT 60.51 5.015 60.68 7.225 ;
      RECT 60.51 7.795 60.68 8.305 ;
      RECT 55.305 5.015 55.475 8.305 ;
      RECT 54.875 5.015 55.045 7.225 ;
      RECT 54.875 7.795 55.045 8.305 ;
      RECT 48.03 7.8 48.2 8.31 ;
      RECT 47.04 0.57 47.21 1.08 ;
      RECT 47.04 2.39 47.21 3.86 ;
      RECT 47.04 5.02 47.21 6.49 ;
      RECT 47.04 7.8 47.21 8.31 ;
      RECT 45.68 0.575 45.85 3.865 ;
      RECT 45.68 5.015 45.85 8.305 ;
      RECT 45.25 0.575 45.42 1.085 ;
      RECT 45.25 1.655 45.42 3.865 ;
      RECT 45.25 5.015 45.42 7.225 ;
      RECT 45.25 7.795 45.42 8.305 ;
      RECT 40.045 5.015 40.215 8.305 ;
      RECT 39.615 5.015 39.785 7.225 ;
      RECT 39.615 7.795 39.785 8.305 ;
      RECT 32.77 7.8 32.94 8.31 ;
      RECT 31.78 0.57 31.95 1.08 ;
      RECT 31.78 2.39 31.95 3.86 ;
      RECT 31.78 5.02 31.95 6.49 ;
      RECT 31.78 7.8 31.95 8.31 ;
      RECT 30.42 0.575 30.59 3.865 ;
      RECT 30.42 5.015 30.59 8.305 ;
      RECT 29.99 0.575 30.16 1.085 ;
      RECT 29.99 1.655 30.16 3.865 ;
      RECT 29.99 5.015 30.16 7.225 ;
      RECT 29.99 7.795 30.16 8.305 ;
      RECT 24.785 5.015 24.955 8.305 ;
      RECT 24.355 5.015 24.525 7.225 ;
      RECT 24.355 7.795 24.525 8.305 ;
      RECT 17.51 7.8 17.68 8.31 ;
      RECT 16.52 0.57 16.69 1.08 ;
      RECT 16.52 2.39 16.69 3.86 ;
      RECT 16.52 5.02 16.69 6.49 ;
      RECT 16.52 7.8 16.69 8.31 ;
      RECT 15.16 0.575 15.33 3.865 ;
      RECT 15.16 5.015 15.33 8.305 ;
      RECT 14.73 0.575 14.9 1.085 ;
      RECT 14.73 1.655 14.9 3.865 ;
      RECT 14.73 5.015 14.9 7.225 ;
      RECT 14.73 7.795 14.9 8.305 ;
      RECT 9.525 5.015 9.695 8.305 ;
      RECT 9.095 5.015 9.265 7.225 ;
      RECT 9.095 7.795 9.265 8.305 ;
      RECT 1.6 5.015 1.77 7.225 ;
      RECT 1.6 7.795 1.77 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r2

END LIBRARY
