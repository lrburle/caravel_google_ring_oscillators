magic
tech sky130A
magscale 1 2
timestamp 1704982549
<< viali >>
rect 301933 492201 301967 492235
rect 294256 472005 294290 472039
rect 296038 471189 296072 471223
rect 299623 471189 299657 471223
rect 303208 471189 303242 471223
rect 306793 471189 306827 471223
rect 310378 471189 310412 471223
rect 302378 471053 302412 471087
rect 295769 449701 295803 449735
rect 299086 449701 299120 449735
rect 302403 449701 302437 449735
rect 299341 429165 299375 429199
rect 293763 408969 293797 409003
rect 297028 408833 297062 408867
rect 298981 408221 299015 408255
rect 305511 408153 305545 408187
rect 294209 388025 294243 388059
rect 309057 388025 309091 388059
rect 303586 387209 303620 387243
rect 295503 366197 295537 366231
rect 307711 366197 307745 366231
rect 293545 346001 293579 346035
rect 299649 346001 299683 346035
rect 295502 345185 295536 345219
rect 307710 345185 307744 345219
rect 301930 323697 301964 323731
rect 310406 303161 310440 303195
rect 292728 262021 292762 262055
rect 299339 261205 299373 261239
rect 309671 261205 309705 261239
rect 293762 241009 293796 241043
rect 297027 240805 297061 240839
rect 298980 240193 299014 240227
rect 305510 240193 305544 240227
rect 297921 219793 297955 219827
rect 303586 218705 303620 218739
rect 295502 198169 295536 198203
rect 307710 198169 307744 198203
rect 296597 178177 296631 178211
rect 295502 177361 295536 177395
rect 307710 177361 307744 177395
<< metal1 >>
rect 301130 493348 301136 493400
rect 301188 493348 301194 493400
rect 301148 492844 301176 493348
rect 296996 492832 297048 492838
rect 289722 492668 289728 492720
rect 289780 492708 289786 492720
rect 292040 492708 292068 492806
rect 301103 492820 301176 492844
rect 301070 492816 301176 492820
rect 301070 492792 301131 492816
rect 304290 492792 304672 492820
rect 296996 492774 297048 492780
rect 289780 492680 292068 492708
rect 304644 492708 304672 492792
rect 308398 492708 308404 492720
rect 304644 492680 308404 492708
rect 289780 492668 289786 492680
rect 308398 492668 308404 492680
rect 308456 492668 308462 492720
rect 292482 492600 292488 492652
rect 292540 492640 292546 492652
rect 296990 492640 296996 492652
rect 292540 492612 296996 492640
rect 292540 492600 292546 492612
rect 296990 492600 296996 492612
rect 297048 492600 297054 492652
rect 301958 492241 301964 492244
rect 301921 492235 301964 492241
rect 301921 492201 301933 492235
rect 301921 492195 301964 492201
rect 301958 492192 301964 492195
rect 302016 492192 302022 492244
rect 309594 492232 309600 492244
rect 307588 492204 309600 492232
rect 307588 492184 307616 492204
rect 309594 492192 309600 492204
rect 309652 492192 309658 492244
rect 291930 492124 291936 492176
rect 291988 492164 291994 492176
rect 291988 492136 294814 492164
rect 307418 492156 307616 492184
rect 291988 492124 291994 492136
rect 295616 491825 295668 491831
rect 295616 491767 295668 491773
rect 298744 491825 298796 491831
rect 298744 491767 298796 491773
rect 305092 491825 305144 491831
rect 305092 491767 305144 491773
rect 308232 491484 308260 491799
rect 313918 491484 313924 491496
rect 308232 491456 313924 491484
rect 313918 491444 313924 491456
rect 313976 491444 313982 491496
rect 305086 488996 305092 489048
rect 305144 489036 305150 489048
rect 312722 489036 312728 489048
rect 305144 489008 312728 489036
rect 305144 488996 305150 489008
rect 312722 488996 312728 489008
rect 312780 488996 312786 489048
rect 301958 488656 301964 488708
rect 302016 488696 302022 488708
rect 312906 488696 312912 488708
rect 302016 488668 312912 488696
rect 302016 488656 302022 488668
rect 312906 488656 312912 488668
rect 312964 488656 312970 488708
rect 298738 488588 298744 488640
rect 298796 488628 298802 488640
rect 367738 488628 367744 488640
rect 298796 488600 367744 488628
rect 298796 488588 298802 488600
rect 367738 488588 367744 488600
rect 367796 488588 367802 488640
rect 295610 488520 295616 488572
rect 295668 488560 295674 488572
rect 404998 488560 405004 488572
rect 295668 488532 405004 488560
rect 295668 488520 295674 488532
rect 404998 488520 405004 488532
rect 405056 488520 405062 488572
rect 296622 473288 296628 473340
rect 296680 473328 296686 473340
rect 298370 473328 298376 473340
rect 296680 473300 298376 473328
rect 296680 473288 296686 473300
rect 298370 473288 298376 473300
rect 298428 473288 298434 473340
rect 298370 472404 298376 472456
rect 298428 472404 298434 472456
rect 302418 472404 302424 472456
rect 302476 472444 302482 472456
rect 302476 472416 303016 472444
rect 302476 472404 302482 472416
rect 298388 472184 298416 472404
rect 302988 472184 303016 472416
rect 298370 472132 298376 472184
rect 298428 472132 298434 472184
rect 302970 472132 302976 472184
rect 303028 472132 303034 472184
rect 291838 471996 291844 472048
rect 291896 472036 291902 472048
rect 294244 472039 294302 472045
rect 294244 472036 294256 472039
rect 291896 472008 294256 472036
rect 291896 471996 291902 472008
rect 294244 472005 294256 472008
rect 294290 472005 294302 472039
rect 294244 471999 294302 472005
rect 289722 471928 289728 471980
rect 289780 471968 289786 471980
rect 289780 471940 292068 471968
rect 289780 471928 289786 471940
rect 292040 471806 292068 471940
rect 298370 471780 298376 471832
rect 298428 471780 298434 471832
rect 310514 471288 310520 471300
rect 306116 471260 310520 471288
rect 295978 471180 295984 471232
rect 296036 471229 296042 471232
rect 296036 471223 296084 471229
rect 296036 471189 296038 471223
rect 296072 471189 296084 471223
rect 296036 471183 296084 471189
rect 296036 471180 296042 471183
rect 299566 471180 299572 471232
rect 299624 471229 299630 471232
rect 299624 471223 299669 471229
rect 299657 471189 299669 471223
rect 299624 471183 299669 471189
rect 299624 471180 299630 471183
rect 303154 471180 303160 471232
rect 303212 471229 303218 471232
rect 303212 471223 303254 471229
rect 303242 471189 303254 471223
rect 303212 471183 303254 471189
rect 306116 471184 306144 471260
rect 310514 471248 310520 471260
rect 310572 471248 310578 471300
rect 303212 471180 303218 471183
rect 306038 471156 306144 471184
rect 306742 471180 306748 471232
rect 306800 471229 306806 471232
rect 306800 471223 306839 471229
rect 306827 471189 306839 471223
rect 306800 471183 306839 471189
rect 310366 471223 310424 471229
rect 310366 471189 310378 471223
rect 310412 471220 310424 471223
rect 312538 471220 312544 471232
rect 310412 471192 312544 471220
rect 310412 471189 310424 471192
rect 310366 471183 310424 471189
rect 306800 471180 306806 471183
rect 312538 471180 312544 471192
rect 312596 471180 312602 471232
rect 302366 471087 302424 471093
rect 302366 471053 302378 471087
rect 302412 471053 302424 471087
rect 302366 471047 302424 471053
rect 302378 471016 302406 471047
rect 302970 471016 302976 471028
rect 302378 470988 302976 471016
rect 302142 470704 302148 470756
rect 302200 470744 302206 470756
rect 302436 470744 302464 470988
rect 302970 470976 302976 470988
rect 303028 470976 303034 471028
rect 302200 470716 302464 470744
rect 302200 470704 302206 470716
rect 306742 469140 306748 469192
rect 306800 469180 306806 469192
rect 306800 469152 311894 469180
rect 306800 469140 306806 469152
rect 311866 469112 311894 469152
rect 314102 469112 314108 469124
rect 311866 469084 314108 469112
rect 314102 469072 314108 469084
rect 314160 469072 314166 469124
rect 296070 468052 296076 468104
rect 296128 468092 296134 468104
rect 296128 468064 296714 468092
rect 296128 468052 296134 468064
rect 296686 468024 296714 468064
rect 338758 468024 338764 468036
rect 296686 467996 338764 468024
rect 338758 467984 338764 467996
rect 338816 467984 338822 468036
rect 303154 467916 303160 467968
rect 303212 467956 303218 467968
rect 363598 467956 363604 467968
rect 303212 467928 363604 467956
rect 303212 467916 303218 467928
rect 363598 467916 363604 467928
rect 363656 467916 363662 467968
rect 299658 467848 299664 467900
rect 299716 467888 299722 467900
rect 388438 467888 388444 467900
rect 299716 467860 388444 467888
rect 299716 467848 299722 467860
rect 388438 467848 388444 467860
rect 388496 467848 388502 467900
rect 338758 451868 338764 451920
rect 338816 451908 338822 451920
rect 515398 451908 515404 451920
rect 338816 451880 515404 451908
rect 338816 451868 338822 451880
rect 515398 451868 515404 451880
rect 515456 451868 515462 451920
rect 289722 450780 289728 450832
rect 289780 450820 289786 450832
rect 289780 450792 292054 450820
rect 289780 450780 289786 450792
rect 309060 449936 309088 450095
rect 314010 449936 314016 449948
rect 309060 449908 314016 449936
rect 314010 449896 314016 449908
rect 314068 449896 314074 449948
rect 305736 449825 305788 449831
rect 305736 449767 305788 449773
rect 295794 449741 295800 449744
rect 295757 449735 295800 449741
rect 295757 449701 295769 449735
rect 295757 449695 295800 449701
rect 295794 449692 295800 449695
rect 295852 449692 295858 449744
rect 299106 449741 299112 449744
rect 299074 449735 299112 449741
rect 299074 449701 299086 449735
rect 299074 449695 299112 449701
rect 299106 449692 299112 449695
rect 299164 449692 299170 449744
rect 302418 449741 302424 449744
rect 302391 449735 302424 449741
rect 302391 449701 302403 449735
rect 302391 449695 302424 449701
rect 302418 449692 302424 449695
rect 302476 449692 302482 449744
rect 305730 447652 305736 447704
rect 305788 447692 305794 447704
rect 314194 447692 314200 447704
rect 305788 447664 314200 447692
rect 305788 447652 305794 447664
rect 314194 447652 314200 447664
rect 314252 447652 314258 447704
rect 295794 447244 295800 447296
rect 295852 447284 295858 447296
rect 295852 447256 296714 447284
rect 295852 447244 295858 447256
rect 296686 447148 296714 447256
rect 299106 447244 299112 447296
rect 299164 447244 299170 447296
rect 302418 447244 302424 447296
rect 302476 447284 302482 447296
rect 370590 447284 370596 447296
rect 302476 447256 370596 447284
rect 302476 447244 302482 447256
rect 370590 447244 370596 447256
rect 370648 447244 370654 447296
rect 299124 447216 299152 447244
rect 406378 447216 406384 447228
rect 299124 447188 406384 447216
rect 406378 447176 406384 447188
rect 406436 447176 406442 447228
rect 443638 447148 443644 447160
rect 296686 447120 443644 447148
rect 443638 447108 443644 447120
rect 443696 447108 443702 447160
rect 296070 430040 296076 430092
rect 296128 430040 296134 430092
rect 292764 429832 292816 429838
rect 289722 429768 289728 429820
rect 289780 429808 289786 429820
rect 289780 429780 292068 429808
rect 296088 429820 296116 430040
rect 296088 429792 296194 429820
rect 289780 429768 289786 429780
rect 292764 429774 292816 429780
rect 299290 429156 299296 429208
rect 299348 429205 299354 429208
rect 299348 429199 299387 429205
rect 299375 429165 299387 429199
rect 299348 429159 299387 429165
rect 299348 429156 299354 429159
rect 308876 428924 308904 429170
rect 309134 428924 309140 428936
rect 308876 428896 309140 428924
rect 309134 428884 309140 428896
rect 309192 428884 309198 428936
rect 302792 428825 302844 428831
rect 295904 428788 295932 428799
rect 296530 428788 296536 428800
rect 295904 428760 296536 428788
rect 296530 428748 296536 428760
rect 296588 428748 296594 428800
rect 302792 428767 302844 428773
rect 306196 428825 306248 428831
rect 309718 428788 310008 428813
rect 312814 428788 312820 428800
rect 309718 428785 312820 428788
rect 306196 428767 306248 428773
rect 309980 428760 312820 428785
rect 312814 428748 312820 428760
rect 312872 428748 312878 428800
rect 306190 425552 306196 425604
rect 306248 425592 306254 425604
rect 314378 425592 314384 425604
rect 306248 425564 314384 425592
rect 306248 425552 306254 425564
rect 314378 425552 314384 425564
rect 314436 425552 314442 425604
rect 299290 425144 299296 425196
rect 299348 425144 299354 425196
rect 302786 425144 302792 425196
rect 302844 425184 302850 425196
rect 391198 425184 391204 425196
rect 302844 425156 391204 425184
rect 302844 425144 302850 425156
rect 391198 425144 391204 425156
rect 391256 425144 391262 425196
rect 299308 425116 299336 425144
rect 427078 425116 427084 425128
rect 299308 425088 427084 425116
rect 427078 425076 427084 425088
rect 427136 425076 427142 425128
rect 404998 422220 405004 422272
rect 405056 422260 405062 422272
rect 514754 422260 514760 422272
rect 405056 422232 514760 422260
rect 405056 422220 405062 422232
rect 514754 422220 514760 422232
rect 514812 422220 514818 422272
rect 524322 421404 524328 421456
rect 524380 421444 524386 421456
rect 527174 421444 527180 421456
rect 524380 421416 527180 421444
rect 524380 421404 524386 421416
rect 527174 421404 527180 421416
rect 527232 421404 527238 421456
rect 517422 421336 517428 421388
rect 517480 421376 517486 421388
rect 518986 421376 518992 421388
rect 517480 421348 518992 421376
rect 517480 421336 517486 421348
rect 518986 421336 518992 421348
rect 519044 421336 519050 421388
rect 526990 421336 526996 421388
rect 527048 421376 527054 421388
rect 529198 421376 529204 421388
rect 527048 421348 529204 421376
rect 527048 421336 527054 421348
rect 529198 421336 529204 421348
rect 529256 421336 529262 421388
rect 443638 419432 443644 419484
rect 443696 419472 443702 419484
rect 514754 419472 514760 419484
rect 443696 419444 514760 419472
rect 443696 419432 443702 419444
rect 514754 419432 514760 419444
rect 514812 419432 514818 419484
rect 296530 418072 296536 418124
rect 296588 418112 296594 418124
rect 514754 418112 514760 418124
rect 296588 418084 514760 418112
rect 296588 418072 296594 418084
rect 514754 418072 514760 418084
rect 514812 418072 514818 418124
rect 291838 409028 291844 409080
rect 291896 409068 291902 409080
rect 291896 409040 293816 409068
rect 291896 409028 291902 409040
rect 293788 409009 293816 409040
rect 293751 409003 293816 409009
rect 293751 408969 293763 409003
rect 293797 408972 293816 409003
rect 293797 408969 293809 408972
rect 293751 408963 293809 408969
rect 297016 408867 297074 408873
rect 297016 408864 297028 408867
rect 296686 408836 297028 408864
rect 292040 408796 292068 408806
rect 289740 408768 292068 408796
rect 289740 408740 289768 408768
rect 289722 408688 289728 408740
rect 289780 408688 289786 408740
rect 291930 408688 291936 408740
rect 291988 408728 291994 408740
rect 296686 408728 296714 408836
rect 297016 408833 297028 408836
rect 297062 408833 297074 408867
rect 297016 408827 297074 408833
rect 291988 408700 296714 408728
rect 291988 408688 291994 408700
rect 298922 408212 298928 408264
rect 298980 408261 298986 408264
rect 298980 408255 299027 408261
rect 298980 408221 298981 408255
rect 299015 408221 299027 408255
rect 298980 408215 299027 408221
rect 298980 408212 298986 408215
rect 305499 408187 305557 408193
rect 305499 408153 305511 408187
rect 305545 408184 305557 408187
rect 305638 408184 305644 408196
rect 305545 408156 305644 408184
rect 305545 408153 305557 408156
rect 305499 408147 305557 408153
rect 305638 408144 305644 408156
rect 305696 408144 305702 408196
rect 309042 408184 309048 408196
rect 307970 408156 309048 408184
rect 309042 408144 309048 408156
rect 309100 408144 309106 408196
rect 295708 407825 295760 407831
rect 295708 407767 295760 407773
rect 302240 407825 302292 407831
rect 302240 407767 302292 407773
rect 308784 407776 308812 407799
rect 311434 407776 311440 407788
rect 308784 407748 311440 407776
rect 311434 407736 311440 407748
rect 311492 407736 311498 407788
rect 312998 407124 313004 407176
rect 313056 407164 313062 407176
rect 514754 407164 514760 407176
rect 313056 407136 514760 407164
rect 313056 407124 313062 407136
rect 514754 407124 514760 407136
rect 514812 407124 514818 407176
rect 311526 405696 311532 405748
rect 311584 405736 311590 405748
rect 514754 405736 514760 405748
rect 311584 405708 514760 405736
rect 311584 405696 311590 405708
rect 514754 405696 514760 405708
rect 514812 405696 514818 405748
rect 295702 405628 295708 405680
rect 295760 405668 295766 405680
rect 515398 405668 515404 405680
rect 295760 405640 515404 405668
rect 295760 405628 295766 405640
rect 515398 405628 515404 405640
rect 515456 405628 515462 405680
rect 302234 405560 302240 405612
rect 302292 405560 302298 405612
rect 305638 405560 305644 405612
rect 305696 405600 305702 405612
rect 314470 405600 314476 405612
rect 305696 405572 314476 405600
rect 305696 405560 305702 405572
rect 314470 405560 314476 405572
rect 314528 405560 314534 405612
rect 302252 405532 302280 405560
rect 313182 405532 313188 405544
rect 302252 405504 313188 405532
rect 313182 405492 313188 405504
rect 313240 405492 313246 405544
rect 298922 404608 298928 404660
rect 298980 404608 298986 404660
rect 298940 404444 298968 404608
rect 446398 404444 446404 404456
rect 298940 404416 446404 404444
rect 446398 404404 446404 404416
rect 446456 404404 446462 404456
rect 311250 404336 311256 404388
rect 311308 404376 311314 404388
rect 514754 404376 514760 404388
rect 311308 404348 514760 404376
rect 311308 404336 311314 404348
rect 514754 404336 514760 404348
rect 514812 404336 514818 404388
rect 311158 402976 311164 403028
rect 311216 403016 311222 403028
rect 514754 403016 514760 403028
rect 311216 402988 514760 403016
rect 311216 402976 311222 402988
rect 514754 402976 514760 402988
rect 514812 402976 514818 403028
rect 312630 401616 312636 401668
rect 312688 401656 312694 401668
rect 514754 401656 514760 401668
rect 312688 401628 514760 401656
rect 312688 401616 312694 401628
rect 514754 401616 514760 401628
rect 514812 401616 514818 401668
rect 289722 388016 289728 388068
rect 289780 388016 289786 388068
rect 291838 388016 291844 388068
rect 291896 388056 291902 388068
rect 294197 388059 294255 388065
rect 294197 388056 294209 388059
rect 291896 388028 294209 388056
rect 291896 388016 291902 388028
rect 294197 388025 294209 388028
rect 294243 388025 294255 388059
rect 294197 388019 294255 388025
rect 309042 388016 309048 388068
rect 309100 388016 309106 388068
rect 289740 387988 289768 388016
rect 289740 387960 292068 387988
rect 292040 387806 292068 387960
rect 302234 387780 302240 387832
rect 302292 387780 302298 387832
rect 306498 387792 306788 387820
rect 306760 387716 306788 387792
rect 311894 387716 311900 387728
rect 306760 387688 311900 387716
rect 311894 387676 311900 387688
rect 311952 387676 311958 387728
rect 303614 387249 303620 387252
rect 303574 387243 303620 387249
rect 303574 387209 303586 387243
rect 303574 387203 303620 387209
rect 303614 387200 303620 387203
rect 303672 387200 303678 387252
rect 314286 386832 314292 386844
rect 296168 386825 296220 386831
rect 296168 386767 296220 386773
rect 299848 386825 299900 386831
rect 299848 386767 299900 386773
rect 307300 386825 307352 386831
rect 310992 386804 314292 386832
rect 310992 386799 311020 386804
rect 314286 386792 314292 386804
rect 314344 386792 314350 386844
rect 307300 386767 307352 386773
rect 296162 384956 296168 385008
rect 296220 384996 296226 385008
rect 515858 384996 515864 385008
rect 296220 384968 515864 384996
rect 296220 384956 296226 384968
rect 515858 384956 515864 384968
rect 515916 384956 515922 385008
rect 299842 384888 299848 384940
rect 299900 384928 299906 384940
rect 300762 384928 300768 384940
rect 299900 384900 300768 384928
rect 299900 384888 299906 384900
rect 300762 384888 300768 384900
rect 300820 384888 300826 384940
rect 303614 384888 303620 384940
rect 303672 384928 303678 384940
rect 308398 384928 308404 384940
rect 303672 384900 308404 384928
rect 303672 384888 303678 384900
rect 308398 384888 308404 384900
rect 308456 384888 308462 384940
rect 307294 384004 307300 384056
rect 307352 384044 307358 384056
rect 307352 384016 311894 384044
rect 307352 384004 307358 384016
rect 311866 383908 311894 384016
rect 311866 383880 316034 383908
rect 316006 383704 316034 383880
rect 393958 383704 393964 383716
rect 316006 383676 393964 383704
rect 393958 383664 393964 383676
rect 394016 383664 394022 383716
rect 367738 382168 367744 382220
rect 367796 382208 367802 382220
rect 514754 382208 514760 382220
rect 367796 382180 514760 382208
rect 367796 382168 367802 382180
rect 514754 382168 514760 382180
rect 514812 382168 514818 382220
rect 388438 380808 388444 380860
rect 388496 380848 388502 380860
rect 514754 380848 514760 380860
rect 388496 380820 514760 380848
rect 388496 380808 388502 380820
rect 514754 380808 514760 380820
rect 514812 380808 514818 380860
rect 406378 379448 406384 379500
rect 406436 379488 406442 379500
rect 514754 379488 514760 379500
rect 406436 379460 514760 379488
rect 406436 379448 406442 379460
rect 514754 379448 514760 379460
rect 514812 379448 514818 379500
rect 427078 378088 427084 378140
rect 427136 378128 427142 378140
rect 514754 378128 514760 378140
rect 427136 378100 514760 378128
rect 427136 378088 427142 378100
rect 514754 378088 514760 378100
rect 514812 378088 514818 378140
rect 446398 376660 446404 376712
rect 446456 376700 446462 376712
rect 514754 376700 514760 376712
rect 446456 376672 514760 376700
rect 446456 376660 446462 376672
rect 514754 376660 514760 376672
rect 514812 376660 514818 376712
rect 300762 375300 300768 375352
rect 300820 375340 300826 375352
rect 514754 375340 514760 375352
rect 300820 375312 514760 375340
rect 300820 375300 300826 375312
rect 514754 375300 514760 375312
rect 514812 375300 514818 375352
rect 373258 367072 373264 367124
rect 373316 367112 373322 367124
rect 514754 367112 514760 367124
rect 373316 367084 514760 367112
rect 373316 367072 373322 367084
rect 514754 367072 514760 367084
rect 514812 367072 514818 367124
rect 289722 367004 289728 367056
rect 289780 367044 289786 367056
rect 289780 367016 292068 367044
rect 289780 367004 289786 367016
rect 292040 366806 292068 367016
rect 307662 366840 307668 366852
rect 294046 366780 294052 366832
rect 294104 366780 294110 366832
rect 300210 366780 300216 366832
rect 300268 366780 300274 366832
rect 307220 366820 307668 366840
rect 306958 366812 307668 366820
rect 306958 366792 307248 366812
rect 307662 366800 307668 366812
rect 307720 366840 307726 366852
rect 308030 366840 308036 366852
rect 307720 366812 308036 366840
rect 307720 366800 307726 366812
rect 308030 366800 308036 366812
rect 308088 366800 308094 366852
rect 295518 366237 295524 366240
rect 295491 366231 295524 366237
rect 295491 366197 295503 366231
rect 295491 366191 295524 366197
rect 295518 366188 295524 366191
rect 295576 366188 295582 366240
rect 307699 366231 307757 366237
rect 307699 366197 307711 366231
rect 307745 366228 307757 366231
rect 307745 366200 316034 366228
rect 307745 366197 307757 366200
rect 307699 366191 307757 366197
rect 298560 365825 298612 365831
rect 298560 365767 298612 365773
rect 301596 365825 301648 365831
rect 301596 365767 301648 365773
rect 304632 365825 304684 365831
rect 316006 365820 316034 366200
rect 370498 365820 370504 365832
rect 316006 365792 370504 365820
rect 370498 365780 370504 365792
rect 370556 365780 370562 365832
rect 304632 365767 304684 365773
rect 313090 365712 313096 365764
rect 313148 365752 313154 365764
rect 514754 365752 514760 365764
rect 313148 365724 514760 365752
rect 313148 365712 313154 365724
rect 514754 365712 514760 365724
rect 514812 365712 514818 365764
rect 359458 364352 359464 364404
rect 359516 364392 359522 364404
rect 514754 364392 514760 364404
rect 359516 364364 514760 364392
rect 359516 364352 359522 364364
rect 514754 364352 514760 364364
rect 514812 364352 514818 364404
rect 295518 364284 295524 364336
rect 295576 364324 295582 364336
rect 515490 364324 515496 364336
rect 295576 364296 515496 364324
rect 295576 364284 295582 364296
rect 515490 364284 515496 364296
rect 515548 364284 515554 364336
rect 298554 364216 298560 364268
rect 298612 364256 298618 364268
rect 515306 364256 515312 364268
rect 298612 364228 515312 364256
rect 298612 364216 298618 364228
rect 515306 364216 515312 364228
rect 515364 364216 515370 364268
rect 301590 364148 301596 364200
rect 301648 364188 301654 364200
rect 308490 364188 308496 364200
rect 301648 364160 308496 364188
rect 301648 364148 301654 364160
rect 308490 364148 308496 364160
rect 308548 364148 308554 364200
rect 304626 363332 304632 363384
rect 304684 363372 304690 363384
rect 314562 363372 314568 363384
rect 304684 363344 314568 363372
rect 304684 363332 304690 363344
rect 314562 363332 314568 363344
rect 314620 363332 314626 363384
rect 311618 362924 311624 362976
rect 311676 362964 311682 362976
rect 514754 362964 514760 362976
rect 311676 362936 514760 362964
rect 311676 362924 311682 362936
rect 514754 362924 514760 362936
rect 514812 362924 514818 362976
rect 311342 361564 311348 361616
rect 311400 361604 311406 361616
rect 514754 361604 514760 361616
rect 311400 361576 514760 361604
rect 311400 361564 311406 361576
rect 514754 361564 514760 361576
rect 514812 361564 514818 361616
rect 299566 346400 299572 346452
rect 299624 346400 299630 346452
rect 299584 346168 299612 346400
rect 299584 346140 299704 346168
rect 291746 346060 291752 346112
rect 291804 346100 291810 346112
rect 291804 346072 293540 346100
rect 291804 346060 291810 346072
rect 289722 345992 289728 346044
rect 289780 346032 289786 346044
rect 293512 346041 293540 346072
rect 293512 346035 293591 346041
rect 289780 346004 292068 346032
rect 293512 346004 293545 346035
rect 289780 345992 289786 346004
rect 292040 345806 292068 346004
rect 293533 346001 293545 346004
rect 293579 346032 293591 346035
rect 294414 346032 294420 346044
rect 293579 346004 294420 346032
rect 293579 346001 293591 346004
rect 293533 345995 293591 346001
rect 294414 345992 294420 346004
rect 294472 345992 294478 346044
rect 299676 346041 299704 346140
rect 299637 346035 299704 346041
rect 299637 346001 299649 346035
rect 299683 346004 299704 346035
rect 299683 346001 299695 346004
rect 299637 345995 299695 346001
rect 307846 345828 307852 345840
rect 307036 345820 307852 345828
rect 306958 345800 307852 345820
rect 306958 345792 307064 345800
rect 307846 345788 307852 345800
rect 307904 345788 307910 345840
rect 313182 345652 313188 345704
rect 313240 345692 313246 345704
rect 515306 345692 515312 345704
rect 313240 345664 515312 345692
rect 313240 345652 313246 345664
rect 515306 345652 515312 345664
rect 515364 345652 515370 345704
rect 295518 345225 295524 345228
rect 295490 345219 295524 345225
rect 295490 345185 295502 345219
rect 295490 345179 295524 345185
rect 295518 345176 295524 345179
rect 295576 345176 295582 345228
rect 307698 345219 307756 345225
rect 307698 345216 307710 345219
rect 307680 345185 307710 345216
rect 307744 345185 307756 345219
rect 307680 345179 307756 345185
rect 307680 345080 307708 345179
rect 307680 345052 307800 345080
rect 307772 344876 307800 345052
rect 313182 344876 313188 344888
rect 307772 344848 313188 344876
rect 313182 344836 313188 344848
rect 313240 344836 313246 344888
rect 298560 344825 298612 344831
rect 304632 344825 304684 344831
rect 302142 344808 302148 344820
rect 301622 344780 302148 344808
rect 298560 344767 298612 344773
rect 302142 344768 302148 344780
rect 302200 344768 302206 344820
rect 304632 344767 304684 344773
rect 295518 342184 295524 342236
rect 295576 342224 295582 342236
rect 515766 342224 515772 342236
rect 295576 342196 515772 342224
rect 295576 342184 295582 342196
rect 515766 342184 515772 342196
rect 515824 342184 515830 342236
rect 298554 342116 298560 342168
rect 298612 342156 298618 342168
rect 516042 342156 516048 342168
rect 298612 342128 516048 342156
rect 298612 342116 298618 342128
rect 516042 342116 516048 342128
rect 516100 342116 516106 342168
rect 312906 342048 312912 342100
rect 312964 342088 312970 342100
rect 514754 342088 514760 342100
rect 312964 342060 514760 342088
rect 312964 342048 312970 342060
rect 514754 342048 514760 342060
rect 514812 342048 514818 342100
rect 304626 341300 304632 341352
rect 304684 341340 304690 341352
rect 304684 341312 306374 341340
rect 304684 341300 304690 341312
rect 306346 341272 306374 341312
rect 309778 341272 309784 341284
rect 306346 341244 309784 341272
rect 309778 341232 309784 341244
rect 309836 341232 309842 341284
rect 363598 340824 363604 340876
rect 363656 340864 363662 340876
rect 514754 340864 514760 340876
rect 363656 340836 514760 340864
rect 363656 340824 363662 340836
rect 514754 340824 514760 340836
rect 514812 340824 514818 340876
rect 370590 339396 370596 339448
rect 370648 339436 370654 339448
rect 514754 339436 514760 339448
rect 370648 339408 514760 339436
rect 370648 339396 370654 339408
rect 514754 339396 514760 339408
rect 514812 339396 514818 339448
rect 391198 338036 391204 338088
rect 391256 338076 391262 338088
rect 514754 338076 514760 338088
rect 391256 338048 514760 338076
rect 391256 338036 391262 338048
rect 514754 338036 514760 338048
rect 514812 338036 514818 338088
rect 308398 335248 308404 335300
rect 308456 335288 308462 335300
rect 514754 335288 514760 335300
rect 308456 335260 514760 335288
rect 308456 335248 308462 335260
rect 514754 335248 514760 335260
rect 514812 335248 514818 335300
rect 308490 333888 308496 333940
rect 308548 333928 308554 333940
rect 514754 333928 514760 333940
rect 308548 333900 514760 333928
rect 308548 333888 308554 333900
rect 514754 333888 514760 333900
rect 514812 333888 514818 333940
rect 302142 332528 302148 332580
rect 302200 332568 302206 332580
rect 514754 332568 514760 332580
rect 302200 332540 514760 332568
rect 302200 332528 302206 332540
rect 514754 332528 514760 332540
rect 514812 332528 514818 332580
rect 363690 327088 363696 327140
rect 363748 327128 363754 327140
rect 514754 327128 514760 327140
rect 363748 327100 514760 327128
rect 363748 327088 363754 327100
rect 514754 327088 514760 327100
rect 514812 327088 514818 327140
rect 363598 325660 363604 325712
rect 363656 325700 363662 325712
rect 514754 325700 514760 325712
rect 363656 325672 514760 325700
rect 363656 325660 363662 325672
rect 514754 325660 514760 325672
rect 514812 325660 514818 325712
rect 294782 325388 294788 325440
rect 294840 325388 294846 325440
rect 307846 325388 307852 325440
rect 307904 325428 307910 325440
rect 308490 325428 308496 325440
rect 307904 325400 308496 325428
rect 307904 325388 307910 325400
rect 308490 325388 308496 325400
rect 308548 325388 308554 325440
rect 294800 325236 294828 325388
rect 294782 325184 294788 325236
rect 294840 325184 294846 325236
rect 308398 324952 308404 324964
rect 301516 324924 308404 324952
rect 296996 324832 297048 324838
rect 289722 324776 289728 324828
rect 289780 324816 289786 324828
rect 289780 324788 292068 324816
rect 289780 324776 289786 324788
rect 301516 324820 301544 324924
rect 308398 324912 308404 324924
rect 308456 324912 308462 324964
rect 301162 324792 301544 324820
rect 308582 324816 308588 324828
rect 307418 324788 308588 324816
rect 296996 324774 297048 324780
rect 308582 324776 308588 324788
rect 308640 324776 308646 324828
rect 291838 324640 291844 324692
rect 291896 324680 291902 324692
rect 296990 324680 296996 324692
rect 291896 324652 296996 324680
rect 291896 324640 291902 324652
rect 296990 324640 296996 324652
rect 297048 324640 297054 324692
rect 377398 324300 377404 324352
rect 377456 324340 377462 324352
rect 514754 324340 514760 324352
rect 377456 324312 514760 324340
rect 377456 324300 377462 324312
rect 514754 324300 514760 324312
rect 514812 324300 514818 324352
rect 308490 324272 308496 324284
rect 304276 324244 308496 324272
rect 294788 324196 294840 324202
rect 304276 324190 304304 324244
rect 308490 324232 308496 324244
rect 308548 324232 308554 324284
rect 294788 324138 294840 324144
rect 292390 323892 292396 323944
rect 292448 323932 292454 323944
rect 294800 323932 294828 324138
rect 292448 323904 294828 323932
rect 292448 323892 292454 323904
rect 295616 323825 295668 323831
rect 295616 323767 295668 323773
rect 298744 323825 298796 323831
rect 298744 323767 298796 323773
rect 305092 323825 305144 323831
rect 305092 323767 305144 323773
rect 301958 323737 301964 323740
rect 301918 323731 301964 323737
rect 301918 323697 301930 323731
rect 301918 323691 301964 323697
rect 301958 323688 301964 323691
rect 302016 323688 302022 323740
rect 308232 323524 308260 323799
rect 311710 323524 311716 323536
rect 308232 323496 311716 323524
rect 311710 323484 311716 323496
rect 311768 323484 311774 323536
rect 364978 322940 364984 322992
rect 365036 322980 365042 322992
rect 514754 322980 514760 322992
rect 365036 322952 514760 322980
rect 365036 322940 365042 322952
rect 514754 322940 514760 322952
rect 514812 322940 514818 322992
rect 362218 321580 362224 321632
rect 362276 321620 362282 321632
rect 514754 321620 514760 321632
rect 362276 321592 514760 321620
rect 362276 321580 362282 321592
rect 514754 321580 514760 321592
rect 514812 321580 514818 321632
rect 295610 321512 295616 321564
rect 295668 321552 295674 321564
rect 515674 321552 515680 321564
rect 295668 321524 515680 321552
rect 295668 321512 295674 321524
rect 515674 321512 515680 321524
rect 515732 321512 515738 321564
rect 298738 321444 298744 321496
rect 298796 321484 298802 321496
rect 515950 321484 515956 321496
rect 298796 321456 515956 321484
rect 298796 321444 298802 321456
rect 515950 321444 515956 321456
rect 516008 321444 516014 321496
rect 301958 321376 301964 321428
rect 302016 321416 302022 321428
rect 516042 321416 516048 321428
rect 302016 321388 516048 321416
rect 302016 321376 302022 321388
rect 516042 321376 516048 321388
rect 516100 321376 516106 321428
rect 345658 320152 345664 320204
rect 345716 320192 345722 320204
rect 514754 320192 514760 320204
rect 345716 320164 514760 320192
rect 345716 320152 345722 320164
rect 514754 320152 514760 320164
rect 514812 320152 514818 320204
rect 305086 318044 305092 318096
rect 305144 318084 305150 318096
rect 366358 318084 366364 318096
rect 305144 318056 366364 318084
rect 305144 318044 305150 318056
rect 366358 318044 366364 318056
rect 366416 318044 366422 318096
rect 294966 304376 294972 304428
rect 295024 304376 295030 304428
rect 298462 304376 298468 304428
rect 298520 304376 298526 304428
rect 302418 304376 302424 304428
rect 302476 304376 302482 304428
rect 306006 304376 306012 304428
rect 306064 304376 306070 304428
rect 309594 304376 309600 304428
rect 309652 304376 309658 304428
rect 309778 304376 309784 304428
rect 309836 304416 309842 304428
rect 309836 304388 316034 304416
rect 309836 304376 309842 304388
rect 294984 304224 295012 304376
rect 298480 304224 298508 304376
rect 302436 304224 302464 304376
rect 306024 304224 306052 304376
rect 309612 304224 309640 304376
rect 316006 304280 316034 304388
rect 515674 304280 515680 304292
rect 316006 304252 515680 304280
rect 515674 304240 515680 304252
rect 515732 304240 515738 304292
rect 294966 304172 294972 304224
rect 295024 304172 295030 304224
rect 298462 304172 298468 304224
rect 298520 304172 298526 304224
rect 302418 304172 302424 304224
rect 302476 304172 302482 304224
rect 306006 304172 306012 304224
rect 306064 304172 306070 304224
rect 309594 304172 309600 304224
rect 309652 304172 309658 304224
rect 289722 303764 289728 303816
rect 289780 303804 289786 303816
rect 291856 303804 292146 303820
rect 289780 303792 292146 303804
rect 289780 303776 291884 303792
rect 289780 303764 289786 303776
rect 310394 303195 310452 303201
rect 310394 303161 310406 303195
rect 310440 303192 310452 303195
rect 312906 303192 312912 303204
rect 310440 303164 312912 303192
rect 310440 303161 310452 303164
rect 310394 303155 310452 303161
rect 312906 303152 312912 303164
rect 312964 303152 312970 303204
rect 314102 303084 314108 303136
rect 314160 303124 314166 303136
rect 515030 303124 515036 303136
rect 314160 303096 515036 303124
rect 314160 303084 314166 303096
rect 515030 303084 515036 303096
rect 515088 303084 515094 303136
rect 314562 303016 314568 303068
rect 314620 303056 314626 303068
rect 515950 303056 515956 303068
rect 314620 303028 515956 303056
rect 314620 303016 314626 303028
rect 515950 303016 515956 303028
rect 516008 303016 516014 303068
rect 314194 302948 314200 303000
rect 314252 302988 314258 303000
rect 514938 302988 514944 303000
rect 314252 302960 514944 302988
rect 314252 302948 314258 302960
rect 514938 302948 514944 302960
rect 514996 302948 515002 303000
rect 312722 302880 312728 302932
rect 312780 302920 312786 302932
rect 514754 302920 514760 302932
rect 312780 302892 514760 302920
rect 312780 302880 312786 302892
rect 514754 302880 514760 302892
rect 514812 302880 514818 302932
rect 296076 302825 296128 302831
rect 296076 302767 296128 302773
rect 299664 302825 299716 302831
rect 306840 302825 306892 302831
rect 299664 302767 299716 302773
rect 303264 302172 303292 302799
rect 306840 302767 306892 302773
rect 515766 302172 515772 302184
rect 303264 302144 515772 302172
rect 515766 302132 515772 302144
rect 515824 302132 515830 302184
rect 517422 301792 517428 301844
rect 517480 301832 517486 301844
rect 518894 301832 518900 301844
rect 517480 301804 518900 301832
rect 517480 301792 517486 301804
rect 518894 301792 518900 301804
rect 518952 301792 518958 301844
rect 296070 300772 296076 300824
rect 296128 300812 296134 300824
rect 515582 300812 515588 300824
rect 296128 300784 515588 300812
rect 296128 300772 296134 300784
rect 515582 300772 515588 300784
rect 515640 300772 515646 300824
rect 299658 300704 299664 300756
rect 299716 300744 299722 300756
rect 515858 300744 515864 300756
rect 299716 300716 515864 300744
rect 299716 300704 299722 300716
rect 515858 300704 515864 300716
rect 515916 300704 515922 300756
rect 306834 299752 306840 299804
rect 306892 299792 306898 299804
rect 307662 299792 307668 299804
rect 306892 299764 307668 299792
rect 306892 299752 306898 299764
rect 307662 299752 307668 299764
rect 307720 299752 307726 299804
rect 314378 298052 314384 298104
rect 314436 298092 314442 298104
rect 514754 298092 514760 298104
rect 314436 298064 514760 298092
rect 314436 298052 314442 298064
rect 514754 298052 514760 298064
rect 514812 298052 514818 298104
rect 314470 296624 314476 296676
rect 314528 296664 314534 296676
rect 514754 296664 514760 296676
rect 314528 296636 514760 296664
rect 314528 296624 314534 296636
rect 514754 296624 514760 296636
rect 514812 296624 514818 296676
rect 393958 295264 393964 295316
rect 394016 295304 394022 295316
rect 514754 295304 514760 295316
rect 394016 295276 514760 295304
rect 394016 295264 394022 295276
rect 514754 295264 514760 295276
rect 514812 295264 514818 295316
rect 366358 291116 366364 291168
rect 366416 291156 366422 291168
rect 514754 291156 514760 291168
rect 366416 291128 514760 291156
rect 366416 291116 366422 291128
rect 514754 291116 514760 291128
rect 514812 291116 514818 291168
rect 307662 289756 307668 289808
rect 307720 289796 307726 289808
rect 514754 289796 514760 289808
rect 307720 289768 514760 289796
rect 307720 289756 307726 289768
rect 514754 289756 514760 289768
rect 514812 289756 514818 289808
rect 366358 284316 366364 284368
rect 366416 284356 366422 284368
rect 514754 284356 514760 284368
rect 366416 284328 514760 284356
rect 366416 284316 366422 284328
rect 514754 284316 514760 284328
rect 514812 284316 514818 284368
rect 291838 282888 291844 282940
rect 291896 282928 291902 282940
rect 291896 282900 292344 282928
rect 291896 282888 291902 282900
rect 292316 282860 292344 282900
rect 292316 282832 292620 282860
rect 292592 282820 292620 282832
rect 291856 282792 292146 282820
rect 292592 282792 292790 282820
rect 296470 282792 296534 282820
rect 289740 282764 291884 282792
rect 296272 282764 296534 282792
rect 289740 282668 289768 282764
rect 289722 282616 289728 282668
rect 289780 282616 289786 282668
rect 291930 282616 291936 282668
rect 291988 282656 291994 282668
rect 296272 282656 296300 282764
rect 291988 282628 296300 282656
rect 291988 282616 291994 282628
rect 309134 282180 309140 282192
rect 308232 282152 309140 282180
rect 309134 282140 309140 282152
rect 309192 282140 309198 282192
rect 371878 281840 371884 281852
rect 295800 281825 295852 281831
rect 295800 281767 295852 281773
rect 299112 281825 299164 281831
rect 299112 281767 299164 281773
rect 302424 281825 302476 281831
rect 302424 281767 302476 281773
rect 305736 281825 305788 281831
rect 309060 281812 371884 281840
rect 309060 281799 309088 281812
rect 371878 281800 371884 281812
rect 371936 281800 371942 281852
rect 305736 281767 305788 281773
rect 295794 280100 295800 280152
rect 295852 280140 295858 280152
rect 295852 280112 296714 280140
rect 295852 280100 295858 280112
rect 296686 279936 296714 280112
rect 299106 280100 299112 280152
rect 299164 280100 299170 280152
rect 305730 280100 305736 280152
rect 305788 280140 305794 280152
rect 515950 280140 515956 280152
rect 305788 280112 515956 280140
rect 305788 280100 305794 280112
rect 515950 280100 515956 280112
rect 516008 280100 516014 280152
rect 299124 280072 299152 280100
rect 373258 280072 373264 280084
rect 299124 280044 373264 280072
rect 373258 280032 373264 280044
rect 373316 280032 373322 280084
rect 302418 279964 302424 280016
rect 302476 280004 302482 280016
rect 363690 280004 363696 280016
rect 302476 279976 363696 280004
rect 302476 279964 302482 279976
rect 363690 279964 363696 279976
rect 363748 279964 363754 280016
rect 312998 279936 313004 279948
rect 296686 279908 313004 279936
rect 312998 279896 313004 279908
rect 313056 279896 313062 279948
rect 313918 262148 313924 262200
rect 313976 262188 313982 262200
rect 514754 262188 514760 262200
rect 313976 262160 514760 262188
rect 313976 262148 313982 262160
rect 514754 262148 514760 262160
rect 514812 262148 514818 262200
rect 291838 262012 291844 262064
rect 291896 262052 291902 262064
rect 292716 262055 292774 262061
rect 292716 262052 292728 262055
rect 291896 262024 292728 262052
rect 291896 262012 291902 262024
rect 292716 262021 292728 262024
rect 292762 262021 292774 262055
rect 292716 262015 292774 262021
rect 289722 261808 289728 261860
rect 289780 261848 289786 261860
rect 289780 261820 292068 261848
rect 289780 261808 289786 261820
rect 292040 261806 292068 261820
rect 295996 261792 296194 261820
rect 291930 261672 291936 261724
rect 291988 261712 291994 261724
rect 295996 261712 296024 261792
rect 291988 261684 296024 261712
rect 291988 261672 291994 261684
rect 299290 261196 299296 261248
rect 299348 261245 299354 261248
rect 299348 261239 299385 261245
rect 299373 261205 299385 261239
rect 299348 261199 299385 261205
rect 309659 261239 309717 261245
rect 309659 261205 309671 261239
rect 309705 261236 309717 261239
rect 312722 261236 312728 261248
rect 309705 261208 312728 261236
rect 309705 261205 309717 261208
rect 309659 261199 309717 261205
rect 299348 261196 299354 261199
rect 312722 261196 312728 261208
rect 312780 261196 312786 261248
rect 308876 260908 308904 261170
rect 308858 260856 308864 260908
rect 308916 260856 308922 260908
rect 295892 260825 295944 260831
rect 295892 260767 295944 260773
rect 302792 260825 302844 260831
rect 302792 260767 302844 260773
rect 306196 260825 306248 260831
rect 312538 260788 312544 260840
rect 312596 260828 312602 260840
rect 514754 260828 514760 260840
rect 312596 260800 514760 260828
rect 312596 260788 312602 260800
rect 514754 260788 514760 260800
rect 514812 260788 514818 260840
rect 306196 260767 306248 260773
rect 314010 259360 314016 259412
rect 314068 259400 314074 259412
rect 514754 259400 514760 259412
rect 314068 259372 514760 259400
rect 314068 259360 314074 259372
rect 514754 259360 514760 259372
rect 514812 259360 514818 259412
rect 302786 259292 302792 259344
rect 302844 259332 302850 259344
rect 363598 259332 363604 259344
rect 302844 259304 363604 259332
rect 302844 259292 302850 259304
rect 363598 259292 363604 259304
rect 363656 259292 363662 259344
rect 306190 258000 306196 258052
rect 306248 258040 306254 258052
rect 515858 258040 515864 258052
rect 306248 258012 515864 258040
rect 306248 258000 306254 258012
rect 515858 258000 515864 258012
rect 515916 258000 515922 258052
rect 295886 257932 295892 257984
rect 295944 257972 295950 257984
rect 311526 257972 311532 257984
rect 295944 257944 311532 257972
rect 295944 257932 295950 257944
rect 311526 257932 311532 257944
rect 311584 257932 311590 257984
rect 312814 257932 312820 257984
rect 312872 257972 312878 257984
rect 514754 257972 514760 257984
rect 312872 257944 514760 257972
rect 312872 257932 312878 257944
rect 514754 257932 514760 257944
rect 514812 257932 514818 257984
rect 299198 257864 299204 257916
rect 299256 257904 299262 257916
rect 313090 257904 313096 257916
rect 299256 257876 313096 257904
rect 299256 257864 299262 257876
rect 313090 257864 313096 257876
rect 313148 257864 313154 257916
rect 311434 256640 311440 256692
rect 311492 256680 311498 256692
rect 514754 256680 514760 256692
rect 311492 256652 514760 256680
rect 311492 256640 311498 256652
rect 514754 256640 514760 256652
rect 514812 256640 514818 256692
rect 314286 255212 314292 255264
rect 314344 255252 314350 255264
rect 514754 255252 514760 255264
rect 314344 255224 514760 255252
rect 314344 255212 314350 255224
rect 514754 255212 514760 255224
rect 514812 255212 514818 255264
rect 370498 253852 370504 253904
rect 370556 253892 370562 253904
rect 514754 253892 514760 253904
rect 370556 253864 514760 253892
rect 370556 253852 370562 253864
rect 514754 253852 514760 253864
rect 514812 253852 514818 253904
rect 313182 252492 313188 252544
rect 313240 252532 313246 252544
rect 514754 252532 514760 252544
rect 313240 252504 514760 252532
rect 313240 252492 313246 252504
rect 514754 252492 514760 252504
rect 514812 252492 514818 252544
rect 311710 251132 311716 251184
rect 311768 251172 311774 251184
rect 514754 251172 514760 251184
rect 311768 251144 514760 251172
rect 311768 251132 311774 251144
rect 514754 251132 514760 251144
rect 514812 251132 514818 251184
rect 312906 249704 312912 249756
rect 312964 249744 312970 249756
rect 514754 249744 514760 249756
rect 312964 249716 514760 249744
rect 312964 249704 312970 249716
rect 514754 249704 514760 249716
rect 514812 249704 514818 249756
rect 371878 248344 371884 248396
rect 371936 248384 371942 248396
rect 514754 248384 514760 248396
rect 371936 248356 514760 248384
rect 371936 248344 371942 248356
rect 514754 248344 514760 248356
rect 514812 248344 514818 248396
rect 312722 246984 312728 247036
rect 312780 247024 312786 247036
rect 514754 247024 514760 247036
rect 312780 246996 514760 247024
rect 312780 246984 312786 246996
rect 514754 246984 514760 246996
rect 514812 246984 514818 247036
rect 313918 242904 313924 242956
rect 313976 242944 313982 242956
rect 514754 242944 514760 242956
rect 313976 242916 514760 242944
rect 313976 242904 313982 242916
rect 514754 242904 514760 242916
rect 514812 242904 514818 242956
rect 289722 241000 289728 241052
rect 289780 241000 289786 241052
rect 291838 241000 291844 241052
rect 291896 241040 291902 241052
rect 293750 241043 293808 241049
rect 293750 241040 293762 241043
rect 291896 241012 293762 241040
rect 291896 241000 291902 241012
rect 293750 241009 293762 241012
rect 293796 241009 293808 241043
rect 293750 241003 293808 241009
rect 289740 240972 289768 241000
rect 289740 240944 292068 240972
rect 292040 240806 292068 240944
rect 307944 240848 307996 240854
rect 297015 240839 297073 240845
rect 297015 240836 297027 240839
rect 296686 240808 297027 240836
rect 291930 240660 291936 240712
rect 291988 240700 291994 240712
rect 296686 240700 296714 240808
rect 297015 240805 297027 240808
rect 297061 240805 297073 240839
rect 297015 240799 297073 240805
rect 308858 240836 308864 240848
rect 307996 240808 308864 240836
rect 308858 240796 308864 240808
rect 308916 240796 308922 240848
rect 307944 240790 307996 240796
rect 291988 240672 296714 240700
rect 291988 240660 291994 240672
rect 298922 240184 298928 240236
rect 298980 240233 298986 240236
rect 298980 240227 299026 240233
rect 299014 240193 299026 240227
rect 298980 240187 299026 240193
rect 298980 240184 298986 240187
rect 305454 240184 305460 240236
rect 305512 240233 305518 240236
rect 305512 240227 305556 240233
rect 305544 240193 305556 240227
rect 305512 240187 305556 240193
rect 305512 240184 305518 240187
rect 295708 239825 295760 239831
rect 295708 239767 295760 239773
rect 302240 239825 302292 239831
rect 514938 239816 514944 239828
rect 308784 239788 514944 239816
rect 514938 239776 514944 239788
rect 514996 239776 515002 239828
rect 302240 239767 302292 239773
rect 299014 238688 299020 238740
rect 299072 238728 299078 238740
rect 359458 238728 359464 238740
rect 299072 238700 359464 238728
rect 299072 238688 299078 238700
rect 359458 238688 359464 238700
rect 359516 238688 359522 238740
rect 295702 237328 295708 237380
rect 295760 237368 295766 237380
rect 295760 237340 296714 237368
rect 295760 237328 295766 237340
rect 296686 237232 296714 237340
rect 302234 237328 302240 237380
rect 302292 237368 302298 237380
rect 377398 237368 377404 237380
rect 302292 237340 377404 237368
rect 302292 237328 302298 237340
rect 377398 237328 377404 237340
rect 377456 237328 377462 237380
rect 305546 237260 305552 237312
rect 305604 237300 305610 237312
rect 366358 237300 366364 237312
rect 305604 237272 366364 237300
rect 305604 237260 305610 237272
rect 366358 237260 366364 237272
rect 366416 237260 366422 237312
rect 311250 237232 311256 237244
rect 296686 237204 311256 237232
rect 311250 237192 311256 237204
rect 311308 237192 311314 237244
rect 289722 219988 289728 220040
rect 289780 220028 289786 220040
rect 289780 220000 292068 220028
rect 289780 219988 289786 220000
rect 292040 219807 292068 220000
rect 297909 219827 297967 219833
rect 297909 219824 297921 219827
rect 296686 219796 297921 219824
rect 291930 219648 291936 219700
rect 291988 219688 291994 219700
rect 296686 219688 296714 219796
rect 297909 219793 297921 219796
rect 297955 219793 297967 219827
rect 297909 219787 297967 219793
rect 291988 219660 296714 219688
rect 291988 219648 291994 219660
rect 313918 219144 313924 219156
rect 310992 219116 313924 219144
rect 310992 219095 311020 219116
rect 313918 219104 313924 219116
rect 313976 219104 313982 219156
rect 296168 218825 296220 218831
rect 296168 218767 296220 218773
rect 299848 218825 299900 218831
rect 299848 218767 299900 218773
rect 307300 218825 307352 218831
rect 307300 218767 307352 218773
rect 303614 218745 303620 218748
rect 303574 218739 303620 218745
rect 303574 218705 303586 218739
rect 303574 218699 303620 218705
rect 303614 218696 303620 218699
rect 303672 218696 303678 218748
rect 296162 216588 296168 216640
rect 296220 216628 296226 216640
rect 296220 216600 296714 216628
rect 296220 216588 296226 216600
rect 296686 216492 296714 216600
rect 303614 216588 303620 216640
rect 303672 216628 303678 216640
rect 303672 216600 306374 216628
rect 303672 216588 303678 216600
rect 306346 216560 306374 216600
rect 307294 216588 307300 216640
rect 307352 216628 307358 216640
rect 515766 216628 515772 216640
rect 307352 216600 515772 216628
rect 307352 216588 307358 216600
rect 515766 216588 515772 216600
rect 515824 216588 515830 216640
rect 364978 216560 364984 216572
rect 306346 216532 364984 216560
rect 364978 216520 364984 216532
rect 365036 216520 365042 216572
rect 311158 216492 311164 216504
rect 296686 216464 311164 216492
rect 311158 216452 311164 216464
rect 311216 216452 311222 216504
rect 299842 216384 299848 216436
rect 299900 216424 299906 216436
rect 311618 216424 311624 216436
rect 299900 216396 311624 216424
rect 299900 216384 299906 216396
rect 311618 216384 311624 216396
rect 311676 216384 311682 216436
rect 289722 206252 289728 206304
rect 289780 206292 289786 206304
rect 580166 206292 580172 206304
rect 289780 206264 580172 206292
rect 289780 206252 289786 206264
rect 580166 206252 580172 206264
rect 580224 206252 580230 206304
rect 297542 199384 297548 199436
rect 297600 199384 297606 199436
rect 300762 199384 300768 199436
rect 300820 199384 300826 199436
rect 304810 199384 304816 199436
rect 304868 199384 304874 199436
rect 297560 199232 297588 199384
rect 300780 199232 300808 199384
rect 297542 199180 297548 199232
rect 297600 199180 297606 199232
rect 300762 199180 300768 199232
rect 300820 199180 300826 199232
rect 304828 198892 304856 199384
rect 304810 198840 304816 198892
rect 304868 198840 304874 198892
rect 289722 198772 289728 198824
rect 289780 198812 289786 198824
rect 289780 198784 292068 198812
rect 289780 198772 289786 198784
rect 293678 198780 293684 198832
rect 293736 198780 293742 198832
rect 295518 198209 295524 198212
rect 295490 198203 295524 198209
rect 295490 198169 295502 198203
rect 295490 198163 295524 198169
rect 295518 198160 295524 198163
rect 295576 198160 295582 198212
rect 307570 198200 307576 198212
rect 307036 198184 307576 198200
rect 306958 198172 307576 198184
rect 306958 198156 307064 198172
rect 307570 198160 307576 198172
rect 307628 198160 307634 198212
rect 307698 198203 307756 198209
rect 307698 198169 307710 198203
rect 307744 198200 307756 198203
rect 307744 198172 316034 198200
rect 307744 198169 307756 198172
rect 307698 198163 307756 198169
rect 298560 197825 298612 197831
rect 304632 197825 304684 197831
rect 298560 197767 298612 197773
rect 301608 197316 301636 197778
rect 304632 197767 304684 197773
rect 316006 197792 316034 198172
rect 515950 197792 515956 197804
rect 316006 197764 515956 197792
rect 515950 197752 515956 197764
rect 516008 197752 516014 197804
rect 362218 197316 362224 197328
rect 301608 197288 362224 197316
rect 362218 197276 362224 197288
rect 362276 197276 362282 197328
rect 295518 195916 295524 195968
rect 295576 195956 295582 195968
rect 295576 195928 296714 195956
rect 295576 195916 295582 195928
rect 296686 195888 296714 195928
rect 304626 195916 304632 195968
rect 304684 195956 304690 195968
rect 515674 195956 515680 195968
rect 304684 195928 515680 195956
rect 304684 195916 304690 195928
rect 515674 195916 515680 195928
rect 515732 195916 515738 195968
rect 312630 195888 312636 195900
rect 296686 195860 312636 195888
rect 312630 195848 312636 195860
rect 312688 195848 312694 195900
rect 298554 195780 298560 195832
rect 298612 195820 298618 195832
rect 311342 195820 311348 195832
rect 298612 195792 311348 195820
rect 298612 195780 298618 195792
rect 311342 195780 311348 195792
rect 311400 195780 311406 195832
rect 296714 178644 296720 178696
rect 296772 178644 296778 178696
rect 293954 178576 293960 178628
rect 294012 178576 294018 178628
rect 293972 178412 294000 178576
rect 294046 178412 294052 178424
rect 293972 178384 294052 178412
rect 294046 178372 294052 178384
rect 294104 178372 294110 178424
rect 296585 178211 296643 178217
rect 296585 178177 296597 178211
rect 296631 178208 296643 178211
rect 296732 178208 296760 178644
rect 300762 178576 300768 178628
rect 300820 178576 300826 178628
rect 304534 178616 304540 178628
rect 303816 178588 304540 178616
rect 300780 178424 300808 178576
rect 303816 178424 303844 178588
rect 304534 178576 304540 178588
rect 304592 178576 304598 178628
rect 306926 178576 306932 178628
rect 306984 178576 306990 178628
rect 300762 178372 300768 178424
rect 300820 178372 300826 178424
rect 303798 178372 303804 178424
rect 303856 178372 303862 178424
rect 306834 178372 306840 178424
rect 306892 178412 306898 178424
rect 306944 178412 306972 178576
rect 306892 178384 306972 178412
rect 306892 178372 306898 178384
rect 296631 178180 296760 178208
rect 296631 178177 296643 178180
rect 296585 178171 296643 178177
rect 289722 177964 289728 178016
rect 289780 178004 289786 178016
rect 292040 178004 292068 178006
rect 289780 177976 292068 178004
rect 294046 177980 294052 178032
rect 294104 177980 294110 178032
rect 289780 177964 289786 177976
rect 295518 177401 295524 177404
rect 295490 177395 295524 177401
rect 295490 177361 295502 177395
rect 295490 177355 295524 177361
rect 295518 177352 295524 177355
rect 295576 177352 295582 177404
rect 307698 177395 307756 177401
rect 307698 177361 307710 177395
rect 307744 177392 307756 177395
rect 307744 177364 316034 177392
rect 307744 177361 307756 177364
rect 307698 177355 307756 177361
rect 298560 177025 298612 177031
rect 298560 176967 298612 176973
rect 301596 177025 301648 177031
rect 301596 176967 301648 176973
rect 304632 177025 304684 177031
rect 304632 176967 304684 176973
rect 316006 176984 316034 177364
rect 515858 176984 515864 176996
rect 316006 176956 515864 176984
rect 515858 176944 515864 176956
rect 515916 176944 515922 176996
rect 295518 175176 295524 175228
rect 295576 175216 295582 175228
rect 515398 175216 515404 175228
rect 295576 175188 515404 175216
rect 295576 175176 295582 175188
rect 515398 175176 515404 175188
rect 515456 175176 515462 175228
rect 298554 175108 298560 175160
rect 298612 175148 298618 175160
rect 515490 175148 515496 175160
rect 298612 175120 515496 175148
rect 298612 175108 298618 175120
rect 515490 175108 515496 175120
rect 515548 175108 515554 175160
rect 301590 175040 301596 175092
rect 301648 175040 301654 175092
rect 304626 175040 304632 175092
rect 304684 175080 304690 175092
rect 515582 175080 515588 175092
rect 304684 175052 515588 175080
rect 304684 175040 304690 175052
rect 515582 175040 515588 175052
rect 515640 175040 515646 175092
rect 301608 175012 301636 175040
rect 345658 175012 345664 175024
rect 301608 174984 345664 175012
rect 345658 174972 345664 174984
rect 345716 174972 345722 175024
<< via1 >>
rect 301136 493348 301188 493400
rect 289728 492668 289780 492720
rect 296996 492780 297048 492832
rect 308404 492668 308456 492720
rect 292488 492600 292540 492652
rect 296996 492600 297048 492652
rect 301964 492235 302016 492244
rect 301964 492201 301967 492235
rect 301967 492201 302016 492235
rect 301964 492192 302016 492201
rect 309600 492192 309652 492244
rect 291936 492124 291988 492176
rect 295616 491773 295668 491825
rect 298744 491773 298796 491825
rect 305092 491773 305144 491825
rect 313924 491444 313976 491496
rect 305092 488996 305144 489048
rect 312728 488996 312780 489048
rect 301964 488656 302016 488708
rect 312912 488656 312964 488708
rect 298744 488588 298796 488640
rect 367744 488588 367796 488640
rect 295616 488520 295668 488572
rect 405004 488520 405056 488572
rect 296628 473288 296680 473340
rect 298376 473288 298428 473340
rect 298376 472404 298428 472456
rect 302424 472404 302476 472456
rect 298376 472132 298428 472184
rect 302976 472132 303028 472184
rect 291844 471996 291896 472048
rect 289728 471928 289780 471980
rect 298376 471780 298428 471832
rect 295984 471180 296036 471232
rect 299572 471223 299624 471232
rect 299572 471189 299623 471223
rect 299623 471189 299624 471223
rect 299572 471180 299624 471189
rect 303160 471223 303212 471232
rect 303160 471189 303208 471223
rect 303208 471189 303212 471223
rect 303160 471180 303212 471189
rect 310520 471248 310572 471300
rect 306748 471223 306800 471232
rect 306748 471189 306793 471223
rect 306793 471189 306800 471223
rect 306748 471180 306800 471189
rect 312544 471180 312596 471232
rect 302148 470704 302200 470756
rect 302976 470976 303028 471028
rect 306748 469140 306800 469192
rect 314108 469072 314160 469124
rect 296076 468052 296128 468104
rect 338764 467984 338816 468036
rect 303160 467916 303212 467968
rect 363604 467916 363656 467968
rect 299664 467848 299716 467900
rect 388444 467848 388496 467900
rect 338764 451868 338816 451920
rect 515404 451868 515456 451920
rect 289728 450780 289780 450832
rect 314016 449896 314068 449948
rect 305736 449773 305788 449825
rect 295800 449735 295852 449744
rect 295800 449701 295803 449735
rect 295803 449701 295852 449735
rect 295800 449692 295852 449701
rect 299112 449735 299164 449744
rect 299112 449701 299120 449735
rect 299120 449701 299164 449735
rect 299112 449692 299164 449701
rect 302424 449735 302476 449744
rect 302424 449701 302437 449735
rect 302437 449701 302476 449735
rect 302424 449692 302476 449701
rect 305736 447652 305788 447704
rect 314200 447652 314252 447704
rect 295800 447244 295852 447296
rect 299112 447244 299164 447296
rect 302424 447244 302476 447296
rect 370596 447244 370648 447296
rect 406384 447176 406436 447228
rect 443644 447108 443696 447160
rect 296076 430040 296128 430092
rect 289728 429768 289780 429820
rect 292764 429780 292816 429832
rect 299296 429199 299348 429208
rect 299296 429165 299341 429199
rect 299341 429165 299348 429199
rect 299296 429156 299348 429165
rect 309140 428884 309192 428936
rect 296536 428748 296588 428800
rect 302792 428773 302844 428825
rect 306196 428773 306248 428825
rect 312820 428748 312872 428800
rect 306196 425552 306248 425604
rect 314384 425552 314436 425604
rect 299296 425144 299348 425196
rect 302792 425144 302844 425196
rect 391204 425144 391256 425196
rect 427084 425076 427136 425128
rect 405004 422220 405056 422272
rect 514760 422220 514812 422272
rect 524328 421404 524380 421456
rect 527180 421404 527232 421456
rect 517428 421336 517480 421388
rect 518992 421336 519044 421388
rect 526996 421336 527048 421388
rect 529204 421336 529256 421388
rect 443644 419432 443696 419484
rect 514760 419432 514812 419484
rect 296536 418072 296588 418124
rect 514760 418072 514812 418124
rect 291844 409028 291896 409080
rect 289728 408688 289780 408740
rect 291936 408688 291988 408740
rect 298928 408212 298980 408264
rect 305644 408144 305696 408196
rect 309048 408144 309100 408196
rect 295708 407773 295760 407825
rect 302240 407773 302292 407825
rect 311440 407736 311492 407788
rect 313004 407124 313056 407176
rect 514760 407124 514812 407176
rect 311532 405696 311584 405748
rect 514760 405696 514812 405748
rect 295708 405628 295760 405680
rect 515404 405628 515456 405680
rect 302240 405560 302292 405612
rect 305644 405560 305696 405612
rect 314476 405560 314528 405612
rect 313188 405492 313240 405544
rect 298928 404608 298980 404660
rect 446404 404404 446456 404456
rect 311256 404336 311308 404388
rect 514760 404336 514812 404388
rect 311164 402976 311216 403028
rect 514760 402976 514812 403028
rect 312636 401616 312688 401668
rect 514760 401616 514812 401668
rect 289728 388016 289780 388068
rect 291844 388016 291896 388068
rect 309048 388059 309100 388068
rect 309048 388025 309057 388059
rect 309057 388025 309091 388059
rect 309091 388025 309100 388059
rect 309048 388016 309100 388025
rect 302240 387780 302292 387832
rect 311900 387676 311952 387728
rect 303620 387200 303672 387252
rect 296168 386773 296220 386825
rect 299848 386773 299900 386825
rect 307300 386773 307352 386825
rect 314292 386792 314344 386844
rect 296168 384956 296220 385008
rect 515864 384956 515916 385008
rect 299848 384888 299900 384940
rect 300768 384888 300820 384940
rect 303620 384888 303672 384940
rect 308404 384888 308456 384940
rect 307300 384004 307352 384056
rect 393964 383664 394016 383716
rect 367744 382168 367796 382220
rect 514760 382168 514812 382220
rect 388444 380808 388496 380860
rect 514760 380808 514812 380860
rect 406384 379448 406436 379500
rect 514760 379448 514812 379500
rect 427084 378088 427136 378140
rect 514760 378088 514812 378140
rect 446404 376660 446456 376712
rect 514760 376660 514812 376712
rect 300768 375300 300820 375352
rect 514760 375300 514812 375352
rect 373264 367072 373316 367124
rect 514760 367072 514812 367124
rect 289728 367004 289780 367056
rect 294052 366780 294104 366832
rect 300216 366780 300268 366832
rect 307668 366800 307720 366852
rect 308036 366800 308088 366852
rect 295524 366231 295576 366240
rect 295524 366197 295537 366231
rect 295537 366197 295576 366231
rect 295524 366188 295576 366197
rect 298560 365773 298612 365825
rect 301596 365773 301648 365825
rect 304632 365773 304684 365825
rect 370504 365780 370556 365832
rect 313096 365712 313148 365764
rect 514760 365712 514812 365764
rect 359464 364352 359516 364404
rect 514760 364352 514812 364404
rect 295524 364284 295576 364336
rect 515496 364284 515548 364336
rect 298560 364216 298612 364268
rect 515312 364216 515364 364268
rect 301596 364148 301648 364200
rect 308496 364148 308548 364200
rect 304632 363332 304684 363384
rect 314568 363332 314620 363384
rect 311624 362924 311676 362976
rect 514760 362924 514812 362976
rect 311348 361564 311400 361616
rect 514760 361564 514812 361616
rect 299572 346400 299624 346452
rect 291752 346060 291804 346112
rect 289728 345992 289780 346044
rect 294420 345992 294472 346044
rect 307852 345788 307904 345840
rect 313188 345652 313240 345704
rect 515312 345652 515364 345704
rect 295524 345219 295576 345228
rect 295524 345185 295536 345219
rect 295536 345185 295576 345219
rect 295524 345176 295576 345185
rect 313188 344836 313240 344888
rect 298560 344773 298612 344825
rect 302148 344768 302200 344820
rect 304632 344773 304684 344825
rect 295524 342184 295576 342236
rect 515772 342184 515824 342236
rect 298560 342116 298612 342168
rect 516048 342116 516100 342168
rect 312912 342048 312964 342100
rect 514760 342048 514812 342100
rect 304632 341300 304684 341352
rect 309784 341232 309836 341284
rect 363604 340824 363656 340876
rect 514760 340824 514812 340876
rect 370596 339396 370648 339448
rect 514760 339396 514812 339448
rect 391204 338036 391256 338088
rect 514760 338036 514812 338088
rect 308404 335248 308456 335300
rect 514760 335248 514812 335300
rect 308496 333888 308548 333940
rect 514760 333888 514812 333940
rect 302148 332528 302200 332580
rect 514760 332528 514812 332580
rect 363696 327088 363748 327140
rect 514760 327088 514812 327140
rect 363604 325660 363656 325712
rect 514760 325660 514812 325712
rect 294788 325388 294840 325440
rect 307852 325388 307904 325440
rect 308496 325388 308548 325440
rect 294788 325184 294840 325236
rect 289728 324776 289780 324828
rect 296996 324780 297048 324832
rect 308404 324912 308456 324964
rect 308588 324776 308640 324828
rect 291844 324640 291896 324692
rect 296996 324640 297048 324692
rect 377404 324300 377456 324352
rect 514760 324300 514812 324352
rect 294788 324144 294840 324196
rect 308496 324232 308548 324284
rect 292396 323892 292448 323944
rect 295616 323773 295668 323825
rect 298744 323773 298796 323825
rect 305092 323773 305144 323825
rect 301964 323688 302016 323740
rect 311716 323484 311768 323536
rect 364984 322940 365036 322992
rect 514760 322940 514812 322992
rect 362224 321580 362276 321632
rect 514760 321580 514812 321632
rect 295616 321512 295668 321564
rect 515680 321512 515732 321564
rect 298744 321444 298796 321496
rect 515956 321444 516008 321496
rect 301964 321376 302016 321428
rect 516048 321376 516100 321428
rect 345664 320152 345716 320204
rect 514760 320152 514812 320204
rect 305092 318044 305144 318096
rect 366364 318044 366416 318096
rect 294972 304376 295024 304428
rect 298468 304376 298520 304428
rect 302424 304376 302476 304428
rect 306012 304376 306064 304428
rect 309600 304376 309652 304428
rect 309784 304376 309836 304428
rect 515680 304240 515732 304292
rect 294972 304172 295024 304224
rect 298468 304172 298520 304224
rect 302424 304172 302476 304224
rect 306012 304172 306064 304224
rect 309600 304172 309652 304224
rect 289728 303764 289780 303816
rect 312912 303152 312964 303204
rect 314108 303084 314160 303136
rect 515036 303084 515088 303136
rect 314568 303016 314620 303068
rect 515956 303016 516008 303068
rect 314200 302948 314252 303000
rect 514944 302948 514996 303000
rect 312728 302880 312780 302932
rect 514760 302880 514812 302932
rect 296076 302773 296128 302825
rect 299664 302773 299716 302825
rect 306840 302773 306892 302825
rect 515772 302132 515824 302184
rect 517428 301792 517480 301844
rect 518900 301792 518952 301844
rect 296076 300772 296128 300824
rect 515588 300772 515640 300824
rect 299664 300704 299716 300756
rect 515864 300704 515916 300756
rect 306840 299752 306892 299804
rect 307668 299752 307720 299804
rect 314384 298052 314436 298104
rect 514760 298052 514812 298104
rect 314476 296624 314528 296676
rect 514760 296624 514812 296676
rect 393964 295264 394016 295316
rect 514760 295264 514812 295316
rect 366364 291116 366416 291168
rect 514760 291116 514812 291168
rect 307668 289756 307720 289808
rect 514760 289756 514812 289808
rect 366364 284316 366416 284368
rect 514760 284316 514812 284368
rect 291844 282888 291896 282940
rect 289728 282616 289780 282668
rect 291936 282616 291988 282668
rect 309140 282140 309192 282192
rect 295800 281773 295852 281825
rect 299112 281773 299164 281825
rect 302424 281773 302476 281825
rect 305736 281773 305788 281825
rect 371884 281800 371936 281852
rect 295800 280100 295852 280152
rect 299112 280100 299164 280152
rect 305736 280100 305788 280152
rect 515956 280100 516008 280152
rect 373264 280032 373316 280084
rect 302424 279964 302476 280016
rect 363696 279964 363748 280016
rect 313004 279896 313056 279948
rect 313924 262148 313976 262200
rect 514760 262148 514812 262200
rect 291844 262012 291896 262064
rect 289728 261808 289780 261860
rect 291936 261672 291988 261724
rect 299296 261239 299348 261248
rect 299296 261205 299339 261239
rect 299339 261205 299348 261239
rect 299296 261196 299348 261205
rect 312728 261196 312780 261248
rect 308864 260856 308916 260908
rect 295892 260773 295944 260825
rect 302792 260773 302844 260825
rect 306196 260773 306248 260825
rect 312544 260788 312596 260840
rect 514760 260788 514812 260840
rect 314016 259360 314068 259412
rect 514760 259360 514812 259412
rect 302792 259292 302844 259344
rect 363604 259292 363656 259344
rect 306196 258000 306248 258052
rect 515864 258000 515916 258052
rect 295892 257932 295944 257984
rect 311532 257932 311584 257984
rect 312820 257932 312872 257984
rect 514760 257932 514812 257984
rect 299204 257864 299256 257916
rect 313096 257864 313148 257916
rect 311440 256640 311492 256692
rect 514760 256640 514812 256692
rect 314292 255212 314344 255264
rect 514760 255212 514812 255264
rect 370504 253852 370556 253904
rect 514760 253852 514812 253904
rect 313188 252492 313240 252544
rect 514760 252492 514812 252544
rect 311716 251132 311768 251184
rect 514760 251132 514812 251184
rect 312912 249704 312964 249756
rect 514760 249704 514812 249756
rect 371884 248344 371936 248396
rect 514760 248344 514812 248396
rect 312728 246984 312780 247036
rect 514760 246984 514812 247036
rect 313924 242904 313976 242956
rect 514760 242904 514812 242956
rect 289728 241000 289780 241052
rect 291844 241000 291896 241052
rect 291936 240660 291988 240712
rect 307944 240796 307996 240848
rect 308864 240796 308916 240848
rect 298928 240184 298980 240236
rect 305460 240227 305512 240236
rect 305460 240193 305510 240227
rect 305510 240193 305512 240227
rect 305460 240184 305512 240193
rect 295708 239773 295760 239825
rect 302240 239773 302292 239825
rect 514944 239776 514996 239828
rect 299020 238688 299072 238740
rect 359464 238688 359516 238740
rect 295708 237328 295760 237380
rect 302240 237328 302292 237380
rect 377404 237328 377456 237380
rect 305552 237260 305604 237312
rect 366364 237260 366416 237312
rect 311256 237192 311308 237244
rect 289728 219988 289780 220040
rect 291936 219648 291988 219700
rect 313924 219104 313976 219156
rect 296168 218773 296220 218825
rect 299848 218773 299900 218825
rect 307300 218773 307352 218825
rect 303620 218696 303672 218748
rect 296168 216588 296220 216640
rect 303620 216588 303672 216640
rect 307300 216588 307352 216640
rect 515772 216588 515824 216640
rect 364984 216520 365036 216572
rect 311164 216452 311216 216504
rect 299848 216384 299900 216436
rect 311624 216384 311676 216436
rect 289728 206252 289780 206304
rect 580172 206252 580224 206304
rect 297548 199384 297600 199436
rect 300768 199384 300820 199436
rect 304816 199384 304868 199436
rect 297548 199180 297600 199232
rect 300768 199180 300820 199232
rect 304816 198840 304868 198892
rect 289728 198772 289780 198824
rect 293684 198780 293736 198832
rect 295524 198203 295576 198212
rect 295524 198169 295536 198203
rect 295536 198169 295576 198203
rect 295524 198160 295576 198169
rect 307576 198160 307628 198212
rect 298560 197773 298612 197825
rect 304632 197773 304684 197825
rect 515956 197752 516008 197804
rect 362224 197276 362276 197328
rect 295524 195916 295576 195968
rect 304632 195916 304684 195968
rect 515680 195916 515732 195968
rect 312636 195848 312688 195900
rect 298560 195780 298612 195832
rect 311348 195780 311400 195832
rect 296720 178644 296772 178696
rect 293960 178576 294012 178628
rect 294052 178372 294104 178424
rect 300768 178576 300820 178628
rect 304540 178576 304592 178628
rect 306932 178576 306984 178628
rect 300768 178372 300820 178424
rect 303804 178372 303856 178424
rect 306840 178372 306892 178424
rect 289728 177964 289780 178016
rect 294052 177980 294104 178032
rect 295524 177395 295576 177404
rect 295524 177361 295536 177395
rect 295536 177361 295576 177395
rect 295524 177352 295576 177361
rect 298560 176973 298612 177025
rect 301596 176973 301648 177025
rect 304632 176973 304684 177025
rect 515864 176944 515916 176996
rect 295524 175176 295576 175228
rect 515404 175176 515456 175228
rect 298560 175108 298612 175160
rect 515496 175108 515548 175160
rect 301596 175040 301648 175092
rect 304632 175040 304684 175092
rect 515588 175040 515640 175092
rect 345664 174972 345716 175024
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 301134 494320 301190 494329
rect 301134 494255 301190 494264
rect 309138 494320 309194 494329
rect 309138 494255 309194 494264
rect 301148 493406 301176 494255
rect 301136 493400 301188 493406
rect 301136 493342 301188 493348
rect 296996 492832 297048 492838
rect 296996 492774 297048 492780
rect 289728 492720 289780 492726
rect 289728 492662 289780 492668
rect 289740 471986 289768 492662
rect 297008 492658 297036 492774
rect 308404 492720 308456 492726
rect 308404 492662 308456 492668
rect 292488 492652 292540 492658
rect 292488 492594 292540 492600
rect 296996 492652 297048 492658
rect 296996 492594 297048 492600
rect 291936 492176 291988 492182
rect 291936 492118 291988 492124
rect 291948 489914 291976 492118
rect 292500 489914 292528 492594
rect 301964 492244 302016 492250
rect 301964 492186 302016 492192
rect 295616 491825 295668 491831
rect 295616 491767 295668 491773
rect 298744 491825 298796 491831
rect 298744 491767 298796 491773
rect 291856 489886 291976 489914
rect 292408 489886 292528 489914
rect 291856 472054 291884 489886
rect 292408 473385 292436 489886
rect 295628 488578 295656 491767
rect 298756 488646 298784 491767
rect 301976 488714 302004 492186
rect 305092 491825 305144 491831
rect 305092 491767 305144 491773
rect 305104 489054 305132 491767
rect 305092 489048 305144 489054
rect 305092 488990 305144 488996
rect 301964 488708 302016 488714
rect 301964 488650 302016 488656
rect 298744 488640 298796 488646
rect 298744 488582 298796 488588
rect 295616 488572 295668 488578
rect 295616 488514 295668 488520
rect 308416 473521 308444 492662
rect 308402 473512 308458 473521
rect 308402 473447 308458 473456
rect 309152 473385 309180 494255
rect 309600 492244 309652 492250
rect 309600 492186 309652 492192
rect 309612 489914 309640 492186
rect 313924 491496 313976 491502
rect 313924 491438 313976 491444
rect 309612 489886 309824 489914
rect 292394 473376 292450 473385
rect 292394 473311 292450 473320
rect 296626 473376 296682 473385
rect 302422 473376 302478 473385
rect 296626 473311 296628 473320
rect 296680 473311 296682 473320
rect 298376 473340 298428 473346
rect 296628 473282 296680 473288
rect 302422 473311 302478 473320
rect 309138 473376 309194 473385
rect 309138 473311 309194 473320
rect 298376 473282 298428 473288
rect 298388 472462 298416 473282
rect 302436 472462 302464 473311
rect 298376 472456 298428 472462
rect 298376 472398 298428 472404
rect 302424 472456 302476 472462
rect 309796 472433 309824 489886
rect 312728 489048 312780 489054
rect 312728 488990 312780 488996
rect 310518 473512 310574 473521
rect 310518 473447 310574 473456
rect 302424 472398 302476 472404
rect 309782 472424 309838 472433
rect 309782 472359 309838 472368
rect 298376 472184 298428 472190
rect 298376 472126 298428 472132
rect 302976 472184 303028 472190
rect 302976 472126 303028 472132
rect 309506 472152 309562 472161
rect 291844 472048 291896 472054
rect 291844 471990 291896 471996
rect 289728 471980 289780 471986
rect 289728 471922 289780 471928
rect 289740 450838 289768 471922
rect 289728 450832 289780 450838
rect 289728 450774 289780 450780
rect 289740 429826 289768 450774
rect 291856 448633 291884 471990
rect 298388 471838 298416 472126
rect 298376 471832 298428 471838
rect 298376 471774 298428 471780
rect 298388 471594 298416 471774
rect 298388 471580 298807 471594
rect 298388 471566 298821 471580
rect 295984 471232 296036 471238
rect 295984 471174 296036 471180
rect 295996 470594 296024 471174
rect 298793 470778 298821 471566
rect 299572 471232 299624 471238
rect 299572 471174 299624 471180
rect 298480 470750 298821 470778
rect 295996 470566 296116 470594
rect 296088 468110 296116 470566
rect 296076 468104 296128 468110
rect 296076 468046 296128 468052
rect 298480 451489 298508 470750
rect 299584 470594 299612 471174
rect 302988 471034 303016 472126
rect 309506 472087 309562 472096
rect 303160 471232 303212 471238
rect 303160 471174 303212 471180
rect 306748 471232 306800 471238
rect 306748 471174 306800 471180
rect 302976 471028 303028 471034
rect 302976 470970 303028 470976
rect 302148 470756 302200 470762
rect 302148 470698 302200 470704
rect 299584 470566 299704 470594
rect 299676 467906 299704 470566
rect 299664 467900 299716 467906
rect 299664 467842 299716 467848
rect 302160 452849 302188 470698
rect 303172 467974 303200 471174
rect 306760 469198 306788 471174
rect 309520 470594 309548 472087
rect 310532 471306 310560 473447
rect 310520 471300 310572 471306
rect 310520 471242 310572 471248
rect 309060 470566 309548 470594
rect 306748 469192 306800 469198
rect 306748 469134 306800 469140
rect 303160 467968 303212 467974
rect 303160 467910 303212 467916
rect 302146 452840 302202 452849
rect 302146 452775 302202 452784
rect 302160 451489 302188 452775
rect 304906 452704 304962 452713
rect 304906 452639 304962 452648
rect 304920 451625 304948 452639
rect 309060 452554 309088 470566
rect 310532 453937 310560 471242
rect 312544 471232 312596 471238
rect 312544 471174 312596 471180
rect 309230 453928 309286 453937
rect 309230 453863 309286 453872
rect 310518 453928 310574 453937
rect 310518 453863 310574 453872
rect 309244 452713 309272 453863
rect 309414 452840 309470 452849
rect 309414 452775 309470 452784
rect 309230 452704 309286 452713
rect 309230 452639 309286 452648
rect 309060 452526 309180 452554
rect 304906 451616 304962 451625
rect 304906 451551 304962 451560
rect 298466 451480 298522 451489
rect 298466 451415 298522 451424
rect 302146 451480 302202 451489
rect 302146 451415 302202 451424
rect 298098 451072 298154 451081
rect 298098 451007 298154 451016
rect 301560 451072 301616 451081
rect 301560 451007 301616 451016
rect 304877 451072 304933 451081
rect 304877 451007 304933 451016
rect 298112 450922 298140 451007
rect 298112 450908 298271 450922
rect 298112 450894 298285 450908
rect 294940 450242 294968 450364
rect 294892 450214 294968 450242
rect 291842 448624 291898 448633
rect 291842 448559 291898 448568
rect 293958 448624 294014 448633
rect 293958 448559 294014 448568
rect 294786 448624 294842 448633
rect 294892 448610 294920 450214
rect 298257 449970 298285 450894
rect 298112 449942 298285 449970
rect 295800 449744 295852 449750
rect 295800 449686 295852 449692
rect 294842 448582 294920 448610
rect 294786 448559 294842 448568
rect 291842 430808 291898 430817
rect 291842 430743 291898 430752
rect 289728 429820 289780 429826
rect 289728 429762 289780 429768
rect 289740 408746 289768 429762
rect 291856 422294 291884 430743
rect 293972 430681 294000 448559
rect 295812 447302 295840 449686
rect 295800 447296 295852 447302
rect 295800 447238 295852 447244
rect 298112 430817 298140 449942
rect 308232 449857 308260 450364
rect 308218 449848 308274 449857
rect 305736 449825 305788 449831
rect 308218 449783 308274 449792
rect 309046 449848 309102 449857
rect 309152 449834 309180 452526
rect 309102 449806 309180 449834
rect 309046 449783 309102 449792
rect 305736 449767 305788 449773
rect 299112 449744 299164 449750
rect 299112 449686 299164 449692
rect 302424 449744 302476 449750
rect 302424 449686 302476 449692
rect 299124 447302 299152 449686
rect 302436 447302 302464 449686
rect 305748 447710 305776 449767
rect 305736 447704 305788 447710
rect 305736 447646 305788 447652
rect 299112 447296 299164 447302
rect 299112 447238 299164 447244
rect 302424 447296 302476 447302
rect 302424 447238 302476 447244
rect 308232 441614 308260 449783
rect 308232 441586 308904 441614
rect 305550 432168 305606 432177
rect 305550 432103 305606 432112
rect 302054 432032 302110 432041
rect 302054 431967 302110 431976
rect 298098 430808 298154 430817
rect 298098 430743 298154 430752
rect 293958 430672 294014 430681
rect 293958 430607 294014 430616
rect 302068 430522 302096 431967
rect 305564 430545 305592 432103
rect 308876 430545 308904 441586
rect 309244 432177 309272 452639
rect 309428 441614 309456 452775
rect 309428 441586 309916 441614
rect 309230 432168 309286 432177
rect 309230 432103 309286 432112
rect 309244 431954 309272 432103
rect 309888 432041 309916 441586
rect 309874 432032 309930 432041
rect 309874 431967 309930 431976
rect 309244 431926 309824 431954
rect 302146 430536 302202 430545
rect 302068 430494 302146 430522
rect 302146 430471 302202 430480
rect 305550 430536 305606 430545
rect 305550 430471 305606 430480
rect 308862 430536 308918 430545
rect 308862 430471 308918 430480
rect 296074 430264 296130 430273
rect 296074 430199 296130 430208
rect 309322 430264 309378 430273
rect 309322 430199 309378 430208
rect 296088 430098 296116 430199
rect 296076 430092 296128 430098
rect 301935 430072 301944 430128
rect 302000 430072 302009 430128
rect 305379 430072 305388 430128
rect 305444 430072 305453 430128
rect 296076 430034 296128 430040
rect 292762 429856 292818 429865
rect 292500 429814 292762 429842
rect 292500 426329 292528 429814
rect 292762 429791 292764 429800
rect 292816 429791 292818 429800
rect 292764 429774 292816 429780
rect 299296 429208 299348 429214
rect 299296 429150 299348 429156
rect 296536 428800 296588 428806
rect 296536 428742 296588 428748
rect 292486 426320 292542 426329
rect 292486 426255 292542 426264
rect 293958 426320 294014 426329
rect 293958 426255 294014 426264
rect 291856 422266 291976 422294
rect 291106 410136 291162 410145
rect 291106 410071 291162 410080
rect 289728 408740 289780 408746
rect 289728 408682 289780 408688
rect 289740 388074 289768 408682
rect 291120 389473 291148 410071
rect 291842 410000 291898 410009
rect 291842 409935 291898 409944
rect 291856 409086 291884 409935
rect 291844 409080 291896 409086
rect 291844 409022 291896 409028
rect 291106 389464 291162 389473
rect 291106 389399 291162 389408
rect 289728 388068 289780 388074
rect 289728 388010 289780 388016
rect 289740 367062 289768 388010
rect 291120 385665 291148 389399
rect 291856 388074 291884 409022
rect 291948 408746 291976 422266
rect 293972 410009 294000 426255
rect 296548 418130 296576 428742
rect 299308 425202 299336 429150
rect 309140 428936 309192 428942
rect 309336 428890 309364 430199
rect 309192 428884 309364 428890
rect 309140 428878 309364 428884
rect 309152 428862 309364 428878
rect 302792 428825 302844 428831
rect 302792 428767 302844 428773
rect 306196 428825 306248 428831
rect 306196 428767 306248 428773
rect 302804 425202 302832 428767
rect 306208 425610 306236 428767
rect 309152 426306 309180 428862
rect 309060 426278 309180 426306
rect 306196 425604 306248 425610
rect 306196 425546 306248 425552
rect 299296 425196 299348 425202
rect 299296 425138 299348 425144
rect 302792 425196 302844 425202
rect 302792 425138 302844 425144
rect 301502 422920 301558 422929
rect 301502 422855 301558 422864
rect 296536 418124 296588 418130
rect 296536 418066 296588 418072
rect 301516 410145 301544 422855
rect 304814 411360 304870 411369
rect 304814 411295 304870 411304
rect 301502 410136 301558 410145
rect 301502 410071 301558 410080
rect 293958 410000 294014 410009
rect 293958 409935 294014 409944
rect 301516 409465 301544 410071
rect 304828 409465 304856 411295
rect 301502 409456 301558 409465
rect 301502 409391 301558 409400
rect 304814 409456 304870 409465
rect 304814 409391 304870 409400
rect 301410 409184 301466 409193
rect 301410 409119 301466 409128
rect 304722 409184 304778 409193
rect 304722 409119 304778 409128
rect 301424 409034 301452 409119
rect 304736 409034 304764 409119
rect 301419 409006 301452 409034
rect 304684 409006 304764 409034
rect 301419 408748 301447 409006
rect 304684 408748 304712 409006
rect 291936 408740 291988 408746
rect 291936 408682 291988 408688
rect 291948 389201 291976 408682
rect 298928 408264 298980 408270
rect 298928 408206 298980 408212
rect 295708 407825 295760 407831
rect 295708 407767 295760 407773
rect 295720 405686 295748 407767
rect 295708 405680 295760 405686
rect 295708 405622 295760 405628
rect 298940 404666 298968 408206
rect 309060 408202 309088 426278
rect 309796 412634 309824 431926
rect 309888 422929 309916 431967
rect 309874 422920 309930 422929
rect 309874 422855 309930 422864
rect 309152 412606 309824 412634
rect 309152 411369 309180 412606
rect 309138 411360 309194 411369
rect 309138 411295 309194 411304
rect 305644 408196 305696 408202
rect 305644 408138 305696 408144
rect 309048 408196 309100 408202
rect 309048 408138 309100 408144
rect 302240 407825 302292 407831
rect 302240 407767 302292 407773
rect 302252 405618 302280 407767
rect 305656 405618 305684 408138
rect 302240 405612 302292 405618
rect 302240 405554 302292 405560
rect 305644 405612 305696 405618
rect 305644 405554 305696 405560
rect 298928 404660 298980 404666
rect 298928 404602 298980 404608
rect 302238 389464 302294 389473
rect 302238 389399 302294 389408
rect 291934 389192 291990 389201
rect 291934 389127 291990 389136
rect 298834 389192 298890 389201
rect 298834 389127 298890 389136
rect 291844 388068 291896 388074
rect 291844 388010 291896 388016
rect 291106 385656 291162 385665
rect 291106 385591 291162 385600
rect 291856 373994 291884 388010
rect 291948 381585 291976 389127
rect 298848 388521 298876 389127
rect 302252 388521 302280 389399
rect 309060 388521 309088 408138
rect 309152 389337 309180 411295
rect 311440 407788 311492 407794
rect 311440 407730 311492 407736
rect 311256 404388 311308 404394
rect 311256 404330 311308 404336
rect 311164 403028 311216 403034
rect 311164 402970 311216 402976
rect 309138 389328 309194 389337
rect 309138 389263 309194 389272
rect 298834 388512 298890 388521
rect 298834 388447 298890 388456
rect 302238 388512 302294 388521
rect 302238 388447 302294 388456
rect 309046 388512 309102 388521
rect 309046 388447 309102 388456
rect 299018 388240 299074 388249
rect 299018 388175 299074 388184
rect 302238 388240 302294 388249
rect 302238 388175 302294 388184
rect 309046 388240 309102 388249
rect 309046 388175 309102 388184
rect 299032 387804 299060 388175
rect 302252 387838 302280 388175
rect 309060 388074 309088 388175
rect 309048 388068 309100 388074
rect 309048 388010 309100 388016
rect 302240 387832 302292 387838
rect 302240 387774 302292 387780
rect 303620 387252 303672 387258
rect 303620 387194 303672 387200
rect 296168 386825 296220 386831
rect 296168 386767 296220 386773
rect 299848 386825 299900 386831
rect 299848 386767 299900 386773
rect 296180 385014 296208 386767
rect 299478 385656 299534 385665
rect 299478 385591 299534 385600
rect 296168 385008 296220 385014
rect 296168 384950 296220 384956
rect 291934 381576 291990 381585
rect 291934 381511 291990 381520
rect 296718 381576 296774 381585
rect 296718 381511 296774 381520
rect 291764 373966 291884 373994
rect 291764 371385 291792 373966
rect 291750 371376 291806 371385
rect 291750 371311 291806 371320
rect 293958 371376 294014 371385
rect 293958 371311 294014 371320
rect 291934 368520 291990 368529
rect 291934 368455 291990 368464
rect 291750 367160 291806 367169
rect 291750 367095 291806 367104
rect 289728 367056 289780 367062
rect 289728 366998 289780 367004
rect 289740 346050 289768 366998
rect 291764 346118 291792 367095
rect 291948 348401 291976 368455
rect 293972 367441 294000 371311
rect 296732 367441 296760 381511
rect 299492 368529 299520 385591
rect 299860 384946 299888 386767
rect 303632 384946 303660 387194
rect 307300 386825 307352 386831
rect 307300 386767 307352 386773
rect 299848 384940 299900 384946
rect 299848 384882 299900 384888
rect 300768 384940 300820 384946
rect 300768 384882 300820 384888
rect 303620 384940 303672 384946
rect 303620 384882 303672 384888
rect 300780 375358 300808 384882
rect 307312 384062 307340 386767
rect 308404 384940 308456 384946
rect 308404 384882 308456 384888
rect 307300 384056 307352 384062
rect 307300 383998 307352 384004
rect 300768 375352 300820 375358
rect 300768 375294 300820 375300
rect 304078 369744 304134 369753
rect 304078 369679 304134 369688
rect 299478 368520 299534 368529
rect 299478 368455 299534 368464
rect 300122 368520 300178 368529
rect 300122 368455 300178 368464
rect 300136 367441 300164 368455
rect 304092 367441 304120 369679
rect 308034 368520 308090 368529
rect 308034 368455 308090 368464
rect 293958 367432 294014 367441
rect 293958 367367 294014 367376
rect 296718 367432 296774 367441
rect 296718 367367 296774 367376
rect 300122 367432 300178 367441
rect 300122 367367 300178 367376
rect 304078 367432 304134 367441
rect 304078 367367 304134 367376
rect 294050 367160 294106 367169
rect 294050 367095 294106 367104
rect 297362 367160 297418 367169
rect 297362 367095 297418 367104
rect 300214 367160 300270 367169
rect 303986 367160 304042 367169
rect 300214 367095 300270 367104
rect 303816 367118 303986 367146
rect 294064 366838 294092 367095
rect 294052 366832 294104 366838
rect 294052 366774 294104 366780
rect 297376 366738 297404 367095
rect 300228 366838 300256 367095
rect 300216 366832 300268 366838
rect 300216 366774 300268 366780
rect 303816 366738 303844 367118
rect 303986 367095 304042 367104
rect 308048 366858 308076 368455
rect 307668 366852 307720 366858
rect 307668 366794 307720 366800
rect 308036 366852 308088 366858
rect 308036 366794 308088 366800
rect 297376 366724 297742 366738
rect 297376 366710 297756 366724
rect 295524 366240 295576 366246
rect 295524 366182 295576 366188
rect 295536 364342 295564 366182
rect 297728 366058 297756 366710
rect 297652 366030 297756 366058
rect 303816 366710 303846 366738
rect 295524 364336 295576 364342
rect 295524 364278 295576 364284
rect 297652 360233 297680 366030
rect 298560 365825 298612 365831
rect 298560 365767 298612 365773
rect 301596 365825 301648 365831
rect 301596 365767 301648 365773
rect 298572 364274 298600 365767
rect 298560 364268 298612 364274
rect 298560 364210 298612 364216
rect 301608 364206 301636 365767
rect 301596 364200 301648 364206
rect 301596 364142 301648 364148
rect 303816 361593 303844 366710
rect 304632 365825 304684 365831
rect 304632 365767 304684 365773
rect 307680 365786 307708 366794
rect 304644 363390 304672 365767
rect 307680 365758 307800 365786
rect 307772 364290 307800 365758
rect 307680 364262 307800 364290
rect 304632 363384 304684 363390
rect 304632 363326 304684 363332
rect 303802 361584 303858 361593
rect 303802 361519 303858 361528
rect 304906 361584 304962 361593
rect 304906 361519 304962 361528
rect 296718 360224 296774 360233
rect 296718 360159 296774 360168
rect 297638 360224 297694 360233
rect 297638 360159 297694 360168
rect 291934 348392 291990 348401
rect 291934 348327 291990 348336
rect 296732 346633 296760 360159
rect 299570 348392 299626 348401
rect 299570 348327 299626 348336
rect 299584 347857 299612 348327
rect 299570 347848 299626 347857
rect 299570 347783 299626 347792
rect 291842 346624 291898 346633
rect 291842 346559 291898 346568
rect 296718 346624 296774 346633
rect 296718 346559 296774 346568
rect 291752 346112 291804 346118
rect 291752 346054 291804 346060
rect 289728 346044 289780 346050
rect 289728 345986 289780 345992
rect 289740 324834 289768 345986
rect 289728 324828 289780 324834
rect 289728 324770 289780 324776
rect 289740 303822 289768 324770
rect 291856 324698 291884 346559
rect 299584 346458 299612 347783
rect 304920 346497 304948 361519
rect 304906 346488 304962 346497
rect 299572 346452 299624 346458
rect 307680 346474 307708 364262
rect 308034 347848 308090 347857
rect 308034 347783 308090 347792
rect 307942 346488 307998 346497
rect 307680 346446 307892 346474
rect 304906 346423 304962 346432
rect 299572 346394 299624 346400
rect 297270 346216 297326 346225
rect 303986 346216 304042 346225
rect 297326 346174 297404 346202
rect 297270 346151 297326 346160
rect 294420 346044 294472 346050
rect 294420 345986 294472 345992
rect 294432 345386 294460 345986
rect 297376 345794 297404 346174
rect 303908 346174 303986 346202
rect 303908 346066 303936 346174
rect 303986 346151 304042 346160
rect 303830 346038 303936 346066
rect 297376 345766 297740 345794
rect 303830 345780 303858 346038
rect 307864 345846 307892 346446
rect 307942 346423 307998 346432
rect 307852 345840 307904 345846
rect 307852 345782 307904 345788
rect 307864 345386 307892 345782
rect 294432 345372 294688 345386
rect 294432 345358 294702 345372
rect 294674 345014 294702 345358
rect 307772 345358 307892 345386
rect 295524 345228 295576 345234
rect 295524 345170 295576 345176
rect 294674 344986 294828 345014
rect 294800 325446 294828 344986
rect 295536 342242 295564 345170
rect 298560 344825 298612 344831
rect 298560 344767 298612 344773
rect 302148 344820 302200 344826
rect 295524 342236 295576 342242
rect 295524 342178 295576 342184
rect 298572 342174 298600 344767
rect 302148 344762 302200 344768
rect 304632 344825 304684 344831
rect 304632 344767 304684 344773
rect 298560 342168 298612 342174
rect 298560 342110 298612 342116
rect 302160 332586 302188 344762
rect 304644 341358 304672 344767
rect 304632 341352 304684 341358
rect 304632 341294 304684 341300
rect 307772 340898 307800 345358
rect 307956 345014 307984 346423
rect 307680 340870 307800 340898
rect 307864 344986 307984 345014
rect 302148 332580 302200 332586
rect 302148 332522 302200 332528
rect 307680 325825 307708 340870
rect 307666 325816 307722 325825
rect 307666 325751 307722 325760
rect 307864 325446 307892 344986
rect 308048 335354 308076 347783
rect 307956 335326 308076 335354
rect 307956 331214 307984 335326
rect 308416 335306 308444 384882
rect 308496 364200 308548 364206
rect 308496 364142 308548 364148
rect 308404 335300 308456 335306
rect 308404 335242 308456 335248
rect 308508 333946 308536 364142
rect 309784 341284 309836 341290
rect 309784 341226 309836 341232
rect 308496 333940 308548 333946
rect 308496 333882 308548 333888
rect 307956 331186 308444 331214
rect 294788 325440 294840 325446
rect 294788 325382 294840 325388
rect 307852 325440 307904 325446
rect 307852 325382 307904 325388
rect 294788 325236 294840 325242
rect 294788 325178 294840 325184
rect 291844 324692 291896 324698
rect 291844 324634 291896 324640
rect 291856 306374 291884 324634
rect 294800 324202 294828 325178
rect 308416 324970 308444 331186
rect 308586 325816 308642 325825
rect 308586 325751 308642 325760
rect 309598 325816 309654 325825
rect 309598 325751 309654 325760
rect 308496 325440 308548 325446
rect 308496 325382 308548 325388
rect 308404 324964 308456 324970
rect 308404 324906 308456 324912
rect 296996 324832 297048 324838
rect 296996 324774 297048 324780
rect 297008 324698 297036 324774
rect 296996 324692 297048 324698
rect 296996 324634 297048 324640
rect 294788 324196 294840 324202
rect 294788 324138 294840 324144
rect 292396 323944 292448 323950
rect 292396 323886 292448 323892
rect 291856 306346 291976 306374
rect 291948 305153 291976 306346
rect 291934 305144 291990 305153
rect 291934 305079 291990 305088
rect 289728 303816 289780 303822
rect 289728 303758 289780 303764
rect 289740 282674 289768 303758
rect 291842 283520 291898 283529
rect 291842 283455 291898 283464
rect 291856 282946 291884 283455
rect 291844 282940 291896 282946
rect 291844 282882 291896 282888
rect 289728 282668 289780 282674
rect 289728 282610 289780 282616
rect 289740 261866 289768 282610
rect 291856 262070 291884 282882
rect 291948 282674 291976 305079
rect 292408 305017 292436 323886
rect 295616 323825 295668 323831
rect 295616 323767 295668 323773
rect 298744 323825 298796 323831
rect 298744 323767 298796 323773
rect 305092 323825 305144 323831
rect 305092 323767 305144 323773
rect 295628 321570 295656 323767
rect 295616 321564 295668 321570
rect 295616 321506 295668 321512
rect 298756 321502 298784 323767
rect 301964 323740 302016 323746
rect 301964 323682 302016 323688
rect 298744 321496 298796 321502
rect 298744 321438 298796 321444
rect 301976 321434 302004 323682
rect 301964 321428 302016 321434
rect 301964 321370 302016 321376
rect 305104 318102 305132 323767
rect 305092 318096 305144 318102
rect 305092 318038 305144 318044
rect 306010 305824 306066 305833
rect 306010 305759 306066 305768
rect 302422 305688 302478 305697
rect 302422 305623 302478 305632
rect 298466 305144 298522 305153
rect 298466 305079 298522 305088
rect 292394 305008 292450 305017
rect 292394 304943 292450 304952
rect 294970 305008 295026 305017
rect 294970 304943 295026 304952
rect 294984 304434 295012 304943
rect 298480 304434 298508 305079
rect 302436 304434 302464 305623
rect 306024 304434 306052 305759
rect 308416 305697 308444 324906
rect 308508 324290 308536 325382
rect 308600 324834 308628 325751
rect 308588 324828 308640 324834
rect 308588 324770 308640 324776
rect 308496 324284 308548 324290
rect 308496 324226 308548 324232
rect 308508 305833 308536 324226
rect 308494 305824 308550 305833
rect 308494 305759 308550 305768
rect 308402 305688 308458 305697
rect 308402 305623 308458 305632
rect 308416 305017 308444 305623
rect 308508 305153 308536 305759
rect 308494 305144 308550 305153
rect 308494 305079 308550 305088
rect 308402 305008 308458 305017
rect 308402 304943 308458 304952
rect 309612 304434 309640 325751
rect 309796 304434 309824 341226
rect 310518 305008 310574 305017
rect 310518 304943 310574 304952
rect 294972 304428 295024 304434
rect 294972 304370 295024 304376
rect 298468 304428 298520 304434
rect 298468 304370 298520 304376
rect 302424 304428 302476 304434
rect 302424 304370 302476 304376
rect 306012 304428 306064 304434
rect 306012 304370 306064 304376
rect 309600 304428 309652 304434
rect 309600 304370 309652 304376
rect 309784 304428 309836 304434
rect 309784 304370 309836 304376
rect 294972 304224 295024 304230
rect 294972 304166 295024 304172
rect 298468 304224 298520 304230
rect 298468 304166 298520 304172
rect 302424 304224 302476 304230
rect 302424 304166 302476 304172
rect 306012 304224 306064 304230
rect 306012 304166 306064 304172
rect 309600 304224 309652 304230
rect 309600 304166 309652 304172
rect 294984 303770 295012 304166
rect 298480 303770 298508 304166
rect 302436 304042 302464 304166
rect 306024 304042 306052 304166
rect 302406 304014 302464 304042
rect 305991 304014 306052 304042
rect 294984 303756 295250 303770
rect 294984 303742 295264 303756
rect 298480 303742 298835 303770
rect 302406 303756 302434 304014
rect 305991 303756 306019 304014
rect 309612 303906 309640 304166
rect 309576 303878 309640 303906
rect 295236 303090 295264 303742
rect 309576 303090 309604 303878
rect 295236 303062 295288 303090
rect 309576 303062 309640 303090
rect 295260 283529 295288 303062
rect 296076 302825 296128 302831
rect 296076 302767 296128 302773
rect 299664 302825 299716 302831
rect 299664 302767 299716 302773
rect 306840 302825 306892 302831
rect 306840 302767 306892 302773
rect 296088 300830 296116 302767
rect 296076 300824 296128 300830
rect 296076 300766 296128 300772
rect 299676 300762 299704 302767
rect 299664 300756 299716 300762
rect 299664 300698 299716 300704
rect 306852 299810 306880 302767
rect 308678 302288 308734 302297
rect 308678 302223 308734 302232
rect 309506 302288 309562 302297
rect 309612 302274 309640 303062
rect 309562 302246 309640 302274
rect 309506 302223 309562 302232
rect 306840 299804 306892 299810
rect 306840 299746 306892 299752
rect 307668 299804 307720 299810
rect 307668 299746 307720 299752
rect 307680 289814 307708 299746
rect 307668 289808 307720 289814
rect 307668 289750 307720 289756
rect 304906 284472 304962 284481
rect 304906 284407 304962 284416
rect 301686 284336 301742 284345
rect 301686 284271 301742 284280
rect 301700 283529 301728 284271
rect 304920 283529 304948 284407
rect 295246 283520 295302 283529
rect 295246 283455 295302 283464
rect 301686 283520 301742 283529
rect 301686 283455 301742 283464
rect 304906 283520 304962 283529
rect 308692 283506 308720 302223
rect 309138 285696 309194 285705
rect 309138 285631 309194 285640
rect 309152 284481 309180 285631
rect 309138 284472 309194 284481
rect 309194 284430 309456 284458
rect 309138 284407 309194 284416
rect 309322 284336 309378 284345
rect 309322 284271 309378 284280
rect 308692 283478 309272 283506
rect 304906 283455 304962 283464
rect 301591 283112 301647 283121
rect 301591 283047 301647 283056
rect 304908 283112 304964 283121
rect 304908 283047 304964 283056
rect 309244 282962 309272 283478
rect 309152 282934 309272 282962
rect 291936 282668 291988 282674
rect 291936 282610 291988 282616
rect 291844 262064 291896 262070
rect 291844 262006 291896 262012
rect 289728 261860 289780 261866
rect 289728 261802 289780 261808
rect 289740 241058 289768 261802
rect 291856 241058 291884 262006
rect 291948 261730 291976 282610
rect 309152 282198 309180 282934
rect 309336 282826 309364 284271
rect 309244 282798 309364 282826
rect 309140 282192 309192 282198
rect 309140 282134 309192 282140
rect 295800 281825 295852 281831
rect 295800 281767 295852 281773
rect 299112 281825 299164 281831
rect 299112 281767 299164 281773
rect 302424 281825 302476 281831
rect 302424 281767 302476 281773
rect 305736 281825 305788 281831
rect 305736 281767 305788 281773
rect 295812 280158 295840 281767
rect 299124 280158 299152 281767
rect 295800 280152 295852 280158
rect 295800 280094 295852 280100
rect 299112 280152 299164 280158
rect 299112 280094 299164 280100
rect 302436 280022 302464 281767
rect 305748 280158 305776 281767
rect 305736 280152 305788 280158
rect 309152 280106 309180 282134
rect 305736 280094 305788 280100
rect 309060 280078 309180 280106
rect 302424 280016 302476 280022
rect 302424 279958 302476 279964
rect 305918 263800 305974 263809
rect 305918 263735 305974 263744
rect 302146 263664 302202 263673
rect 302146 263599 302202 263608
rect 302160 262585 302188 263599
rect 305932 262585 305960 263735
rect 309060 262585 309088 280078
rect 309244 263673 309272 282798
rect 309428 277394 309456 284430
rect 310532 284345 310560 304943
rect 310518 284336 310574 284345
rect 310518 284271 310574 284280
rect 309336 277366 309456 277394
rect 309336 263809 309364 277366
rect 309322 263800 309378 263809
rect 309322 263735 309378 263744
rect 309230 263664 309286 263673
rect 309230 263599 309286 263608
rect 309336 262585 309364 263735
rect 309874 263664 309930 263673
rect 309874 263599 309930 263608
rect 302146 262576 302202 262585
rect 302146 262511 302202 262520
rect 305918 262576 305974 262585
rect 305918 262511 305974 262520
rect 309046 262576 309102 262585
rect 309046 262511 309102 262520
rect 309322 262576 309378 262585
rect 309322 262511 309378 262520
rect 309322 262168 309378 262177
rect 301933 262112 301942 262168
rect 301998 262112 302007 262168
rect 305377 262112 305386 262168
rect 305442 262112 305451 262168
rect 309322 262103 309378 262112
rect 308830 262032 308886 262041
rect 308830 261967 308886 261976
rect 291936 261724 291988 261730
rect 291936 261666 291988 261672
rect 289728 241052 289780 241058
rect 289728 240994 289780 241000
rect 291844 241052 291896 241058
rect 291844 240994 291896 241000
rect 289740 220046 289768 240994
rect 289728 220040 289780 220046
rect 289728 219982 289780 219988
rect 289740 206310 289768 219982
rect 291856 218521 291884 240994
rect 291948 240718 291976 261666
rect 299296 261248 299348 261254
rect 299296 261190 299348 261196
rect 295892 260825 295944 260831
rect 295892 260767 295944 260773
rect 295904 257990 295932 260767
rect 299308 258074 299336 261190
rect 308864 260908 308916 260914
rect 308864 260850 308916 260856
rect 302792 260825 302844 260831
rect 302792 260767 302844 260773
rect 306196 260825 306248 260831
rect 306196 260767 306248 260773
rect 302804 259350 302832 260767
rect 302792 259344 302844 259350
rect 302792 259286 302844 259292
rect 299216 258046 299336 258074
rect 306208 258058 306236 260767
rect 306196 258052 306248 258058
rect 295892 257984 295944 257990
rect 295892 257926 295944 257932
rect 299216 257922 299244 258046
rect 306196 257994 306248 258000
rect 299204 257916 299256 257922
rect 299204 257858 299256 257864
rect 304906 250472 304962 250481
rect 304906 250407 304962 250416
rect 304920 248414 304948 250407
rect 304828 248386 304948 248414
rect 301502 242992 301558 243001
rect 301502 242927 301558 242936
rect 301516 241505 301544 242927
rect 304828 241505 304856 248386
rect 301502 241496 301558 241505
rect 301502 241431 301558 241440
rect 304814 241496 304870 241505
rect 304814 241431 304870 241440
rect 301410 241224 301466 241233
rect 301410 241159 301466 241168
rect 304722 241224 304778 241233
rect 304722 241159 304778 241168
rect 301424 240788 301452 241159
rect 304736 241074 304764 241159
rect 304683 241046 304764 241074
rect 304683 240788 304711 241046
rect 308876 240854 308904 260850
rect 309336 253934 309364 262103
rect 309244 253906 309364 253934
rect 309244 250481 309272 253906
rect 309230 250472 309286 250481
rect 309230 250407 309286 250416
rect 309138 242992 309194 243001
rect 309138 242927 309194 242936
rect 307944 240848 307996 240854
rect 307944 240790 307996 240796
rect 308864 240848 308916 240854
rect 308864 240790 308916 240796
rect 291936 240712 291988 240718
rect 291936 240654 291988 240660
rect 291948 219706 291976 240654
rect 298928 240236 298980 240242
rect 298928 240178 298980 240184
rect 305460 240236 305512 240242
rect 305460 240178 305512 240184
rect 295708 239825 295760 239831
rect 295708 239767 295760 239773
rect 295720 237386 295748 239767
rect 298940 238754 298968 240178
rect 302240 239825 302292 239831
rect 302240 239767 302292 239773
rect 298940 238746 299060 238754
rect 298940 238740 299072 238746
rect 298940 238726 299020 238740
rect 299020 238682 299072 238688
rect 302252 237386 302280 239767
rect 305472 238754 305500 240178
rect 305472 238726 305592 238754
rect 295708 237380 295760 237386
rect 295708 237322 295760 237328
rect 302240 237380 302292 237386
rect 302240 237322 302292 237328
rect 305564 237318 305592 238726
rect 305552 237312 305604 237318
rect 305552 237254 305604 237260
rect 306838 223544 306894 223553
rect 306838 223479 306894 223488
rect 302790 222864 302846 222873
rect 302790 222799 302846 222808
rect 302804 220425 302832 222799
rect 306852 220425 306880 223479
rect 307956 222737 307984 240790
rect 309152 222873 309180 242927
rect 309244 223553 309272 250407
rect 309888 243001 309916 263599
rect 309874 242992 309930 243001
rect 309874 242927 309930 242936
rect 309230 223544 309286 223553
rect 309230 223479 309286 223488
rect 309138 222864 309194 222873
rect 309138 222799 309194 222808
rect 307942 222728 307998 222737
rect 307942 222663 307998 222672
rect 309690 222728 309746 222737
rect 309690 222663 309746 222672
rect 309704 220425 309732 222663
rect 302790 220416 302846 220425
rect 302790 220351 302846 220360
rect 306838 220416 306894 220425
rect 306838 220351 306894 220360
rect 309690 220416 309746 220425
rect 309690 220351 309746 220360
rect 306746 220144 306802 220153
rect 306484 220102 306746 220130
rect 302745 220008 302801 220017
rect 302745 219943 302801 219952
rect 302759 219708 302787 219943
rect 291936 219700 291988 219706
rect 291936 219642 291988 219648
rect 291842 218512 291898 218521
rect 291842 218447 291898 218456
rect 291948 209774 291976 219642
rect 306484 219178 306512 220102
rect 306746 220079 306802 220088
rect 309782 220144 309838 220153
rect 309838 220102 309916 220130
rect 309782 220079 309838 220088
rect 309888 219722 309916 220102
rect 309888 219708 310197 219722
rect 309888 219694 310211 219708
rect 310183 219178 310211 219694
rect 294708 219150 295349 219178
rect 306392 219164 306512 219178
rect 310178 219164 310211 219178
rect 306392 219150 306498 219164
rect 310164 219150 310197 219164
rect 294708 218521 294736 219150
rect 296168 218825 296220 218831
rect 296168 218767 296220 218773
rect 299848 218825 299900 218831
rect 299848 218767 299900 218773
rect 294694 218512 294750 218521
rect 294694 218447 294750 218456
rect 291764 209746 291976 209774
rect 289728 206304 289780 206310
rect 289728 206246 289780 206252
rect 289740 198830 289768 206246
rect 291764 200161 291792 209746
rect 291842 200288 291898 200297
rect 291842 200223 291898 200232
rect 291750 200152 291806 200161
rect 291750 200087 291806 200096
rect 289728 198824 289780 198830
rect 289728 198766 289780 198772
rect 289740 178022 289768 198766
rect 291764 180305 291792 200087
rect 291750 180296 291806 180305
rect 291750 180231 291806 180240
rect 291856 180033 291884 200223
rect 294708 199481 294736 218447
rect 296180 216646 296208 218767
rect 296168 216640 296220 216646
rect 296168 216582 296220 216588
rect 299860 216442 299888 218767
rect 303620 218748 303672 218754
rect 303620 218690 303672 218696
rect 303632 216646 303660 218690
rect 306392 217841 306420 219150
rect 307300 218825 307352 218831
rect 307300 218767 307352 218773
rect 304906 217832 304962 217841
rect 304906 217767 304962 217776
rect 306378 217832 306434 217841
rect 306378 217767 306434 217776
rect 306930 217832 306986 217841
rect 306930 217767 306986 217776
rect 303620 216640 303672 216646
rect 303620 216582 303672 216588
rect 299848 216436 299900 216442
rect 299848 216378 299900 216384
rect 300766 200696 300822 200705
rect 300766 200631 300822 200640
rect 300780 200297 300808 200631
rect 300766 200288 300822 200297
rect 300766 200223 300822 200232
rect 297546 200152 297602 200161
rect 297546 200087 297602 200096
rect 294694 199472 294750 199481
rect 297560 199442 297588 200087
rect 300780 199442 300808 200223
rect 304920 200114 304948 217767
rect 304828 200086 304948 200114
rect 304828 199442 304856 200086
rect 306944 199481 306972 217767
rect 307312 216646 307340 218767
rect 310164 217841 310192 219150
rect 310150 217832 310206 217841
rect 310150 217767 310206 217776
rect 307300 216640 307352 216646
rect 307300 216582 307352 216588
rect 311176 216510 311204 402970
rect 311268 237250 311296 404330
rect 311346 388240 311402 388249
rect 311346 388175 311402 388184
rect 311360 368529 311388 388175
rect 311346 368520 311402 368529
rect 311346 368455 311402 368464
rect 311348 361616 311400 361622
rect 311348 361558 311400 361564
rect 311256 237244 311308 237250
rect 311256 237186 311308 237192
rect 311164 216504 311216 216510
rect 311164 216446 311216 216452
rect 306930 199472 306986 199481
rect 294694 199407 294750 199416
rect 297548 199436 297600 199442
rect 297548 199378 297600 199384
rect 300768 199436 300820 199442
rect 300768 199378 300820 199384
rect 304816 199436 304868 199442
rect 306930 199407 306986 199416
rect 304816 199378 304868 199384
rect 297548 199232 297600 199238
rect 297548 199174 297600 199180
rect 300768 199232 300820 199238
rect 300768 199174 300820 199180
rect 307574 199200 307630 199209
rect 293684 198832 293736 198838
rect 292486 198792 292542 198801
rect 292486 198727 292542 198736
rect 293682 198792 293684 198801
rect 293736 198792 293738 198801
rect 297560 198778 297588 199174
rect 300780 199050 300808 199174
rect 307574 199135 307630 199144
rect 300779 199022 300808 199050
rect 297560 198750 297741 198778
rect 300779 198764 300807 199022
rect 304816 198892 304868 198898
rect 304816 198834 304868 198840
rect 293682 198727 293738 198736
rect 291842 180024 291898 180033
rect 291842 179959 291898 179968
rect 292500 179489 292528 198727
rect 295524 198212 295576 198218
rect 295524 198154 295576 198160
rect 295536 195974 295564 198154
rect 303831 197962 303859 198220
rect 303831 197934 303936 197962
rect 298560 197825 298612 197831
rect 298560 197767 298612 197773
rect 295524 195968 295576 195974
rect 295524 195910 295576 195916
rect 298572 195838 298600 197767
rect 303908 197418 303936 197934
rect 304632 197825 304684 197831
rect 304632 197767 304684 197773
rect 303986 197432 304042 197441
rect 303908 197390 303986 197418
rect 303986 197367 304042 197376
rect 304644 195974 304672 197767
rect 304828 197441 304856 198834
rect 307588 198218 307616 199135
rect 307576 198212 307628 198218
rect 307576 198154 307628 198160
rect 307588 198098 307616 198154
rect 307588 198070 307800 198098
rect 304814 197432 304870 197441
rect 304814 197367 304870 197376
rect 304632 195968 304684 195974
rect 304632 195910 304684 195916
rect 298560 195832 298612 195838
rect 298560 195774 298612 195780
rect 304828 180794 304856 197367
rect 304552 180766 304856 180794
rect 296718 180296 296774 180305
rect 296718 180231 296774 180240
rect 298006 180296 298062 180305
rect 298006 180231 298062 180240
rect 292486 179480 292542 179489
rect 292486 179415 292542 179424
rect 293958 179480 294014 179489
rect 293958 179415 294014 179424
rect 293972 178634 294000 179415
rect 296732 178702 296760 180231
rect 298020 179625 298048 180231
rect 304552 179897 304580 180766
rect 307772 180033 307800 198070
rect 311360 195838 311388 361558
rect 311452 256698 311480 407730
rect 311532 405748 311584 405754
rect 311532 405690 311584 405696
rect 311544 257990 311572 405690
rect 311898 389328 311954 389337
rect 311898 389263 311954 389272
rect 311912 387734 311940 389263
rect 311900 387728 311952 387734
rect 311900 387670 311952 387676
rect 311912 369753 311940 387670
rect 311898 369744 311954 369753
rect 311898 369679 311954 369688
rect 311624 362976 311676 362982
rect 311624 362918 311676 362924
rect 311532 257984 311584 257990
rect 311532 257926 311584 257932
rect 311440 256692 311492 256698
rect 311440 256634 311492 256640
rect 311636 216442 311664 362918
rect 311716 323536 311768 323542
rect 311716 323478 311768 323484
rect 311728 251190 311756 323478
rect 311898 305144 311954 305153
rect 311898 305079 311954 305088
rect 311912 285705 311940 305079
rect 311898 285696 311954 285705
rect 311898 285631 311954 285640
rect 312556 260846 312584 471174
rect 312636 401668 312688 401674
rect 312636 401610 312688 401616
rect 312544 260840 312596 260846
rect 312544 260782 312596 260788
rect 311716 251184 311768 251190
rect 311716 251126 311768 251132
rect 311898 222864 311954 222873
rect 311898 222799 311954 222808
rect 311624 216436 311676 216442
rect 311624 216378 311676 216384
rect 311912 200705 311940 222799
rect 311898 200696 311954 200705
rect 311898 200631 311954 200640
rect 312648 195906 312676 401610
rect 312740 302938 312768 488990
rect 312912 488708 312964 488714
rect 312912 488650 312964 488656
rect 312820 428800 312872 428806
rect 312820 428742 312872 428748
rect 312728 302932 312780 302938
rect 312728 302874 312780 302880
rect 312728 261248 312780 261254
rect 312728 261190 312780 261196
rect 312740 247042 312768 261190
rect 312832 257990 312860 428742
rect 312924 342106 312952 488650
rect 313004 407176 313056 407182
rect 313004 407118 313056 407124
rect 312912 342100 312964 342106
rect 312912 342042 312964 342048
rect 312912 303204 312964 303210
rect 312912 303146 312964 303152
rect 312820 257984 312872 257990
rect 312820 257926 312872 257932
rect 312924 249762 312952 303146
rect 313016 279954 313044 407118
rect 313188 405544 313240 405550
rect 313188 405486 313240 405492
rect 313096 365764 313148 365770
rect 313096 365706 313148 365712
rect 313004 279948 313056 279954
rect 313004 279890 313056 279896
rect 313108 257922 313136 365706
rect 313200 345710 313228 405486
rect 313188 345704 313240 345710
rect 313188 345646 313240 345652
rect 313188 344888 313240 344894
rect 313188 344830 313240 344836
rect 313096 257916 313148 257922
rect 313096 257858 313148 257864
rect 313200 252550 313228 344830
rect 313936 262206 313964 491438
rect 367744 488640 367796 488646
rect 367744 488582 367796 488588
rect 314108 469124 314160 469130
rect 314108 469066 314160 469072
rect 314016 449948 314068 449954
rect 314016 449890 314068 449896
rect 313924 262200 313976 262206
rect 313924 262142 313976 262148
rect 314028 259418 314056 449890
rect 314120 303142 314148 469066
rect 338764 468036 338816 468042
rect 338764 467978 338816 467984
rect 338776 451926 338804 467978
rect 363604 467968 363656 467974
rect 363604 467910 363656 467916
rect 338764 451920 338816 451926
rect 338764 451862 338816 451868
rect 314200 447704 314252 447710
rect 314200 447646 314252 447652
rect 314108 303136 314160 303142
rect 314108 303078 314160 303084
rect 314212 303006 314240 447646
rect 314384 425604 314436 425610
rect 314384 425546 314436 425552
rect 314292 386844 314344 386850
rect 314292 386786 314344 386792
rect 314200 303000 314252 303006
rect 314200 302942 314252 302948
rect 314016 259412 314068 259418
rect 314016 259354 314068 259360
rect 314304 255270 314332 386786
rect 314396 298110 314424 425546
rect 314476 405612 314528 405618
rect 314476 405554 314528 405560
rect 314384 298104 314436 298110
rect 314384 298046 314436 298052
rect 314488 296682 314516 405554
rect 359464 364404 359516 364410
rect 359464 364346 359516 364352
rect 314568 363384 314620 363390
rect 314568 363326 314620 363332
rect 314580 303074 314608 363326
rect 345664 320204 345716 320210
rect 345664 320146 345716 320152
rect 314568 303068 314620 303074
rect 314568 303010 314620 303016
rect 314476 296676 314528 296682
rect 314476 296618 314528 296624
rect 314292 255264 314344 255270
rect 314292 255206 314344 255212
rect 313188 252544 313240 252550
rect 313188 252486 313240 252492
rect 312912 249756 312964 249762
rect 312912 249698 312964 249704
rect 312728 247036 312780 247042
rect 312728 246978 312780 246984
rect 313924 242956 313976 242962
rect 313924 242898 313976 242904
rect 313936 219162 313964 242898
rect 313924 219156 313976 219162
rect 313924 219098 313976 219104
rect 312636 195900 312688 195906
rect 312636 195842 312688 195848
rect 311348 195832 311400 195838
rect 311348 195774 311400 195780
rect 306930 180024 306986 180033
rect 306930 179959 306986 179968
rect 307758 180024 307814 180033
rect 307758 179959 307814 179968
rect 304538 179888 304594 179897
rect 304538 179823 304594 179832
rect 300766 179752 300822 179761
rect 300766 179687 300822 179696
rect 298006 179616 298062 179625
rect 298006 179551 298062 179560
rect 296720 178696 296772 178702
rect 296720 178638 296772 178644
rect 300780 178634 300808 179687
rect 304552 178634 304580 179823
rect 306944 178634 306972 179959
rect 308770 179752 308826 179761
rect 308770 179687 308826 179696
rect 308586 179616 308642 179625
rect 308586 179551 308642 179560
rect 308402 179480 308458 179489
rect 308402 179415 308458 179424
rect 293960 178628 294012 178634
rect 293960 178570 294012 178576
rect 300768 178628 300820 178634
rect 300768 178570 300820 178576
rect 304540 178628 304592 178634
rect 304540 178570 304592 178576
rect 306932 178628 306984 178634
rect 306932 178570 306984 178576
rect 294052 178424 294104 178430
rect 294052 178366 294104 178372
rect 300768 178424 300820 178430
rect 300768 178366 300820 178372
rect 303804 178424 303856 178430
rect 303804 178366 303856 178372
rect 306840 178424 306892 178430
rect 306840 178366 306892 178372
rect 294064 178038 294092 178366
rect 300780 178242 300808 178366
rect 300778 178214 300808 178242
rect 303816 178242 303844 178366
rect 303816 178214 303858 178242
rect 294052 178032 294104 178038
rect 289728 178016 289780 178022
rect 294052 177974 294104 177980
rect 289728 177958 289780 177964
rect 300778 177956 300806 178214
rect 303830 177956 303858 178214
rect 306852 178106 306880 178366
rect 306852 178078 306910 178106
rect 306882 177956 306910 178078
rect 295524 177404 295576 177410
rect 295524 177346 295576 177352
rect 295536 175234 295564 177346
rect 298560 177025 298612 177031
rect 298560 176967 298612 176973
rect 301596 177025 301648 177031
rect 301596 176967 301648 176973
rect 304632 177025 304684 177031
rect 304632 176967 304684 176973
rect 295524 175228 295576 175234
rect 295524 175170 295576 175176
rect 298572 175166 298600 176967
rect 298560 175160 298612 175166
rect 298560 175102 298612 175108
rect 301608 175098 301636 176967
rect 304644 175098 304672 176967
rect 301596 175092 301648 175098
rect 301596 175034 301648 175040
rect 304632 175092 304684 175098
rect 304632 175034 304684 175040
rect 308416 6633 308444 179415
rect 308600 46345 308628 179551
rect 308784 86193 308812 179687
rect 345676 175030 345704 320146
rect 359476 238746 359504 364346
rect 363616 340882 363644 467910
rect 367756 382226 367784 488582
rect 405004 488572 405056 488578
rect 405004 488514 405056 488520
rect 388444 467900 388496 467906
rect 388444 467842 388496 467848
rect 370596 447296 370648 447302
rect 370596 447238 370648 447244
rect 367744 382220 367796 382226
rect 367744 382162 367796 382168
rect 370504 365832 370556 365838
rect 370504 365774 370556 365780
rect 363604 340876 363656 340882
rect 363604 340818 363656 340824
rect 363696 327140 363748 327146
rect 363696 327082 363748 327088
rect 363604 325712 363656 325718
rect 363604 325654 363656 325660
rect 362224 321632 362276 321638
rect 362224 321574 362276 321580
rect 359464 238740 359516 238746
rect 359464 238682 359516 238688
rect 362236 197334 362264 321574
rect 363616 259350 363644 325654
rect 363708 280022 363736 327082
rect 364984 322992 365036 322998
rect 364984 322934 365036 322940
rect 363696 280016 363748 280022
rect 363696 279958 363748 279964
rect 363604 259344 363656 259350
rect 363604 259286 363656 259292
rect 364996 216578 365024 322934
rect 366364 318096 366416 318102
rect 366364 318038 366416 318044
rect 366376 291174 366404 318038
rect 366364 291168 366416 291174
rect 366364 291110 366416 291116
rect 366364 284368 366416 284374
rect 366364 284310 366416 284316
rect 366376 237318 366404 284310
rect 370516 253910 370544 365774
rect 370608 339454 370636 447238
rect 388456 380866 388484 467842
rect 391204 425196 391256 425202
rect 391204 425138 391256 425144
rect 388444 380860 388496 380866
rect 388444 380802 388496 380808
rect 373264 367124 373316 367130
rect 373264 367066 373316 367072
rect 370596 339448 370648 339454
rect 370596 339390 370648 339396
rect 371884 281852 371936 281858
rect 371884 281794 371936 281800
rect 370504 253904 370556 253910
rect 370504 253846 370556 253852
rect 371896 248402 371924 281794
rect 373276 280090 373304 367066
rect 391216 338094 391244 425138
rect 405016 422278 405044 488514
rect 515404 451920 515456 451926
rect 515404 451862 515456 451868
rect 406384 447228 406436 447234
rect 406384 447170 406436 447176
rect 405004 422272 405056 422278
rect 405004 422214 405056 422220
rect 393964 383716 394016 383722
rect 393964 383658 394016 383664
rect 391204 338088 391256 338094
rect 391204 338030 391256 338036
rect 377404 324352 377456 324358
rect 377404 324294 377456 324300
rect 373264 280084 373316 280090
rect 373264 280026 373316 280032
rect 371884 248396 371936 248402
rect 371884 248338 371936 248344
rect 377416 237386 377444 324294
rect 393976 295322 394004 383658
rect 406396 379506 406424 447170
rect 443644 447160 443696 447166
rect 443644 447102 443696 447108
rect 427084 425128 427136 425134
rect 427084 425070 427136 425076
rect 406384 379500 406436 379506
rect 406384 379442 406436 379448
rect 427096 378146 427124 425070
rect 443656 419490 443684 447102
rect 514760 422272 514812 422278
rect 514760 422214 514812 422220
rect 514772 421025 514800 422214
rect 514758 421016 514814 421025
rect 514758 420951 514814 420960
rect 515416 419665 515444 451862
rect 518622 423872 518678 423881
rect 518622 423807 518678 423816
rect 521658 423872 521714 423881
rect 521658 423807 521714 423816
rect 517428 421388 517480 421394
rect 517428 421330 517480 421336
rect 515402 419656 515458 419665
rect 515402 419591 515458 419600
rect 443644 419484 443696 419490
rect 443644 419426 443696 419432
rect 514760 419484 514812 419490
rect 514760 419426 514812 419432
rect 514772 418305 514800 419426
rect 514758 418296 514814 418305
rect 514758 418231 514814 418240
rect 514760 418124 514812 418130
rect 514760 418066 514812 418072
rect 514772 416945 514800 418066
rect 514758 416936 514814 416945
rect 514758 416871 514814 416880
rect 515402 415576 515458 415585
rect 515402 415511 515458 415520
rect 514758 407416 514814 407425
rect 514758 407351 514814 407360
rect 514772 407182 514800 407351
rect 514760 407176 514812 407182
rect 514760 407118 514812 407124
rect 514758 406056 514814 406065
rect 514758 405991 514814 406000
rect 514772 405754 514800 405991
rect 514760 405748 514812 405754
rect 514760 405690 514812 405696
rect 515416 405686 515444 415511
rect 515862 414216 515918 414225
rect 515862 414151 515918 414160
rect 515494 412856 515550 412865
rect 515494 412791 515550 412800
rect 515404 405680 515456 405686
rect 515404 405622 515456 405628
rect 514758 404696 514814 404705
rect 514758 404631 514814 404640
rect 446404 404456 446456 404462
rect 446404 404398 446456 404404
rect 427084 378140 427136 378146
rect 427084 378082 427136 378088
rect 446416 376718 446444 404398
rect 514772 404394 514800 404631
rect 514760 404388 514812 404394
rect 514760 404330 514812 404336
rect 514758 403336 514814 403345
rect 514758 403271 514814 403280
rect 514772 403034 514800 403271
rect 514760 403028 514812 403034
rect 514760 402970 514812 402976
rect 514758 401976 514814 401985
rect 514758 401911 514814 401920
rect 514772 401674 514800 401911
rect 514760 401668 514812 401674
rect 514760 401610 514812 401616
rect 515402 400616 515458 400625
rect 515402 400551 515458 400560
rect 514760 382220 514812 382226
rect 514760 382162 514812 382168
rect 514772 381041 514800 382162
rect 514758 381032 514814 381041
rect 514758 380967 514814 380976
rect 514760 380860 514812 380866
rect 514760 380802 514812 380808
rect 514772 379681 514800 380802
rect 514758 379672 514814 379681
rect 514758 379607 514814 379616
rect 514760 379500 514812 379506
rect 514760 379442 514812 379448
rect 514772 378321 514800 379442
rect 514758 378312 514814 378321
rect 514758 378247 514814 378256
rect 514760 378140 514812 378146
rect 514760 378082 514812 378088
rect 514772 376961 514800 378082
rect 514758 376952 514814 376961
rect 514758 376887 514814 376896
rect 446404 376712 446456 376718
rect 446404 376654 446456 376660
rect 514760 376712 514812 376718
rect 514760 376654 514812 376660
rect 514772 375601 514800 376654
rect 514758 375592 514814 375601
rect 514758 375527 514814 375536
rect 514760 375352 514812 375358
rect 514760 375294 514812 375300
rect 514772 374241 514800 375294
rect 514758 374232 514814 374241
rect 514758 374167 514814 374176
rect 515310 372872 515366 372881
rect 515310 372807 515366 372816
rect 514758 367432 514814 367441
rect 514758 367367 514814 367376
rect 514772 367130 514800 367367
rect 514760 367124 514812 367130
rect 514760 367066 514812 367072
rect 514758 366072 514814 366081
rect 514758 366007 514814 366016
rect 514772 365770 514800 366007
rect 514760 365764 514812 365770
rect 514760 365706 514812 365712
rect 514758 364712 514814 364721
rect 514758 364647 514814 364656
rect 514772 364410 514800 364647
rect 514760 364404 514812 364410
rect 514760 364346 514812 364352
rect 515324 364274 515352 372807
rect 515312 364268 515364 364274
rect 515312 364210 515364 364216
rect 514758 363352 514814 363361
rect 514758 363287 514814 363296
rect 514772 362982 514800 363287
rect 514760 362976 514812 362982
rect 514760 362918 514812 362924
rect 514758 361992 514814 362001
rect 514758 361927 514814 361936
rect 514772 361622 514800 361927
rect 514760 361616 514812 361622
rect 514760 361558 514812 361564
rect 515312 345704 515364 345710
rect 515312 345646 515364 345652
rect 514760 342100 514812 342106
rect 514760 342042 514812 342048
rect 514772 341057 514800 342042
rect 514758 341048 514814 341057
rect 514758 340983 514814 340992
rect 514760 340876 514812 340882
rect 514760 340818 514812 340824
rect 514772 339697 514800 340818
rect 514758 339688 514814 339697
rect 514758 339623 514814 339632
rect 514760 339448 514812 339454
rect 514760 339390 514812 339396
rect 514772 338337 514800 339390
rect 514758 338328 514814 338337
rect 514758 338263 514814 338272
rect 514760 338088 514812 338094
rect 514760 338030 514812 338036
rect 514772 336977 514800 338030
rect 514758 336968 514814 336977
rect 514758 336903 514814 336912
rect 515324 335617 515352 345646
rect 515310 335608 515366 335617
rect 515310 335543 515366 335552
rect 514760 335300 514812 335306
rect 514760 335242 514812 335248
rect 514772 334257 514800 335242
rect 514758 334248 514814 334257
rect 514758 334183 514814 334192
rect 514760 333940 514812 333946
rect 514760 333882 514812 333888
rect 514772 332897 514800 333882
rect 514758 332888 514814 332897
rect 514758 332823 514814 332832
rect 514760 332580 514812 332586
rect 514760 332522 514812 332528
rect 514772 331537 514800 332522
rect 514758 331528 514814 331537
rect 514758 331463 514814 331472
rect 514758 327448 514814 327457
rect 514758 327383 514814 327392
rect 514772 327146 514800 327383
rect 514760 327140 514812 327146
rect 514760 327082 514812 327088
rect 514758 326088 514814 326097
rect 514758 326023 514814 326032
rect 514772 325718 514800 326023
rect 514760 325712 514812 325718
rect 514760 325654 514812 325660
rect 514758 324728 514814 324737
rect 514758 324663 514814 324672
rect 514772 324358 514800 324663
rect 514760 324352 514812 324358
rect 514760 324294 514812 324300
rect 514758 323368 514814 323377
rect 514758 323303 514814 323312
rect 514772 322998 514800 323303
rect 514760 322992 514812 322998
rect 514760 322934 514812 322940
rect 514758 322008 514814 322017
rect 514758 321943 514814 321952
rect 514772 321638 514800 321943
rect 514760 321632 514812 321638
rect 514760 321574 514812 321580
rect 514758 320648 514814 320657
rect 514758 320583 514814 320592
rect 514772 320210 514800 320583
rect 514760 320204 514812 320210
rect 514760 320146 514812 320152
rect 515036 303136 515088 303142
rect 515036 303078 515088 303084
rect 514944 303000 514996 303006
rect 514944 302942 514996 302948
rect 514760 302932 514812 302938
rect 514760 302874 514812 302880
rect 514772 301073 514800 302874
rect 514758 301064 514814 301073
rect 514758 300999 514814 301008
rect 514956 298353 514984 302942
rect 515048 299713 515076 303078
rect 515034 299704 515090 299713
rect 515034 299639 515090 299648
rect 514942 298344 514998 298353
rect 514942 298279 514998 298288
rect 514760 298104 514812 298110
rect 514760 298046 514812 298052
rect 514772 296993 514800 298046
rect 514758 296984 514814 296993
rect 514758 296919 514814 296928
rect 514760 296676 514812 296682
rect 514760 296618 514812 296624
rect 514772 295633 514800 296618
rect 514758 295624 514814 295633
rect 514758 295559 514814 295568
rect 393964 295316 394016 295322
rect 393964 295258 394016 295264
rect 514760 295316 514812 295322
rect 514760 295258 514812 295264
rect 514772 294273 514800 295258
rect 514758 294264 514814 294273
rect 514758 294199 514814 294208
rect 514760 291168 514812 291174
rect 514760 291110 514812 291116
rect 514772 290193 514800 291110
rect 514758 290184 514814 290193
rect 514758 290119 514814 290128
rect 514760 289808 514812 289814
rect 514760 289750 514812 289756
rect 514772 288833 514800 289750
rect 514758 288824 514814 288833
rect 514758 288759 514814 288768
rect 514758 284744 514814 284753
rect 514758 284679 514814 284688
rect 514772 284374 514800 284679
rect 514760 284368 514812 284374
rect 514760 284310 514812 284316
rect 514760 262200 514812 262206
rect 514760 262142 514812 262148
rect 514772 261089 514800 262142
rect 514758 261080 514814 261089
rect 514758 261015 514814 261024
rect 514760 260840 514812 260846
rect 514760 260782 514812 260788
rect 514772 259729 514800 260782
rect 514758 259720 514814 259729
rect 514758 259655 514814 259664
rect 514760 259412 514812 259418
rect 514760 259354 514812 259360
rect 514772 258369 514800 259354
rect 514758 258360 514814 258369
rect 514758 258295 514814 258304
rect 514760 257984 514812 257990
rect 514760 257926 514812 257932
rect 514772 257009 514800 257926
rect 514758 257000 514814 257009
rect 514758 256935 514814 256944
rect 514760 256692 514812 256698
rect 514760 256634 514812 256640
rect 514772 255649 514800 256634
rect 514758 255640 514814 255649
rect 514758 255575 514814 255584
rect 514760 255264 514812 255270
rect 514760 255206 514812 255212
rect 514772 254289 514800 255206
rect 514758 254280 514814 254289
rect 514758 254215 514814 254224
rect 514760 253904 514812 253910
rect 514760 253846 514812 253852
rect 514772 252929 514800 253846
rect 514758 252920 514814 252929
rect 514758 252855 514814 252864
rect 514760 252544 514812 252550
rect 514760 252486 514812 252492
rect 514772 251569 514800 252486
rect 514758 251560 514814 251569
rect 514758 251495 514814 251504
rect 514760 251184 514812 251190
rect 514760 251126 514812 251132
rect 514772 250209 514800 251126
rect 514758 250200 514814 250209
rect 514758 250135 514814 250144
rect 514760 249756 514812 249762
rect 514760 249698 514812 249704
rect 514772 248849 514800 249698
rect 514758 248840 514814 248849
rect 514758 248775 514814 248784
rect 514760 248396 514812 248402
rect 514760 248338 514812 248344
rect 514772 247489 514800 248338
rect 514758 247480 514814 247489
rect 514758 247415 514814 247424
rect 514760 247036 514812 247042
rect 514760 246978 514812 246984
rect 514772 246129 514800 246978
rect 514758 246120 514814 246129
rect 514758 246055 514814 246064
rect 514942 244760 514998 244769
rect 514942 244695 514998 244704
rect 514758 243400 514814 243409
rect 514758 243335 514814 243344
rect 514772 242962 514800 243335
rect 514760 242956 514812 242962
rect 514760 242898 514812 242904
rect 514956 239834 514984 244695
rect 514944 239828 514996 239834
rect 514944 239770 514996 239776
rect 377404 237380 377456 237386
rect 377404 237322 377456 237328
rect 366364 237312 366416 237318
rect 366364 237254 366416 237260
rect 364984 216572 365036 216578
rect 364984 216514 365036 216520
rect 362224 197328 362276 197334
rect 362224 197270 362276 197276
rect 367742 180024 367798 180033
rect 367742 179959 367798 179968
rect 364982 179888 365038 179897
rect 364982 179823 365038 179832
rect 345664 175024 345716 175030
rect 345664 174966 345716 174972
rect 364996 126041 365024 179823
rect 367756 165889 367784 179959
rect 515416 175234 515444 400551
rect 515508 364342 515536 412791
rect 515770 411496 515826 411505
rect 515770 411431 515826 411440
rect 515678 410136 515734 410145
rect 515678 410071 515734 410080
rect 515586 408776 515642 408785
rect 515586 408711 515642 408720
rect 515496 364336 515548 364342
rect 515496 364278 515548 364284
rect 515494 360632 515550 360641
rect 515494 360567 515550 360576
rect 515404 175228 515456 175234
rect 515404 175170 515456 175176
rect 515508 175166 515536 360567
rect 515600 300830 515628 408711
rect 515692 321570 515720 410071
rect 515784 342242 515812 411431
rect 515876 385014 515904 414151
rect 517440 400217 517468 421330
rect 517426 400208 517482 400217
rect 517426 400143 517482 400152
rect 518636 399537 518664 423807
rect 521672 421954 521700 423807
rect 521672 421926 521732 421954
rect 524328 421456 524380 421462
rect 519004 421394 519248 421410
rect 518992 421388 519248 421394
rect 519044 421382 519248 421388
rect 524216 421404 524328 421410
rect 527180 421456 527232 421462
rect 524216 421398 524380 421404
rect 524216 421382 524368 421398
rect 526700 421394 527036 421410
rect 527180 421398 527232 421404
rect 526700 421388 527048 421394
rect 526700 421382 526996 421388
rect 518992 421330 519044 421336
rect 526996 421330 527048 421336
rect 527192 412634 527220 421398
rect 529204 421388 529256 421394
rect 529204 421330 529256 421336
rect 527192 412606 527312 412634
rect 518898 400208 518954 400217
rect 518898 400143 518954 400152
rect 518622 399528 518678 399537
rect 518622 399463 518678 399472
rect 515864 385008 515916 385014
rect 515864 384950 515916 384956
rect 517426 383888 517482 383897
rect 517426 383823 517482 383832
rect 516046 371512 516102 371521
rect 516046 371447 516102 371456
rect 515954 370152 516010 370161
rect 515954 370087 516010 370096
rect 515862 368792 515918 368801
rect 515862 368727 515918 368736
rect 515772 342236 515824 342242
rect 515772 342178 515824 342184
rect 515770 328808 515826 328817
rect 515770 328743 515826 328752
rect 515680 321564 515732 321570
rect 515680 321506 515732 321512
rect 515680 304292 515732 304298
rect 515680 304234 515732 304240
rect 515588 300824 515640 300830
rect 515588 300766 515640 300772
rect 515692 291553 515720 304234
rect 515784 302190 515812 328743
rect 515772 302184 515824 302190
rect 515772 302126 515824 302132
rect 515876 300762 515904 368727
rect 515968 321502 515996 370087
rect 516060 342174 516088 371447
rect 517440 359417 517468 383823
rect 518912 381970 518940 400143
rect 521658 399528 521714 399537
rect 521658 399463 521714 399472
rect 521672 383897 521700 399463
rect 527284 398857 527312 412606
rect 529216 404977 529244 421330
rect 529938 410952 529994 410961
rect 529938 410887 529994 410896
rect 529202 404968 529258 404977
rect 529202 404903 529258 404912
rect 529216 402974 529244 404903
rect 529216 402946 529428 402974
rect 524326 398848 524382 398857
rect 524326 398783 524382 398792
rect 527270 398848 527326 398857
rect 527270 398783 527326 398792
rect 524340 383897 524368 398783
rect 521658 383888 521714 383897
rect 521658 383823 521714 383832
rect 524326 383888 524382 383897
rect 524326 383823 524382 383832
rect 529202 383888 529258 383897
rect 529202 383823 529258 383832
rect 521672 381970 521700 383823
rect 524340 381970 524368 383823
rect 527086 383752 527142 383761
rect 527086 383687 527142 383696
rect 528558 383752 528614 383761
rect 528558 383687 528614 383696
rect 527100 381970 527128 383687
rect 518912 381942 519248 381970
rect 521672 381942 521732 381970
rect 524216 381942 524368 381970
rect 526700 381942 527128 381970
rect 518912 381426 518940 381942
rect 518636 381398 518940 381426
rect 518636 360074 518664 381398
rect 518636 360046 518940 360074
rect 517426 359408 517482 359417
rect 517426 359343 517482 359352
rect 518438 343904 518494 343913
rect 518438 343839 518494 343848
rect 516048 342168 516100 342174
rect 516048 342110 516100 342116
rect 516046 330168 516102 330177
rect 516046 330103 516102 330112
rect 515956 321496 516008 321502
rect 515956 321438 516008 321444
rect 516060 321434 516088 330103
rect 516048 321428 516100 321434
rect 516048 321370 516100 321376
rect 518452 319433 518480 343839
rect 518912 341986 518940 360046
rect 521658 359408 521714 359417
rect 521658 359343 521714 359352
rect 521672 343913 521700 359343
rect 521658 343904 521714 343913
rect 521658 343839 521714 343848
rect 524326 343904 524382 343913
rect 524326 343839 524382 343848
rect 527270 343904 527326 343913
rect 527270 343839 527326 343848
rect 521672 341986 521700 343839
rect 524340 341986 524368 343839
rect 527086 343768 527142 343777
rect 527086 343703 527142 343712
rect 527100 341986 527128 343703
rect 518636 341958 519248 341986
rect 521672 341958 521732 341986
rect 524216 341958 524368 341986
rect 526700 341958 527128 341986
rect 518438 319424 518494 319433
rect 518438 319359 518494 319368
rect 518636 318794 518664 341958
rect 522302 319424 522358 319433
rect 522302 319359 522358 319368
rect 518636 318766 518940 318794
rect 515956 303068 516008 303074
rect 515956 303010 516008 303016
rect 515864 300756 515916 300762
rect 515864 300698 515916 300704
rect 515968 292913 515996 303010
rect 518912 301866 518940 318766
rect 522316 306374 522344 319359
rect 522132 306346 522344 306374
rect 522132 302297 522160 306346
rect 527086 303784 527142 303793
rect 527086 303719 527142 303728
rect 524326 303648 524382 303657
rect 524326 303583 524382 303592
rect 522118 302288 522174 302297
rect 522118 302223 522174 302232
rect 522132 301866 522160 302223
rect 524340 301866 524368 303583
rect 527100 301866 527128 303719
rect 527284 303657 527312 343839
rect 528572 343777 528600 383687
rect 529216 351937 529244 383823
rect 529400 383761 529428 402946
rect 529386 383752 529442 383761
rect 529386 383687 529442 383696
rect 529952 370977 529980 410887
rect 529938 370968 529994 370977
rect 529938 370903 529994 370912
rect 529202 351928 529258 351937
rect 529202 351863 529258 351872
rect 529216 343913 529244 351863
rect 529202 343904 529258 343913
rect 529202 343839 529258 343848
rect 528558 343768 528614 343777
rect 528558 343703 528614 343712
rect 528572 303793 528600 343703
rect 529952 330993 529980 370903
rect 529938 330984 529994 330993
rect 529938 330919 529994 330928
rect 528558 303784 528614 303793
rect 528558 303719 528614 303728
rect 527270 303648 527326 303657
rect 527270 303583 527326 303592
rect 518912 301850 519248 301866
rect 517428 301844 517480 301850
rect 517428 301786 517480 301792
rect 518900 301844 519248 301850
rect 518952 301838 519248 301844
rect 521732 301838 522160 301866
rect 524216 301838 524368 301866
rect 526700 301838 527128 301866
rect 518900 301786 518952 301792
rect 515954 292904 516010 292913
rect 515954 292839 516010 292848
rect 515678 291544 515734 291553
rect 515678 291479 515734 291488
rect 515954 287464 516010 287473
rect 515954 287399 516010 287408
rect 515862 286104 515918 286113
rect 515862 286039 515918 286048
rect 515770 283384 515826 283393
rect 515770 283319 515826 283328
rect 515678 282024 515734 282033
rect 515678 281959 515734 281968
rect 515586 280664 515642 280673
rect 515586 280599 515642 280608
rect 515496 175160 515548 175166
rect 515496 175102 515548 175108
rect 515600 175098 515628 280599
rect 515692 195974 515720 281959
rect 515784 216646 515812 283319
rect 515876 258058 515904 286039
rect 515968 280158 515996 287399
rect 515956 280152 516008 280158
rect 515956 280094 516008 280100
rect 517440 278905 517468 301786
rect 517426 278896 517482 278905
rect 517426 278831 517482 278840
rect 519542 278896 519598 278905
rect 519542 278831 519598 278840
rect 519556 267734 519584 278831
rect 519556 267706 519676 267734
rect 519648 263673 519676 267706
rect 527086 264888 527142 264897
rect 527086 264823 527142 264832
rect 524326 264616 524382 264625
rect 524326 264551 524382 264560
rect 522118 264480 522174 264489
rect 522118 264415 522174 264424
rect 519634 263664 519690 263673
rect 519634 263599 519690 263608
rect 519648 261882 519676 263599
rect 522132 261882 522160 264415
rect 524340 261882 524368 264551
rect 527100 261882 527128 264823
rect 527284 264625 527312 303583
rect 528572 264897 528600 303719
rect 528650 302288 528706 302297
rect 528650 302223 528706 302232
rect 528558 264888 528614 264897
rect 528558 264823 528614 264832
rect 527270 264616 527326 264625
rect 527270 264551 527326 264560
rect 528664 264489 528692 302223
rect 529952 291009 529980 330919
rect 580170 302288 580226 302297
rect 580170 302223 580226 302232
rect 580184 298761 580212 302223
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 529938 291000 529994 291009
rect 529938 290935 529994 290944
rect 528650 264480 528706 264489
rect 528650 264415 528706 264424
rect 527822 263664 527878 263673
rect 527822 263599 527878 263608
rect 519248 261854 519676 261882
rect 521732 261854 522160 261882
rect 524216 261854 524368 261882
rect 526700 261854 527128 261882
rect 515864 258052 515916 258058
rect 515864 257994 515916 258000
rect 527836 245585 527864 263599
rect 529952 251025 529980 290935
rect 529938 251016 529994 251025
rect 529938 250951 529994 250960
rect 530582 251016 530638 251025
rect 530582 250951 530638 250960
rect 527822 245576 527878 245585
rect 527822 245511 527878 245520
rect 515954 242040 516010 242049
rect 515954 241975 516010 241984
rect 515862 240680 515918 240689
rect 515862 240615 515918 240624
rect 515772 216640 515824 216646
rect 515772 216582 515824 216588
rect 515680 195968 515732 195974
rect 515680 195910 515732 195916
rect 515876 177002 515904 240615
rect 515968 197810 515996 241975
rect 515956 197804 516008 197810
rect 515956 197746 516008 197752
rect 515864 176996 515916 177002
rect 515864 176938 515916 176944
rect 515588 175092 515640 175098
rect 515588 175034 515640 175040
rect 367742 165880 367798 165889
rect 367742 165815 367798 165824
rect 364982 126032 365038 126041
rect 364982 125967 365038 125976
rect 308770 86184 308826 86193
rect 308770 86119 308826 86128
rect 308586 46336 308642 46345
rect 308586 46271 308642 46280
rect 530596 19825 530624 250951
rect 580172 206304 580224 206310
rect 580172 206246 580224 206252
rect 580184 205737 580212 206246
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 530582 19816 530638 19825
rect 530582 19751 530638 19760
rect 308402 6624 308458 6633
rect 308402 6559 308458 6568
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
<< via2 >>
rect 301134 494264 301190 494320
rect 309138 494264 309194 494320
rect 308402 473456 308458 473512
rect 292394 473320 292450 473376
rect 296626 473340 296682 473376
rect 296626 473320 296628 473340
rect 296628 473320 296680 473340
rect 296680 473320 296682 473340
rect 302422 473320 302478 473376
rect 309138 473320 309194 473376
rect 310518 473456 310574 473512
rect 309782 472368 309838 472424
rect 309506 472096 309562 472152
rect 302146 452784 302202 452840
rect 304906 452648 304962 452704
rect 309230 453872 309286 453928
rect 310518 453872 310574 453928
rect 309414 452784 309470 452840
rect 309230 452648 309286 452704
rect 304906 451560 304962 451616
rect 298466 451424 298522 451480
rect 302146 451424 302202 451480
rect 298098 451016 298154 451072
rect 301560 451016 301616 451072
rect 304877 451016 304933 451072
rect 291842 448568 291898 448624
rect 293958 448568 294014 448624
rect 294786 448568 294842 448624
rect 291842 430752 291898 430808
rect 308218 449792 308274 449848
rect 309046 449792 309102 449848
rect 305550 432112 305606 432168
rect 302054 431976 302110 432032
rect 298098 430752 298154 430808
rect 293958 430616 294014 430672
rect 309230 432112 309286 432168
rect 309874 431976 309930 432032
rect 302146 430480 302202 430536
rect 305550 430480 305606 430536
rect 308862 430480 308918 430536
rect 296074 430208 296130 430264
rect 309322 430208 309378 430264
rect 301944 430072 302000 430128
rect 305388 430072 305444 430128
rect 292762 429832 292818 429856
rect 292762 429800 292764 429832
rect 292764 429800 292816 429832
rect 292816 429800 292818 429832
rect 292486 426264 292542 426320
rect 293958 426264 294014 426320
rect 291106 410080 291162 410136
rect 291842 409944 291898 410000
rect 291106 389408 291162 389464
rect 301502 422864 301558 422920
rect 304814 411304 304870 411360
rect 301502 410080 301558 410136
rect 293958 409944 294014 410000
rect 301502 409400 301558 409456
rect 304814 409400 304870 409456
rect 301410 409128 301466 409184
rect 304722 409128 304778 409184
rect 309874 422864 309930 422920
rect 309138 411304 309194 411360
rect 302238 389408 302294 389464
rect 291934 389136 291990 389192
rect 298834 389136 298890 389192
rect 291106 385600 291162 385656
rect 309138 389272 309194 389328
rect 298834 388456 298890 388512
rect 302238 388456 302294 388512
rect 309046 388456 309102 388512
rect 299018 388184 299074 388240
rect 302238 388184 302294 388240
rect 309046 388184 309102 388240
rect 299478 385600 299534 385656
rect 291934 381520 291990 381576
rect 296718 381520 296774 381576
rect 291750 371320 291806 371376
rect 293958 371320 294014 371376
rect 291934 368464 291990 368520
rect 291750 367104 291806 367160
rect 304078 369688 304134 369744
rect 299478 368464 299534 368520
rect 300122 368464 300178 368520
rect 308034 368464 308090 368520
rect 293958 367376 294014 367432
rect 296718 367376 296774 367432
rect 300122 367376 300178 367432
rect 304078 367376 304134 367432
rect 294050 367104 294106 367160
rect 297362 367104 297418 367160
rect 300214 367104 300270 367160
rect 303986 367104 304042 367160
rect 303802 361528 303858 361584
rect 304906 361528 304962 361584
rect 296718 360168 296774 360224
rect 297638 360168 297694 360224
rect 291934 348336 291990 348392
rect 299570 348336 299626 348392
rect 299570 347792 299626 347848
rect 291842 346568 291898 346624
rect 296718 346568 296774 346624
rect 304906 346432 304962 346488
rect 308034 347792 308090 347848
rect 297270 346160 297326 346216
rect 303986 346160 304042 346216
rect 307942 346432 307998 346488
rect 307666 325760 307722 325816
rect 308586 325760 308642 325816
rect 309598 325760 309654 325816
rect 291934 305088 291990 305144
rect 291842 283464 291898 283520
rect 306010 305768 306066 305824
rect 302422 305632 302478 305688
rect 298466 305088 298522 305144
rect 292394 304952 292450 305008
rect 294970 304952 295026 305008
rect 308494 305768 308550 305824
rect 308402 305632 308458 305688
rect 308494 305088 308550 305144
rect 308402 304952 308458 305008
rect 310518 304952 310574 305008
rect 308678 302232 308734 302288
rect 309506 302232 309562 302288
rect 304906 284416 304962 284472
rect 301686 284280 301742 284336
rect 295246 283464 295302 283520
rect 301686 283464 301742 283520
rect 304906 283464 304962 283520
rect 309138 285640 309194 285696
rect 309138 284416 309194 284472
rect 309322 284280 309378 284336
rect 301591 283056 301647 283112
rect 304908 283056 304964 283112
rect 305918 263744 305974 263800
rect 302146 263608 302202 263664
rect 310518 284280 310574 284336
rect 309322 263744 309378 263800
rect 309230 263608 309286 263664
rect 309874 263608 309930 263664
rect 302146 262520 302202 262576
rect 305918 262520 305974 262576
rect 309046 262520 309102 262576
rect 309322 262520 309378 262576
rect 301942 262112 301998 262168
rect 305386 262112 305442 262168
rect 309322 262112 309378 262168
rect 308830 261976 308886 262032
rect 304906 250416 304962 250472
rect 301502 242936 301558 242992
rect 301502 241440 301558 241496
rect 304814 241440 304870 241496
rect 301410 241168 301466 241224
rect 304722 241168 304778 241224
rect 309230 250416 309286 250472
rect 309138 242936 309194 242992
rect 306838 223488 306894 223544
rect 302790 222808 302846 222864
rect 309874 242936 309930 242992
rect 309230 223488 309286 223544
rect 309138 222808 309194 222864
rect 307942 222672 307998 222728
rect 309690 222672 309746 222728
rect 302790 220360 302846 220416
rect 306838 220360 306894 220416
rect 309690 220360 309746 220416
rect 302745 219952 302801 220008
rect 291842 218456 291898 218512
rect 306746 220088 306802 220144
rect 309782 220088 309838 220144
rect 294694 218456 294750 218512
rect 291842 200232 291898 200288
rect 291750 200096 291806 200152
rect 291750 180240 291806 180296
rect 304906 217776 304962 217832
rect 306378 217776 306434 217832
rect 306930 217776 306986 217832
rect 300766 200640 300822 200696
rect 300766 200232 300822 200288
rect 297546 200096 297602 200152
rect 294694 199416 294750 199472
rect 310150 217776 310206 217832
rect 311346 388184 311402 388240
rect 311346 368464 311402 368520
rect 306930 199416 306986 199472
rect 292486 198736 292542 198792
rect 293682 198780 293684 198792
rect 293684 198780 293736 198792
rect 293736 198780 293738 198792
rect 293682 198736 293738 198780
rect 307574 199144 307630 199200
rect 291842 179968 291898 180024
rect 303986 197376 304042 197432
rect 304814 197376 304870 197432
rect 296718 180240 296774 180296
rect 298006 180240 298062 180296
rect 292486 179424 292542 179480
rect 293958 179424 294014 179480
rect 311898 389272 311954 389328
rect 311898 369688 311954 369744
rect 311898 305088 311954 305144
rect 311898 285640 311954 285696
rect 311898 222808 311954 222864
rect 311898 200640 311954 200696
rect 306930 179968 306986 180024
rect 307758 179968 307814 180024
rect 304538 179832 304594 179888
rect 300766 179696 300822 179752
rect 298006 179560 298062 179616
rect 308770 179696 308826 179752
rect 308586 179560 308642 179616
rect 308402 179424 308458 179480
rect 514758 420960 514814 421016
rect 518622 423816 518678 423872
rect 521658 423816 521714 423872
rect 515402 419600 515458 419656
rect 514758 418240 514814 418296
rect 514758 416880 514814 416936
rect 515402 415520 515458 415576
rect 514758 407360 514814 407416
rect 514758 406000 514814 406056
rect 515862 414160 515918 414216
rect 515494 412800 515550 412856
rect 514758 404640 514814 404696
rect 514758 403280 514814 403336
rect 514758 401920 514814 401976
rect 515402 400560 515458 400616
rect 514758 380976 514814 381032
rect 514758 379616 514814 379672
rect 514758 378256 514814 378312
rect 514758 376896 514814 376952
rect 514758 375536 514814 375592
rect 514758 374176 514814 374232
rect 515310 372816 515366 372872
rect 514758 367376 514814 367432
rect 514758 366016 514814 366072
rect 514758 364656 514814 364712
rect 514758 363296 514814 363352
rect 514758 361936 514814 361992
rect 514758 340992 514814 341048
rect 514758 339632 514814 339688
rect 514758 338272 514814 338328
rect 514758 336912 514814 336968
rect 515310 335552 515366 335608
rect 514758 334192 514814 334248
rect 514758 332832 514814 332888
rect 514758 331472 514814 331528
rect 514758 327392 514814 327448
rect 514758 326032 514814 326088
rect 514758 324672 514814 324728
rect 514758 323312 514814 323368
rect 514758 321952 514814 322008
rect 514758 320592 514814 320648
rect 514758 301008 514814 301064
rect 515034 299648 515090 299704
rect 514942 298288 514998 298344
rect 514758 296928 514814 296984
rect 514758 295568 514814 295624
rect 514758 294208 514814 294264
rect 514758 290128 514814 290184
rect 514758 288768 514814 288824
rect 514758 284688 514814 284744
rect 514758 261024 514814 261080
rect 514758 259664 514814 259720
rect 514758 258304 514814 258360
rect 514758 256944 514814 257000
rect 514758 255584 514814 255640
rect 514758 254224 514814 254280
rect 514758 252864 514814 252920
rect 514758 251504 514814 251560
rect 514758 250144 514814 250200
rect 514758 248784 514814 248840
rect 514758 247424 514814 247480
rect 514758 246064 514814 246120
rect 514942 244704 514998 244760
rect 514758 243344 514814 243400
rect 367742 179968 367798 180024
rect 364982 179832 365038 179888
rect 515770 411440 515826 411496
rect 515678 410080 515734 410136
rect 515586 408720 515642 408776
rect 515494 360576 515550 360632
rect 517426 400152 517482 400208
rect 518898 400152 518954 400208
rect 518622 399472 518678 399528
rect 517426 383832 517482 383888
rect 516046 371456 516102 371512
rect 515954 370096 516010 370152
rect 515862 368736 515918 368792
rect 515770 328752 515826 328808
rect 521658 399472 521714 399528
rect 529938 410896 529994 410952
rect 529202 404912 529258 404968
rect 524326 398792 524382 398848
rect 527270 398792 527326 398848
rect 521658 383832 521714 383888
rect 524326 383832 524382 383888
rect 529202 383832 529258 383888
rect 527086 383696 527142 383752
rect 528558 383696 528614 383752
rect 517426 359352 517482 359408
rect 518438 343848 518494 343904
rect 516046 330112 516102 330168
rect 521658 359352 521714 359408
rect 521658 343848 521714 343904
rect 524326 343848 524382 343904
rect 527270 343848 527326 343904
rect 527086 343712 527142 343768
rect 518438 319368 518494 319424
rect 522302 319368 522358 319424
rect 527086 303728 527142 303784
rect 524326 303592 524382 303648
rect 522118 302232 522174 302288
rect 529386 383696 529442 383752
rect 529938 370912 529994 370968
rect 529202 351872 529258 351928
rect 529202 343848 529258 343904
rect 528558 343712 528614 343768
rect 529938 330928 529994 330984
rect 528558 303728 528614 303784
rect 527270 303592 527326 303648
rect 515954 292848 516010 292904
rect 515678 291488 515734 291544
rect 515954 287408 516010 287464
rect 515862 286048 515918 286104
rect 515770 283328 515826 283384
rect 515678 281968 515734 282024
rect 515586 280608 515642 280664
rect 517426 278840 517482 278896
rect 519542 278840 519598 278896
rect 527086 264832 527142 264888
rect 524326 264560 524382 264616
rect 522118 264424 522174 264480
rect 519634 263608 519690 263664
rect 528650 302232 528706 302288
rect 528558 264832 528614 264888
rect 527270 264560 527326 264616
rect 580170 302232 580226 302288
rect 580170 298696 580226 298752
rect 529938 290944 529994 291000
rect 528650 264424 528706 264480
rect 527822 263608 527878 263664
rect 529938 250960 529994 251016
rect 530582 250960 530638 251016
rect 527822 245520 527878 245576
rect 515954 241984 516010 242040
rect 515862 240624 515918 240680
rect 367742 165824 367798 165880
rect 364982 125976 365038 126032
rect 308770 86128 308826 86184
rect 308586 46280 308642 46336
rect 580170 205672 580226 205728
rect 530582 19760 530638 19816
rect 308402 6568 308458 6624
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect 301129 494322 301195 494325
rect 309133 494322 309199 494325
rect 301129 494320 309199 494322
rect 301129 494264 301134 494320
rect 301190 494264 309138 494320
rect 309194 494264 309199 494320
rect 301129 494262 309199 494264
rect 301129 494259 301195 494262
rect 309133 494259 309199 494262
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 308397 473514 308463 473517
rect 310513 473514 310579 473517
rect 308397 473512 310579 473514
rect 308397 473456 308402 473512
rect 308458 473456 310518 473512
rect 310574 473456 310579 473512
rect 308397 473454 310579 473456
rect 308397 473451 308463 473454
rect 310513 473451 310579 473454
rect 292389 473378 292455 473381
rect 296621 473378 296687 473381
rect 292389 473376 296687 473378
rect 292389 473320 292394 473376
rect 292450 473320 296626 473376
rect 296682 473320 296687 473376
rect 292389 473318 296687 473320
rect 292389 473315 292455 473318
rect 296621 473315 296687 473318
rect 302417 473378 302483 473381
rect 309133 473378 309199 473381
rect 302417 473376 309199 473378
rect 302417 473320 302422 473376
rect 302478 473320 309138 473376
rect 309194 473320 309199 473376
rect 302417 473318 309199 473320
rect 302417 473315 302483 473318
rect 309133 473315 309199 473318
rect 309777 472426 309843 472429
rect 309734 472424 309843 472426
rect 309734 472368 309782 472424
rect 309838 472368 309843 472424
rect 309734 472363 309843 472368
rect 309501 472154 309567 472157
rect 309734 472154 309794 472363
rect 309501 472152 309794 472154
rect 309501 472096 309506 472152
rect 309562 472096 309794 472152
rect 309501 472094 309794 472096
rect 309501 472091 309567 472094
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect 309225 453930 309291 453933
rect 310513 453930 310579 453933
rect 309225 453928 310579 453930
rect 309225 453872 309230 453928
rect 309286 453872 310518 453928
rect 310574 453872 310579 453928
rect 309225 453870 310579 453872
rect 309225 453867 309291 453870
rect 310513 453867 310579 453870
rect 302141 452842 302207 452845
rect 309409 452842 309475 452845
rect 302141 452840 309475 452842
rect 302141 452784 302146 452840
rect 302202 452784 309414 452840
rect 309470 452784 309475 452840
rect 302141 452782 309475 452784
rect 302141 452779 302207 452782
rect 309409 452779 309475 452782
rect 304901 452706 304967 452709
rect 309225 452706 309291 452709
rect 304901 452704 309291 452706
rect 304901 452648 304906 452704
rect 304962 452648 309230 452704
rect 309286 452648 309291 452704
rect 304901 452646 309291 452648
rect 304901 452643 304967 452646
rect 309225 452643 309291 452646
rect 304901 451616 304967 451621
rect 304901 451560 304906 451616
rect 304962 451560 304967 451616
rect 304901 451555 304967 451560
rect 298461 451482 298527 451485
rect 302141 451482 302207 451485
rect 298142 451480 298527 451482
rect 298142 451424 298466 451480
rect 298522 451424 298527 451480
rect 298142 451422 298527 451424
rect 298142 451077 298202 451422
rect 298461 451419 298527 451422
rect 301684 451480 302207 451482
rect 301684 451424 302146 451480
rect 302202 451424 302207 451480
rect 301684 451422 302207 451424
rect 298093 451072 298202 451077
rect 298093 451016 298098 451072
rect 298154 451016 298202 451072
rect 298093 451014 298202 451016
rect 301555 451074 301621 451077
rect 301684 451074 301744 451422
rect 302141 451419 302207 451422
rect 304904 451077 304964 451555
rect 301555 451072 301744 451074
rect 301555 451016 301560 451072
rect 301616 451016 301744 451072
rect 301555 451014 301744 451016
rect 304872 451072 304964 451077
rect 304872 451016 304877 451072
rect 304933 451016 304964 451072
rect 304872 451014 304964 451016
rect 298093 451011 298159 451014
rect 301555 451011 301621 451014
rect 304872 451011 304938 451014
rect 308213 449850 308279 449853
rect 309041 449850 309107 449853
rect 308213 449848 309107 449850
rect 308213 449792 308218 449848
rect 308274 449792 309046 449848
rect 309102 449792 309107 449848
rect 308213 449790 309107 449792
rect 308213 449787 308279 449790
rect 309041 449787 309107 449790
rect -960 449428 480 449668
rect 291837 448626 291903 448629
rect 293953 448626 294019 448629
rect 294781 448626 294847 448629
rect 291837 448624 294847 448626
rect 291837 448568 291842 448624
rect 291898 448568 293958 448624
rect 294014 448568 294786 448624
rect 294842 448568 294847 448624
rect 291837 448566 294847 448568
rect 291837 448563 291903 448566
rect 293953 448563 294019 448566
rect 294781 448563 294847 448566
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 305545 432170 305611 432173
rect 309225 432170 309291 432173
rect 305545 432168 309291 432170
rect 305545 432112 305550 432168
rect 305606 432112 309230 432168
rect 309286 432112 309291 432168
rect 305545 432110 309291 432112
rect 305545 432107 305611 432110
rect 309225 432107 309291 432110
rect 302049 432034 302115 432037
rect 309869 432034 309935 432037
rect 302049 432032 309935 432034
rect 302049 431976 302054 432032
rect 302110 431976 309874 432032
rect 309930 431976 309935 432032
rect 302049 431974 309935 431976
rect 302049 431971 302115 431974
rect 309869 431971 309935 431974
rect 583520 431476 584960 431716
rect 291837 430810 291903 430813
rect 298093 430810 298159 430813
rect 291837 430808 298159 430810
rect 291837 430752 291842 430808
rect 291898 430752 298098 430808
rect 298154 430752 298159 430808
rect 291837 430750 298159 430752
rect 291837 430747 291903 430750
rect 293953 430674 294019 430677
rect 292806 430672 294019 430674
rect 292806 430616 293958 430672
rect 294014 430616 294019 430672
rect 292806 430614 294019 430616
rect 292806 429861 292866 430614
rect 293953 430611 294019 430614
rect 296118 430269 296178 430750
rect 298093 430747 298159 430750
rect 302141 430538 302207 430541
rect 302141 430536 302250 430538
rect 302141 430480 302146 430536
rect 302202 430480 302250 430536
rect 302141 430475 302250 430480
rect 305545 430536 305611 430541
rect 305545 430480 305550 430536
rect 305606 430480 305611 430536
rect 305545 430475 305611 430480
rect 308857 430538 308923 430541
rect 308857 430536 309058 430538
rect 308857 430480 308862 430536
rect 308918 430480 309058 430536
rect 308857 430478 309058 430480
rect 308857 430475 308923 430478
rect 296069 430264 296178 430269
rect 296069 430208 296074 430264
rect 296130 430208 296178 430264
rect 296069 430206 296178 430208
rect 296069 430203 296135 430206
rect 301939 430130 302005 430133
rect 302190 430130 302250 430475
rect 301939 430128 302250 430130
rect 301939 430072 301944 430128
rect 302000 430072 302250 430128
rect 301939 430070 302250 430072
rect 305383 430130 305449 430133
rect 305548 430130 305608 430475
rect 308998 430266 309058 430478
rect 309317 430266 309383 430269
rect 308998 430264 309383 430266
rect 308998 430208 309322 430264
rect 309378 430208 309383 430264
rect 308998 430206 309383 430208
rect 309317 430203 309383 430206
rect 305383 430128 305608 430130
rect 305383 430072 305388 430128
rect 305444 430072 305608 430128
rect 305383 430070 305608 430072
rect 301939 430067 302005 430070
rect 305383 430067 305449 430070
rect 292757 429856 292866 429861
rect 292757 429800 292762 429856
rect 292818 429800 292866 429856
rect 292757 429798 292866 429800
rect 292757 429795 292823 429798
rect 292481 426322 292547 426325
rect 293953 426322 294019 426325
rect 292481 426320 294019 426322
rect 292481 426264 292486 426320
rect 292542 426264 293958 426320
rect 294014 426264 294019 426320
rect 292481 426262 294019 426264
rect 292481 426259 292547 426262
rect 293953 426259 294019 426262
rect 518617 423874 518683 423877
rect 521653 423874 521719 423877
rect 518617 423872 521719 423874
rect 518617 423816 518622 423872
rect 518678 423816 521658 423872
rect 521714 423816 521719 423872
rect 518617 423814 521719 423816
rect 518617 423811 518683 423814
rect 521653 423811 521719 423814
rect -960 423452 480 423692
rect 301497 422922 301563 422925
rect 309869 422922 309935 422925
rect 301497 422920 309935 422922
rect 301497 422864 301502 422920
rect 301558 422864 309874 422920
rect 309930 422864 309935 422920
rect 301497 422862 309935 422864
rect 301497 422859 301563 422862
rect 309869 422859 309935 422862
rect 514753 421018 514819 421021
rect 514753 421016 518052 421018
rect 514753 420960 514758 421016
rect 514814 420960 518052 421016
rect 514753 420958 518052 420960
rect 514753 420955 514819 420958
rect 515397 419658 515463 419661
rect 515397 419656 518052 419658
rect 515397 419600 515402 419656
rect 515458 419600 518052 419656
rect 515397 419598 518052 419600
rect 515397 419595 515463 419598
rect 514753 418298 514819 418301
rect 514753 418296 518052 418298
rect 514753 418240 514758 418296
rect 514814 418240 518052 418296
rect 514753 418238 518052 418240
rect 514753 418235 514819 418238
rect 583520 418148 584960 418388
rect 514753 416938 514819 416941
rect 514753 416936 518052 416938
rect 514753 416880 514758 416936
rect 514814 416880 518052 416936
rect 514753 416878 518052 416880
rect 514753 416875 514819 416878
rect 515397 415578 515463 415581
rect 515397 415576 518052 415578
rect 515397 415520 515402 415576
rect 515458 415520 518052 415576
rect 515397 415518 518052 415520
rect 515397 415515 515463 415518
rect 515857 414218 515923 414221
rect 515857 414216 518052 414218
rect 515857 414160 515862 414216
rect 515918 414160 518052 414216
rect 515857 414158 518052 414160
rect 515857 414155 515923 414158
rect 515489 412858 515555 412861
rect 515489 412856 518052 412858
rect 515489 412800 515494 412856
rect 515550 412800 518052 412856
rect 515489 412798 518052 412800
rect 515489 412795 515555 412798
rect 515765 411498 515831 411501
rect 515765 411496 518052 411498
rect 515765 411440 515770 411496
rect 515826 411440 518052 411496
rect 515765 411438 518052 411440
rect 515765 411435 515831 411438
rect 304809 411362 304875 411365
rect 309133 411362 309199 411365
rect 304809 411360 309199 411362
rect 304809 411304 304814 411360
rect 304870 411304 309138 411360
rect 309194 411304 309199 411360
rect 304809 411302 309199 411304
rect 304809 411299 304875 411302
rect 309133 411299 309199 411302
rect 529933 410954 529999 410957
rect 527804 410952 529999 410954
rect 527804 410896 529938 410952
rect 529994 410896 529999 410952
rect 527804 410894 529999 410896
rect 529933 410891 529999 410894
rect -960 410396 480 410636
rect 291101 410138 291167 410141
rect 301497 410138 301563 410141
rect 291101 410136 301563 410138
rect 291101 410080 291106 410136
rect 291162 410080 301502 410136
rect 301558 410080 301563 410136
rect 291101 410078 301563 410080
rect 291101 410075 291167 410078
rect 301497 410075 301563 410078
rect 515673 410138 515739 410141
rect 515673 410136 518052 410138
rect 515673 410080 515678 410136
rect 515734 410080 518052 410136
rect 515673 410078 518052 410080
rect 515673 410075 515739 410078
rect 291837 410002 291903 410005
rect 293953 410002 294019 410005
rect 291837 410000 294019 410002
rect 291837 409944 291842 410000
rect 291898 409944 293958 410000
rect 294014 409944 294019 410000
rect 291837 409942 294019 409944
rect 291837 409939 291903 409942
rect 293953 409939 294019 409942
rect 301497 409458 301563 409461
rect 304809 409458 304875 409461
rect 301454 409456 301563 409458
rect 301454 409400 301502 409456
rect 301558 409400 301563 409456
rect 301454 409395 301563 409400
rect 304766 409456 304875 409458
rect 304766 409400 304814 409456
rect 304870 409400 304875 409456
rect 304766 409395 304875 409400
rect 301454 409189 301514 409395
rect 304766 409189 304826 409395
rect 301405 409184 301514 409189
rect 301405 409128 301410 409184
rect 301466 409128 301514 409184
rect 301405 409126 301514 409128
rect 304717 409184 304826 409189
rect 304717 409128 304722 409184
rect 304778 409128 304826 409184
rect 304717 409126 304826 409128
rect 301405 409123 301471 409126
rect 304717 409123 304783 409126
rect 515581 408778 515647 408781
rect 515581 408776 518052 408778
rect 515581 408720 515586 408776
rect 515642 408720 518052 408776
rect 515581 408718 518052 408720
rect 515581 408715 515647 408718
rect 514753 407418 514819 407421
rect 514753 407416 518052 407418
rect 514753 407360 514758 407416
rect 514814 407360 518052 407416
rect 514753 407358 518052 407360
rect 514753 407355 514819 407358
rect 514753 406058 514819 406061
rect 514753 406056 518052 406058
rect 514753 406000 514758 406056
rect 514814 406000 518052 406056
rect 514753 405998 518052 406000
rect 514753 405995 514819 405998
rect 529197 404970 529263 404973
rect 583520 404970 584960 405060
rect 529197 404968 584960 404970
rect 529197 404912 529202 404968
rect 529258 404912 584960 404968
rect 529197 404910 584960 404912
rect 529197 404907 529263 404910
rect 583520 404820 584960 404910
rect 514753 404698 514819 404701
rect 514753 404696 518052 404698
rect 514753 404640 514758 404696
rect 514814 404640 518052 404696
rect 514753 404638 518052 404640
rect 514753 404635 514819 404638
rect 514753 403338 514819 403341
rect 514753 403336 518052 403338
rect 514753 403280 514758 403336
rect 514814 403280 518052 403336
rect 514753 403278 518052 403280
rect 514753 403275 514819 403278
rect 514753 401978 514819 401981
rect 514753 401976 518052 401978
rect 514753 401920 514758 401976
rect 514814 401920 518052 401976
rect 514753 401918 518052 401920
rect 514753 401915 514819 401918
rect 515397 400618 515463 400621
rect 515397 400616 518052 400618
rect 515397 400560 515402 400616
rect 515458 400560 518052 400616
rect 515397 400558 518052 400560
rect 515397 400555 515463 400558
rect 517421 400210 517487 400213
rect 518893 400210 518959 400213
rect 517421 400208 518959 400210
rect 517421 400152 517426 400208
rect 517482 400152 518898 400208
rect 518954 400152 518959 400208
rect 517421 400150 518959 400152
rect 517421 400147 517487 400150
rect 518893 400147 518959 400150
rect 518617 399530 518683 399533
rect 521653 399530 521719 399533
rect 518617 399528 521719 399530
rect 518617 399472 518622 399528
rect 518678 399472 521658 399528
rect 521714 399472 521719 399528
rect 518617 399470 521719 399472
rect 518617 399467 518683 399470
rect 521653 399467 521719 399470
rect 524321 398850 524387 398853
rect 527265 398850 527331 398853
rect 524321 398848 527331 398850
rect 524321 398792 524326 398848
rect 524382 398792 527270 398848
rect 527326 398792 527331 398848
rect 524321 398790 527331 398792
rect 524321 398787 524387 398790
rect 527265 398787 527331 398790
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect 291101 389466 291167 389469
rect 302233 389466 302299 389469
rect 291101 389464 302299 389466
rect 291101 389408 291106 389464
rect 291162 389408 302238 389464
rect 302294 389408 302299 389464
rect 291101 389406 302299 389408
rect 291101 389403 291167 389406
rect 302233 389403 302299 389406
rect 309133 389330 309199 389333
rect 311893 389330 311959 389333
rect 309133 389328 311959 389330
rect 309133 389272 309138 389328
rect 309194 389272 311898 389328
rect 311954 389272 311959 389328
rect 309133 389270 311959 389272
rect 309133 389267 309199 389270
rect 311893 389267 311959 389270
rect 291929 389194 291995 389197
rect 298829 389194 298895 389197
rect 291929 389192 298895 389194
rect 291929 389136 291934 389192
rect 291990 389136 298834 389192
rect 298890 389136 298895 389192
rect 291929 389134 298895 389136
rect 291929 389131 291995 389134
rect 298829 389131 298895 389134
rect 298829 388514 298895 388517
rect 298829 388512 298938 388514
rect 298829 388456 298834 388512
rect 298890 388456 298938 388512
rect 298829 388451 298938 388456
rect 302233 388512 302299 388517
rect 309041 388514 309107 388517
rect 302233 388456 302238 388512
rect 302294 388456 302299 388512
rect 302233 388451 302299 388456
rect 308998 388512 309107 388514
rect 308998 388456 309046 388512
rect 309102 388456 309107 388512
rect 308998 388451 309107 388456
rect 298878 388242 298938 388451
rect 302236 388245 302296 388451
rect 308998 388245 309058 388451
rect 299013 388242 299079 388245
rect 298878 388240 299079 388242
rect 298878 388184 299018 388240
rect 299074 388184 299079 388240
rect 298878 388182 299079 388184
rect 299013 388179 299079 388182
rect 302233 388240 302299 388245
rect 302233 388184 302238 388240
rect 302294 388184 302299 388240
rect 302233 388179 302299 388184
rect 308998 388242 309107 388245
rect 311341 388242 311407 388245
rect 308998 388240 311407 388242
rect 308998 388184 309046 388240
rect 309102 388184 311346 388240
rect 311402 388184 311407 388240
rect 308998 388182 311407 388184
rect 309041 388179 309107 388182
rect 311341 388179 311407 388182
rect 291101 385658 291167 385661
rect 299473 385658 299539 385661
rect 291101 385656 299539 385658
rect 291101 385600 291106 385656
rect 291162 385600 299478 385656
rect 299534 385600 299539 385656
rect 291101 385598 299539 385600
rect 291101 385595 291167 385598
rect 299473 385595 299539 385598
rect -960 384284 480 384524
rect 517421 383890 517487 383893
rect 521653 383890 521719 383893
rect 517421 383888 521719 383890
rect 517421 383832 517426 383888
rect 517482 383832 521658 383888
rect 521714 383832 521719 383888
rect 517421 383830 521719 383832
rect 517421 383827 517487 383830
rect 521653 383827 521719 383830
rect 524321 383890 524387 383893
rect 529197 383890 529263 383893
rect 524321 383888 529263 383890
rect 524321 383832 524326 383888
rect 524382 383832 529202 383888
rect 529258 383832 529263 383888
rect 524321 383830 529263 383832
rect 524321 383827 524387 383830
rect 529197 383827 529263 383830
rect 527081 383754 527147 383757
rect 528553 383754 528619 383757
rect 529381 383754 529447 383757
rect 527081 383752 529447 383754
rect 527081 383696 527086 383752
rect 527142 383696 528558 383752
rect 528614 383696 529386 383752
rect 529442 383696 529447 383752
rect 527081 383694 529447 383696
rect 527081 383691 527147 383694
rect 528553 383691 528619 383694
rect 529381 383691 529447 383694
rect 291929 381578 291995 381581
rect 296713 381578 296779 381581
rect 291929 381576 296779 381578
rect 291929 381520 291934 381576
rect 291990 381520 296718 381576
rect 296774 381520 296779 381576
rect 291929 381518 296779 381520
rect 291929 381515 291995 381518
rect 296713 381515 296779 381518
rect 514753 381034 514819 381037
rect 514753 381032 518052 381034
rect 514753 380976 514758 381032
rect 514814 380976 518052 381032
rect 514753 380974 518052 380976
rect 514753 380971 514819 380974
rect 514753 379674 514819 379677
rect 514753 379672 518052 379674
rect 514753 379616 514758 379672
rect 514814 379616 518052 379672
rect 514753 379614 518052 379616
rect 514753 379611 514819 379614
rect 514753 378314 514819 378317
rect 514753 378312 518052 378314
rect 514753 378256 514758 378312
rect 514814 378256 518052 378312
rect 583520 378300 584960 378540
rect 514753 378254 518052 378256
rect 514753 378251 514819 378254
rect 514753 376954 514819 376957
rect 514753 376952 518052 376954
rect 514753 376896 514758 376952
rect 514814 376896 518052 376952
rect 514753 376894 518052 376896
rect 514753 376891 514819 376894
rect 514753 375594 514819 375597
rect 514753 375592 518052 375594
rect 514753 375536 514758 375592
rect 514814 375536 518052 375592
rect 514753 375534 518052 375536
rect 514753 375531 514819 375534
rect 514753 374234 514819 374237
rect 514753 374232 518052 374234
rect 514753 374176 514758 374232
rect 514814 374176 518052 374232
rect 514753 374174 518052 374176
rect 514753 374171 514819 374174
rect 515305 372874 515371 372877
rect 515305 372872 518052 372874
rect 515305 372816 515310 372872
rect 515366 372816 518052 372872
rect 515305 372814 518052 372816
rect 515305 372811 515371 372814
rect 516041 371514 516107 371517
rect 516041 371512 518052 371514
rect -960 371228 480 371468
rect 516041 371456 516046 371512
rect 516102 371456 518052 371512
rect 516041 371454 518052 371456
rect 516041 371451 516107 371454
rect 291745 371378 291811 371381
rect 293953 371378 294019 371381
rect 291745 371376 294019 371378
rect 291745 371320 291750 371376
rect 291806 371320 293958 371376
rect 294014 371320 294019 371376
rect 291745 371318 294019 371320
rect 291745 371315 291811 371318
rect 293953 371315 294019 371318
rect 529933 370970 529999 370973
rect 527804 370968 529999 370970
rect 527804 370912 529938 370968
rect 529994 370912 529999 370968
rect 527804 370910 529999 370912
rect 529933 370907 529999 370910
rect 515949 370154 516015 370157
rect 515949 370152 518052 370154
rect 515949 370096 515954 370152
rect 516010 370096 518052 370152
rect 515949 370094 518052 370096
rect 515949 370091 516015 370094
rect 304073 369746 304139 369749
rect 311893 369746 311959 369749
rect 304073 369744 311959 369746
rect 304073 369688 304078 369744
rect 304134 369688 311898 369744
rect 311954 369688 311959 369744
rect 304073 369686 311959 369688
rect 304073 369683 304139 369686
rect 311893 369683 311959 369686
rect 515857 368794 515923 368797
rect 515857 368792 518052 368794
rect 515857 368736 515862 368792
rect 515918 368736 518052 368792
rect 515857 368734 518052 368736
rect 515857 368731 515923 368734
rect 291929 368522 291995 368525
rect 299473 368522 299539 368525
rect 300117 368522 300183 368525
rect 291929 368520 300183 368522
rect 291929 368464 291934 368520
rect 291990 368464 299478 368520
rect 299534 368464 300122 368520
rect 300178 368464 300183 368520
rect 291929 368462 300183 368464
rect 291929 368459 291995 368462
rect 299473 368459 299539 368462
rect 300117 368459 300183 368462
rect 308029 368522 308095 368525
rect 311341 368522 311407 368525
rect 308029 368520 311407 368522
rect 308029 368464 308034 368520
rect 308090 368464 311346 368520
rect 311402 368464 311407 368520
rect 308029 368462 311407 368464
rect 308029 368459 308095 368462
rect 311341 368459 311407 368462
rect 293953 367434 294019 367437
rect 296713 367434 296779 367437
rect 300117 367434 300183 367437
rect 304073 367434 304139 367437
rect 293953 367432 294154 367434
rect 293953 367376 293958 367432
rect 294014 367376 294154 367432
rect 293953 367374 294154 367376
rect 293953 367371 294019 367374
rect 294094 367298 294154 367374
rect 296713 367432 297282 367434
rect 296713 367376 296718 367432
rect 296774 367376 297282 367432
rect 296713 367374 297282 367376
rect 296713 367371 296779 367374
rect 292254 367238 294154 367298
rect 291745 367162 291811 367165
rect 292254 367162 292314 367238
rect 294094 367165 294154 367238
rect 291745 367160 292314 367162
rect 291745 367104 291750 367160
rect 291806 367104 292314 367160
rect 291745 367102 292314 367104
rect 294045 367160 294154 367165
rect 294045 367104 294050 367160
rect 294106 367104 294154 367160
rect 294045 367102 294154 367104
rect 297222 367162 297282 367374
rect 300117 367432 300226 367434
rect 300117 367376 300122 367432
rect 300178 367376 300226 367432
rect 300117 367371 300226 367376
rect 300166 367165 300226 367371
rect 304030 367432 304139 367434
rect 304030 367376 304078 367432
rect 304134 367376 304139 367432
rect 304030 367371 304139 367376
rect 514753 367434 514819 367437
rect 514753 367432 518052 367434
rect 514753 367376 514758 367432
rect 514814 367376 518052 367432
rect 514753 367374 518052 367376
rect 514753 367371 514819 367374
rect 304030 367165 304090 367371
rect 297357 367162 297423 367165
rect 297222 367160 297423 367162
rect 297222 367104 297362 367160
rect 297418 367104 297423 367160
rect 297222 367102 297423 367104
rect 300166 367160 300275 367165
rect 300166 367104 300214 367160
rect 300270 367104 300275 367160
rect 300166 367102 300275 367104
rect 291745 367099 291811 367102
rect 294045 367099 294111 367102
rect 297357 367099 297423 367102
rect 300209 367099 300275 367102
rect 303981 367160 304090 367165
rect 303981 367104 303986 367160
rect 304042 367104 304090 367160
rect 303981 367102 304090 367104
rect 303981 367099 304047 367102
rect 514753 366074 514819 366077
rect 514753 366072 518052 366074
rect 514753 366016 514758 366072
rect 514814 366016 518052 366072
rect 514753 366014 518052 366016
rect 514753 366011 514819 366014
rect 583520 364972 584960 365212
rect 514753 364714 514819 364717
rect 514753 364712 518052 364714
rect 514753 364656 514758 364712
rect 514814 364656 518052 364712
rect 514753 364654 518052 364656
rect 514753 364651 514819 364654
rect 514753 363354 514819 363357
rect 514753 363352 518052 363354
rect 514753 363296 514758 363352
rect 514814 363296 518052 363352
rect 514753 363294 518052 363296
rect 514753 363291 514819 363294
rect 514753 361994 514819 361997
rect 514753 361992 518052 361994
rect 514753 361936 514758 361992
rect 514814 361936 518052 361992
rect 514753 361934 518052 361936
rect 514753 361931 514819 361934
rect 303797 361586 303863 361589
rect 304901 361586 304967 361589
rect 303797 361584 304967 361586
rect 303797 361528 303802 361584
rect 303858 361528 304906 361584
rect 304962 361528 304967 361584
rect 303797 361526 304967 361528
rect 303797 361523 303863 361526
rect 304901 361523 304967 361526
rect 515489 360634 515555 360637
rect 515489 360632 518052 360634
rect 515489 360576 515494 360632
rect 515550 360576 518052 360632
rect 515489 360574 518052 360576
rect 515489 360571 515555 360574
rect 296713 360226 296779 360229
rect 297633 360226 297699 360229
rect 296713 360224 297699 360226
rect 296713 360168 296718 360224
rect 296774 360168 297638 360224
rect 297694 360168 297699 360224
rect 296713 360166 297699 360168
rect 296713 360163 296779 360166
rect 297633 360163 297699 360166
rect 517421 359410 517487 359413
rect 521653 359410 521719 359413
rect 517421 359408 521719 359410
rect 517421 359352 517426 359408
rect 517482 359352 521658 359408
rect 521714 359352 521719 359408
rect 517421 359350 521719 359352
rect 517421 359347 517487 359350
rect 521653 359347 521719 359350
rect -960 358308 480 358548
rect 529197 351930 529263 351933
rect 583520 351930 584960 352020
rect 529197 351928 584960 351930
rect 529197 351872 529202 351928
rect 529258 351872 584960 351928
rect 529197 351870 584960 351872
rect 529197 351867 529263 351870
rect 583520 351780 584960 351870
rect 291929 348394 291995 348397
rect 299565 348394 299631 348397
rect 291929 348392 299631 348394
rect 291929 348336 291934 348392
rect 291990 348336 299570 348392
rect 299626 348336 299631 348392
rect 291929 348334 299631 348336
rect 291929 348331 291995 348334
rect 299565 348331 299631 348334
rect 299565 347850 299631 347853
rect 308029 347850 308095 347853
rect 299565 347848 308095 347850
rect 299565 347792 299570 347848
rect 299626 347792 308034 347848
rect 308090 347792 308095 347848
rect 299565 347790 308095 347792
rect 299565 347787 299631 347790
rect 308029 347787 308095 347790
rect 291837 346626 291903 346629
rect 296713 346626 296779 346629
rect 291837 346624 297282 346626
rect 291837 346568 291842 346624
rect 291898 346568 296718 346624
rect 296774 346568 297282 346624
rect 291837 346566 297282 346568
rect 291837 346563 291903 346566
rect 296713 346563 296779 346566
rect 297222 346221 297282 346566
rect 304901 346490 304967 346493
rect 307937 346490 308003 346493
rect 304030 346488 308003 346490
rect 304030 346432 304906 346488
rect 304962 346432 307942 346488
rect 307998 346432 308003 346488
rect 304030 346430 308003 346432
rect 304030 346221 304090 346430
rect 304901 346427 304967 346430
rect 307937 346427 308003 346430
rect 297222 346216 297331 346221
rect 297222 346160 297270 346216
rect 297326 346160 297331 346216
rect 297222 346158 297331 346160
rect 297265 346155 297331 346158
rect 303981 346216 304090 346221
rect 303981 346160 303986 346216
rect 304042 346160 304090 346216
rect 303981 346158 304090 346160
rect 303981 346155 304047 346158
rect -960 345252 480 345492
rect 518433 343906 518499 343909
rect 521653 343906 521719 343909
rect 518433 343904 521719 343906
rect 518433 343848 518438 343904
rect 518494 343848 521658 343904
rect 521714 343848 521719 343904
rect 518433 343846 521719 343848
rect 518433 343843 518499 343846
rect 521653 343843 521719 343846
rect 524321 343906 524387 343909
rect 527265 343906 527331 343909
rect 529197 343906 529263 343909
rect 524321 343904 529263 343906
rect 524321 343848 524326 343904
rect 524382 343848 527270 343904
rect 527326 343848 529202 343904
rect 529258 343848 529263 343904
rect 524321 343846 529263 343848
rect 524321 343843 524387 343846
rect 527265 343843 527331 343846
rect 529197 343843 529263 343846
rect 527081 343770 527147 343773
rect 528553 343770 528619 343773
rect 527081 343768 528619 343770
rect 527081 343712 527086 343768
rect 527142 343712 528558 343768
rect 528614 343712 528619 343768
rect 527081 343710 528619 343712
rect 527081 343707 527147 343710
rect 528553 343707 528619 343710
rect 514753 341050 514819 341053
rect 514753 341048 518052 341050
rect 514753 340992 514758 341048
rect 514814 340992 518052 341048
rect 514753 340990 518052 340992
rect 514753 340987 514819 340990
rect 514753 339690 514819 339693
rect 514753 339688 518052 339690
rect 514753 339632 514758 339688
rect 514814 339632 518052 339688
rect 514753 339630 518052 339632
rect 514753 339627 514819 339630
rect 583520 338452 584960 338692
rect 514753 338330 514819 338333
rect 514753 338328 518052 338330
rect 514753 338272 514758 338328
rect 514814 338272 518052 338328
rect 514753 338270 518052 338272
rect 514753 338267 514819 338270
rect 514753 336970 514819 336973
rect 514753 336968 518052 336970
rect 514753 336912 514758 336968
rect 514814 336912 518052 336968
rect 514753 336910 518052 336912
rect 514753 336907 514819 336910
rect 515305 335610 515371 335613
rect 515305 335608 518052 335610
rect 515305 335552 515310 335608
rect 515366 335552 518052 335608
rect 515305 335550 518052 335552
rect 515305 335547 515371 335550
rect 514753 334250 514819 334253
rect 514753 334248 518052 334250
rect 514753 334192 514758 334248
rect 514814 334192 518052 334248
rect 514753 334190 518052 334192
rect 514753 334187 514819 334190
rect 514753 332890 514819 332893
rect 514753 332888 518052 332890
rect 514753 332832 514758 332888
rect 514814 332832 518052 332888
rect 514753 332830 518052 332832
rect 514753 332827 514819 332830
rect -960 332196 480 332436
rect 514753 331530 514819 331533
rect 514753 331528 518052 331530
rect 514753 331472 514758 331528
rect 514814 331472 518052 331528
rect 514753 331470 518052 331472
rect 514753 331467 514819 331470
rect 529933 330986 529999 330989
rect 527804 330984 529999 330986
rect 527804 330928 529938 330984
rect 529994 330928 529999 330984
rect 527804 330926 529999 330928
rect 529933 330923 529999 330926
rect 516041 330170 516107 330173
rect 516041 330168 518052 330170
rect 516041 330112 516046 330168
rect 516102 330112 518052 330168
rect 516041 330110 518052 330112
rect 516041 330107 516107 330110
rect 515765 328810 515831 328813
rect 515765 328808 518052 328810
rect 515765 328752 515770 328808
rect 515826 328752 518052 328808
rect 515765 328750 518052 328752
rect 515765 328747 515831 328750
rect 514753 327450 514819 327453
rect 514753 327448 518052 327450
rect 514753 327392 514758 327448
rect 514814 327392 518052 327448
rect 514753 327390 518052 327392
rect 514753 327387 514819 327390
rect 514753 326090 514819 326093
rect 514753 326088 518052 326090
rect 514753 326032 514758 326088
rect 514814 326032 518052 326088
rect 514753 326030 518052 326032
rect 514753 326027 514819 326030
rect 307661 325818 307727 325821
rect 308581 325818 308647 325821
rect 309593 325818 309659 325821
rect 307661 325816 309659 325818
rect 307661 325760 307666 325816
rect 307722 325760 308586 325816
rect 308642 325760 309598 325816
rect 309654 325760 309659 325816
rect 307661 325758 309659 325760
rect 307661 325755 307727 325758
rect 308581 325755 308647 325758
rect 309593 325755 309659 325758
rect 583520 325124 584960 325364
rect 514753 324730 514819 324733
rect 514753 324728 518052 324730
rect 514753 324672 514758 324728
rect 514814 324672 518052 324728
rect 514753 324670 518052 324672
rect 514753 324667 514819 324670
rect 514753 323370 514819 323373
rect 514753 323368 518052 323370
rect 514753 323312 514758 323368
rect 514814 323312 518052 323368
rect 514753 323310 518052 323312
rect 514753 323307 514819 323310
rect 514753 322010 514819 322013
rect 514753 322008 518052 322010
rect 514753 321952 514758 322008
rect 514814 321952 518052 322008
rect 514753 321950 518052 321952
rect 514753 321947 514819 321950
rect 514753 320650 514819 320653
rect 514753 320648 518052 320650
rect 514753 320592 514758 320648
rect 514814 320592 518052 320648
rect 514753 320590 518052 320592
rect 514753 320587 514819 320590
rect 518433 319426 518499 319429
rect 522297 319426 522363 319429
rect 518433 319424 522363 319426
rect -960 319140 480 319380
rect 518433 319368 518438 319424
rect 518494 319368 522302 319424
rect 522358 319368 522363 319424
rect 518433 319366 522363 319368
rect 518433 319363 518499 319366
rect 522297 319363 522363 319366
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 306005 305826 306071 305829
rect 308489 305826 308555 305829
rect 306005 305824 308555 305826
rect 306005 305768 306010 305824
rect 306066 305768 308494 305824
rect 308550 305768 308555 305824
rect 306005 305766 308555 305768
rect 306005 305763 306071 305766
rect 308489 305763 308555 305766
rect 302417 305690 302483 305693
rect 308397 305690 308463 305693
rect 302417 305688 308463 305690
rect 302417 305632 302422 305688
rect 302478 305632 308402 305688
rect 308458 305632 308463 305688
rect 302417 305630 308463 305632
rect 302417 305627 302483 305630
rect 308397 305627 308463 305630
rect 291929 305146 291995 305149
rect 298461 305146 298527 305149
rect 291929 305144 298527 305146
rect 291929 305088 291934 305144
rect 291990 305088 298466 305144
rect 298522 305088 298527 305144
rect 291929 305086 298527 305088
rect 291929 305083 291995 305086
rect 298461 305083 298527 305086
rect 308489 305146 308555 305149
rect 311893 305146 311959 305149
rect 308489 305144 311959 305146
rect 308489 305088 308494 305144
rect 308550 305088 311898 305144
rect 311954 305088 311959 305144
rect 308489 305086 311959 305088
rect 308489 305083 308555 305086
rect 311893 305083 311959 305086
rect 292389 305010 292455 305013
rect 294965 305010 295031 305013
rect 292389 305008 295031 305010
rect 292389 304952 292394 305008
rect 292450 304952 294970 305008
rect 295026 304952 295031 305008
rect 292389 304950 295031 304952
rect 292389 304947 292455 304950
rect 294965 304947 295031 304950
rect 308397 305010 308463 305013
rect 310513 305010 310579 305013
rect 308397 305008 310579 305010
rect 308397 304952 308402 305008
rect 308458 304952 310518 305008
rect 310574 304952 310579 305008
rect 308397 304950 310579 304952
rect 308397 304947 308463 304950
rect 310513 304947 310579 304950
rect 527081 303786 527147 303789
rect 528553 303786 528619 303789
rect 527081 303784 528619 303786
rect 527081 303728 527086 303784
rect 527142 303728 528558 303784
rect 528614 303728 528619 303784
rect 527081 303726 528619 303728
rect 527081 303723 527147 303726
rect 528553 303723 528619 303726
rect 524321 303650 524387 303653
rect 527265 303650 527331 303653
rect 524321 303648 527331 303650
rect 524321 303592 524326 303648
rect 524382 303592 527270 303648
rect 527326 303592 527331 303648
rect 524321 303590 527331 303592
rect 524321 303587 524387 303590
rect 527265 303587 527331 303590
rect 308673 302290 308739 302293
rect 309501 302290 309567 302293
rect 308673 302288 309567 302290
rect 308673 302232 308678 302288
rect 308734 302232 309506 302288
rect 309562 302232 309567 302288
rect 308673 302230 309567 302232
rect 308673 302227 308739 302230
rect 309501 302227 309567 302230
rect 522113 302290 522179 302293
rect 528645 302290 528711 302293
rect 580165 302290 580231 302293
rect 522113 302288 580231 302290
rect 522113 302232 522118 302288
rect 522174 302232 528650 302288
rect 528706 302232 580170 302288
rect 580226 302232 580231 302288
rect 522113 302230 580231 302232
rect 522113 302227 522179 302230
rect 528645 302227 528711 302230
rect 580165 302227 580231 302230
rect 514753 301066 514819 301069
rect 514753 301064 518052 301066
rect 514753 301008 514758 301064
rect 514814 301008 518052 301064
rect 514753 301006 518052 301008
rect 514753 301003 514819 301006
rect 515029 299706 515095 299709
rect 515029 299704 518052 299706
rect 515029 299648 515034 299704
rect 515090 299648 518052 299704
rect 515029 299646 518052 299648
rect 515029 299643 515095 299646
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 514937 298346 515003 298349
rect 514937 298344 518052 298346
rect 514937 298288 514942 298344
rect 514998 298288 518052 298344
rect 514937 298286 518052 298288
rect 514937 298283 515003 298286
rect 514753 296986 514819 296989
rect 514753 296984 518052 296986
rect 514753 296928 514758 296984
rect 514814 296928 518052 296984
rect 514753 296926 518052 296928
rect 514753 296923 514819 296926
rect 514753 295626 514819 295629
rect 514753 295624 518052 295626
rect 514753 295568 514758 295624
rect 514814 295568 518052 295624
rect 514753 295566 518052 295568
rect 514753 295563 514819 295566
rect 514753 294266 514819 294269
rect 514753 294264 518052 294266
rect 514753 294208 514758 294264
rect 514814 294208 518052 294264
rect 514753 294206 518052 294208
rect 514753 294203 514819 294206
rect -960 293028 480 293268
rect 515949 292906 516015 292909
rect 515949 292904 518052 292906
rect 515949 292848 515954 292904
rect 516010 292848 518052 292904
rect 515949 292846 518052 292848
rect 515949 292843 516015 292846
rect 515673 291546 515739 291549
rect 515673 291544 518052 291546
rect 515673 291488 515678 291544
rect 515734 291488 518052 291544
rect 515673 291486 518052 291488
rect 515673 291483 515739 291486
rect 529933 291002 529999 291005
rect 527804 291000 529999 291002
rect 527804 290944 529938 291000
rect 529994 290944 529999 291000
rect 527804 290942 529999 290944
rect 529933 290939 529999 290942
rect 514753 290186 514819 290189
rect 514753 290184 518052 290186
rect 514753 290128 514758 290184
rect 514814 290128 518052 290184
rect 514753 290126 518052 290128
rect 514753 290123 514819 290126
rect 514753 288826 514819 288829
rect 514753 288824 518052 288826
rect 514753 288768 514758 288824
rect 514814 288768 518052 288824
rect 514753 288766 518052 288768
rect 514753 288763 514819 288766
rect 515949 287466 516015 287469
rect 515949 287464 518052 287466
rect 515949 287408 515954 287464
rect 516010 287408 518052 287464
rect 515949 287406 518052 287408
rect 515949 287403 516015 287406
rect 515857 286106 515923 286109
rect 515857 286104 518052 286106
rect 515857 286048 515862 286104
rect 515918 286048 518052 286104
rect 515857 286046 518052 286048
rect 515857 286043 515923 286046
rect 309133 285698 309199 285701
rect 311893 285698 311959 285701
rect 309133 285696 311959 285698
rect 309133 285640 309138 285696
rect 309194 285640 311898 285696
rect 311954 285640 311959 285696
rect 309133 285638 311959 285640
rect 309133 285635 309199 285638
rect 311893 285635 311959 285638
rect 583520 285276 584960 285516
rect 514753 284746 514819 284749
rect 514753 284744 518052 284746
rect 514753 284688 514758 284744
rect 514814 284688 518052 284744
rect 514753 284686 518052 284688
rect 514753 284683 514819 284686
rect 304901 284474 304967 284477
rect 309133 284474 309199 284477
rect 304901 284472 309199 284474
rect 304901 284416 304906 284472
rect 304962 284416 309138 284472
rect 309194 284416 309199 284472
rect 304901 284414 309199 284416
rect 304901 284411 304967 284414
rect 309133 284411 309199 284414
rect 301681 284338 301747 284341
rect 309317 284338 309383 284341
rect 310513 284338 310579 284341
rect 301681 284336 310579 284338
rect 301681 284280 301686 284336
rect 301742 284280 309322 284336
rect 309378 284280 310518 284336
rect 310574 284280 310579 284336
rect 301681 284278 310579 284280
rect 301681 284275 301747 284278
rect 309317 284275 309383 284278
rect 310513 284275 310579 284278
rect 291837 283522 291903 283525
rect 295241 283522 295307 283525
rect 301681 283522 301747 283525
rect 291837 283520 295307 283522
rect 291837 283464 291842 283520
rect 291898 283464 295246 283520
rect 295302 283464 295307 283520
rect 291837 283462 295307 283464
rect 291837 283459 291903 283462
rect 295241 283459 295307 283462
rect 301638 283520 301747 283522
rect 301638 283464 301686 283520
rect 301742 283464 301747 283520
rect 301638 283459 301747 283464
rect 304901 283522 304967 283525
rect 304901 283520 305010 283522
rect 304901 283464 304906 283520
rect 304962 283464 305010 283520
rect 304901 283459 305010 283464
rect 301638 283117 301698 283459
rect 304950 283117 305010 283459
rect 515765 283386 515831 283389
rect 515765 283384 518052 283386
rect 515765 283328 515770 283384
rect 515826 283328 518052 283384
rect 515765 283326 518052 283328
rect 515765 283323 515831 283326
rect 301586 283112 301698 283117
rect 301586 283056 301591 283112
rect 301647 283056 301698 283112
rect 301586 283054 301698 283056
rect 304903 283112 305010 283117
rect 304903 283056 304908 283112
rect 304964 283056 305010 283112
rect 304903 283054 305010 283056
rect 301586 283051 301652 283054
rect 304903 283051 304969 283054
rect 515673 282026 515739 282029
rect 515673 282024 518052 282026
rect 515673 281968 515678 282024
rect 515734 281968 518052 282024
rect 515673 281966 518052 281968
rect 515673 281963 515739 281966
rect 515581 280666 515647 280669
rect 515581 280664 518052 280666
rect 515581 280608 515586 280664
rect 515642 280608 518052 280664
rect 515581 280606 518052 280608
rect 515581 280603 515647 280606
rect -960 279972 480 280212
rect 517421 278898 517487 278901
rect 519537 278898 519603 278901
rect 517421 278896 519603 278898
rect 517421 278840 517426 278896
rect 517482 278840 519542 278896
rect 519598 278840 519603 278896
rect 517421 278838 519603 278840
rect 517421 278835 517487 278838
rect 519537 278835 519603 278838
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 527081 264890 527147 264893
rect 528553 264890 528619 264893
rect 527081 264888 528619 264890
rect 527081 264832 527086 264888
rect 527142 264832 528558 264888
rect 528614 264832 528619 264888
rect 527081 264830 528619 264832
rect 527081 264827 527147 264830
rect 528553 264827 528619 264830
rect 524321 264618 524387 264621
rect 527265 264618 527331 264621
rect 524321 264616 527331 264618
rect 524321 264560 524326 264616
rect 524382 264560 527270 264616
rect 527326 264560 527331 264616
rect 524321 264558 527331 264560
rect 524321 264555 524387 264558
rect 527265 264555 527331 264558
rect 522113 264482 522179 264485
rect 528645 264482 528711 264485
rect 522113 264480 528711 264482
rect 522113 264424 522118 264480
rect 522174 264424 528650 264480
rect 528706 264424 528711 264480
rect 522113 264422 528711 264424
rect 522113 264419 522179 264422
rect 528645 264419 528711 264422
rect 305913 263802 305979 263805
rect 309317 263802 309383 263805
rect 305913 263800 309383 263802
rect 305913 263744 305918 263800
rect 305974 263744 309322 263800
rect 309378 263744 309383 263800
rect 305913 263742 309383 263744
rect 305913 263739 305979 263742
rect 309317 263739 309383 263742
rect 302141 263666 302207 263669
rect 309225 263666 309291 263669
rect 309869 263666 309935 263669
rect 302141 263664 309935 263666
rect 302141 263608 302146 263664
rect 302202 263608 309230 263664
rect 309286 263608 309874 263664
rect 309930 263608 309935 263664
rect 302141 263606 309935 263608
rect 302141 263603 302207 263606
rect 309225 263603 309291 263606
rect 309869 263603 309935 263606
rect 519629 263666 519695 263669
rect 527817 263666 527883 263669
rect 519629 263664 527883 263666
rect 519629 263608 519634 263664
rect 519690 263608 527822 263664
rect 527878 263608 527883 263664
rect 519629 263606 527883 263608
rect 519629 263603 519695 263606
rect 527817 263603 527883 263606
rect 302141 262578 302207 262581
rect 302141 262576 302250 262578
rect 302141 262520 302146 262576
rect 302202 262520 302250 262576
rect 302141 262515 302250 262520
rect 305913 262576 305979 262581
rect 309041 262578 309107 262581
rect 305913 262520 305918 262576
rect 305974 262520 305979 262576
rect 305913 262515 305979 262520
rect 308998 262576 309107 262578
rect 308998 262520 309046 262576
rect 309102 262520 309107 262576
rect 308998 262515 309107 262520
rect 309317 262578 309383 262581
rect 309317 262576 309426 262578
rect 309317 262520 309322 262576
rect 309378 262520 309426 262576
rect 309317 262515 309426 262520
rect 301937 262170 302003 262173
rect 302190 262170 302250 262515
rect 301937 262168 302250 262170
rect 301937 262112 301942 262168
rect 301998 262112 302250 262168
rect 301937 262110 302250 262112
rect 305381 262170 305447 262173
rect 305916 262170 305976 262515
rect 305381 262168 305976 262170
rect 305381 262112 305386 262168
rect 305442 262112 305976 262168
rect 305381 262110 305976 262112
rect 301937 262107 302003 262110
rect 305381 262107 305447 262110
rect 308825 262034 308891 262037
rect 308998 262034 309058 262515
rect 309366 262173 309426 262515
rect 309317 262168 309426 262173
rect 309317 262112 309322 262168
rect 309378 262112 309426 262168
rect 309317 262110 309426 262112
rect 309317 262107 309383 262110
rect 308825 262032 309058 262034
rect 308825 261976 308830 262032
rect 308886 261976 309058 262032
rect 308825 261974 309058 261976
rect 308825 261971 308891 261974
rect 514753 261082 514819 261085
rect 514753 261080 518052 261082
rect 514753 261024 514758 261080
rect 514814 261024 518052 261080
rect 514753 261022 518052 261024
rect 514753 261019 514819 261022
rect 514753 259722 514819 259725
rect 514753 259720 518052 259722
rect 514753 259664 514758 259720
rect 514814 259664 518052 259720
rect 514753 259662 518052 259664
rect 514753 259659 514819 259662
rect 583520 258756 584960 258996
rect 514753 258362 514819 258365
rect 514753 258360 518052 258362
rect 514753 258304 514758 258360
rect 514814 258304 518052 258360
rect 514753 258302 518052 258304
rect 514753 258299 514819 258302
rect 514753 257002 514819 257005
rect 514753 257000 518052 257002
rect 514753 256944 514758 257000
rect 514814 256944 518052 257000
rect 514753 256942 518052 256944
rect 514753 256939 514819 256942
rect 514753 255642 514819 255645
rect 514753 255640 518052 255642
rect 514753 255584 514758 255640
rect 514814 255584 518052 255640
rect 514753 255582 518052 255584
rect 514753 255579 514819 255582
rect 514753 254282 514819 254285
rect 514753 254280 518052 254282
rect -960 253996 480 254236
rect 514753 254224 514758 254280
rect 514814 254224 518052 254280
rect 514753 254222 518052 254224
rect 514753 254219 514819 254222
rect 514753 252922 514819 252925
rect 514753 252920 518052 252922
rect 514753 252864 514758 252920
rect 514814 252864 518052 252920
rect 514753 252862 518052 252864
rect 514753 252859 514819 252862
rect 514753 251562 514819 251565
rect 514753 251560 518052 251562
rect 514753 251504 514758 251560
rect 514814 251504 518052 251560
rect 514753 251502 518052 251504
rect 514753 251499 514819 251502
rect 529933 251018 529999 251021
rect 530577 251018 530643 251021
rect 527804 251016 530643 251018
rect 527804 250960 529938 251016
rect 529994 250960 530582 251016
rect 530638 250960 530643 251016
rect 527804 250958 530643 250960
rect 529933 250955 529999 250958
rect 530577 250955 530643 250958
rect 304901 250474 304967 250477
rect 309225 250474 309291 250477
rect 304901 250472 309291 250474
rect 304901 250416 304906 250472
rect 304962 250416 309230 250472
rect 309286 250416 309291 250472
rect 304901 250414 309291 250416
rect 304901 250411 304967 250414
rect 309225 250411 309291 250414
rect 514753 250202 514819 250205
rect 514753 250200 518052 250202
rect 514753 250144 514758 250200
rect 514814 250144 518052 250200
rect 514753 250142 518052 250144
rect 514753 250139 514819 250142
rect 514753 248842 514819 248845
rect 514753 248840 518052 248842
rect 514753 248784 514758 248840
rect 514814 248784 518052 248840
rect 514753 248782 518052 248784
rect 514753 248779 514819 248782
rect 514753 247482 514819 247485
rect 514753 247480 518052 247482
rect 514753 247424 514758 247480
rect 514814 247424 518052 247480
rect 514753 247422 518052 247424
rect 514753 247419 514819 247422
rect 514753 246122 514819 246125
rect 514753 246120 518052 246122
rect 514753 246064 514758 246120
rect 514814 246064 518052 246120
rect 514753 246062 518052 246064
rect 514753 246059 514819 246062
rect 527817 245578 527883 245581
rect 583520 245578 584960 245668
rect 527817 245576 584960 245578
rect 527817 245520 527822 245576
rect 527878 245520 584960 245576
rect 527817 245518 584960 245520
rect 527817 245515 527883 245518
rect 583520 245428 584960 245518
rect 514937 244762 515003 244765
rect 514937 244760 518052 244762
rect 514937 244704 514942 244760
rect 514998 244704 518052 244760
rect 514937 244702 518052 244704
rect 514937 244699 515003 244702
rect 514753 243402 514819 243405
rect 514753 243400 518052 243402
rect 514753 243344 514758 243400
rect 514814 243344 518052 243400
rect 514753 243342 518052 243344
rect 514753 243339 514819 243342
rect 301497 242994 301563 242997
rect 309133 242994 309199 242997
rect 309869 242994 309935 242997
rect 301497 242992 309935 242994
rect 301497 242936 301502 242992
rect 301558 242936 309138 242992
rect 309194 242936 309874 242992
rect 309930 242936 309935 242992
rect 301497 242934 309935 242936
rect 301497 242931 301563 242934
rect 309133 242931 309199 242934
rect 309869 242931 309935 242934
rect 515949 242042 516015 242045
rect 515949 242040 518052 242042
rect 515949 241984 515954 242040
rect 516010 241984 518052 242040
rect 515949 241982 518052 241984
rect 515949 241979 516015 241982
rect 301497 241498 301563 241501
rect 304809 241498 304875 241501
rect 301454 241496 301563 241498
rect 301454 241440 301502 241496
rect 301558 241440 301563 241496
rect 301454 241435 301563 241440
rect 304766 241496 304875 241498
rect 304766 241440 304814 241496
rect 304870 241440 304875 241496
rect 304766 241435 304875 241440
rect 301454 241229 301514 241435
rect 304766 241229 304826 241435
rect 301405 241224 301514 241229
rect -960 240940 480 241180
rect 301405 241168 301410 241224
rect 301466 241168 301514 241224
rect 301405 241166 301514 241168
rect 304717 241224 304826 241229
rect 304717 241168 304722 241224
rect 304778 241168 304826 241224
rect 304717 241166 304826 241168
rect 301405 241163 301471 241166
rect 304717 241163 304783 241166
rect 515857 240682 515923 240685
rect 515857 240680 518052 240682
rect 515857 240624 515862 240680
rect 515918 240624 518052 240680
rect 515857 240622 518052 240624
rect 515857 240619 515923 240622
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 306833 223546 306899 223549
rect 309225 223546 309291 223549
rect 306833 223544 309291 223546
rect 306833 223488 306838 223544
rect 306894 223488 309230 223544
rect 309286 223488 309291 223544
rect 306833 223486 309291 223488
rect 306833 223483 306899 223486
rect 309225 223483 309291 223486
rect 302785 222866 302851 222869
rect 309133 222866 309199 222869
rect 311893 222866 311959 222869
rect 302785 222864 311959 222866
rect 302785 222808 302790 222864
rect 302846 222808 309138 222864
rect 309194 222808 311898 222864
rect 311954 222808 311959 222864
rect 302785 222806 311959 222808
rect 302785 222803 302851 222806
rect 309133 222803 309199 222806
rect 311893 222803 311959 222806
rect 307937 222730 308003 222733
rect 309685 222730 309751 222733
rect 307937 222728 309751 222730
rect 307937 222672 307942 222728
rect 307998 222672 309690 222728
rect 309746 222672 309751 222728
rect 307937 222670 309751 222672
rect 307937 222667 308003 222670
rect 309685 222667 309751 222670
rect 302785 220418 302851 220421
rect 306833 220418 306899 220421
rect 302742 220416 302851 220418
rect 302742 220360 302790 220416
rect 302846 220360 302851 220416
rect 302742 220355 302851 220360
rect 306790 220416 306899 220418
rect 306790 220360 306838 220416
rect 306894 220360 306899 220416
rect 306790 220355 306899 220360
rect 309685 220418 309751 220421
rect 309685 220416 309794 220418
rect 309685 220360 309690 220416
rect 309746 220360 309794 220416
rect 309685 220355 309794 220360
rect 302742 220013 302802 220355
rect 306790 220149 306850 220355
rect 306741 220144 306850 220149
rect 306741 220088 306746 220144
rect 306802 220088 306850 220144
rect 306741 220086 306850 220088
rect 309734 220149 309794 220355
rect 309734 220144 309843 220149
rect 309734 220088 309782 220144
rect 309838 220088 309843 220144
rect 309734 220086 309843 220088
rect 306741 220083 306807 220086
rect 309777 220083 309843 220086
rect 302740 220008 302806 220013
rect 302740 219952 302745 220008
rect 302801 219952 302806 220008
rect 302740 219947 302806 219952
rect 583520 218908 584960 219148
rect 291837 218514 291903 218517
rect 294689 218514 294755 218517
rect 291837 218512 294755 218514
rect 291837 218456 291842 218512
rect 291898 218456 294694 218512
rect 294750 218456 294755 218512
rect 291837 218454 294755 218456
rect 291837 218451 291903 218454
rect 294689 218451 294755 218454
rect 304901 217834 304967 217837
rect 306373 217834 306439 217837
rect 304901 217832 306439 217834
rect 304901 217776 304906 217832
rect 304962 217776 306378 217832
rect 306434 217776 306439 217832
rect 304901 217774 306439 217776
rect 304901 217771 304967 217774
rect 306373 217771 306439 217774
rect 306925 217834 306991 217837
rect 310145 217834 310211 217837
rect 306925 217832 310211 217834
rect 306925 217776 306930 217832
rect 306986 217776 310150 217832
rect 310206 217776 310211 217832
rect 306925 217774 310211 217776
rect 306925 217771 306991 217774
rect 310145 217771 310211 217774
rect -960 214828 480 215068
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 300761 200698 300827 200701
rect 311893 200698 311959 200701
rect 300761 200696 311959 200698
rect 300761 200640 300766 200696
rect 300822 200640 311898 200696
rect 311954 200640 311959 200696
rect 300761 200638 311959 200640
rect 300761 200635 300827 200638
rect 311893 200635 311959 200638
rect 291837 200290 291903 200293
rect 300761 200290 300827 200293
rect 291837 200288 300827 200290
rect 291837 200232 291842 200288
rect 291898 200232 300766 200288
rect 300822 200232 300827 200288
rect 291837 200230 300827 200232
rect 291837 200227 291903 200230
rect 300761 200227 300827 200230
rect 291745 200154 291811 200157
rect 297541 200154 297607 200157
rect 291745 200152 297607 200154
rect 291745 200096 291750 200152
rect 291806 200096 297546 200152
rect 297602 200096 297607 200152
rect 291745 200094 297607 200096
rect 291745 200091 291811 200094
rect 297541 200091 297607 200094
rect 294689 199474 294755 199477
rect 293542 199472 294755 199474
rect 293542 199416 294694 199472
rect 294750 199416 294755 199472
rect 293542 199414 294755 199416
rect 292481 198794 292547 198797
rect 293542 198794 293602 199414
rect 294689 199411 294755 199414
rect 306925 199474 306991 199477
rect 306925 199472 307034 199474
rect 306925 199416 306930 199472
rect 306986 199416 307034 199472
rect 306925 199411 307034 199416
rect 306974 199202 307034 199411
rect 307569 199202 307635 199205
rect 306974 199200 307635 199202
rect 306974 199144 307574 199200
rect 307630 199144 307635 199200
rect 306974 199142 307635 199144
rect 307569 199139 307635 199142
rect 293677 198794 293743 198797
rect 292481 198792 293743 198794
rect 292481 198736 292486 198792
rect 292542 198736 293682 198792
rect 293738 198736 293743 198792
rect 292481 198734 293743 198736
rect 292481 198731 292547 198734
rect 293677 198731 293743 198734
rect 303981 197434 304047 197437
rect 304809 197434 304875 197437
rect 303981 197432 304875 197434
rect 303981 197376 303986 197432
rect 304042 197376 304814 197432
rect 304870 197376 304875 197432
rect 303981 197374 304875 197376
rect 303981 197371 304047 197374
rect 304809 197371 304875 197374
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 291745 180298 291811 180301
rect 296713 180298 296779 180301
rect 298001 180298 298067 180301
rect 291745 180296 298067 180298
rect 291745 180240 291750 180296
rect 291806 180240 296718 180296
rect 296774 180240 298006 180296
rect 298062 180240 298067 180296
rect 291745 180238 298067 180240
rect 291745 180235 291811 180238
rect 296713 180235 296779 180238
rect 298001 180235 298067 180238
rect 291837 180026 291903 180029
rect 306925 180026 306991 180029
rect 307753 180026 307819 180029
rect 367737 180026 367803 180029
rect 291837 180024 300778 180026
rect 291837 179968 291842 180024
rect 291898 179968 300778 180024
rect 291837 179966 300778 179968
rect 291837 179963 291903 179966
rect 300718 179757 300778 179966
rect 306925 180024 367803 180026
rect 306925 179968 306930 180024
rect 306986 179968 307758 180024
rect 307814 179968 367742 180024
rect 367798 179968 367803 180024
rect 306925 179966 367803 179968
rect 306925 179963 306991 179966
rect 307753 179963 307819 179966
rect 367737 179963 367803 179966
rect 304533 179890 304599 179893
rect 364977 179890 365043 179893
rect 304533 179888 365043 179890
rect 304533 179832 304538 179888
rect 304594 179832 364982 179888
rect 365038 179832 365043 179888
rect 304533 179830 365043 179832
rect 304533 179827 304599 179830
rect 364977 179827 365043 179830
rect 300718 179754 300827 179757
rect 308765 179754 308831 179757
rect 300718 179752 308831 179754
rect 300718 179696 300766 179752
rect 300822 179696 308770 179752
rect 308826 179696 308831 179752
rect 300718 179694 308831 179696
rect 300761 179691 300827 179694
rect 308765 179691 308831 179694
rect 298001 179618 298067 179621
rect 308581 179618 308647 179621
rect 298001 179616 308647 179618
rect 298001 179560 298006 179616
rect 298062 179560 308586 179616
rect 308642 179560 308647 179616
rect 298001 179558 308647 179560
rect 298001 179555 298067 179558
rect 308581 179555 308647 179558
rect 292481 179482 292547 179485
rect 293953 179482 294019 179485
rect 308397 179482 308463 179485
rect 292481 179480 308463 179482
rect 292481 179424 292486 179480
rect 292542 179424 293958 179480
rect 294014 179424 308402 179480
rect 308458 179424 308463 179480
rect 292481 179422 308463 179424
rect 292481 179419 292547 179422
rect 293953 179419 294019 179422
rect 308397 179419 308463 179422
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 367737 165882 367803 165885
rect 583520 165882 584960 165972
rect 367737 165880 584960 165882
rect 367737 165824 367742 165880
rect 367798 165824 584960 165880
rect 367737 165822 584960 165824
rect 367737 165819 367803 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 364977 126034 365043 126037
rect 583520 126034 584960 126124
rect 364977 126032 584960 126034
rect 364977 125976 364982 126032
rect 365038 125976 584960 126032
rect 364977 125974 584960 125976
rect 364977 125971 365043 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 308765 86186 308831 86189
rect 583520 86186 584960 86276
rect 308765 86184 584960 86186
rect 308765 86128 308770 86184
rect 308826 86128 584960 86184
rect 308765 86126 584960 86128
rect 308765 86123 308831 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 308581 46338 308647 46341
rect 583520 46338 584960 46428
rect 308581 46336 584960 46338
rect 308581 46280 308586 46336
rect 308642 46280 584960 46336
rect 308581 46278 584960 46280
rect 308581 46275 308647 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 530577 19818 530643 19821
rect 583520 19818 584960 19908
rect 530577 19816 584960 19818
rect 530577 19760 530582 19816
rect 530638 19760 584960 19816
rect 530577 19758 584960 19760
rect 530577 19755 530643 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect 308397 6626 308463 6629
rect 583520 6626 584960 6716
rect 308397 6624 584960 6626
rect -960 6340 480 6580
rect 308397 6568 308402 6624
rect 308458 6568 584960 6624
rect 308397 6566 584960 6568
rect 308397 6563 308463 6566
rect 583520 6476 584960 6566
<< metal4 >>
rect -4950 696434 -3538 707814
rect -4950 696198 -4842 696434
rect -4606 696198 -4522 696434
rect -4286 696198 -4202 696434
rect -3966 696198 -3882 696434
rect -3646 696198 -3538 696434
rect -4950 689434 -3538 696198
rect -4950 689198 -4842 689434
rect -4606 689198 -4522 689434
rect -4286 689198 -4202 689434
rect -3966 689198 -3882 689434
rect -3646 689198 -3538 689434
rect -4950 682434 -3538 689198
rect -4950 682198 -4842 682434
rect -4606 682198 -4522 682434
rect -4286 682198 -4202 682434
rect -3966 682198 -3882 682434
rect -3646 682198 -3538 682434
rect -4950 675434 -3538 682198
rect -4950 675198 -4842 675434
rect -4606 675198 -4522 675434
rect -4286 675198 -4202 675434
rect -3966 675198 -3882 675434
rect -3646 675198 -3538 675434
rect -4950 668434 -3538 675198
rect -4950 668198 -4842 668434
rect -4606 668198 -4522 668434
rect -4286 668198 -4202 668434
rect -3966 668198 -3882 668434
rect -3646 668198 -3538 668434
rect -4950 661434 -3538 668198
rect -4950 661198 -4842 661434
rect -4606 661198 -4522 661434
rect -4286 661198 -4202 661434
rect -3966 661198 -3882 661434
rect -3646 661198 -3538 661434
rect -4950 654434 -3538 661198
rect -4950 654198 -4842 654434
rect -4606 654198 -4522 654434
rect -4286 654198 -4202 654434
rect -3966 654198 -3882 654434
rect -3646 654198 -3538 654434
rect -4950 647434 -3538 654198
rect -4950 647198 -4842 647434
rect -4606 647198 -4522 647434
rect -4286 647198 -4202 647434
rect -3966 647198 -3882 647434
rect -3646 647198 -3538 647434
rect -4950 640434 -3538 647198
rect -4950 640198 -4842 640434
rect -4606 640198 -4522 640434
rect -4286 640198 -4202 640434
rect -3966 640198 -3882 640434
rect -3646 640198 -3538 640434
rect -4950 633434 -3538 640198
rect -4950 633198 -4842 633434
rect -4606 633198 -4522 633434
rect -4286 633198 -4202 633434
rect -3966 633198 -3882 633434
rect -3646 633198 -3538 633434
rect -4950 626434 -3538 633198
rect -4950 626198 -4842 626434
rect -4606 626198 -4522 626434
rect -4286 626198 -4202 626434
rect -3966 626198 -3882 626434
rect -3646 626198 -3538 626434
rect -4950 619434 -3538 626198
rect -4950 619198 -4842 619434
rect -4606 619198 -4522 619434
rect -4286 619198 -4202 619434
rect -3966 619198 -3882 619434
rect -3646 619198 -3538 619434
rect -4950 612434 -3538 619198
rect -4950 612198 -4842 612434
rect -4606 612198 -4522 612434
rect -4286 612198 -4202 612434
rect -3966 612198 -3882 612434
rect -3646 612198 -3538 612434
rect -4950 605434 -3538 612198
rect -4950 605198 -4842 605434
rect -4606 605198 -4522 605434
rect -4286 605198 -4202 605434
rect -3966 605198 -3882 605434
rect -3646 605198 -3538 605434
rect -4950 598434 -3538 605198
rect -4950 598198 -4842 598434
rect -4606 598198 -4522 598434
rect -4286 598198 -4202 598434
rect -3966 598198 -3882 598434
rect -3646 598198 -3538 598434
rect -4950 591434 -3538 598198
rect -4950 591198 -4842 591434
rect -4606 591198 -4522 591434
rect -4286 591198 -4202 591434
rect -3966 591198 -3882 591434
rect -3646 591198 -3538 591434
rect -4950 584434 -3538 591198
rect -4950 584198 -4842 584434
rect -4606 584198 -4522 584434
rect -4286 584198 -4202 584434
rect -3966 584198 -3882 584434
rect -3646 584198 -3538 584434
rect -4950 577434 -3538 584198
rect -4950 577198 -4842 577434
rect -4606 577198 -4522 577434
rect -4286 577198 -4202 577434
rect -3966 577198 -3882 577434
rect -3646 577198 -3538 577434
rect -4950 570434 -3538 577198
rect -4950 570198 -4842 570434
rect -4606 570198 -4522 570434
rect -4286 570198 -4202 570434
rect -3966 570198 -3882 570434
rect -3646 570198 -3538 570434
rect -4950 563434 -3538 570198
rect -4950 563198 -4842 563434
rect -4606 563198 -4522 563434
rect -4286 563198 -4202 563434
rect -3966 563198 -3882 563434
rect -3646 563198 -3538 563434
rect -4950 556434 -3538 563198
rect -4950 556198 -4842 556434
rect -4606 556198 -4522 556434
rect -4286 556198 -4202 556434
rect -3966 556198 -3882 556434
rect -3646 556198 -3538 556434
rect -4950 549434 -3538 556198
rect -4950 549198 -4842 549434
rect -4606 549198 -4522 549434
rect -4286 549198 -4202 549434
rect -3966 549198 -3882 549434
rect -3646 549198 -3538 549434
rect -4950 542434 -3538 549198
rect -4950 542198 -4842 542434
rect -4606 542198 -4522 542434
rect -4286 542198 -4202 542434
rect -3966 542198 -3882 542434
rect -3646 542198 -3538 542434
rect -4950 535434 -3538 542198
rect -4950 535198 -4842 535434
rect -4606 535198 -4522 535434
rect -4286 535198 -4202 535434
rect -3966 535198 -3882 535434
rect -3646 535198 -3538 535434
rect -4950 528434 -3538 535198
rect -4950 528198 -4842 528434
rect -4606 528198 -4522 528434
rect -4286 528198 -4202 528434
rect -3966 528198 -3882 528434
rect -3646 528198 -3538 528434
rect -4950 521434 -3538 528198
rect -4950 521198 -4842 521434
rect -4606 521198 -4522 521434
rect -4286 521198 -4202 521434
rect -3966 521198 -3882 521434
rect -3646 521198 -3538 521434
rect -4950 514434 -3538 521198
rect -4950 514198 -4842 514434
rect -4606 514198 -4522 514434
rect -4286 514198 -4202 514434
rect -3966 514198 -3882 514434
rect -3646 514198 -3538 514434
rect -4950 507434 -3538 514198
rect -4950 507198 -4842 507434
rect -4606 507198 -4522 507434
rect -4286 507198 -4202 507434
rect -3966 507198 -3882 507434
rect -3646 507198 -3538 507434
rect -4950 500434 -3538 507198
rect -4950 500198 -4842 500434
rect -4606 500198 -4522 500434
rect -4286 500198 -4202 500434
rect -3966 500198 -3882 500434
rect -3646 500198 -3538 500434
rect -4950 493434 -3538 500198
rect -4950 493198 -4842 493434
rect -4606 493198 -4522 493434
rect -4286 493198 -4202 493434
rect -3966 493198 -3882 493434
rect -3646 493198 -3538 493434
rect -4950 486434 -3538 493198
rect -4950 486198 -4842 486434
rect -4606 486198 -4522 486434
rect -4286 486198 -4202 486434
rect -3966 486198 -3882 486434
rect -3646 486198 -3538 486434
rect -4950 479434 -3538 486198
rect -4950 479198 -4842 479434
rect -4606 479198 -4522 479434
rect -4286 479198 -4202 479434
rect -3966 479198 -3882 479434
rect -3646 479198 -3538 479434
rect -4950 472434 -3538 479198
rect -4950 472198 -4842 472434
rect -4606 472198 -4522 472434
rect -4286 472198 -4202 472434
rect -3966 472198 -3882 472434
rect -3646 472198 -3538 472434
rect -4950 465434 -3538 472198
rect -4950 465198 -4842 465434
rect -4606 465198 -4522 465434
rect -4286 465198 -4202 465434
rect -3966 465198 -3882 465434
rect -3646 465198 -3538 465434
rect -4950 458434 -3538 465198
rect -4950 458198 -4842 458434
rect -4606 458198 -4522 458434
rect -4286 458198 -4202 458434
rect -3966 458198 -3882 458434
rect -3646 458198 -3538 458434
rect -4950 451434 -3538 458198
rect -4950 451198 -4842 451434
rect -4606 451198 -4522 451434
rect -4286 451198 -4202 451434
rect -3966 451198 -3882 451434
rect -3646 451198 -3538 451434
rect -4950 444434 -3538 451198
rect -4950 444198 -4842 444434
rect -4606 444198 -4522 444434
rect -4286 444198 -4202 444434
rect -3966 444198 -3882 444434
rect -3646 444198 -3538 444434
rect -4950 437434 -3538 444198
rect -4950 437198 -4842 437434
rect -4606 437198 -4522 437434
rect -4286 437198 -4202 437434
rect -3966 437198 -3882 437434
rect -3646 437198 -3538 437434
rect -4950 430434 -3538 437198
rect -4950 430198 -4842 430434
rect -4606 430198 -4522 430434
rect -4286 430198 -4202 430434
rect -3966 430198 -3882 430434
rect -3646 430198 -3538 430434
rect -4950 423434 -3538 430198
rect -4950 423198 -4842 423434
rect -4606 423198 -4522 423434
rect -4286 423198 -4202 423434
rect -3966 423198 -3882 423434
rect -3646 423198 -3538 423434
rect -4950 416434 -3538 423198
rect -4950 416198 -4842 416434
rect -4606 416198 -4522 416434
rect -4286 416198 -4202 416434
rect -3966 416198 -3882 416434
rect -3646 416198 -3538 416434
rect -4950 409434 -3538 416198
rect -4950 409198 -4842 409434
rect -4606 409198 -4522 409434
rect -4286 409198 -4202 409434
rect -3966 409198 -3882 409434
rect -3646 409198 -3538 409434
rect -4950 402434 -3538 409198
rect -4950 402198 -4842 402434
rect -4606 402198 -4522 402434
rect -4286 402198 -4202 402434
rect -3966 402198 -3882 402434
rect -3646 402198 -3538 402434
rect -4950 395434 -3538 402198
rect -4950 395198 -4842 395434
rect -4606 395198 -4522 395434
rect -4286 395198 -4202 395434
rect -3966 395198 -3882 395434
rect -3646 395198 -3538 395434
rect -4950 388434 -3538 395198
rect -4950 388198 -4842 388434
rect -4606 388198 -4522 388434
rect -4286 388198 -4202 388434
rect -3966 388198 -3882 388434
rect -3646 388198 -3538 388434
rect -4950 381434 -3538 388198
rect -4950 381198 -4842 381434
rect -4606 381198 -4522 381434
rect -4286 381198 -4202 381434
rect -3966 381198 -3882 381434
rect -3646 381198 -3538 381434
rect -4950 374434 -3538 381198
rect -4950 374198 -4842 374434
rect -4606 374198 -4522 374434
rect -4286 374198 -4202 374434
rect -3966 374198 -3882 374434
rect -3646 374198 -3538 374434
rect -4950 367434 -3538 374198
rect -4950 367198 -4842 367434
rect -4606 367198 -4522 367434
rect -4286 367198 -4202 367434
rect -3966 367198 -3882 367434
rect -3646 367198 -3538 367434
rect -4950 360434 -3538 367198
rect -4950 360198 -4842 360434
rect -4606 360198 -4522 360434
rect -4286 360198 -4202 360434
rect -3966 360198 -3882 360434
rect -3646 360198 -3538 360434
rect -4950 353434 -3538 360198
rect -4950 353198 -4842 353434
rect -4606 353198 -4522 353434
rect -4286 353198 -4202 353434
rect -3966 353198 -3882 353434
rect -3646 353198 -3538 353434
rect -4950 346434 -3538 353198
rect -4950 346198 -4842 346434
rect -4606 346198 -4522 346434
rect -4286 346198 -4202 346434
rect -3966 346198 -3882 346434
rect -3646 346198 -3538 346434
rect -4950 339434 -3538 346198
rect -4950 339198 -4842 339434
rect -4606 339198 -4522 339434
rect -4286 339198 -4202 339434
rect -3966 339198 -3882 339434
rect -3646 339198 -3538 339434
rect -4950 332434 -3538 339198
rect -4950 332198 -4842 332434
rect -4606 332198 -4522 332434
rect -4286 332198 -4202 332434
rect -3966 332198 -3882 332434
rect -3646 332198 -3538 332434
rect -4950 325434 -3538 332198
rect -4950 325198 -4842 325434
rect -4606 325198 -4522 325434
rect -4286 325198 -4202 325434
rect -3966 325198 -3882 325434
rect -3646 325198 -3538 325434
rect -4950 318434 -3538 325198
rect -4950 318198 -4842 318434
rect -4606 318198 -4522 318434
rect -4286 318198 -4202 318434
rect -3966 318198 -3882 318434
rect -3646 318198 -3538 318434
rect -4950 311434 -3538 318198
rect -4950 311198 -4842 311434
rect -4606 311198 -4522 311434
rect -4286 311198 -4202 311434
rect -3966 311198 -3882 311434
rect -3646 311198 -3538 311434
rect -4950 304434 -3538 311198
rect -4950 304198 -4842 304434
rect -4606 304198 -4522 304434
rect -4286 304198 -4202 304434
rect -3966 304198 -3882 304434
rect -3646 304198 -3538 304434
rect -4950 297434 -3538 304198
rect -4950 297198 -4842 297434
rect -4606 297198 -4522 297434
rect -4286 297198 -4202 297434
rect -3966 297198 -3882 297434
rect -3646 297198 -3538 297434
rect -4950 290434 -3538 297198
rect -4950 290198 -4842 290434
rect -4606 290198 -4522 290434
rect -4286 290198 -4202 290434
rect -3966 290198 -3882 290434
rect -3646 290198 -3538 290434
rect -4950 283434 -3538 290198
rect -4950 283198 -4842 283434
rect -4606 283198 -4522 283434
rect -4286 283198 -4202 283434
rect -3966 283198 -3882 283434
rect -3646 283198 -3538 283434
rect -4950 276434 -3538 283198
rect -4950 276198 -4842 276434
rect -4606 276198 -4522 276434
rect -4286 276198 -4202 276434
rect -3966 276198 -3882 276434
rect -3646 276198 -3538 276434
rect -4950 269434 -3538 276198
rect -4950 269198 -4842 269434
rect -4606 269198 -4522 269434
rect -4286 269198 -4202 269434
rect -3966 269198 -3882 269434
rect -3646 269198 -3538 269434
rect -4950 262434 -3538 269198
rect -4950 262198 -4842 262434
rect -4606 262198 -4522 262434
rect -4286 262198 -4202 262434
rect -3966 262198 -3882 262434
rect -3646 262198 -3538 262434
rect -4950 255434 -3538 262198
rect -4950 255198 -4842 255434
rect -4606 255198 -4522 255434
rect -4286 255198 -4202 255434
rect -3966 255198 -3882 255434
rect -3646 255198 -3538 255434
rect -4950 248434 -3538 255198
rect -4950 248198 -4842 248434
rect -4606 248198 -4522 248434
rect -4286 248198 -4202 248434
rect -3966 248198 -3882 248434
rect -3646 248198 -3538 248434
rect -4950 241434 -3538 248198
rect -4950 241198 -4842 241434
rect -4606 241198 -4522 241434
rect -4286 241198 -4202 241434
rect -3966 241198 -3882 241434
rect -3646 241198 -3538 241434
rect -4950 234434 -3538 241198
rect -4950 234198 -4842 234434
rect -4606 234198 -4522 234434
rect -4286 234198 -4202 234434
rect -3966 234198 -3882 234434
rect -3646 234198 -3538 234434
rect -4950 227434 -3538 234198
rect -4950 227198 -4842 227434
rect -4606 227198 -4522 227434
rect -4286 227198 -4202 227434
rect -3966 227198 -3882 227434
rect -3646 227198 -3538 227434
rect -4950 220434 -3538 227198
rect -4950 220198 -4842 220434
rect -4606 220198 -4522 220434
rect -4286 220198 -4202 220434
rect -3966 220198 -3882 220434
rect -3646 220198 -3538 220434
rect -4950 213434 -3538 220198
rect -4950 213198 -4842 213434
rect -4606 213198 -4522 213434
rect -4286 213198 -4202 213434
rect -3966 213198 -3882 213434
rect -3646 213198 -3538 213434
rect -4950 206434 -3538 213198
rect -4950 206198 -4842 206434
rect -4606 206198 -4522 206434
rect -4286 206198 -4202 206434
rect -3966 206198 -3882 206434
rect -3646 206198 -3538 206434
rect -4950 199434 -3538 206198
rect -4950 199198 -4842 199434
rect -4606 199198 -4522 199434
rect -4286 199198 -4202 199434
rect -3966 199198 -3882 199434
rect -3646 199198 -3538 199434
rect -4950 192434 -3538 199198
rect -4950 192198 -4842 192434
rect -4606 192198 -4522 192434
rect -4286 192198 -4202 192434
rect -3966 192198 -3882 192434
rect -3646 192198 -3538 192434
rect -4950 185434 -3538 192198
rect -4950 185198 -4842 185434
rect -4606 185198 -4522 185434
rect -4286 185198 -4202 185434
rect -3966 185198 -3882 185434
rect -3646 185198 -3538 185434
rect -4950 178434 -3538 185198
rect -4950 178198 -4842 178434
rect -4606 178198 -4522 178434
rect -4286 178198 -4202 178434
rect -3966 178198 -3882 178434
rect -3646 178198 -3538 178434
rect -4950 171434 -3538 178198
rect -4950 171198 -4842 171434
rect -4606 171198 -4522 171434
rect -4286 171198 -4202 171434
rect -3966 171198 -3882 171434
rect -3646 171198 -3538 171434
rect -4950 164434 -3538 171198
rect -4950 164198 -4842 164434
rect -4606 164198 -4522 164434
rect -4286 164198 -4202 164434
rect -3966 164198 -3882 164434
rect -3646 164198 -3538 164434
rect -4950 157434 -3538 164198
rect -4950 157198 -4842 157434
rect -4606 157198 -4522 157434
rect -4286 157198 -4202 157434
rect -3966 157198 -3882 157434
rect -3646 157198 -3538 157434
rect -4950 150434 -3538 157198
rect -4950 150198 -4842 150434
rect -4606 150198 -4522 150434
rect -4286 150198 -4202 150434
rect -3966 150198 -3882 150434
rect -3646 150198 -3538 150434
rect -4950 143434 -3538 150198
rect -4950 143198 -4842 143434
rect -4606 143198 -4522 143434
rect -4286 143198 -4202 143434
rect -3966 143198 -3882 143434
rect -3646 143198 -3538 143434
rect -4950 136434 -3538 143198
rect -4950 136198 -4842 136434
rect -4606 136198 -4522 136434
rect -4286 136198 -4202 136434
rect -3966 136198 -3882 136434
rect -3646 136198 -3538 136434
rect -4950 129434 -3538 136198
rect -4950 129198 -4842 129434
rect -4606 129198 -4522 129434
rect -4286 129198 -4202 129434
rect -3966 129198 -3882 129434
rect -3646 129198 -3538 129434
rect -4950 122434 -3538 129198
rect -4950 122198 -4842 122434
rect -4606 122198 -4522 122434
rect -4286 122198 -4202 122434
rect -3966 122198 -3882 122434
rect -3646 122198 -3538 122434
rect -4950 115434 -3538 122198
rect -4950 115198 -4842 115434
rect -4606 115198 -4522 115434
rect -4286 115198 -4202 115434
rect -3966 115198 -3882 115434
rect -3646 115198 -3538 115434
rect -4950 108434 -3538 115198
rect -4950 108198 -4842 108434
rect -4606 108198 -4522 108434
rect -4286 108198 -4202 108434
rect -3966 108198 -3882 108434
rect -3646 108198 -3538 108434
rect -4950 101434 -3538 108198
rect -4950 101198 -4842 101434
rect -4606 101198 -4522 101434
rect -4286 101198 -4202 101434
rect -3966 101198 -3882 101434
rect -3646 101198 -3538 101434
rect -4950 94434 -3538 101198
rect -4950 94198 -4842 94434
rect -4606 94198 -4522 94434
rect -4286 94198 -4202 94434
rect -3966 94198 -3882 94434
rect -3646 94198 -3538 94434
rect -4950 87434 -3538 94198
rect -4950 87198 -4842 87434
rect -4606 87198 -4522 87434
rect -4286 87198 -4202 87434
rect -3966 87198 -3882 87434
rect -3646 87198 -3538 87434
rect -4950 80434 -3538 87198
rect -4950 80198 -4842 80434
rect -4606 80198 -4522 80434
rect -4286 80198 -4202 80434
rect -3966 80198 -3882 80434
rect -3646 80198 -3538 80434
rect -4950 73434 -3538 80198
rect -4950 73198 -4842 73434
rect -4606 73198 -4522 73434
rect -4286 73198 -4202 73434
rect -3966 73198 -3882 73434
rect -3646 73198 -3538 73434
rect -4950 66434 -3538 73198
rect -4950 66198 -4842 66434
rect -4606 66198 -4522 66434
rect -4286 66198 -4202 66434
rect -3966 66198 -3882 66434
rect -3646 66198 -3538 66434
rect -4950 59434 -3538 66198
rect -4950 59198 -4842 59434
rect -4606 59198 -4522 59434
rect -4286 59198 -4202 59434
rect -3966 59198 -3882 59434
rect -3646 59198 -3538 59434
rect -4950 52434 -3538 59198
rect -4950 52198 -4842 52434
rect -4606 52198 -4522 52434
rect -4286 52198 -4202 52434
rect -3966 52198 -3882 52434
rect -3646 52198 -3538 52434
rect -4950 45434 -3538 52198
rect -4950 45198 -4842 45434
rect -4606 45198 -4522 45434
rect -4286 45198 -4202 45434
rect -3966 45198 -3882 45434
rect -3646 45198 -3538 45434
rect -4950 38434 -3538 45198
rect -4950 38198 -4842 38434
rect -4606 38198 -4522 38434
rect -4286 38198 -4202 38434
rect -3966 38198 -3882 38434
rect -3646 38198 -3538 38434
rect -4950 31434 -3538 38198
rect -4950 31198 -4842 31434
rect -4606 31198 -4522 31434
rect -4286 31198 -4202 31434
rect -3966 31198 -3882 31434
rect -3646 31198 -3538 31434
rect -4950 24434 -3538 31198
rect -4950 24198 -4842 24434
rect -4606 24198 -4522 24434
rect -4286 24198 -4202 24434
rect -3966 24198 -3882 24434
rect -3646 24198 -3538 24434
rect -4950 17434 -3538 24198
rect -4950 17198 -4842 17434
rect -4606 17198 -4522 17434
rect -4286 17198 -4202 17434
rect -3966 17198 -3882 17434
rect -3646 17198 -3538 17434
rect -4950 10434 -3538 17198
rect -4950 10198 -4842 10434
rect -4606 10198 -4522 10434
rect -4286 10198 -4202 10434
rect -3966 10198 -3882 10434
rect -3646 10198 -3538 10434
rect -4950 3434 -3538 10198
rect -4950 3198 -4842 3434
rect -4606 3198 -4522 3434
rect -4286 3198 -4202 3434
rect -3966 3198 -3882 3434
rect -3646 3198 -3538 3434
rect -4950 -3878 -3538 3198
rect -3198 705238 -1786 706062
rect -3198 705002 -2374 705238
rect -2138 705002 -2054 705238
rect -1818 705002 -1786 705238
rect -3198 704918 -1786 705002
rect -3198 704682 -2374 704918
rect -2138 704682 -2054 704918
rect -1818 704682 -1786 704918
rect -3198 695494 -1786 704682
rect -3198 695258 -3090 695494
rect -2854 695258 -2770 695494
rect -2534 695258 -2450 695494
rect -2214 695258 -2130 695494
rect -1894 695258 -1786 695494
rect -3198 688494 -1786 695258
rect -3198 688258 -3090 688494
rect -2854 688258 -2770 688494
rect -2534 688258 -2450 688494
rect -2214 688258 -2130 688494
rect -1894 688258 -1786 688494
rect -3198 681494 -1786 688258
rect -3198 681258 -3090 681494
rect -2854 681258 -2770 681494
rect -2534 681258 -2450 681494
rect -2214 681258 -2130 681494
rect -1894 681258 -1786 681494
rect -3198 674494 -1786 681258
rect -3198 674258 -3090 674494
rect -2854 674258 -2770 674494
rect -2534 674258 -2450 674494
rect -2214 674258 -2130 674494
rect -1894 674258 -1786 674494
rect -3198 667494 -1786 674258
rect -3198 667258 -3090 667494
rect -2854 667258 -2770 667494
rect -2534 667258 -2450 667494
rect -2214 667258 -2130 667494
rect -1894 667258 -1786 667494
rect -3198 660494 -1786 667258
rect -3198 660258 -3090 660494
rect -2854 660258 -2770 660494
rect -2534 660258 -2450 660494
rect -2214 660258 -2130 660494
rect -1894 660258 -1786 660494
rect -3198 653494 -1786 660258
rect -3198 653258 -3090 653494
rect -2854 653258 -2770 653494
rect -2534 653258 -2450 653494
rect -2214 653258 -2130 653494
rect -1894 653258 -1786 653494
rect -3198 646494 -1786 653258
rect -3198 646258 -3090 646494
rect -2854 646258 -2770 646494
rect -2534 646258 -2450 646494
rect -2214 646258 -2130 646494
rect -1894 646258 -1786 646494
rect -3198 639494 -1786 646258
rect -3198 639258 -3090 639494
rect -2854 639258 -2770 639494
rect -2534 639258 -2450 639494
rect -2214 639258 -2130 639494
rect -1894 639258 -1786 639494
rect -3198 632494 -1786 639258
rect -3198 632258 -3090 632494
rect -2854 632258 -2770 632494
rect -2534 632258 -2450 632494
rect -2214 632258 -2130 632494
rect -1894 632258 -1786 632494
rect -3198 625494 -1786 632258
rect -3198 625258 -3090 625494
rect -2854 625258 -2770 625494
rect -2534 625258 -2450 625494
rect -2214 625258 -2130 625494
rect -1894 625258 -1786 625494
rect -3198 618494 -1786 625258
rect -3198 618258 -3090 618494
rect -2854 618258 -2770 618494
rect -2534 618258 -2450 618494
rect -2214 618258 -2130 618494
rect -1894 618258 -1786 618494
rect -3198 611494 -1786 618258
rect -3198 611258 -3090 611494
rect -2854 611258 -2770 611494
rect -2534 611258 -2450 611494
rect -2214 611258 -2130 611494
rect -1894 611258 -1786 611494
rect -3198 604494 -1786 611258
rect -3198 604258 -3090 604494
rect -2854 604258 -2770 604494
rect -2534 604258 -2450 604494
rect -2214 604258 -2130 604494
rect -1894 604258 -1786 604494
rect -3198 597494 -1786 604258
rect -3198 597258 -3090 597494
rect -2854 597258 -2770 597494
rect -2534 597258 -2450 597494
rect -2214 597258 -2130 597494
rect -1894 597258 -1786 597494
rect -3198 590494 -1786 597258
rect -3198 590258 -3090 590494
rect -2854 590258 -2770 590494
rect -2534 590258 -2450 590494
rect -2214 590258 -2130 590494
rect -1894 590258 -1786 590494
rect -3198 583494 -1786 590258
rect -3198 583258 -3090 583494
rect -2854 583258 -2770 583494
rect -2534 583258 -2450 583494
rect -2214 583258 -2130 583494
rect -1894 583258 -1786 583494
rect -3198 576494 -1786 583258
rect -3198 576258 -3090 576494
rect -2854 576258 -2770 576494
rect -2534 576258 -2450 576494
rect -2214 576258 -2130 576494
rect -1894 576258 -1786 576494
rect -3198 569494 -1786 576258
rect -3198 569258 -3090 569494
rect -2854 569258 -2770 569494
rect -2534 569258 -2450 569494
rect -2214 569258 -2130 569494
rect -1894 569258 -1786 569494
rect -3198 562494 -1786 569258
rect -3198 562258 -3090 562494
rect -2854 562258 -2770 562494
rect -2534 562258 -2450 562494
rect -2214 562258 -2130 562494
rect -1894 562258 -1786 562494
rect -3198 555494 -1786 562258
rect -3198 555258 -3090 555494
rect -2854 555258 -2770 555494
rect -2534 555258 -2450 555494
rect -2214 555258 -2130 555494
rect -1894 555258 -1786 555494
rect -3198 548494 -1786 555258
rect -3198 548258 -3090 548494
rect -2854 548258 -2770 548494
rect -2534 548258 -2450 548494
rect -2214 548258 -2130 548494
rect -1894 548258 -1786 548494
rect -3198 541494 -1786 548258
rect -3198 541258 -3090 541494
rect -2854 541258 -2770 541494
rect -2534 541258 -2450 541494
rect -2214 541258 -2130 541494
rect -1894 541258 -1786 541494
rect -3198 534494 -1786 541258
rect -3198 534258 -3090 534494
rect -2854 534258 -2770 534494
rect -2534 534258 -2450 534494
rect -2214 534258 -2130 534494
rect -1894 534258 -1786 534494
rect -3198 527494 -1786 534258
rect -3198 527258 -3090 527494
rect -2854 527258 -2770 527494
rect -2534 527258 -2450 527494
rect -2214 527258 -2130 527494
rect -1894 527258 -1786 527494
rect -3198 520494 -1786 527258
rect -3198 520258 -3090 520494
rect -2854 520258 -2770 520494
rect -2534 520258 -2450 520494
rect -2214 520258 -2130 520494
rect -1894 520258 -1786 520494
rect -3198 513494 -1786 520258
rect -3198 513258 -3090 513494
rect -2854 513258 -2770 513494
rect -2534 513258 -2450 513494
rect -2214 513258 -2130 513494
rect -1894 513258 -1786 513494
rect -3198 506494 -1786 513258
rect -3198 506258 -3090 506494
rect -2854 506258 -2770 506494
rect -2534 506258 -2450 506494
rect -2214 506258 -2130 506494
rect -1894 506258 -1786 506494
rect -3198 499494 -1786 506258
rect -3198 499258 -3090 499494
rect -2854 499258 -2770 499494
rect -2534 499258 -2450 499494
rect -2214 499258 -2130 499494
rect -1894 499258 -1786 499494
rect -3198 492494 -1786 499258
rect -3198 492258 -3090 492494
rect -2854 492258 -2770 492494
rect -2534 492258 -2450 492494
rect -2214 492258 -2130 492494
rect -1894 492258 -1786 492494
rect -3198 485494 -1786 492258
rect -3198 485258 -3090 485494
rect -2854 485258 -2770 485494
rect -2534 485258 -2450 485494
rect -2214 485258 -2130 485494
rect -1894 485258 -1786 485494
rect -3198 478494 -1786 485258
rect -3198 478258 -3090 478494
rect -2854 478258 -2770 478494
rect -2534 478258 -2450 478494
rect -2214 478258 -2130 478494
rect -1894 478258 -1786 478494
rect -3198 471494 -1786 478258
rect -3198 471258 -3090 471494
rect -2854 471258 -2770 471494
rect -2534 471258 -2450 471494
rect -2214 471258 -2130 471494
rect -1894 471258 -1786 471494
rect -3198 464494 -1786 471258
rect -3198 464258 -3090 464494
rect -2854 464258 -2770 464494
rect -2534 464258 -2450 464494
rect -2214 464258 -2130 464494
rect -1894 464258 -1786 464494
rect -3198 457494 -1786 464258
rect -3198 457258 -3090 457494
rect -2854 457258 -2770 457494
rect -2534 457258 -2450 457494
rect -2214 457258 -2130 457494
rect -1894 457258 -1786 457494
rect -3198 450494 -1786 457258
rect -3198 450258 -3090 450494
rect -2854 450258 -2770 450494
rect -2534 450258 -2450 450494
rect -2214 450258 -2130 450494
rect -1894 450258 -1786 450494
rect -3198 443494 -1786 450258
rect -3198 443258 -3090 443494
rect -2854 443258 -2770 443494
rect -2534 443258 -2450 443494
rect -2214 443258 -2130 443494
rect -1894 443258 -1786 443494
rect -3198 436494 -1786 443258
rect -3198 436258 -3090 436494
rect -2854 436258 -2770 436494
rect -2534 436258 -2450 436494
rect -2214 436258 -2130 436494
rect -1894 436258 -1786 436494
rect -3198 429494 -1786 436258
rect -3198 429258 -3090 429494
rect -2854 429258 -2770 429494
rect -2534 429258 -2450 429494
rect -2214 429258 -2130 429494
rect -1894 429258 -1786 429494
rect -3198 422494 -1786 429258
rect -3198 422258 -3090 422494
rect -2854 422258 -2770 422494
rect -2534 422258 -2450 422494
rect -2214 422258 -2130 422494
rect -1894 422258 -1786 422494
rect -3198 415494 -1786 422258
rect -3198 415258 -3090 415494
rect -2854 415258 -2770 415494
rect -2534 415258 -2450 415494
rect -2214 415258 -2130 415494
rect -1894 415258 -1786 415494
rect -3198 408494 -1786 415258
rect -3198 408258 -3090 408494
rect -2854 408258 -2770 408494
rect -2534 408258 -2450 408494
rect -2214 408258 -2130 408494
rect -1894 408258 -1786 408494
rect -3198 401494 -1786 408258
rect -3198 401258 -3090 401494
rect -2854 401258 -2770 401494
rect -2534 401258 -2450 401494
rect -2214 401258 -2130 401494
rect -1894 401258 -1786 401494
rect -3198 394494 -1786 401258
rect -3198 394258 -3090 394494
rect -2854 394258 -2770 394494
rect -2534 394258 -2450 394494
rect -2214 394258 -2130 394494
rect -1894 394258 -1786 394494
rect -3198 387494 -1786 394258
rect -3198 387258 -3090 387494
rect -2854 387258 -2770 387494
rect -2534 387258 -2450 387494
rect -2214 387258 -2130 387494
rect -1894 387258 -1786 387494
rect -3198 380494 -1786 387258
rect -3198 380258 -3090 380494
rect -2854 380258 -2770 380494
rect -2534 380258 -2450 380494
rect -2214 380258 -2130 380494
rect -1894 380258 -1786 380494
rect -3198 373494 -1786 380258
rect -3198 373258 -3090 373494
rect -2854 373258 -2770 373494
rect -2534 373258 -2450 373494
rect -2214 373258 -2130 373494
rect -1894 373258 -1786 373494
rect -3198 366494 -1786 373258
rect -3198 366258 -3090 366494
rect -2854 366258 -2770 366494
rect -2534 366258 -2450 366494
rect -2214 366258 -2130 366494
rect -1894 366258 -1786 366494
rect -3198 359494 -1786 366258
rect -3198 359258 -3090 359494
rect -2854 359258 -2770 359494
rect -2534 359258 -2450 359494
rect -2214 359258 -2130 359494
rect -1894 359258 -1786 359494
rect -3198 352494 -1786 359258
rect -3198 352258 -3090 352494
rect -2854 352258 -2770 352494
rect -2534 352258 -2450 352494
rect -2214 352258 -2130 352494
rect -1894 352258 -1786 352494
rect -3198 345494 -1786 352258
rect -3198 345258 -3090 345494
rect -2854 345258 -2770 345494
rect -2534 345258 -2450 345494
rect -2214 345258 -2130 345494
rect -1894 345258 -1786 345494
rect -3198 338494 -1786 345258
rect -3198 338258 -3090 338494
rect -2854 338258 -2770 338494
rect -2534 338258 -2450 338494
rect -2214 338258 -2130 338494
rect -1894 338258 -1786 338494
rect -3198 331494 -1786 338258
rect -3198 331258 -3090 331494
rect -2854 331258 -2770 331494
rect -2534 331258 -2450 331494
rect -2214 331258 -2130 331494
rect -1894 331258 -1786 331494
rect -3198 324494 -1786 331258
rect -3198 324258 -3090 324494
rect -2854 324258 -2770 324494
rect -2534 324258 -2450 324494
rect -2214 324258 -2130 324494
rect -1894 324258 -1786 324494
rect -3198 317494 -1786 324258
rect -3198 317258 -3090 317494
rect -2854 317258 -2770 317494
rect -2534 317258 -2450 317494
rect -2214 317258 -2130 317494
rect -1894 317258 -1786 317494
rect -3198 310494 -1786 317258
rect -3198 310258 -3090 310494
rect -2854 310258 -2770 310494
rect -2534 310258 -2450 310494
rect -2214 310258 -2130 310494
rect -1894 310258 -1786 310494
rect -3198 303494 -1786 310258
rect -3198 303258 -3090 303494
rect -2854 303258 -2770 303494
rect -2534 303258 -2450 303494
rect -2214 303258 -2130 303494
rect -1894 303258 -1786 303494
rect -3198 296494 -1786 303258
rect -3198 296258 -3090 296494
rect -2854 296258 -2770 296494
rect -2534 296258 -2450 296494
rect -2214 296258 -2130 296494
rect -1894 296258 -1786 296494
rect -3198 289494 -1786 296258
rect -3198 289258 -3090 289494
rect -2854 289258 -2770 289494
rect -2534 289258 -2450 289494
rect -2214 289258 -2130 289494
rect -1894 289258 -1786 289494
rect -3198 282494 -1786 289258
rect -3198 282258 -3090 282494
rect -2854 282258 -2770 282494
rect -2534 282258 -2450 282494
rect -2214 282258 -2130 282494
rect -1894 282258 -1786 282494
rect -3198 275494 -1786 282258
rect -3198 275258 -3090 275494
rect -2854 275258 -2770 275494
rect -2534 275258 -2450 275494
rect -2214 275258 -2130 275494
rect -1894 275258 -1786 275494
rect -3198 268494 -1786 275258
rect -3198 268258 -3090 268494
rect -2854 268258 -2770 268494
rect -2534 268258 -2450 268494
rect -2214 268258 -2130 268494
rect -1894 268258 -1786 268494
rect -3198 261494 -1786 268258
rect -3198 261258 -3090 261494
rect -2854 261258 -2770 261494
rect -2534 261258 -2450 261494
rect -2214 261258 -2130 261494
rect -1894 261258 -1786 261494
rect -3198 254494 -1786 261258
rect -3198 254258 -3090 254494
rect -2854 254258 -2770 254494
rect -2534 254258 -2450 254494
rect -2214 254258 -2130 254494
rect -1894 254258 -1786 254494
rect -3198 247494 -1786 254258
rect -3198 247258 -3090 247494
rect -2854 247258 -2770 247494
rect -2534 247258 -2450 247494
rect -2214 247258 -2130 247494
rect -1894 247258 -1786 247494
rect -3198 240494 -1786 247258
rect -3198 240258 -3090 240494
rect -2854 240258 -2770 240494
rect -2534 240258 -2450 240494
rect -2214 240258 -2130 240494
rect -1894 240258 -1786 240494
rect -3198 233494 -1786 240258
rect -3198 233258 -3090 233494
rect -2854 233258 -2770 233494
rect -2534 233258 -2450 233494
rect -2214 233258 -2130 233494
rect -1894 233258 -1786 233494
rect -3198 226494 -1786 233258
rect -3198 226258 -3090 226494
rect -2854 226258 -2770 226494
rect -2534 226258 -2450 226494
rect -2214 226258 -2130 226494
rect -1894 226258 -1786 226494
rect -3198 219494 -1786 226258
rect -3198 219258 -3090 219494
rect -2854 219258 -2770 219494
rect -2534 219258 -2450 219494
rect -2214 219258 -2130 219494
rect -1894 219258 -1786 219494
rect -3198 212494 -1786 219258
rect -3198 212258 -3090 212494
rect -2854 212258 -2770 212494
rect -2534 212258 -2450 212494
rect -2214 212258 -2130 212494
rect -1894 212258 -1786 212494
rect -3198 205494 -1786 212258
rect -3198 205258 -3090 205494
rect -2854 205258 -2770 205494
rect -2534 205258 -2450 205494
rect -2214 205258 -2130 205494
rect -1894 205258 -1786 205494
rect -3198 198494 -1786 205258
rect -3198 198258 -3090 198494
rect -2854 198258 -2770 198494
rect -2534 198258 -2450 198494
rect -2214 198258 -2130 198494
rect -1894 198258 -1786 198494
rect -3198 191494 -1786 198258
rect -3198 191258 -3090 191494
rect -2854 191258 -2770 191494
rect -2534 191258 -2450 191494
rect -2214 191258 -2130 191494
rect -1894 191258 -1786 191494
rect -3198 184494 -1786 191258
rect -3198 184258 -3090 184494
rect -2854 184258 -2770 184494
rect -2534 184258 -2450 184494
rect -2214 184258 -2130 184494
rect -1894 184258 -1786 184494
rect -3198 177494 -1786 184258
rect -3198 177258 -3090 177494
rect -2854 177258 -2770 177494
rect -2534 177258 -2450 177494
rect -2214 177258 -2130 177494
rect -1894 177258 -1786 177494
rect -3198 170494 -1786 177258
rect -3198 170258 -3090 170494
rect -2854 170258 -2770 170494
rect -2534 170258 -2450 170494
rect -2214 170258 -2130 170494
rect -1894 170258 -1786 170494
rect -3198 163494 -1786 170258
rect -3198 163258 -3090 163494
rect -2854 163258 -2770 163494
rect -2534 163258 -2450 163494
rect -2214 163258 -2130 163494
rect -1894 163258 -1786 163494
rect -3198 156494 -1786 163258
rect -3198 156258 -3090 156494
rect -2854 156258 -2770 156494
rect -2534 156258 -2450 156494
rect -2214 156258 -2130 156494
rect -1894 156258 -1786 156494
rect -3198 149494 -1786 156258
rect -3198 149258 -3090 149494
rect -2854 149258 -2770 149494
rect -2534 149258 -2450 149494
rect -2214 149258 -2130 149494
rect -1894 149258 -1786 149494
rect -3198 142494 -1786 149258
rect -3198 142258 -3090 142494
rect -2854 142258 -2770 142494
rect -2534 142258 -2450 142494
rect -2214 142258 -2130 142494
rect -1894 142258 -1786 142494
rect -3198 135494 -1786 142258
rect -3198 135258 -3090 135494
rect -2854 135258 -2770 135494
rect -2534 135258 -2450 135494
rect -2214 135258 -2130 135494
rect -1894 135258 -1786 135494
rect -3198 128494 -1786 135258
rect -3198 128258 -3090 128494
rect -2854 128258 -2770 128494
rect -2534 128258 -2450 128494
rect -2214 128258 -2130 128494
rect -1894 128258 -1786 128494
rect -3198 121494 -1786 128258
rect -3198 121258 -3090 121494
rect -2854 121258 -2770 121494
rect -2534 121258 -2450 121494
rect -2214 121258 -2130 121494
rect -1894 121258 -1786 121494
rect -3198 114494 -1786 121258
rect -3198 114258 -3090 114494
rect -2854 114258 -2770 114494
rect -2534 114258 -2450 114494
rect -2214 114258 -2130 114494
rect -1894 114258 -1786 114494
rect -3198 107494 -1786 114258
rect -3198 107258 -3090 107494
rect -2854 107258 -2770 107494
rect -2534 107258 -2450 107494
rect -2214 107258 -2130 107494
rect -1894 107258 -1786 107494
rect -3198 100494 -1786 107258
rect -3198 100258 -3090 100494
rect -2854 100258 -2770 100494
rect -2534 100258 -2450 100494
rect -2214 100258 -2130 100494
rect -1894 100258 -1786 100494
rect -3198 93494 -1786 100258
rect -3198 93258 -3090 93494
rect -2854 93258 -2770 93494
rect -2534 93258 -2450 93494
rect -2214 93258 -2130 93494
rect -1894 93258 -1786 93494
rect -3198 86494 -1786 93258
rect -3198 86258 -3090 86494
rect -2854 86258 -2770 86494
rect -2534 86258 -2450 86494
rect -2214 86258 -2130 86494
rect -1894 86258 -1786 86494
rect -3198 79494 -1786 86258
rect -3198 79258 -3090 79494
rect -2854 79258 -2770 79494
rect -2534 79258 -2450 79494
rect -2214 79258 -2130 79494
rect -1894 79258 -1786 79494
rect -3198 72494 -1786 79258
rect -3198 72258 -3090 72494
rect -2854 72258 -2770 72494
rect -2534 72258 -2450 72494
rect -2214 72258 -2130 72494
rect -1894 72258 -1786 72494
rect -3198 65494 -1786 72258
rect -3198 65258 -3090 65494
rect -2854 65258 -2770 65494
rect -2534 65258 -2450 65494
rect -2214 65258 -2130 65494
rect -1894 65258 -1786 65494
rect -3198 58494 -1786 65258
rect -3198 58258 -3090 58494
rect -2854 58258 -2770 58494
rect -2534 58258 -2450 58494
rect -2214 58258 -2130 58494
rect -1894 58258 -1786 58494
rect -3198 51494 -1786 58258
rect -3198 51258 -3090 51494
rect -2854 51258 -2770 51494
rect -2534 51258 -2450 51494
rect -2214 51258 -2130 51494
rect -1894 51258 -1786 51494
rect -3198 44494 -1786 51258
rect -3198 44258 -3090 44494
rect -2854 44258 -2770 44494
rect -2534 44258 -2450 44494
rect -2214 44258 -2130 44494
rect -1894 44258 -1786 44494
rect -3198 37494 -1786 44258
rect -3198 37258 -3090 37494
rect -2854 37258 -2770 37494
rect -2534 37258 -2450 37494
rect -2214 37258 -2130 37494
rect -1894 37258 -1786 37494
rect -3198 30494 -1786 37258
rect -3198 30258 -3090 30494
rect -2854 30258 -2770 30494
rect -2534 30258 -2450 30494
rect -2214 30258 -2130 30494
rect -1894 30258 -1786 30494
rect -3198 23494 -1786 30258
rect -3198 23258 -3090 23494
rect -2854 23258 -2770 23494
rect -2534 23258 -2450 23494
rect -2214 23258 -2130 23494
rect -1894 23258 -1786 23494
rect -3198 16494 -1786 23258
rect -3198 16258 -3090 16494
rect -2854 16258 -2770 16494
rect -2534 16258 -2450 16494
rect -2214 16258 -2130 16494
rect -1894 16258 -1786 16494
rect -3198 9494 -1786 16258
rect -3198 9258 -3090 9494
rect -2854 9258 -2770 9494
rect -2534 9258 -2450 9494
rect -2214 9258 -2130 9494
rect -1894 9258 -1786 9494
rect -3198 2494 -1786 9258
rect -3198 2258 -3090 2494
rect -2854 2258 -2770 2494
rect -2534 2258 -2450 2494
rect -2214 2258 -2130 2494
rect -1894 2258 -1786 2494
rect -3198 -746 -1786 2258
rect -3198 -982 -2374 -746
rect -2138 -982 -2054 -746
rect -1818 -982 -1786 -746
rect -3198 -1066 -1786 -982
rect -3198 -1302 -2374 -1066
rect -2138 -1302 -2054 -1066
rect -1818 -1302 -1786 -1066
rect -3198 -2126 -1786 -1302
rect 1144 705238 1464 706230
rect 1144 705002 1186 705238
rect 1422 705002 1464 705238
rect 1144 704918 1464 705002
rect 1144 704682 1186 704918
rect 1422 704682 1464 704918
rect 1144 695494 1464 704682
rect 1144 695258 1186 695494
rect 1422 695258 1464 695494
rect 1144 688494 1464 695258
rect 1144 688258 1186 688494
rect 1422 688258 1464 688494
rect 1144 681494 1464 688258
rect 1144 681258 1186 681494
rect 1422 681258 1464 681494
rect 1144 674494 1464 681258
rect 1144 674258 1186 674494
rect 1422 674258 1464 674494
rect 1144 667494 1464 674258
rect 1144 667258 1186 667494
rect 1422 667258 1464 667494
rect 1144 660494 1464 667258
rect 1144 660258 1186 660494
rect 1422 660258 1464 660494
rect 1144 653494 1464 660258
rect 1144 653258 1186 653494
rect 1422 653258 1464 653494
rect 1144 646494 1464 653258
rect 1144 646258 1186 646494
rect 1422 646258 1464 646494
rect 1144 639494 1464 646258
rect 1144 639258 1186 639494
rect 1422 639258 1464 639494
rect 1144 632494 1464 639258
rect 1144 632258 1186 632494
rect 1422 632258 1464 632494
rect 1144 625494 1464 632258
rect 1144 625258 1186 625494
rect 1422 625258 1464 625494
rect 1144 618494 1464 625258
rect 1144 618258 1186 618494
rect 1422 618258 1464 618494
rect 1144 611494 1464 618258
rect 1144 611258 1186 611494
rect 1422 611258 1464 611494
rect 1144 604494 1464 611258
rect 1144 604258 1186 604494
rect 1422 604258 1464 604494
rect 1144 597494 1464 604258
rect 1144 597258 1186 597494
rect 1422 597258 1464 597494
rect 1144 590494 1464 597258
rect 1144 590258 1186 590494
rect 1422 590258 1464 590494
rect 1144 583494 1464 590258
rect 1144 583258 1186 583494
rect 1422 583258 1464 583494
rect 1144 576494 1464 583258
rect 1144 576258 1186 576494
rect 1422 576258 1464 576494
rect 1144 569494 1464 576258
rect 1144 569258 1186 569494
rect 1422 569258 1464 569494
rect 1144 562494 1464 569258
rect 1144 562258 1186 562494
rect 1422 562258 1464 562494
rect 1144 555494 1464 562258
rect 1144 555258 1186 555494
rect 1422 555258 1464 555494
rect 1144 548494 1464 555258
rect 1144 548258 1186 548494
rect 1422 548258 1464 548494
rect 1144 541494 1464 548258
rect 1144 541258 1186 541494
rect 1422 541258 1464 541494
rect 1144 534494 1464 541258
rect 1144 534258 1186 534494
rect 1422 534258 1464 534494
rect 1144 527494 1464 534258
rect 1144 527258 1186 527494
rect 1422 527258 1464 527494
rect 1144 520494 1464 527258
rect 1144 520258 1186 520494
rect 1422 520258 1464 520494
rect 1144 513494 1464 520258
rect 1144 513258 1186 513494
rect 1422 513258 1464 513494
rect 1144 506494 1464 513258
rect 1144 506258 1186 506494
rect 1422 506258 1464 506494
rect 1144 499494 1464 506258
rect 1144 499258 1186 499494
rect 1422 499258 1464 499494
rect 1144 492494 1464 499258
rect 1144 492258 1186 492494
rect 1422 492258 1464 492494
rect 1144 485494 1464 492258
rect 1144 485258 1186 485494
rect 1422 485258 1464 485494
rect 1144 478494 1464 485258
rect 1144 478258 1186 478494
rect 1422 478258 1464 478494
rect 1144 471494 1464 478258
rect 1144 471258 1186 471494
rect 1422 471258 1464 471494
rect 1144 464494 1464 471258
rect 1144 464258 1186 464494
rect 1422 464258 1464 464494
rect 1144 457494 1464 464258
rect 1144 457258 1186 457494
rect 1422 457258 1464 457494
rect 1144 450494 1464 457258
rect 1144 450258 1186 450494
rect 1422 450258 1464 450494
rect 1144 443494 1464 450258
rect 1144 443258 1186 443494
rect 1422 443258 1464 443494
rect 1144 436494 1464 443258
rect 1144 436258 1186 436494
rect 1422 436258 1464 436494
rect 1144 429494 1464 436258
rect 1144 429258 1186 429494
rect 1422 429258 1464 429494
rect 1144 422494 1464 429258
rect 1144 422258 1186 422494
rect 1422 422258 1464 422494
rect 1144 415494 1464 422258
rect 1144 415258 1186 415494
rect 1422 415258 1464 415494
rect 1144 408494 1464 415258
rect 1144 408258 1186 408494
rect 1422 408258 1464 408494
rect 1144 401494 1464 408258
rect 1144 401258 1186 401494
rect 1422 401258 1464 401494
rect 1144 394494 1464 401258
rect 1144 394258 1186 394494
rect 1422 394258 1464 394494
rect 1144 387494 1464 394258
rect 1144 387258 1186 387494
rect 1422 387258 1464 387494
rect 1144 380494 1464 387258
rect 1144 380258 1186 380494
rect 1422 380258 1464 380494
rect 1144 373494 1464 380258
rect 1144 373258 1186 373494
rect 1422 373258 1464 373494
rect 1144 366494 1464 373258
rect 1144 366258 1186 366494
rect 1422 366258 1464 366494
rect 1144 359494 1464 366258
rect 1144 359258 1186 359494
rect 1422 359258 1464 359494
rect 1144 352494 1464 359258
rect 1144 352258 1186 352494
rect 1422 352258 1464 352494
rect 1144 345494 1464 352258
rect 1144 345258 1186 345494
rect 1422 345258 1464 345494
rect 1144 338494 1464 345258
rect 1144 338258 1186 338494
rect 1422 338258 1464 338494
rect 1144 331494 1464 338258
rect 1144 331258 1186 331494
rect 1422 331258 1464 331494
rect 1144 324494 1464 331258
rect 1144 324258 1186 324494
rect 1422 324258 1464 324494
rect 1144 317494 1464 324258
rect 1144 317258 1186 317494
rect 1422 317258 1464 317494
rect 1144 310494 1464 317258
rect 1144 310258 1186 310494
rect 1422 310258 1464 310494
rect 1144 303494 1464 310258
rect 1144 303258 1186 303494
rect 1422 303258 1464 303494
rect 1144 296494 1464 303258
rect 1144 296258 1186 296494
rect 1422 296258 1464 296494
rect 1144 289494 1464 296258
rect 1144 289258 1186 289494
rect 1422 289258 1464 289494
rect 1144 282494 1464 289258
rect 1144 282258 1186 282494
rect 1422 282258 1464 282494
rect 1144 275494 1464 282258
rect 1144 275258 1186 275494
rect 1422 275258 1464 275494
rect 1144 268494 1464 275258
rect 1144 268258 1186 268494
rect 1422 268258 1464 268494
rect 1144 261494 1464 268258
rect 1144 261258 1186 261494
rect 1422 261258 1464 261494
rect 1144 254494 1464 261258
rect 1144 254258 1186 254494
rect 1422 254258 1464 254494
rect 1144 247494 1464 254258
rect 1144 247258 1186 247494
rect 1422 247258 1464 247494
rect 1144 240494 1464 247258
rect 1144 240258 1186 240494
rect 1422 240258 1464 240494
rect 1144 233494 1464 240258
rect 1144 233258 1186 233494
rect 1422 233258 1464 233494
rect 1144 226494 1464 233258
rect 1144 226258 1186 226494
rect 1422 226258 1464 226494
rect 1144 219494 1464 226258
rect 1144 219258 1186 219494
rect 1422 219258 1464 219494
rect 1144 212494 1464 219258
rect 1144 212258 1186 212494
rect 1422 212258 1464 212494
rect 1144 205494 1464 212258
rect 1144 205258 1186 205494
rect 1422 205258 1464 205494
rect 1144 198494 1464 205258
rect 1144 198258 1186 198494
rect 1422 198258 1464 198494
rect 1144 191494 1464 198258
rect 1144 191258 1186 191494
rect 1422 191258 1464 191494
rect 1144 184494 1464 191258
rect 1144 184258 1186 184494
rect 1422 184258 1464 184494
rect 1144 177494 1464 184258
rect 1144 177258 1186 177494
rect 1422 177258 1464 177494
rect 1144 170494 1464 177258
rect 1144 170258 1186 170494
rect 1422 170258 1464 170494
rect 1144 163494 1464 170258
rect 1144 163258 1186 163494
rect 1422 163258 1464 163494
rect 1144 156494 1464 163258
rect 1144 156258 1186 156494
rect 1422 156258 1464 156494
rect 1144 149494 1464 156258
rect 1144 149258 1186 149494
rect 1422 149258 1464 149494
rect 1144 142494 1464 149258
rect 1144 142258 1186 142494
rect 1422 142258 1464 142494
rect 1144 135494 1464 142258
rect 1144 135258 1186 135494
rect 1422 135258 1464 135494
rect 1144 128494 1464 135258
rect 1144 128258 1186 128494
rect 1422 128258 1464 128494
rect 1144 121494 1464 128258
rect 1144 121258 1186 121494
rect 1422 121258 1464 121494
rect 1144 114494 1464 121258
rect 1144 114258 1186 114494
rect 1422 114258 1464 114494
rect 1144 107494 1464 114258
rect 1144 107258 1186 107494
rect 1422 107258 1464 107494
rect 1144 100494 1464 107258
rect 1144 100258 1186 100494
rect 1422 100258 1464 100494
rect 1144 93494 1464 100258
rect 1144 93258 1186 93494
rect 1422 93258 1464 93494
rect 1144 86494 1464 93258
rect 1144 86258 1186 86494
rect 1422 86258 1464 86494
rect 1144 79494 1464 86258
rect 1144 79258 1186 79494
rect 1422 79258 1464 79494
rect 1144 72494 1464 79258
rect 1144 72258 1186 72494
rect 1422 72258 1464 72494
rect 1144 65494 1464 72258
rect 1144 65258 1186 65494
rect 1422 65258 1464 65494
rect 1144 58494 1464 65258
rect 1144 58258 1186 58494
rect 1422 58258 1464 58494
rect 1144 51494 1464 58258
rect 1144 51258 1186 51494
rect 1422 51258 1464 51494
rect 1144 44494 1464 51258
rect 1144 44258 1186 44494
rect 1422 44258 1464 44494
rect 1144 37494 1464 44258
rect 1144 37258 1186 37494
rect 1422 37258 1464 37494
rect 1144 30494 1464 37258
rect 1144 30258 1186 30494
rect 1422 30258 1464 30494
rect 1144 23494 1464 30258
rect 1144 23258 1186 23494
rect 1422 23258 1464 23494
rect 1144 16494 1464 23258
rect 1144 16258 1186 16494
rect 1422 16258 1464 16494
rect 1144 9494 1464 16258
rect 1144 9258 1186 9494
rect 1422 9258 1464 9494
rect 1144 2494 1464 9258
rect 1144 2258 1186 2494
rect 1422 2258 1464 2494
rect 1144 -746 1464 2258
rect 1144 -982 1186 -746
rect 1422 -982 1464 -746
rect 1144 -1066 1464 -982
rect 1144 -1302 1186 -1066
rect 1422 -1302 1464 -1066
rect 1144 -2294 1464 -1302
rect 2876 706198 3196 706230
rect 2876 705962 2918 706198
rect 3154 705962 3196 706198
rect 2876 705878 3196 705962
rect 2876 705642 2918 705878
rect 3154 705642 3196 705878
rect 2876 696434 3196 705642
rect 2876 696198 2918 696434
rect 3154 696198 3196 696434
rect 2876 689434 3196 696198
rect 2876 689198 2918 689434
rect 3154 689198 3196 689434
rect 2876 682434 3196 689198
rect 2876 682198 2918 682434
rect 3154 682198 3196 682434
rect 2876 675434 3196 682198
rect 2876 675198 2918 675434
rect 3154 675198 3196 675434
rect 2876 668434 3196 675198
rect 2876 668198 2918 668434
rect 3154 668198 3196 668434
rect 2876 661434 3196 668198
rect 2876 661198 2918 661434
rect 3154 661198 3196 661434
rect 2876 654434 3196 661198
rect 2876 654198 2918 654434
rect 3154 654198 3196 654434
rect 2876 647434 3196 654198
rect 2876 647198 2918 647434
rect 3154 647198 3196 647434
rect 2876 640434 3196 647198
rect 2876 640198 2918 640434
rect 3154 640198 3196 640434
rect 2876 633434 3196 640198
rect 2876 633198 2918 633434
rect 3154 633198 3196 633434
rect 2876 626434 3196 633198
rect 2876 626198 2918 626434
rect 3154 626198 3196 626434
rect 2876 619434 3196 626198
rect 2876 619198 2918 619434
rect 3154 619198 3196 619434
rect 2876 612434 3196 619198
rect 2876 612198 2918 612434
rect 3154 612198 3196 612434
rect 2876 605434 3196 612198
rect 2876 605198 2918 605434
rect 3154 605198 3196 605434
rect 2876 598434 3196 605198
rect 2876 598198 2918 598434
rect 3154 598198 3196 598434
rect 2876 591434 3196 598198
rect 2876 591198 2918 591434
rect 3154 591198 3196 591434
rect 2876 584434 3196 591198
rect 2876 584198 2918 584434
rect 3154 584198 3196 584434
rect 2876 577434 3196 584198
rect 2876 577198 2918 577434
rect 3154 577198 3196 577434
rect 2876 570434 3196 577198
rect 2876 570198 2918 570434
rect 3154 570198 3196 570434
rect 2876 563434 3196 570198
rect 2876 563198 2918 563434
rect 3154 563198 3196 563434
rect 2876 556434 3196 563198
rect 2876 556198 2918 556434
rect 3154 556198 3196 556434
rect 2876 549434 3196 556198
rect 2876 549198 2918 549434
rect 3154 549198 3196 549434
rect 2876 542434 3196 549198
rect 2876 542198 2918 542434
rect 3154 542198 3196 542434
rect 2876 535434 3196 542198
rect 2876 535198 2918 535434
rect 3154 535198 3196 535434
rect 2876 528434 3196 535198
rect 2876 528198 2918 528434
rect 3154 528198 3196 528434
rect 2876 521434 3196 528198
rect 2876 521198 2918 521434
rect 3154 521198 3196 521434
rect 2876 514434 3196 521198
rect 2876 514198 2918 514434
rect 3154 514198 3196 514434
rect 2876 507434 3196 514198
rect 2876 507198 2918 507434
rect 3154 507198 3196 507434
rect 2876 500434 3196 507198
rect 2876 500198 2918 500434
rect 3154 500198 3196 500434
rect 2876 493434 3196 500198
rect 2876 493198 2918 493434
rect 3154 493198 3196 493434
rect 2876 486434 3196 493198
rect 2876 486198 2918 486434
rect 3154 486198 3196 486434
rect 2876 479434 3196 486198
rect 2876 479198 2918 479434
rect 3154 479198 3196 479434
rect 2876 472434 3196 479198
rect 2876 472198 2918 472434
rect 3154 472198 3196 472434
rect 2876 465434 3196 472198
rect 2876 465198 2918 465434
rect 3154 465198 3196 465434
rect 2876 458434 3196 465198
rect 2876 458198 2918 458434
rect 3154 458198 3196 458434
rect 2876 451434 3196 458198
rect 2876 451198 2918 451434
rect 3154 451198 3196 451434
rect 2876 444434 3196 451198
rect 2876 444198 2918 444434
rect 3154 444198 3196 444434
rect 2876 437434 3196 444198
rect 2876 437198 2918 437434
rect 3154 437198 3196 437434
rect 2876 430434 3196 437198
rect 2876 430198 2918 430434
rect 3154 430198 3196 430434
rect 2876 423434 3196 430198
rect 2876 423198 2918 423434
rect 3154 423198 3196 423434
rect 2876 416434 3196 423198
rect 2876 416198 2918 416434
rect 3154 416198 3196 416434
rect 2876 409434 3196 416198
rect 2876 409198 2918 409434
rect 3154 409198 3196 409434
rect 2876 402434 3196 409198
rect 2876 402198 2918 402434
rect 3154 402198 3196 402434
rect 2876 395434 3196 402198
rect 2876 395198 2918 395434
rect 3154 395198 3196 395434
rect 2876 388434 3196 395198
rect 2876 388198 2918 388434
rect 3154 388198 3196 388434
rect 2876 381434 3196 388198
rect 2876 381198 2918 381434
rect 3154 381198 3196 381434
rect 2876 374434 3196 381198
rect 2876 374198 2918 374434
rect 3154 374198 3196 374434
rect 2876 367434 3196 374198
rect 2876 367198 2918 367434
rect 3154 367198 3196 367434
rect 2876 360434 3196 367198
rect 2876 360198 2918 360434
rect 3154 360198 3196 360434
rect 2876 353434 3196 360198
rect 2876 353198 2918 353434
rect 3154 353198 3196 353434
rect 2876 346434 3196 353198
rect 2876 346198 2918 346434
rect 3154 346198 3196 346434
rect 2876 339434 3196 346198
rect 2876 339198 2918 339434
rect 3154 339198 3196 339434
rect 2876 332434 3196 339198
rect 2876 332198 2918 332434
rect 3154 332198 3196 332434
rect 2876 325434 3196 332198
rect 2876 325198 2918 325434
rect 3154 325198 3196 325434
rect 2876 318434 3196 325198
rect 2876 318198 2918 318434
rect 3154 318198 3196 318434
rect 2876 311434 3196 318198
rect 2876 311198 2918 311434
rect 3154 311198 3196 311434
rect 2876 304434 3196 311198
rect 2876 304198 2918 304434
rect 3154 304198 3196 304434
rect 2876 297434 3196 304198
rect 2876 297198 2918 297434
rect 3154 297198 3196 297434
rect 2876 290434 3196 297198
rect 2876 290198 2918 290434
rect 3154 290198 3196 290434
rect 2876 283434 3196 290198
rect 2876 283198 2918 283434
rect 3154 283198 3196 283434
rect 2876 276434 3196 283198
rect 2876 276198 2918 276434
rect 3154 276198 3196 276434
rect 2876 269434 3196 276198
rect 2876 269198 2918 269434
rect 3154 269198 3196 269434
rect 2876 262434 3196 269198
rect 2876 262198 2918 262434
rect 3154 262198 3196 262434
rect 2876 255434 3196 262198
rect 2876 255198 2918 255434
rect 3154 255198 3196 255434
rect 2876 248434 3196 255198
rect 2876 248198 2918 248434
rect 3154 248198 3196 248434
rect 2876 241434 3196 248198
rect 2876 241198 2918 241434
rect 3154 241198 3196 241434
rect 2876 234434 3196 241198
rect 2876 234198 2918 234434
rect 3154 234198 3196 234434
rect 2876 227434 3196 234198
rect 2876 227198 2918 227434
rect 3154 227198 3196 227434
rect 2876 220434 3196 227198
rect 2876 220198 2918 220434
rect 3154 220198 3196 220434
rect 2876 213434 3196 220198
rect 2876 213198 2918 213434
rect 3154 213198 3196 213434
rect 2876 206434 3196 213198
rect 2876 206198 2918 206434
rect 3154 206198 3196 206434
rect 2876 199434 3196 206198
rect 2876 199198 2918 199434
rect 3154 199198 3196 199434
rect 2876 192434 3196 199198
rect 2876 192198 2918 192434
rect 3154 192198 3196 192434
rect 2876 185434 3196 192198
rect 2876 185198 2918 185434
rect 3154 185198 3196 185434
rect 2876 178434 3196 185198
rect 2876 178198 2918 178434
rect 3154 178198 3196 178434
rect 2876 171434 3196 178198
rect 2876 171198 2918 171434
rect 3154 171198 3196 171434
rect 2876 164434 3196 171198
rect 2876 164198 2918 164434
rect 3154 164198 3196 164434
rect 2876 157434 3196 164198
rect 2876 157198 2918 157434
rect 3154 157198 3196 157434
rect 2876 150434 3196 157198
rect 2876 150198 2918 150434
rect 3154 150198 3196 150434
rect 2876 143434 3196 150198
rect 2876 143198 2918 143434
rect 3154 143198 3196 143434
rect 2876 136434 3196 143198
rect 2876 136198 2918 136434
rect 3154 136198 3196 136434
rect 2876 129434 3196 136198
rect 2876 129198 2918 129434
rect 3154 129198 3196 129434
rect 2876 122434 3196 129198
rect 2876 122198 2918 122434
rect 3154 122198 3196 122434
rect 2876 115434 3196 122198
rect 2876 115198 2918 115434
rect 3154 115198 3196 115434
rect 2876 108434 3196 115198
rect 2876 108198 2918 108434
rect 3154 108198 3196 108434
rect 2876 101434 3196 108198
rect 2876 101198 2918 101434
rect 3154 101198 3196 101434
rect 2876 94434 3196 101198
rect 2876 94198 2918 94434
rect 3154 94198 3196 94434
rect 2876 87434 3196 94198
rect 2876 87198 2918 87434
rect 3154 87198 3196 87434
rect 2876 80434 3196 87198
rect 2876 80198 2918 80434
rect 3154 80198 3196 80434
rect 2876 73434 3196 80198
rect 2876 73198 2918 73434
rect 3154 73198 3196 73434
rect 2876 66434 3196 73198
rect 2876 66198 2918 66434
rect 3154 66198 3196 66434
rect 2876 59434 3196 66198
rect 2876 59198 2918 59434
rect 3154 59198 3196 59434
rect 2876 52434 3196 59198
rect 2876 52198 2918 52434
rect 3154 52198 3196 52434
rect 2876 45434 3196 52198
rect 2876 45198 2918 45434
rect 3154 45198 3196 45434
rect 2876 38434 3196 45198
rect 2876 38198 2918 38434
rect 3154 38198 3196 38434
rect 2876 31434 3196 38198
rect 2876 31198 2918 31434
rect 3154 31198 3196 31434
rect 2876 24434 3196 31198
rect 2876 24198 2918 24434
rect 3154 24198 3196 24434
rect 2876 17434 3196 24198
rect 2876 17198 2918 17434
rect 3154 17198 3196 17434
rect 2876 10434 3196 17198
rect 2876 10198 2918 10434
rect 3154 10198 3196 10434
rect 2876 3434 3196 10198
rect 2876 3198 2918 3434
rect 3154 3198 3196 3434
rect 2876 -1706 3196 3198
rect 2876 -1942 2918 -1706
rect 3154 -1942 3196 -1706
rect 2876 -2026 3196 -1942
rect 2876 -2262 2918 -2026
rect 3154 -2262 3196 -2026
rect 2876 -2294 3196 -2262
rect 8144 705238 8464 706230
rect 8144 705002 8186 705238
rect 8422 705002 8464 705238
rect 8144 704918 8464 705002
rect 8144 704682 8186 704918
rect 8422 704682 8464 704918
rect 8144 695494 8464 704682
rect 8144 695258 8186 695494
rect 8422 695258 8464 695494
rect 8144 688494 8464 695258
rect 8144 688258 8186 688494
rect 8422 688258 8464 688494
rect 8144 681494 8464 688258
rect 8144 681258 8186 681494
rect 8422 681258 8464 681494
rect 8144 674494 8464 681258
rect 8144 674258 8186 674494
rect 8422 674258 8464 674494
rect 8144 667494 8464 674258
rect 8144 667258 8186 667494
rect 8422 667258 8464 667494
rect 8144 660494 8464 667258
rect 8144 660258 8186 660494
rect 8422 660258 8464 660494
rect 8144 653494 8464 660258
rect 8144 653258 8186 653494
rect 8422 653258 8464 653494
rect 8144 646494 8464 653258
rect 8144 646258 8186 646494
rect 8422 646258 8464 646494
rect 8144 639494 8464 646258
rect 8144 639258 8186 639494
rect 8422 639258 8464 639494
rect 8144 632494 8464 639258
rect 8144 632258 8186 632494
rect 8422 632258 8464 632494
rect 8144 625494 8464 632258
rect 8144 625258 8186 625494
rect 8422 625258 8464 625494
rect 8144 618494 8464 625258
rect 8144 618258 8186 618494
rect 8422 618258 8464 618494
rect 8144 611494 8464 618258
rect 8144 611258 8186 611494
rect 8422 611258 8464 611494
rect 8144 604494 8464 611258
rect 8144 604258 8186 604494
rect 8422 604258 8464 604494
rect 8144 597494 8464 604258
rect 8144 597258 8186 597494
rect 8422 597258 8464 597494
rect 8144 590494 8464 597258
rect 8144 590258 8186 590494
rect 8422 590258 8464 590494
rect 8144 583494 8464 590258
rect 8144 583258 8186 583494
rect 8422 583258 8464 583494
rect 8144 576494 8464 583258
rect 8144 576258 8186 576494
rect 8422 576258 8464 576494
rect 8144 569494 8464 576258
rect 8144 569258 8186 569494
rect 8422 569258 8464 569494
rect 8144 562494 8464 569258
rect 8144 562258 8186 562494
rect 8422 562258 8464 562494
rect 8144 555494 8464 562258
rect 8144 555258 8186 555494
rect 8422 555258 8464 555494
rect 8144 548494 8464 555258
rect 8144 548258 8186 548494
rect 8422 548258 8464 548494
rect 8144 541494 8464 548258
rect 8144 541258 8186 541494
rect 8422 541258 8464 541494
rect 8144 534494 8464 541258
rect 8144 534258 8186 534494
rect 8422 534258 8464 534494
rect 8144 527494 8464 534258
rect 8144 527258 8186 527494
rect 8422 527258 8464 527494
rect 8144 520494 8464 527258
rect 8144 520258 8186 520494
rect 8422 520258 8464 520494
rect 8144 513494 8464 520258
rect 8144 513258 8186 513494
rect 8422 513258 8464 513494
rect 8144 506494 8464 513258
rect 8144 506258 8186 506494
rect 8422 506258 8464 506494
rect 8144 499494 8464 506258
rect 8144 499258 8186 499494
rect 8422 499258 8464 499494
rect 8144 492494 8464 499258
rect 8144 492258 8186 492494
rect 8422 492258 8464 492494
rect 8144 485494 8464 492258
rect 8144 485258 8186 485494
rect 8422 485258 8464 485494
rect 8144 478494 8464 485258
rect 8144 478258 8186 478494
rect 8422 478258 8464 478494
rect 8144 471494 8464 478258
rect 8144 471258 8186 471494
rect 8422 471258 8464 471494
rect 8144 464494 8464 471258
rect 8144 464258 8186 464494
rect 8422 464258 8464 464494
rect 8144 457494 8464 464258
rect 8144 457258 8186 457494
rect 8422 457258 8464 457494
rect 8144 450494 8464 457258
rect 8144 450258 8186 450494
rect 8422 450258 8464 450494
rect 8144 443494 8464 450258
rect 8144 443258 8186 443494
rect 8422 443258 8464 443494
rect 8144 436494 8464 443258
rect 8144 436258 8186 436494
rect 8422 436258 8464 436494
rect 8144 429494 8464 436258
rect 8144 429258 8186 429494
rect 8422 429258 8464 429494
rect 8144 422494 8464 429258
rect 8144 422258 8186 422494
rect 8422 422258 8464 422494
rect 8144 415494 8464 422258
rect 8144 415258 8186 415494
rect 8422 415258 8464 415494
rect 8144 408494 8464 415258
rect 8144 408258 8186 408494
rect 8422 408258 8464 408494
rect 8144 401494 8464 408258
rect 8144 401258 8186 401494
rect 8422 401258 8464 401494
rect 8144 394494 8464 401258
rect 8144 394258 8186 394494
rect 8422 394258 8464 394494
rect 8144 387494 8464 394258
rect 8144 387258 8186 387494
rect 8422 387258 8464 387494
rect 8144 380494 8464 387258
rect 8144 380258 8186 380494
rect 8422 380258 8464 380494
rect 8144 373494 8464 380258
rect 8144 373258 8186 373494
rect 8422 373258 8464 373494
rect 8144 366494 8464 373258
rect 8144 366258 8186 366494
rect 8422 366258 8464 366494
rect 8144 359494 8464 366258
rect 8144 359258 8186 359494
rect 8422 359258 8464 359494
rect 8144 352494 8464 359258
rect 8144 352258 8186 352494
rect 8422 352258 8464 352494
rect 8144 345494 8464 352258
rect 8144 345258 8186 345494
rect 8422 345258 8464 345494
rect 8144 338494 8464 345258
rect 8144 338258 8186 338494
rect 8422 338258 8464 338494
rect 8144 331494 8464 338258
rect 8144 331258 8186 331494
rect 8422 331258 8464 331494
rect 8144 324494 8464 331258
rect 8144 324258 8186 324494
rect 8422 324258 8464 324494
rect 8144 317494 8464 324258
rect 8144 317258 8186 317494
rect 8422 317258 8464 317494
rect 8144 310494 8464 317258
rect 8144 310258 8186 310494
rect 8422 310258 8464 310494
rect 8144 303494 8464 310258
rect 8144 303258 8186 303494
rect 8422 303258 8464 303494
rect 8144 296494 8464 303258
rect 8144 296258 8186 296494
rect 8422 296258 8464 296494
rect 8144 289494 8464 296258
rect 8144 289258 8186 289494
rect 8422 289258 8464 289494
rect 8144 282494 8464 289258
rect 8144 282258 8186 282494
rect 8422 282258 8464 282494
rect 8144 275494 8464 282258
rect 8144 275258 8186 275494
rect 8422 275258 8464 275494
rect 8144 268494 8464 275258
rect 8144 268258 8186 268494
rect 8422 268258 8464 268494
rect 8144 261494 8464 268258
rect 8144 261258 8186 261494
rect 8422 261258 8464 261494
rect 8144 254494 8464 261258
rect 8144 254258 8186 254494
rect 8422 254258 8464 254494
rect 8144 247494 8464 254258
rect 8144 247258 8186 247494
rect 8422 247258 8464 247494
rect 8144 240494 8464 247258
rect 8144 240258 8186 240494
rect 8422 240258 8464 240494
rect 8144 233494 8464 240258
rect 8144 233258 8186 233494
rect 8422 233258 8464 233494
rect 8144 226494 8464 233258
rect 8144 226258 8186 226494
rect 8422 226258 8464 226494
rect 8144 219494 8464 226258
rect 8144 219258 8186 219494
rect 8422 219258 8464 219494
rect 8144 212494 8464 219258
rect 8144 212258 8186 212494
rect 8422 212258 8464 212494
rect 8144 205494 8464 212258
rect 8144 205258 8186 205494
rect 8422 205258 8464 205494
rect 8144 198494 8464 205258
rect 8144 198258 8186 198494
rect 8422 198258 8464 198494
rect 8144 191494 8464 198258
rect 8144 191258 8186 191494
rect 8422 191258 8464 191494
rect 8144 184494 8464 191258
rect 8144 184258 8186 184494
rect 8422 184258 8464 184494
rect 8144 177494 8464 184258
rect 8144 177258 8186 177494
rect 8422 177258 8464 177494
rect 8144 170494 8464 177258
rect 8144 170258 8186 170494
rect 8422 170258 8464 170494
rect 8144 163494 8464 170258
rect 8144 163258 8186 163494
rect 8422 163258 8464 163494
rect 8144 156494 8464 163258
rect 8144 156258 8186 156494
rect 8422 156258 8464 156494
rect 8144 149494 8464 156258
rect 8144 149258 8186 149494
rect 8422 149258 8464 149494
rect 8144 142494 8464 149258
rect 8144 142258 8186 142494
rect 8422 142258 8464 142494
rect 8144 135494 8464 142258
rect 8144 135258 8186 135494
rect 8422 135258 8464 135494
rect 8144 128494 8464 135258
rect 8144 128258 8186 128494
rect 8422 128258 8464 128494
rect 8144 121494 8464 128258
rect 8144 121258 8186 121494
rect 8422 121258 8464 121494
rect 8144 114494 8464 121258
rect 8144 114258 8186 114494
rect 8422 114258 8464 114494
rect 8144 107494 8464 114258
rect 8144 107258 8186 107494
rect 8422 107258 8464 107494
rect 8144 100494 8464 107258
rect 8144 100258 8186 100494
rect 8422 100258 8464 100494
rect 8144 93494 8464 100258
rect 8144 93258 8186 93494
rect 8422 93258 8464 93494
rect 8144 86494 8464 93258
rect 8144 86258 8186 86494
rect 8422 86258 8464 86494
rect 8144 79494 8464 86258
rect 8144 79258 8186 79494
rect 8422 79258 8464 79494
rect 8144 72494 8464 79258
rect 8144 72258 8186 72494
rect 8422 72258 8464 72494
rect 8144 65494 8464 72258
rect 8144 65258 8186 65494
rect 8422 65258 8464 65494
rect 8144 58494 8464 65258
rect 8144 58258 8186 58494
rect 8422 58258 8464 58494
rect 8144 51494 8464 58258
rect 8144 51258 8186 51494
rect 8422 51258 8464 51494
rect 8144 44494 8464 51258
rect 8144 44258 8186 44494
rect 8422 44258 8464 44494
rect 8144 37494 8464 44258
rect 8144 37258 8186 37494
rect 8422 37258 8464 37494
rect 8144 30494 8464 37258
rect 8144 30258 8186 30494
rect 8422 30258 8464 30494
rect 8144 23494 8464 30258
rect 8144 23258 8186 23494
rect 8422 23258 8464 23494
rect 8144 16494 8464 23258
rect 8144 16258 8186 16494
rect 8422 16258 8464 16494
rect 8144 9494 8464 16258
rect 8144 9258 8186 9494
rect 8422 9258 8464 9494
rect 8144 2494 8464 9258
rect 8144 2258 8186 2494
rect 8422 2258 8464 2494
rect 8144 -746 8464 2258
rect 8144 -982 8186 -746
rect 8422 -982 8464 -746
rect 8144 -1066 8464 -982
rect 8144 -1302 8186 -1066
rect 8422 -1302 8464 -1066
rect 8144 -2294 8464 -1302
rect 9876 706198 10196 706230
rect 9876 705962 9918 706198
rect 10154 705962 10196 706198
rect 9876 705878 10196 705962
rect 9876 705642 9918 705878
rect 10154 705642 10196 705878
rect 9876 696434 10196 705642
rect 9876 696198 9918 696434
rect 10154 696198 10196 696434
rect 9876 689434 10196 696198
rect 9876 689198 9918 689434
rect 10154 689198 10196 689434
rect 9876 682434 10196 689198
rect 9876 682198 9918 682434
rect 10154 682198 10196 682434
rect 9876 675434 10196 682198
rect 9876 675198 9918 675434
rect 10154 675198 10196 675434
rect 9876 668434 10196 675198
rect 9876 668198 9918 668434
rect 10154 668198 10196 668434
rect 9876 661434 10196 668198
rect 9876 661198 9918 661434
rect 10154 661198 10196 661434
rect 9876 654434 10196 661198
rect 9876 654198 9918 654434
rect 10154 654198 10196 654434
rect 9876 647434 10196 654198
rect 9876 647198 9918 647434
rect 10154 647198 10196 647434
rect 9876 640434 10196 647198
rect 9876 640198 9918 640434
rect 10154 640198 10196 640434
rect 9876 633434 10196 640198
rect 9876 633198 9918 633434
rect 10154 633198 10196 633434
rect 9876 626434 10196 633198
rect 9876 626198 9918 626434
rect 10154 626198 10196 626434
rect 9876 619434 10196 626198
rect 9876 619198 9918 619434
rect 10154 619198 10196 619434
rect 9876 612434 10196 619198
rect 9876 612198 9918 612434
rect 10154 612198 10196 612434
rect 9876 605434 10196 612198
rect 9876 605198 9918 605434
rect 10154 605198 10196 605434
rect 9876 598434 10196 605198
rect 9876 598198 9918 598434
rect 10154 598198 10196 598434
rect 9876 591434 10196 598198
rect 9876 591198 9918 591434
rect 10154 591198 10196 591434
rect 9876 584434 10196 591198
rect 9876 584198 9918 584434
rect 10154 584198 10196 584434
rect 9876 577434 10196 584198
rect 9876 577198 9918 577434
rect 10154 577198 10196 577434
rect 9876 570434 10196 577198
rect 9876 570198 9918 570434
rect 10154 570198 10196 570434
rect 9876 563434 10196 570198
rect 9876 563198 9918 563434
rect 10154 563198 10196 563434
rect 9876 556434 10196 563198
rect 9876 556198 9918 556434
rect 10154 556198 10196 556434
rect 9876 549434 10196 556198
rect 9876 549198 9918 549434
rect 10154 549198 10196 549434
rect 9876 542434 10196 549198
rect 9876 542198 9918 542434
rect 10154 542198 10196 542434
rect 9876 535434 10196 542198
rect 9876 535198 9918 535434
rect 10154 535198 10196 535434
rect 9876 528434 10196 535198
rect 9876 528198 9918 528434
rect 10154 528198 10196 528434
rect 9876 521434 10196 528198
rect 9876 521198 9918 521434
rect 10154 521198 10196 521434
rect 9876 514434 10196 521198
rect 9876 514198 9918 514434
rect 10154 514198 10196 514434
rect 9876 507434 10196 514198
rect 9876 507198 9918 507434
rect 10154 507198 10196 507434
rect 9876 500434 10196 507198
rect 9876 500198 9918 500434
rect 10154 500198 10196 500434
rect 9876 493434 10196 500198
rect 9876 493198 9918 493434
rect 10154 493198 10196 493434
rect 9876 486434 10196 493198
rect 9876 486198 9918 486434
rect 10154 486198 10196 486434
rect 9876 479434 10196 486198
rect 9876 479198 9918 479434
rect 10154 479198 10196 479434
rect 9876 472434 10196 479198
rect 9876 472198 9918 472434
rect 10154 472198 10196 472434
rect 9876 465434 10196 472198
rect 9876 465198 9918 465434
rect 10154 465198 10196 465434
rect 9876 458434 10196 465198
rect 9876 458198 9918 458434
rect 10154 458198 10196 458434
rect 9876 451434 10196 458198
rect 9876 451198 9918 451434
rect 10154 451198 10196 451434
rect 9876 444434 10196 451198
rect 9876 444198 9918 444434
rect 10154 444198 10196 444434
rect 9876 437434 10196 444198
rect 9876 437198 9918 437434
rect 10154 437198 10196 437434
rect 9876 430434 10196 437198
rect 9876 430198 9918 430434
rect 10154 430198 10196 430434
rect 9876 423434 10196 430198
rect 9876 423198 9918 423434
rect 10154 423198 10196 423434
rect 9876 416434 10196 423198
rect 9876 416198 9918 416434
rect 10154 416198 10196 416434
rect 9876 409434 10196 416198
rect 9876 409198 9918 409434
rect 10154 409198 10196 409434
rect 9876 402434 10196 409198
rect 9876 402198 9918 402434
rect 10154 402198 10196 402434
rect 9876 395434 10196 402198
rect 9876 395198 9918 395434
rect 10154 395198 10196 395434
rect 9876 388434 10196 395198
rect 9876 388198 9918 388434
rect 10154 388198 10196 388434
rect 9876 381434 10196 388198
rect 9876 381198 9918 381434
rect 10154 381198 10196 381434
rect 9876 374434 10196 381198
rect 9876 374198 9918 374434
rect 10154 374198 10196 374434
rect 9876 367434 10196 374198
rect 9876 367198 9918 367434
rect 10154 367198 10196 367434
rect 9876 360434 10196 367198
rect 9876 360198 9918 360434
rect 10154 360198 10196 360434
rect 9876 353434 10196 360198
rect 9876 353198 9918 353434
rect 10154 353198 10196 353434
rect 9876 346434 10196 353198
rect 9876 346198 9918 346434
rect 10154 346198 10196 346434
rect 9876 339434 10196 346198
rect 9876 339198 9918 339434
rect 10154 339198 10196 339434
rect 9876 332434 10196 339198
rect 9876 332198 9918 332434
rect 10154 332198 10196 332434
rect 9876 325434 10196 332198
rect 9876 325198 9918 325434
rect 10154 325198 10196 325434
rect 9876 318434 10196 325198
rect 9876 318198 9918 318434
rect 10154 318198 10196 318434
rect 9876 311434 10196 318198
rect 9876 311198 9918 311434
rect 10154 311198 10196 311434
rect 9876 304434 10196 311198
rect 9876 304198 9918 304434
rect 10154 304198 10196 304434
rect 9876 297434 10196 304198
rect 9876 297198 9918 297434
rect 10154 297198 10196 297434
rect 9876 290434 10196 297198
rect 9876 290198 9918 290434
rect 10154 290198 10196 290434
rect 9876 283434 10196 290198
rect 9876 283198 9918 283434
rect 10154 283198 10196 283434
rect 9876 276434 10196 283198
rect 9876 276198 9918 276434
rect 10154 276198 10196 276434
rect 9876 269434 10196 276198
rect 9876 269198 9918 269434
rect 10154 269198 10196 269434
rect 9876 262434 10196 269198
rect 9876 262198 9918 262434
rect 10154 262198 10196 262434
rect 9876 255434 10196 262198
rect 9876 255198 9918 255434
rect 10154 255198 10196 255434
rect 9876 248434 10196 255198
rect 9876 248198 9918 248434
rect 10154 248198 10196 248434
rect 9876 241434 10196 248198
rect 9876 241198 9918 241434
rect 10154 241198 10196 241434
rect 9876 234434 10196 241198
rect 9876 234198 9918 234434
rect 10154 234198 10196 234434
rect 9876 227434 10196 234198
rect 9876 227198 9918 227434
rect 10154 227198 10196 227434
rect 9876 220434 10196 227198
rect 9876 220198 9918 220434
rect 10154 220198 10196 220434
rect 9876 213434 10196 220198
rect 9876 213198 9918 213434
rect 10154 213198 10196 213434
rect 9876 206434 10196 213198
rect 9876 206198 9918 206434
rect 10154 206198 10196 206434
rect 9876 199434 10196 206198
rect 9876 199198 9918 199434
rect 10154 199198 10196 199434
rect 9876 192434 10196 199198
rect 9876 192198 9918 192434
rect 10154 192198 10196 192434
rect 9876 185434 10196 192198
rect 9876 185198 9918 185434
rect 10154 185198 10196 185434
rect 9876 178434 10196 185198
rect 9876 178198 9918 178434
rect 10154 178198 10196 178434
rect 9876 171434 10196 178198
rect 9876 171198 9918 171434
rect 10154 171198 10196 171434
rect 9876 164434 10196 171198
rect 9876 164198 9918 164434
rect 10154 164198 10196 164434
rect 9876 157434 10196 164198
rect 9876 157198 9918 157434
rect 10154 157198 10196 157434
rect 9876 150434 10196 157198
rect 9876 150198 9918 150434
rect 10154 150198 10196 150434
rect 9876 143434 10196 150198
rect 9876 143198 9918 143434
rect 10154 143198 10196 143434
rect 9876 136434 10196 143198
rect 9876 136198 9918 136434
rect 10154 136198 10196 136434
rect 9876 129434 10196 136198
rect 9876 129198 9918 129434
rect 10154 129198 10196 129434
rect 9876 122434 10196 129198
rect 9876 122198 9918 122434
rect 10154 122198 10196 122434
rect 9876 115434 10196 122198
rect 9876 115198 9918 115434
rect 10154 115198 10196 115434
rect 9876 108434 10196 115198
rect 9876 108198 9918 108434
rect 10154 108198 10196 108434
rect 9876 101434 10196 108198
rect 9876 101198 9918 101434
rect 10154 101198 10196 101434
rect 9876 94434 10196 101198
rect 9876 94198 9918 94434
rect 10154 94198 10196 94434
rect 9876 87434 10196 94198
rect 9876 87198 9918 87434
rect 10154 87198 10196 87434
rect 9876 80434 10196 87198
rect 9876 80198 9918 80434
rect 10154 80198 10196 80434
rect 9876 73434 10196 80198
rect 9876 73198 9918 73434
rect 10154 73198 10196 73434
rect 9876 66434 10196 73198
rect 9876 66198 9918 66434
rect 10154 66198 10196 66434
rect 9876 59434 10196 66198
rect 9876 59198 9918 59434
rect 10154 59198 10196 59434
rect 9876 52434 10196 59198
rect 9876 52198 9918 52434
rect 10154 52198 10196 52434
rect 9876 45434 10196 52198
rect 9876 45198 9918 45434
rect 10154 45198 10196 45434
rect 9876 38434 10196 45198
rect 9876 38198 9918 38434
rect 10154 38198 10196 38434
rect 9876 31434 10196 38198
rect 9876 31198 9918 31434
rect 10154 31198 10196 31434
rect 9876 24434 10196 31198
rect 9876 24198 9918 24434
rect 10154 24198 10196 24434
rect 9876 17434 10196 24198
rect 9876 17198 9918 17434
rect 10154 17198 10196 17434
rect 9876 10434 10196 17198
rect 9876 10198 9918 10434
rect 10154 10198 10196 10434
rect 9876 3434 10196 10198
rect 9876 3198 9918 3434
rect 10154 3198 10196 3434
rect 9876 -1706 10196 3198
rect 9876 -1942 9918 -1706
rect 10154 -1942 10196 -1706
rect 9876 -2026 10196 -1942
rect 9876 -2262 9918 -2026
rect 10154 -2262 10196 -2026
rect 9876 -2294 10196 -2262
rect 15144 705238 15464 706230
rect 15144 705002 15186 705238
rect 15422 705002 15464 705238
rect 15144 704918 15464 705002
rect 15144 704682 15186 704918
rect 15422 704682 15464 704918
rect 15144 695494 15464 704682
rect 15144 695258 15186 695494
rect 15422 695258 15464 695494
rect 15144 688494 15464 695258
rect 15144 688258 15186 688494
rect 15422 688258 15464 688494
rect 15144 681494 15464 688258
rect 15144 681258 15186 681494
rect 15422 681258 15464 681494
rect 15144 674494 15464 681258
rect 15144 674258 15186 674494
rect 15422 674258 15464 674494
rect 15144 667494 15464 674258
rect 15144 667258 15186 667494
rect 15422 667258 15464 667494
rect 15144 660494 15464 667258
rect 15144 660258 15186 660494
rect 15422 660258 15464 660494
rect 15144 653494 15464 660258
rect 15144 653258 15186 653494
rect 15422 653258 15464 653494
rect 15144 646494 15464 653258
rect 15144 646258 15186 646494
rect 15422 646258 15464 646494
rect 15144 639494 15464 646258
rect 15144 639258 15186 639494
rect 15422 639258 15464 639494
rect 15144 632494 15464 639258
rect 15144 632258 15186 632494
rect 15422 632258 15464 632494
rect 15144 625494 15464 632258
rect 15144 625258 15186 625494
rect 15422 625258 15464 625494
rect 15144 618494 15464 625258
rect 15144 618258 15186 618494
rect 15422 618258 15464 618494
rect 15144 611494 15464 618258
rect 15144 611258 15186 611494
rect 15422 611258 15464 611494
rect 15144 604494 15464 611258
rect 15144 604258 15186 604494
rect 15422 604258 15464 604494
rect 15144 597494 15464 604258
rect 15144 597258 15186 597494
rect 15422 597258 15464 597494
rect 15144 590494 15464 597258
rect 15144 590258 15186 590494
rect 15422 590258 15464 590494
rect 15144 583494 15464 590258
rect 15144 583258 15186 583494
rect 15422 583258 15464 583494
rect 15144 576494 15464 583258
rect 15144 576258 15186 576494
rect 15422 576258 15464 576494
rect 15144 569494 15464 576258
rect 15144 569258 15186 569494
rect 15422 569258 15464 569494
rect 15144 562494 15464 569258
rect 15144 562258 15186 562494
rect 15422 562258 15464 562494
rect 15144 555494 15464 562258
rect 15144 555258 15186 555494
rect 15422 555258 15464 555494
rect 15144 548494 15464 555258
rect 15144 548258 15186 548494
rect 15422 548258 15464 548494
rect 15144 541494 15464 548258
rect 15144 541258 15186 541494
rect 15422 541258 15464 541494
rect 15144 534494 15464 541258
rect 15144 534258 15186 534494
rect 15422 534258 15464 534494
rect 15144 527494 15464 534258
rect 15144 527258 15186 527494
rect 15422 527258 15464 527494
rect 15144 520494 15464 527258
rect 15144 520258 15186 520494
rect 15422 520258 15464 520494
rect 15144 513494 15464 520258
rect 15144 513258 15186 513494
rect 15422 513258 15464 513494
rect 15144 506494 15464 513258
rect 15144 506258 15186 506494
rect 15422 506258 15464 506494
rect 15144 499494 15464 506258
rect 15144 499258 15186 499494
rect 15422 499258 15464 499494
rect 15144 492494 15464 499258
rect 15144 492258 15186 492494
rect 15422 492258 15464 492494
rect 15144 485494 15464 492258
rect 15144 485258 15186 485494
rect 15422 485258 15464 485494
rect 15144 478494 15464 485258
rect 15144 478258 15186 478494
rect 15422 478258 15464 478494
rect 15144 471494 15464 478258
rect 15144 471258 15186 471494
rect 15422 471258 15464 471494
rect 15144 464494 15464 471258
rect 15144 464258 15186 464494
rect 15422 464258 15464 464494
rect 15144 457494 15464 464258
rect 15144 457258 15186 457494
rect 15422 457258 15464 457494
rect 15144 450494 15464 457258
rect 15144 450258 15186 450494
rect 15422 450258 15464 450494
rect 15144 443494 15464 450258
rect 15144 443258 15186 443494
rect 15422 443258 15464 443494
rect 15144 436494 15464 443258
rect 15144 436258 15186 436494
rect 15422 436258 15464 436494
rect 15144 429494 15464 436258
rect 15144 429258 15186 429494
rect 15422 429258 15464 429494
rect 15144 422494 15464 429258
rect 15144 422258 15186 422494
rect 15422 422258 15464 422494
rect 15144 415494 15464 422258
rect 15144 415258 15186 415494
rect 15422 415258 15464 415494
rect 15144 408494 15464 415258
rect 15144 408258 15186 408494
rect 15422 408258 15464 408494
rect 15144 401494 15464 408258
rect 15144 401258 15186 401494
rect 15422 401258 15464 401494
rect 15144 394494 15464 401258
rect 15144 394258 15186 394494
rect 15422 394258 15464 394494
rect 15144 387494 15464 394258
rect 15144 387258 15186 387494
rect 15422 387258 15464 387494
rect 15144 380494 15464 387258
rect 15144 380258 15186 380494
rect 15422 380258 15464 380494
rect 15144 373494 15464 380258
rect 15144 373258 15186 373494
rect 15422 373258 15464 373494
rect 15144 366494 15464 373258
rect 15144 366258 15186 366494
rect 15422 366258 15464 366494
rect 15144 359494 15464 366258
rect 15144 359258 15186 359494
rect 15422 359258 15464 359494
rect 15144 352494 15464 359258
rect 15144 352258 15186 352494
rect 15422 352258 15464 352494
rect 15144 345494 15464 352258
rect 15144 345258 15186 345494
rect 15422 345258 15464 345494
rect 15144 338494 15464 345258
rect 15144 338258 15186 338494
rect 15422 338258 15464 338494
rect 15144 331494 15464 338258
rect 15144 331258 15186 331494
rect 15422 331258 15464 331494
rect 15144 324494 15464 331258
rect 15144 324258 15186 324494
rect 15422 324258 15464 324494
rect 15144 317494 15464 324258
rect 15144 317258 15186 317494
rect 15422 317258 15464 317494
rect 15144 310494 15464 317258
rect 15144 310258 15186 310494
rect 15422 310258 15464 310494
rect 15144 303494 15464 310258
rect 15144 303258 15186 303494
rect 15422 303258 15464 303494
rect 15144 296494 15464 303258
rect 15144 296258 15186 296494
rect 15422 296258 15464 296494
rect 15144 289494 15464 296258
rect 15144 289258 15186 289494
rect 15422 289258 15464 289494
rect 15144 282494 15464 289258
rect 15144 282258 15186 282494
rect 15422 282258 15464 282494
rect 15144 275494 15464 282258
rect 15144 275258 15186 275494
rect 15422 275258 15464 275494
rect 15144 268494 15464 275258
rect 15144 268258 15186 268494
rect 15422 268258 15464 268494
rect 15144 261494 15464 268258
rect 15144 261258 15186 261494
rect 15422 261258 15464 261494
rect 15144 254494 15464 261258
rect 15144 254258 15186 254494
rect 15422 254258 15464 254494
rect 15144 247494 15464 254258
rect 15144 247258 15186 247494
rect 15422 247258 15464 247494
rect 15144 240494 15464 247258
rect 15144 240258 15186 240494
rect 15422 240258 15464 240494
rect 15144 233494 15464 240258
rect 15144 233258 15186 233494
rect 15422 233258 15464 233494
rect 15144 226494 15464 233258
rect 15144 226258 15186 226494
rect 15422 226258 15464 226494
rect 15144 219494 15464 226258
rect 15144 219258 15186 219494
rect 15422 219258 15464 219494
rect 15144 212494 15464 219258
rect 15144 212258 15186 212494
rect 15422 212258 15464 212494
rect 15144 205494 15464 212258
rect 15144 205258 15186 205494
rect 15422 205258 15464 205494
rect 15144 198494 15464 205258
rect 15144 198258 15186 198494
rect 15422 198258 15464 198494
rect 15144 191494 15464 198258
rect 15144 191258 15186 191494
rect 15422 191258 15464 191494
rect 15144 184494 15464 191258
rect 15144 184258 15186 184494
rect 15422 184258 15464 184494
rect 15144 177494 15464 184258
rect 15144 177258 15186 177494
rect 15422 177258 15464 177494
rect 15144 170494 15464 177258
rect 15144 170258 15186 170494
rect 15422 170258 15464 170494
rect 15144 163494 15464 170258
rect 15144 163258 15186 163494
rect 15422 163258 15464 163494
rect 15144 156494 15464 163258
rect 15144 156258 15186 156494
rect 15422 156258 15464 156494
rect 15144 149494 15464 156258
rect 15144 149258 15186 149494
rect 15422 149258 15464 149494
rect 15144 142494 15464 149258
rect 15144 142258 15186 142494
rect 15422 142258 15464 142494
rect 15144 135494 15464 142258
rect 15144 135258 15186 135494
rect 15422 135258 15464 135494
rect 15144 128494 15464 135258
rect 15144 128258 15186 128494
rect 15422 128258 15464 128494
rect 15144 121494 15464 128258
rect 15144 121258 15186 121494
rect 15422 121258 15464 121494
rect 15144 114494 15464 121258
rect 15144 114258 15186 114494
rect 15422 114258 15464 114494
rect 15144 107494 15464 114258
rect 15144 107258 15186 107494
rect 15422 107258 15464 107494
rect 15144 100494 15464 107258
rect 15144 100258 15186 100494
rect 15422 100258 15464 100494
rect 15144 93494 15464 100258
rect 15144 93258 15186 93494
rect 15422 93258 15464 93494
rect 15144 86494 15464 93258
rect 15144 86258 15186 86494
rect 15422 86258 15464 86494
rect 15144 79494 15464 86258
rect 15144 79258 15186 79494
rect 15422 79258 15464 79494
rect 15144 72494 15464 79258
rect 15144 72258 15186 72494
rect 15422 72258 15464 72494
rect 15144 65494 15464 72258
rect 15144 65258 15186 65494
rect 15422 65258 15464 65494
rect 15144 58494 15464 65258
rect 15144 58258 15186 58494
rect 15422 58258 15464 58494
rect 15144 51494 15464 58258
rect 15144 51258 15186 51494
rect 15422 51258 15464 51494
rect 15144 44494 15464 51258
rect 15144 44258 15186 44494
rect 15422 44258 15464 44494
rect 15144 37494 15464 44258
rect 15144 37258 15186 37494
rect 15422 37258 15464 37494
rect 15144 30494 15464 37258
rect 15144 30258 15186 30494
rect 15422 30258 15464 30494
rect 15144 23494 15464 30258
rect 15144 23258 15186 23494
rect 15422 23258 15464 23494
rect 15144 16494 15464 23258
rect 15144 16258 15186 16494
rect 15422 16258 15464 16494
rect 15144 9494 15464 16258
rect 15144 9258 15186 9494
rect 15422 9258 15464 9494
rect 15144 2494 15464 9258
rect 15144 2258 15186 2494
rect 15422 2258 15464 2494
rect 15144 -746 15464 2258
rect 15144 -982 15186 -746
rect 15422 -982 15464 -746
rect 15144 -1066 15464 -982
rect 15144 -1302 15186 -1066
rect 15422 -1302 15464 -1066
rect 15144 -2294 15464 -1302
rect 16876 706198 17196 706230
rect 16876 705962 16918 706198
rect 17154 705962 17196 706198
rect 16876 705878 17196 705962
rect 16876 705642 16918 705878
rect 17154 705642 17196 705878
rect 16876 696434 17196 705642
rect 16876 696198 16918 696434
rect 17154 696198 17196 696434
rect 16876 689434 17196 696198
rect 16876 689198 16918 689434
rect 17154 689198 17196 689434
rect 16876 682434 17196 689198
rect 16876 682198 16918 682434
rect 17154 682198 17196 682434
rect 16876 675434 17196 682198
rect 16876 675198 16918 675434
rect 17154 675198 17196 675434
rect 16876 668434 17196 675198
rect 16876 668198 16918 668434
rect 17154 668198 17196 668434
rect 16876 661434 17196 668198
rect 16876 661198 16918 661434
rect 17154 661198 17196 661434
rect 16876 654434 17196 661198
rect 16876 654198 16918 654434
rect 17154 654198 17196 654434
rect 16876 647434 17196 654198
rect 16876 647198 16918 647434
rect 17154 647198 17196 647434
rect 16876 640434 17196 647198
rect 16876 640198 16918 640434
rect 17154 640198 17196 640434
rect 16876 633434 17196 640198
rect 16876 633198 16918 633434
rect 17154 633198 17196 633434
rect 16876 626434 17196 633198
rect 16876 626198 16918 626434
rect 17154 626198 17196 626434
rect 16876 619434 17196 626198
rect 16876 619198 16918 619434
rect 17154 619198 17196 619434
rect 16876 612434 17196 619198
rect 16876 612198 16918 612434
rect 17154 612198 17196 612434
rect 16876 605434 17196 612198
rect 16876 605198 16918 605434
rect 17154 605198 17196 605434
rect 16876 598434 17196 605198
rect 16876 598198 16918 598434
rect 17154 598198 17196 598434
rect 16876 591434 17196 598198
rect 16876 591198 16918 591434
rect 17154 591198 17196 591434
rect 16876 584434 17196 591198
rect 16876 584198 16918 584434
rect 17154 584198 17196 584434
rect 16876 577434 17196 584198
rect 16876 577198 16918 577434
rect 17154 577198 17196 577434
rect 16876 570434 17196 577198
rect 16876 570198 16918 570434
rect 17154 570198 17196 570434
rect 16876 563434 17196 570198
rect 16876 563198 16918 563434
rect 17154 563198 17196 563434
rect 16876 556434 17196 563198
rect 16876 556198 16918 556434
rect 17154 556198 17196 556434
rect 16876 549434 17196 556198
rect 16876 549198 16918 549434
rect 17154 549198 17196 549434
rect 16876 542434 17196 549198
rect 16876 542198 16918 542434
rect 17154 542198 17196 542434
rect 16876 535434 17196 542198
rect 16876 535198 16918 535434
rect 17154 535198 17196 535434
rect 16876 528434 17196 535198
rect 16876 528198 16918 528434
rect 17154 528198 17196 528434
rect 16876 521434 17196 528198
rect 16876 521198 16918 521434
rect 17154 521198 17196 521434
rect 16876 514434 17196 521198
rect 16876 514198 16918 514434
rect 17154 514198 17196 514434
rect 16876 507434 17196 514198
rect 16876 507198 16918 507434
rect 17154 507198 17196 507434
rect 16876 500434 17196 507198
rect 16876 500198 16918 500434
rect 17154 500198 17196 500434
rect 16876 493434 17196 500198
rect 16876 493198 16918 493434
rect 17154 493198 17196 493434
rect 16876 486434 17196 493198
rect 16876 486198 16918 486434
rect 17154 486198 17196 486434
rect 16876 479434 17196 486198
rect 16876 479198 16918 479434
rect 17154 479198 17196 479434
rect 16876 472434 17196 479198
rect 16876 472198 16918 472434
rect 17154 472198 17196 472434
rect 16876 465434 17196 472198
rect 16876 465198 16918 465434
rect 17154 465198 17196 465434
rect 16876 458434 17196 465198
rect 16876 458198 16918 458434
rect 17154 458198 17196 458434
rect 16876 451434 17196 458198
rect 16876 451198 16918 451434
rect 17154 451198 17196 451434
rect 16876 444434 17196 451198
rect 16876 444198 16918 444434
rect 17154 444198 17196 444434
rect 16876 437434 17196 444198
rect 16876 437198 16918 437434
rect 17154 437198 17196 437434
rect 16876 430434 17196 437198
rect 16876 430198 16918 430434
rect 17154 430198 17196 430434
rect 16876 423434 17196 430198
rect 16876 423198 16918 423434
rect 17154 423198 17196 423434
rect 16876 416434 17196 423198
rect 16876 416198 16918 416434
rect 17154 416198 17196 416434
rect 16876 409434 17196 416198
rect 16876 409198 16918 409434
rect 17154 409198 17196 409434
rect 16876 402434 17196 409198
rect 16876 402198 16918 402434
rect 17154 402198 17196 402434
rect 16876 395434 17196 402198
rect 16876 395198 16918 395434
rect 17154 395198 17196 395434
rect 16876 388434 17196 395198
rect 16876 388198 16918 388434
rect 17154 388198 17196 388434
rect 16876 381434 17196 388198
rect 16876 381198 16918 381434
rect 17154 381198 17196 381434
rect 16876 374434 17196 381198
rect 16876 374198 16918 374434
rect 17154 374198 17196 374434
rect 16876 367434 17196 374198
rect 16876 367198 16918 367434
rect 17154 367198 17196 367434
rect 16876 360434 17196 367198
rect 16876 360198 16918 360434
rect 17154 360198 17196 360434
rect 16876 353434 17196 360198
rect 16876 353198 16918 353434
rect 17154 353198 17196 353434
rect 16876 346434 17196 353198
rect 16876 346198 16918 346434
rect 17154 346198 17196 346434
rect 16876 339434 17196 346198
rect 16876 339198 16918 339434
rect 17154 339198 17196 339434
rect 16876 332434 17196 339198
rect 16876 332198 16918 332434
rect 17154 332198 17196 332434
rect 16876 325434 17196 332198
rect 16876 325198 16918 325434
rect 17154 325198 17196 325434
rect 16876 318434 17196 325198
rect 16876 318198 16918 318434
rect 17154 318198 17196 318434
rect 16876 311434 17196 318198
rect 16876 311198 16918 311434
rect 17154 311198 17196 311434
rect 16876 304434 17196 311198
rect 16876 304198 16918 304434
rect 17154 304198 17196 304434
rect 16876 297434 17196 304198
rect 16876 297198 16918 297434
rect 17154 297198 17196 297434
rect 16876 290434 17196 297198
rect 16876 290198 16918 290434
rect 17154 290198 17196 290434
rect 16876 283434 17196 290198
rect 16876 283198 16918 283434
rect 17154 283198 17196 283434
rect 16876 276434 17196 283198
rect 16876 276198 16918 276434
rect 17154 276198 17196 276434
rect 16876 269434 17196 276198
rect 16876 269198 16918 269434
rect 17154 269198 17196 269434
rect 16876 262434 17196 269198
rect 16876 262198 16918 262434
rect 17154 262198 17196 262434
rect 16876 255434 17196 262198
rect 16876 255198 16918 255434
rect 17154 255198 17196 255434
rect 16876 248434 17196 255198
rect 16876 248198 16918 248434
rect 17154 248198 17196 248434
rect 16876 241434 17196 248198
rect 16876 241198 16918 241434
rect 17154 241198 17196 241434
rect 16876 234434 17196 241198
rect 16876 234198 16918 234434
rect 17154 234198 17196 234434
rect 16876 227434 17196 234198
rect 16876 227198 16918 227434
rect 17154 227198 17196 227434
rect 16876 220434 17196 227198
rect 16876 220198 16918 220434
rect 17154 220198 17196 220434
rect 16876 213434 17196 220198
rect 16876 213198 16918 213434
rect 17154 213198 17196 213434
rect 16876 206434 17196 213198
rect 16876 206198 16918 206434
rect 17154 206198 17196 206434
rect 16876 199434 17196 206198
rect 16876 199198 16918 199434
rect 17154 199198 17196 199434
rect 16876 192434 17196 199198
rect 16876 192198 16918 192434
rect 17154 192198 17196 192434
rect 16876 185434 17196 192198
rect 16876 185198 16918 185434
rect 17154 185198 17196 185434
rect 16876 178434 17196 185198
rect 16876 178198 16918 178434
rect 17154 178198 17196 178434
rect 16876 171434 17196 178198
rect 16876 171198 16918 171434
rect 17154 171198 17196 171434
rect 16876 164434 17196 171198
rect 16876 164198 16918 164434
rect 17154 164198 17196 164434
rect 16876 157434 17196 164198
rect 16876 157198 16918 157434
rect 17154 157198 17196 157434
rect 16876 150434 17196 157198
rect 16876 150198 16918 150434
rect 17154 150198 17196 150434
rect 16876 143434 17196 150198
rect 16876 143198 16918 143434
rect 17154 143198 17196 143434
rect 16876 136434 17196 143198
rect 16876 136198 16918 136434
rect 17154 136198 17196 136434
rect 16876 129434 17196 136198
rect 16876 129198 16918 129434
rect 17154 129198 17196 129434
rect 16876 122434 17196 129198
rect 16876 122198 16918 122434
rect 17154 122198 17196 122434
rect 16876 115434 17196 122198
rect 16876 115198 16918 115434
rect 17154 115198 17196 115434
rect 16876 108434 17196 115198
rect 16876 108198 16918 108434
rect 17154 108198 17196 108434
rect 16876 101434 17196 108198
rect 16876 101198 16918 101434
rect 17154 101198 17196 101434
rect 16876 94434 17196 101198
rect 16876 94198 16918 94434
rect 17154 94198 17196 94434
rect 16876 87434 17196 94198
rect 16876 87198 16918 87434
rect 17154 87198 17196 87434
rect 16876 80434 17196 87198
rect 16876 80198 16918 80434
rect 17154 80198 17196 80434
rect 16876 73434 17196 80198
rect 16876 73198 16918 73434
rect 17154 73198 17196 73434
rect 16876 66434 17196 73198
rect 16876 66198 16918 66434
rect 17154 66198 17196 66434
rect 16876 59434 17196 66198
rect 16876 59198 16918 59434
rect 17154 59198 17196 59434
rect 16876 52434 17196 59198
rect 16876 52198 16918 52434
rect 17154 52198 17196 52434
rect 16876 45434 17196 52198
rect 16876 45198 16918 45434
rect 17154 45198 17196 45434
rect 16876 38434 17196 45198
rect 16876 38198 16918 38434
rect 17154 38198 17196 38434
rect 16876 31434 17196 38198
rect 16876 31198 16918 31434
rect 17154 31198 17196 31434
rect 16876 24434 17196 31198
rect 16876 24198 16918 24434
rect 17154 24198 17196 24434
rect 16876 17434 17196 24198
rect 16876 17198 16918 17434
rect 17154 17198 17196 17434
rect 16876 10434 17196 17198
rect 16876 10198 16918 10434
rect 17154 10198 17196 10434
rect 16876 3434 17196 10198
rect 16876 3198 16918 3434
rect 17154 3198 17196 3434
rect 16876 -1706 17196 3198
rect 16876 -1942 16918 -1706
rect 17154 -1942 17196 -1706
rect 16876 -2026 17196 -1942
rect 16876 -2262 16918 -2026
rect 17154 -2262 17196 -2026
rect 16876 -2294 17196 -2262
rect 22144 705238 22464 706230
rect 22144 705002 22186 705238
rect 22422 705002 22464 705238
rect 22144 704918 22464 705002
rect 22144 704682 22186 704918
rect 22422 704682 22464 704918
rect 22144 695494 22464 704682
rect 22144 695258 22186 695494
rect 22422 695258 22464 695494
rect 22144 688494 22464 695258
rect 22144 688258 22186 688494
rect 22422 688258 22464 688494
rect 22144 681494 22464 688258
rect 22144 681258 22186 681494
rect 22422 681258 22464 681494
rect 22144 674494 22464 681258
rect 22144 674258 22186 674494
rect 22422 674258 22464 674494
rect 22144 667494 22464 674258
rect 22144 667258 22186 667494
rect 22422 667258 22464 667494
rect 22144 660494 22464 667258
rect 22144 660258 22186 660494
rect 22422 660258 22464 660494
rect 22144 653494 22464 660258
rect 22144 653258 22186 653494
rect 22422 653258 22464 653494
rect 22144 646494 22464 653258
rect 22144 646258 22186 646494
rect 22422 646258 22464 646494
rect 22144 639494 22464 646258
rect 22144 639258 22186 639494
rect 22422 639258 22464 639494
rect 22144 632494 22464 639258
rect 22144 632258 22186 632494
rect 22422 632258 22464 632494
rect 22144 625494 22464 632258
rect 22144 625258 22186 625494
rect 22422 625258 22464 625494
rect 22144 618494 22464 625258
rect 22144 618258 22186 618494
rect 22422 618258 22464 618494
rect 22144 611494 22464 618258
rect 22144 611258 22186 611494
rect 22422 611258 22464 611494
rect 22144 604494 22464 611258
rect 22144 604258 22186 604494
rect 22422 604258 22464 604494
rect 22144 597494 22464 604258
rect 22144 597258 22186 597494
rect 22422 597258 22464 597494
rect 22144 590494 22464 597258
rect 22144 590258 22186 590494
rect 22422 590258 22464 590494
rect 22144 583494 22464 590258
rect 22144 583258 22186 583494
rect 22422 583258 22464 583494
rect 22144 576494 22464 583258
rect 22144 576258 22186 576494
rect 22422 576258 22464 576494
rect 22144 569494 22464 576258
rect 22144 569258 22186 569494
rect 22422 569258 22464 569494
rect 22144 562494 22464 569258
rect 22144 562258 22186 562494
rect 22422 562258 22464 562494
rect 22144 555494 22464 562258
rect 22144 555258 22186 555494
rect 22422 555258 22464 555494
rect 22144 548494 22464 555258
rect 22144 548258 22186 548494
rect 22422 548258 22464 548494
rect 22144 541494 22464 548258
rect 22144 541258 22186 541494
rect 22422 541258 22464 541494
rect 22144 534494 22464 541258
rect 22144 534258 22186 534494
rect 22422 534258 22464 534494
rect 22144 527494 22464 534258
rect 22144 527258 22186 527494
rect 22422 527258 22464 527494
rect 22144 520494 22464 527258
rect 22144 520258 22186 520494
rect 22422 520258 22464 520494
rect 22144 513494 22464 520258
rect 22144 513258 22186 513494
rect 22422 513258 22464 513494
rect 22144 506494 22464 513258
rect 22144 506258 22186 506494
rect 22422 506258 22464 506494
rect 22144 499494 22464 506258
rect 22144 499258 22186 499494
rect 22422 499258 22464 499494
rect 22144 492494 22464 499258
rect 22144 492258 22186 492494
rect 22422 492258 22464 492494
rect 22144 485494 22464 492258
rect 22144 485258 22186 485494
rect 22422 485258 22464 485494
rect 22144 478494 22464 485258
rect 22144 478258 22186 478494
rect 22422 478258 22464 478494
rect 22144 471494 22464 478258
rect 22144 471258 22186 471494
rect 22422 471258 22464 471494
rect 22144 464494 22464 471258
rect 22144 464258 22186 464494
rect 22422 464258 22464 464494
rect 22144 457494 22464 464258
rect 22144 457258 22186 457494
rect 22422 457258 22464 457494
rect 22144 450494 22464 457258
rect 22144 450258 22186 450494
rect 22422 450258 22464 450494
rect 22144 443494 22464 450258
rect 22144 443258 22186 443494
rect 22422 443258 22464 443494
rect 22144 436494 22464 443258
rect 22144 436258 22186 436494
rect 22422 436258 22464 436494
rect 22144 429494 22464 436258
rect 22144 429258 22186 429494
rect 22422 429258 22464 429494
rect 22144 422494 22464 429258
rect 22144 422258 22186 422494
rect 22422 422258 22464 422494
rect 22144 415494 22464 422258
rect 22144 415258 22186 415494
rect 22422 415258 22464 415494
rect 22144 408494 22464 415258
rect 22144 408258 22186 408494
rect 22422 408258 22464 408494
rect 22144 401494 22464 408258
rect 22144 401258 22186 401494
rect 22422 401258 22464 401494
rect 22144 394494 22464 401258
rect 22144 394258 22186 394494
rect 22422 394258 22464 394494
rect 22144 387494 22464 394258
rect 22144 387258 22186 387494
rect 22422 387258 22464 387494
rect 22144 380494 22464 387258
rect 22144 380258 22186 380494
rect 22422 380258 22464 380494
rect 22144 373494 22464 380258
rect 22144 373258 22186 373494
rect 22422 373258 22464 373494
rect 22144 366494 22464 373258
rect 22144 366258 22186 366494
rect 22422 366258 22464 366494
rect 22144 359494 22464 366258
rect 22144 359258 22186 359494
rect 22422 359258 22464 359494
rect 22144 352494 22464 359258
rect 22144 352258 22186 352494
rect 22422 352258 22464 352494
rect 22144 345494 22464 352258
rect 22144 345258 22186 345494
rect 22422 345258 22464 345494
rect 22144 338494 22464 345258
rect 22144 338258 22186 338494
rect 22422 338258 22464 338494
rect 22144 331494 22464 338258
rect 22144 331258 22186 331494
rect 22422 331258 22464 331494
rect 22144 324494 22464 331258
rect 22144 324258 22186 324494
rect 22422 324258 22464 324494
rect 22144 317494 22464 324258
rect 22144 317258 22186 317494
rect 22422 317258 22464 317494
rect 22144 310494 22464 317258
rect 22144 310258 22186 310494
rect 22422 310258 22464 310494
rect 22144 303494 22464 310258
rect 22144 303258 22186 303494
rect 22422 303258 22464 303494
rect 22144 296494 22464 303258
rect 22144 296258 22186 296494
rect 22422 296258 22464 296494
rect 22144 289494 22464 296258
rect 22144 289258 22186 289494
rect 22422 289258 22464 289494
rect 22144 282494 22464 289258
rect 22144 282258 22186 282494
rect 22422 282258 22464 282494
rect 22144 275494 22464 282258
rect 22144 275258 22186 275494
rect 22422 275258 22464 275494
rect 22144 268494 22464 275258
rect 22144 268258 22186 268494
rect 22422 268258 22464 268494
rect 22144 261494 22464 268258
rect 22144 261258 22186 261494
rect 22422 261258 22464 261494
rect 22144 254494 22464 261258
rect 22144 254258 22186 254494
rect 22422 254258 22464 254494
rect 22144 247494 22464 254258
rect 22144 247258 22186 247494
rect 22422 247258 22464 247494
rect 22144 240494 22464 247258
rect 22144 240258 22186 240494
rect 22422 240258 22464 240494
rect 22144 233494 22464 240258
rect 22144 233258 22186 233494
rect 22422 233258 22464 233494
rect 22144 226494 22464 233258
rect 22144 226258 22186 226494
rect 22422 226258 22464 226494
rect 22144 219494 22464 226258
rect 22144 219258 22186 219494
rect 22422 219258 22464 219494
rect 22144 212494 22464 219258
rect 22144 212258 22186 212494
rect 22422 212258 22464 212494
rect 22144 205494 22464 212258
rect 22144 205258 22186 205494
rect 22422 205258 22464 205494
rect 22144 198494 22464 205258
rect 22144 198258 22186 198494
rect 22422 198258 22464 198494
rect 22144 191494 22464 198258
rect 22144 191258 22186 191494
rect 22422 191258 22464 191494
rect 22144 184494 22464 191258
rect 22144 184258 22186 184494
rect 22422 184258 22464 184494
rect 22144 177494 22464 184258
rect 22144 177258 22186 177494
rect 22422 177258 22464 177494
rect 22144 170494 22464 177258
rect 22144 170258 22186 170494
rect 22422 170258 22464 170494
rect 22144 163494 22464 170258
rect 22144 163258 22186 163494
rect 22422 163258 22464 163494
rect 22144 156494 22464 163258
rect 22144 156258 22186 156494
rect 22422 156258 22464 156494
rect 22144 149494 22464 156258
rect 22144 149258 22186 149494
rect 22422 149258 22464 149494
rect 22144 142494 22464 149258
rect 22144 142258 22186 142494
rect 22422 142258 22464 142494
rect 22144 135494 22464 142258
rect 22144 135258 22186 135494
rect 22422 135258 22464 135494
rect 22144 128494 22464 135258
rect 22144 128258 22186 128494
rect 22422 128258 22464 128494
rect 22144 121494 22464 128258
rect 22144 121258 22186 121494
rect 22422 121258 22464 121494
rect 22144 114494 22464 121258
rect 22144 114258 22186 114494
rect 22422 114258 22464 114494
rect 22144 107494 22464 114258
rect 22144 107258 22186 107494
rect 22422 107258 22464 107494
rect 22144 100494 22464 107258
rect 22144 100258 22186 100494
rect 22422 100258 22464 100494
rect 22144 93494 22464 100258
rect 22144 93258 22186 93494
rect 22422 93258 22464 93494
rect 22144 86494 22464 93258
rect 22144 86258 22186 86494
rect 22422 86258 22464 86494
rect 22144 79494 22464 86258
rect 22144 79258 22186 79494
rect 22422 79258 22464 79494
rect 22144 72494 22464 79258
rect 22144 72258 22186 72494
rect 22422 72258 22464 72494
rect 22144 65494 22464 72258
rect 22144 65258 22186 65494
rect 22422 65258 22464 65494
rect 22144 58494 22464 65258
rect 22144 58258 22186 58494
rect 22422 58258 22464 58494
rect 22144 51494 22464 58258
rect 22144 51258 22186 51494
rect 22422 51258 22464 51494
rect 22144 44494 22464 51258
rect 22144 44258 22186 44494
rect 22422 44258 22464 44494
rect 22144 37494 22464 44258
rect 22144 37258 22186 37494
rect 22422 37258 22464 37494
rect 22144 30494 22464 37258
rect 22144 30258 22186 30494
rect 22422 30258 22464 30494
rect 22144 23494 22464 30258
rect 22144 23258 22186 23494
rect 22422 23258 22464 23494
rect 22144 16494 22464 23258
rect 22144 16258 22186 16494
rect 22422 16258 22464 16494
rect 22144 9494 22464 16258
rect 22144 9258 22186 9494
rect 22422 9258 22464 9494
rect 22144 2494 22464 9258
rect 22144 2258 22186 2494
rect 22422 2258 22464 2494
rect 22144 -746 22464 2258
rect 22144 -982 22186 -746
rect 22422 -982 22464 -746
rect 22144 -1066 22464 -982
rect 22144 -1302 22186 -1066
rect 22422 -1302 22464 -1066
rect 22144 -2294 22464 -1302
rect 23876 706198 24196 706230
rect 23876 705962 23918 706198
rect 24154 705962 24196 706198
rect 23876 705878 24196 705962
rect 23876 705642 23918 705878
rect 24154 705642 24196 705878
rect 23876 696434 24196 705642
rect 23876 696198 23918 696434
rect 24154 696198 24196 696434
rect 23876 689434 24196 696198
rect 23876 689198 23918 689434
rect 24154 689198 24196 689434
rect 23876 682434 24196 689198
rect 23876 682198 23918 682434
rect 24154 682198 24196 682434
rect 23876 675434 24196 682198
rect 23876 675198 23918 675434
rect 24154 675198 24196 675434
rect 23876 668434 24196 675198
rect 23876 668198 23918 668434
rect 24154 668198 24196 668434
rect 23876 661434 24196 668198
rect 23876 661198 23918 661434
rect 24154 661198 24196 661434
rect 23876 654434 24196 661198
rect 23876 654198 23918 654434
rect 24154 654198 24196 654434
rect 23876 647434 24196 654198
rect 23876 647198 23918 647434
rect 24154 647198 24196 647434
rect 23876 640434 24196 647198
rect 23876 640198 23918 640434
rect 24154 640198 24196 640434
rect 23876 633434 24196 640198
rect 23876 633198 23918 633434
rect 24154 633198 24196 633434
rect 23876 626434 24196 633198
rect 23876 626198 23918 626434
rect 24154 626198 24196 626434
rect 23876 619434 24196 626198
rect 23876 619198 23918 619434
rect 24154 619198 24196 619434
rect 23876 612434 24196 619198
rect 23876 612198 23918 612434
rect 24154 612198 24196 612434
rect 23876 605434 24196 612198
rect 23876 605198 23918 605434
rect 24154 605198 24196 605434
rect 23876 598434 24196 605198
rect 23876 598198 23918 598434
rect 24154 598198 24196 598434
rect 23876 591434 24196 598198
rect 23876 591198 23918 591434
rect 24154 591198 24196 591434
rect 23876 584434 24196 591198
rect 23876 584198 23918 584434
rect 24154 584198 24196 584434
rect 23876 577434 24196 584198
rect 23876 577198 23918 577434
rect 24154 577198 24196 577434
rect 23876 570434 24196 577198
rect 23876 570198 23918 570434
rect 24154 570198 24196 570434
rect 23876 563434 24196 570198
rect 23876 563198 23918 563434
rect 24154 563198 24196 563434
rect 23876 556434 24196 563198
rect 23876 556198 23918 556434
rect 24154 556198 24196 556434
rect 23876 549434 24196 556198
rect 23876 549198 23918 549434
rect 24154 549198 24196 549434
rect 23876 542434 24196 549198
rect 23876 542198 23918 542434
rect 24154 542198 24196 542434
rect 23876 535434 24196 542198
rect 23876 535198 23918 535434
rect 24154 535198 24196 535434
rect 23876 528434 24196 535198
rect 23876 528198 23918 528434
rect 24154 528198 24196 528434
rect 23876 521434 24196 528198
rect 23876 521198 23918 521434
rect 24154 521198 24196 521434
rect 23876 514434 24196 521198
rect 23876 514198 23918 514434
rect 24154 514198 24196 514434
rect 23876 507434 24196 514198
rect 23876 507198 23918 507434
rect 24154 507198 24196 507434
rect 23876 500434 24196 507198
rect 23876 500198 23918 500434
rect 24154 500198 24196 500434
rect 23876 493434 24196 500198
rect 23876 493198 23918 493434
rect 24154 493198 24196 493434
rect 23876 486434 24196 493198
rect 23876 486198 23918 486434
rect 24154 486198 24196 486434
rect 23876 479434 24196 486198
rect 23876 479198 23918 479434
rect 24154 479198 24196 479434
rect 23876 472434 24196 479198
rect 23876 472198 23918 472434
rect 24154 472198 24196 472434
rect 23876 465434 24196 472198
rect 23876 465198 23918 465434
rect 24154 465198 24196 465434
rect 23876 458434 24196 465198
rect 23876 458198 23918 458434
rect 24154 458198 24196 458434
rect 23876 451434 24196 458198
rect 23876 451198 23918 451434
rect 24154 451198 24196 451434
rect 23876 444434 24196 451198
rect 23876 444198 23918 444434
rect 24154 444198 24196 444434
rect 23876 437434 24196 444198
rect 23876 437198 23918 437434
rect 24154 437198 24196 437434
rect 23876 430434 24196 437198
rect 23876 430198 23918 430434
rect 24154 430198 24196 430434
rect 23876 423434 24196 430198
rect 23876 423198 23918 423434
rect 24154 423198 24196 423434
rect 23876 416434 24196 423198
rect 23876 416198 23918 416434
rect 24154 416198 24196 416434
rect 23876 409434 24196 416198
rect 23876 409198 23918 409434
rect 24154 409198 24196 409434
rect 23876 402434 24196 409198
rect 23876 402198 23918 402434
rect 24154 402198 24196 402434
rect 23876 395434 24196 402198
rect 23876 395198 23918 395434
rect 24154 395198 24196 395434
rect 23876 388434 24196 395198
rect 23876 388198 23918 388434
rect 24154 388198 24196 388434
rect 23876 381434 24196 388198
rect 23876 381198 23918 381434
rect 24154 381198 24196 381434
rect 23876 374434 24196 381198
rect 23876 374198 23918 374434
rect 24154 374198 24196 374434
rect 23876 367434 24196 374198
rect 23876 367198 23918 367434
rect 24154 367198 24196 367434
rect 23876 360434 24196 367198
rect 23876 360198 23918 360434
rect 24154 360198 24196 360434
rect 23876 353434 24196 360198
rect 23876 353198 23918 353434
rect 24154 353198 24196 353434
rect 23876 346434 24196 353198
rect 23876 346198 23918 346434
rect 24154 346198 24196 346434
rect 23876 339434 24196 346198
rect 23876 339198 23918 339434
rect 24154 339198 24196 339434
rect 23876 332434 24196 339198
rect 23876 332198 23918 332434
rect 24154 332198 24196 332434
rect 23876 325434 24196 332198
rect 23876 325198 23918 325434
rect 24154 325198 24196 325434
rect 23876 318434 24196 325198
rect 23876 318198 23918 318434
rect 24154 318198 24196 318434
rect 23876 311434 24196 318198
rect 23876 311198 23918 311434
rect 24154 311198 24196 311434
rect 23876 304434 24196 311198
rect 23876 304198 23918 304434
rect 24154 304198 24196 304434
rect 23876 297434 24196 304198
rect 23876 297198 23918 297434
rect 24154 297198 24196 297434
rect 23876 290434 24196 297198
rect 23876 290198 23918 290434
rect 24154 290198 24196 290434
rect 23876 283434 24196 290198
rect 23876 283198 23918 283434
rect 24154 283198 24196 283434
rect 23876 276434 24196 283198
rect 23876 276198 23918 276434
rect 24154 276198 24196 276434
rect 23876 269434 24196 276198
rect 23876 269198 23918 269434
rect 24154 269198 24196 269434
rect 23876 262434 24196 269198
rect 23876 262198 23918 262434
rect 24154 262198 24196 262434
rect 23876 255434 24196 262198
rect 23876 255198 23918 255434
rect 24154 255198 24196 255434
rect 23876 248434 24196 255198
rect 23876 248198 23918 248434
rect 24154 248198 24196 248434
rect 23876 241434 24196 248198
rect 23876 241198 23918 241434
rect 24154 241198 24196 241434
rect 23876 234434 24196 241198
rect 23876 234198 23918 234434
rect 24154 234198 24196 234434
rect 23876 227434 24196 234198
rect 23876 227198 23918 227434
rect 24154 227198 24196 227434
rect 23876 220434 24196 227198
rect 23876 220198 23918 220434
rect 24154 220198 24196 220434
rect 23876 213434 24196 220198
rect 23876 213198 23918 213434
rect 24154 213198 24196 213434
rect 23876 206434 24196 213198
rect 23876 206198 23918 206434
rect 24154 206198 24196 206434
rect 23876 199434 24196 206198
rect 23876 199198 23918 199434
rect 24154 199198 24196 199434
rect 23876 192434 24196 199198
rect 23876 192198 23918 192434
rect 24154 192198 24196 192434
rect 23876 185434 24196 192198
rect 23876 185198 23918 185434
rect 24154 185198 24196 185434
rect 23876 178434 24196 185198
rect 23876 178198 23918 178434
rect 24154 178198 24196 178434
rect 23876 171434 24196 178198
rect 23876 171198 23918 171434
rect 24154 171198 24196 171434
rect 23876 164434 24196 171198
rect 23876 164198 23918 164434
rect 24154 164198 24196 164434
rect 23876 157434 24196 164198
rect 23876 157198 23918 157434
rect 24154 157198 24196 157434
rect 23876 150434 24196 157198
rect 23876 150198 23918 150434
rect 24154 150198 24196 150434
rect 23876 143434 24196 150198
rect 23876 143198 23918 143434
rect 24154 143198 24196 143434
rect 23876 136434 24196 143198
rect 23876 136198 23918 136434
rect 24154 136198 24196 136434
rect 23876 129434 24196 136198
rect 23876 129198 23918 129434
rect 24154 129198 24196 129434
rect 23876 122434 24196 129198
rect 23876 122198 23918 122434
rect 24154 122198 24196 122434
rect 23876 115434 24196 122198
rect 23876 115198 23918 115434
rect 24154 115198 24196 115434
rect 23876 108434 24196 115198
rect 23876 108198 23918 108434
rect 24154 108198 24196 108434
rect 23876 101434 24196 108198
rect 23876 101198 23918 101434
rect 24154 101198 24196 101434
rect 23876 94434 24196 101198
rect 23876 94198 23918 94434
rect 24154 94198 24196 94434
rect 23876 87434 24196 94198
rect 23876 87198 23918 87434
rect 24154 87198 24196 87434
rect 23876 80434 24196 87198
rect 23876 80198 23918 80434
rect 24154 80198 24196 80434
rect 23876 73434 24196 80198
rect 23876 73198 23918 73434
rect 24154 73198 24196 73434
rect 23876 66434 24196 73198
rect 23876 66198 23918 66434
rect 24154 66198 24196 66434
rect 23876 59434 24196 66198
rect 23876 59198 23918 59434
rect 24154 59198 24196 59434
rect 23876 52434 24196 59198
rect 23876 52198 23918 52434
rect 24154 52198 24196 52434
rect 23876 45434 24196 52198
rect 23876 45198 23918 45434
rect 24154 45198 24196 45434
rect 23876 38434 24196 45198
rect 23876 38198 23918 38434
rect 24154 38198 24196 38434
rect 23876 31434 24196 38198
rect 23876 31198 23918 31434
rect 24154 31198 24196 31434
rect 23876 24434 24196 31198
rect 23876 24198 23918 24434
rect 24154 24198 24196 24434
rect 23876 17434 24196 24198
rect 23876 17198 23918 17434
rect 24154 17198 24196 17434
rect 23876 10434 24196 17198
rect 23876 10198 23918 10434
rect 24154 10198 24196 10434
rect 23876 3434 24196 10198
rect 23876 3198 23918 3434
rect 24154 3198 24196 3434
rect 23876 -1706 24196 3198
rect 23876 -1942 23918 -1706
rect 24154 -1942 24196 -1706
rect 23876 -2026 24196 -1942
rect 23876 -2262 23918 -2026
rect 24154 -2262 24196 -2026
rect 23876 -2294 24196 -2262
rect 29144 705238 29464 706230
rect 29144 705002 29186 705238
rect 29422 705002 29464 705238
rect 29144 704918 29464 705002
rect 29144 704682 29186 704918
rect 29422 704682 29464 704918
rect 29144 695494 29464 704682
rect 29144 695258 29186 695494
rect 29422 695258 29464 695494
rect 29144 688494 29464 695258
rect 29144 688258 29186 688494
rect 29422 688258 29464 688494
rect 29144 681494 29464 688258
rect 29144 681258 29186 681494
rect 29422 681258 29464 681494
rect 29144 674494 29464 681258
rect 29144 674258 29186 674494
rect 29422 674258 29464 674494
rect 29144 667494 29464 674258
rect 29144 667258 29186 667494
rect 29422 667258 29464 667494
rect 29144 660494 29464 667258
rect 29144 660258 29186 660494
rect 29422 660258 29464 660494
rect 29144 653494 29464 660258
rect 29144 653258 29186 653494
rect 29422 653258 29464 653494
rect 29144 646494 29464 653258
rect 29144 646258 29186 646494
rect 29422 646258 29464 646494
rect 29144 639494 29464 646258
rect 29144 639258 29186 639494
rect 29422 639258 29464 639494
rect 29144 632494 29464 639258
rect 29144 632258 29186 632494
rect 29422 632258 29464 632494
rect 29144 625494 29464 632258
rect 29144 625258 29186 625494
rect 29422 625258 29464 625494
rect 29144 618494 29464 625258
rect 29144 618258 29186 618494
rect 29422 618258 29464 618494
rect 29144 611494 29464 618258
rect 29144 611258 29186 611494
rect 29422 611258 29464 611494
rect 29144 604494 29464 611258
rect 29144 604258 29186 604494
rect 29422 604258 29464 604494
rect 29144 597494 29464 604258
rect 29144 597258 29186 597494
rect 29422 597258 29464 597494
rect 29144 590494 29464 597258
rect 29144 590258 29186 590494
rect 29422 590258 29464 590494
rect 29144 583494 29464 590258
rect 29144 583258 29186 583494
rect 29422 583258 29464 583494
rect 29144 576494 29464 583258
rect 29144 576258 29186 576494
rect 29422 576258 29464 576494
rect 29144 569494 29464 576258
rect 29144 569258 29186 569494
rect 29422 569258 29464 569494
rect 29144 562494 29464 569258
rect 29144 562258 29186 562494
rect 29422 562258 29464 562494
rect 29144 555494 29464 562258
rect 29144 555258 29186 555494
rect 29422 555258 29464 555494
rect 29144 548494 29464 555258
rect 29144 548258 29186 548494
rect 29422 548258 29464 548494
rect 29144 541494 29464 548258
rect 29144 541258 29186 541494
rect 29422 541258 29464 541494
rect 29144 534494 29464 541258
rect 29144 534258 29186 534494
rect 29422 534258 29464 534494
rect 29144 527494 29464 534258
rect 29144 527258 29186 527494
rect 29422 527258 29464 527494
rect 29144 520494 29464 527258
rect 29144 520258 29186 520494
rect 29422 520258 29464 520494
rect 29144 513494 29464 520258
rect 29144 513258 29186 513494
rect 29422 513258 29464 513494
rect 29144 506494 29464 513258
rect 29144 506258 29186 506494
rect 29422 506258 29464 506494
rect 29144 499494 29464 506258
rect 29144 499258 29186 499494
rect 29422 499258 29464 499494
rect 29144 492494 29464 499258
rect 29144 492258 29186 492494
rect 29422 492258 29464 492494
rect 29144 485494 29464 492258
rect 29144 485258 29186 485494
rect 29422 485258 29464 485494
rect 29144 478494 29464 485258
rect 29144 478258 29186 478494
rect 29422 478258 29464 478494
rect 29144 471494 29464 478258
rect 29144 471258 29186 471494
rect 29422 471258 29464 471494
rect 29144 464494 29464 471258
rect 29144 464258 29186 464494
rect 29422 464258 29464 464494
rect 29144 457494 29464 464258
rect 29144 457258 29186 457494
rect 29422 457258 29464 457494
rect 29144 450494 29464 457258
rect 29144 450258 29186 450494
rect 29422 450258 29464 450494
rect 29144 443494 29464 450258
rect 29144 443258 29186 443494
rect 29422 443258 29464 443494
rect 29144 436494 29464 443258
rect 29144 436258 29186 436494
rect 29422 436258 29464 436494
rect 29144 429494 29464 436258
rect 29144 429258 29186 429494
rect 29422 429258 29464 429494
rect 29144 422494 29464 429258
rect 29144 422258 29186 422494
rect 29422 422258 29464 422494
rect 29144 415494 29464 422258
rect 29144 415258 29186 415494
rect 29422 415258 29464 415494
rect 29144 408494 29464 415258
rect 29144 408258 29186 408494
rect 29422 408258 29464 408494
rect 29144 401494 29464 408258
rect 29144 401258 29186 401494
rect 29422 401258 29464 401494
rect 29144 394494 29464 401258
rect 29144 394258 29186 394494
rect 29422 394258 29464 394494
rect 29144 387494 29464 394258
rect 29144 387258 29186 387494
rect 29422 387258 29464 387494
rect 29144 380494 29464 387258
rect 29144 380258 29186 380494
rect 29422 380258 29464 380494
rect 29144 373494 29464 380258
rect 29144 373258 29186 373494
rect 29422 373258 29464 373494
rect 29144 366494 29464 373258
rect 29144 366258 29186 366494
rect 29422 366258 29464 366494
rect 29144 359494 29464 366258
rect 29144 359258 29186 359494
rect 29422 359258 29464 359494
rect 29144 352494 29464 359258
rect 29144 352258 29186 352494
rect 29422 352258 29464 352494
rect 29144 345494 29464 352258
rect 29144 345258 29186 345494
rect 29422 345258 29464 345494
rect 29144 338494 29464 345258
rect 29144 338258 29186 338494
rect 29422 338258 29464 338494
rect 29144 331494 29464 338258
rect 29144 331258 29186 331494
rect 29422 331258 29464 331494
rect 29144 324494 29464 331258
rect 29144 324258 29186 324494
rect 29422 324258 29464 324494
rect 29144 317494 29464 324258
rect 29144 317258 29186 317494
rect 29422 317258 29464 317494
rect 29144 310494 29464 317258
rect 29144 310258 29186 310494
rect 29422 310258 29464 310494
rect 29144 303494 29464 310258
rect 29144 303258 29186 303494
rect 29422 303258 29464 303494
rect 29144 296494 29464 303258
rect 29144 296258 29186 296494
rect 29422 296258 29464 296494
rect 29144 289494 29464 296258
rect 29144 289258 29186 289494
rect 29422 289258 29464 289494
rect 29144 282494 29464 289258
rect 29144 282258 29186 282494
rect 29422 282258 29464 282494
rect 29144 275494 29464 282258
rect 29144 275258 29186 275494
rect 29422 275258 29464 275494
rect 29144 268494 29464 275258
rect 29144 268258 29186 268494
rect 29422 268258 29464 268494
rect 29144 261494 29464 268258
rect 29144 261258 29186 261494
rect 29422 261258 29464 261494
rect 29144 254494 29464 261258
rect 29144 254258 29186 254494
rect 29422 254258 29464 254494
rect 29144 247494 29464 254258
rect 29144 247258 29186 247494
rect 29422 247258 29464 247494
rect 29144 240494 29464 247258
rect 29144 240258 29186 240494
rect 29422 240258 29464 240494
rect 29144 233494 29464 240258
rect 29144 233258 29186 233494
rect 29422 233258 29464 233494
rect 29144 226494 29464 233258
rect 29144 226258 29186 226494
rect 29422 226258 29464 226494
rect 29144 219494 29464 226258
rect 29144 219258 29186 219494
rect 29422 219258 29464 219494
rect 29144 212494 29464 219258
rect 29144 212258 29186 212494
rect 29422 212258 29464 212494
rect 29144 205494 29464 212258
rect 29144 205258 29186 205494
rect 29422 205258 29464 205494
rect 29144 198494 29464 205258
rect 29144 198258 29186 198494
rect 29422 198258 29464 198494
rect 29144 191494 29464 198258
rect 29144 191258 29186 191494
rect 29422 191258 29464 191494
rect 29144 184494 29464 191258
rect 29144 184258 29186 184494
rect 29422 184258 29464 184494
rect 29144 177494 29464 184258
rect 29144 177258 29186 177494
rect 29422 177258 29464 177494
rect 29144 170494 29464 177258
rect 29144 170258 29186 170494
rect 29422 170258 29464 170494
rect 29144 163494 29464 170258
rect 29144 163258 29186 163494
rect 29422 163258 29464 163494
rect 29144 156494 29464 163258
rect 29144 156258 29186 156494
rect 29422 156258 29464 156494
rect 29144 149494 29464 156258
rect 29144 149258 29186 149494
rect 29422 149258 29464 149494
rect 29144 142494 29464 149258
rect 29144 142258 29186 142494
rect 29422 142258 29464 142494
rect 29144 135494 29464 142258
rect 29144 135258 29186 135494
rect 29422 135258 29464 135494
rect 29144 128494 29464 135258
rect 29144 128258 29186 128494
rect 29422 128258 29464 128494
rect 29144 121494 29464 128258
rect 29144 121258 29186 121494
rect 29422 121258 29464 121494
rect 29144 114494 29464 121258
rect 29144 114258 29186 114494
rect 29422 114258 29464 114494
rect 29144 107494 29464 114258
rect 29144 107258 29186 107494
rect 29422 107258 29464 107494
rect 29144 100494 29464 107258
rect 29144 100258 29186 100494
rect 29422 100258 29464 100494
rect 29144 93494 29464 100258
rect 29144 93258 29186 93494
rect 29422 93258 29464 93494
rect 29144 86494 29464 93258
rect 29144 86258 29186 86494
rect 29422 86258 29464 86494
rect 29144 79494 29464 86258
rect 29144 79258 29186 79494
rect 29422 79258 29464 79494
rect 29144 72494 29464 79258
rect 29144 72258 29186 72494
rect 29422 72258 29464 72494
rect 29144 65494 29464 72258
rect 29144 65258 29186 65494
rect 29422 65258 29464 65494
rect 29144 58494 29464 65258
rect 29144 58258 29186 58494
rect 29422 58258 29464 58494
rect 29144 51494 29464 58258
rect 29144 51258 29186 51494
rect 29422 51258 29464 51494
rect 29144 44494 29464 51258
rect 29144 44258 29186 44494
rect 29422 44258 29464 44494
rect 29144 37494 29464 44258
rect 29144 37258 29186 37494
rect 29422 37258 29464 37494
rect 29144 30494 29464 37258
rect 29144 30258 29186 30494
rect 29422 30258 29464 30494
rect 29144 23494 29464 30258
rect 29144 23258 29186 23494
rect 29422 23258 29464 23494
rect 29144 16494 29464 23258
rect 29144 16258 29186 16494
rect 29422 16258 29464 16494
rect 29144 9494 29464 16258
rect 29144 9258 29186 9494
rect 29422 9258 29464 9494
rect 29144 2494 29464 9258
rect 29144 2258 29186 2494
rect 29422 2258 29464 2494
rect 29144 -746 29464 2258
rect 29144 -982 29186 -746
rect 29422 -982 29464 -746
rect 29144 -1066 29464 -982
rect 29144 -1302 29186 -1066
rect 29422 -1302 29464 -1066
rect 29144 -2294 29464 -1302
rect 30876 706198 31196 706230
rect 30876 705962 30918 706198
rect 31154 705962 31196 706198
rect 30876 705878 31196 705962
rect 30876 705642 30918 705878
rect 31154 705642 31196 705878
rect 30876 696434 31196 705642
rect 30876 696198 30918 696434
rect 31154 696198 31196 696434
rect 30876 689434 31196 696198
rect 30876 689198 30918 689434
rect 31154 689198 31196 689434
rect 30876 682434 31196 689198
rect 30876 682198 30918 682434
rect 31154 682198 31196 682434
rect 30876 675434 31196 682198
rect 30876 675198 30918 675434
rect 31154 675198 31196 675434
rect 30876 668434 31196 675198
rect 30876 668198 30918 668434
rect 31154 668198 31196 668434
rect 30876 661434 31196 668198
rect 30876 661198 30918 661434
rect 31154 661198 31196 661434
rect 30876 654434 31196 661198
rect 30876 654198 30918 654434
rect 31154 654198 31196 654434
rect 30876 647434 31196 654198
rect 30876 647198 30918 647434
rect 31154 647198 31196 647434
rect 30876 640434 31196 647198
rect 30876 640198 30918 640434
rect 31154 640198 31196 640434
rect 30876 633434 31196 640198
rect 30876 633198 30918 633434
rect 31154 633198 31196 633434
rect 30876 626434 31196 633198
rect 30876 626198 30918 626434
rect 31154 626198 31196 626434
rect 30876 619434 31196 626198
rect 30876 619198 30918 619434
rect 31154 619198 31196 619434
rect 30876 612434 31196 619198
rect 30876 612198 30918 612434
rect 31154 612198 31196 612434
rect 30876 605434 31196 612198
rect 30876 605198 30918 605434
rect 31154 605198 31196 605434
rect 30876 598434 31196 605198
rect 30876 598198 30918 598434
rect 31154 598198 31196 598434
rect 30876 591434 31196 598198
rect 30876 591198 30918 591434
rect 31154 591198 31196 591434
rect 30876 584434 31196 591198
rect 30876 584198 30918 584434
rect 31154 584198 31196 584434
rect 30876 577434 31196 584198
rect 30876 577198 30918 577434
rect 31154 577198 31196 577434
rect 30876 570434 31196 577198
rect 30876 570198 30918 570434
rect 31154 570198 31196 570434
rect 30876 563434 31196 570198
rect 30876 563198 30918 563434
rect 31154 563198 31196 563434
rect 30876 556434 31196 563198
rect 30876 556198 30918 556434
rect 31154 556198 31196 556434
rect 30876 549434 31196 556198
rect 30876 549198 30918 549434
rect 31154 549198 31196 549434
rect 30876 542434 31196 549198
rect 30876 542198 30918 542434
rect 31154 542198 31196 542434
rect 30876 535434 31196 542198
rect 30876 535198 30918 535434
rect 31154 535198 31196 535434
rect 30876 528434 31196 535198
rect 30876 528198 30918 528434
rect 31154 528198 31196 528434
rect 30876 521434 31196 528198
rect 30876 521198 30918 521434
rect 31154 521198 31196 521434
rect 30876 514434 31196 521198
rect 30876 514198 30918 514434
rect 31154 514198 31196 514434
rect 30876 507434 31196 514198
rect 30876 507198 30918 507434
rect 31154 507198 31196 507434
rect 30876 500434 31196 507198
rect 30876 500198 30918 500434
rect 31154 500198 31196 500434
rect 30876 493434 31196 500198
rect 30876 493198 30918 493434
rect 31154 493198 31196 493434
rect 30876 486434 31196 493198
rect 30876 486198 30918 486434
rect 31154 486198 31196 486434
rect 30876 479434 31196 486198
rect 30876 479198 30918 479434
rect 31154 479198 31196 479434
rect 30876 472434 31196 479198
rect 30876 472198 30918 472434
rect 31154 472198 31196 472434
rect 30876 465434 31196 472198
rect 30876 465198 30918 465434
rect 31154 465198 31196 465434
rect 30876 458434 31196 465198
rect 30876 458198 30918 458434
rect 31154 458198 31196 458434
rect 30876 451434 31196 458198
rect 30876 451198 30918 451434
rect 31154 451198 31196 451434
rect 30876 444434 31196 451198
rect 30876 444198 30918 444434
rect 31154 444198 31196 444434
rect 30876 437434 31196 444198
rect 30876 437198 30918 437434
rect 31154 437198 31196 437434
rect 30876 430434 31196 437198
rect 30876 430198 30918 430434
rect 31154 430198 31196 430434
rect 30876 423434 31196 430198
rect 30876 423198 30918 423434
rect 31154 423198 31196 423434
rect 30876 416434 31196 423198
rect 30876 416198 30918 416434
rect 31154 416198 31196 416434
rect 30876 409434 31196 416198
rect 30876 409198 30918 409434
rect 31154 409198 31196 409434
rect 30876 402434 31196 409198
rect 30876 402198 30918 402434
rect 31154 402198 31196 402434
rect 30876 395434 31196 402198
rect 30876 395198 30918 395434
rect 31154 395198 31196 395434
rect 30876 388434 31196 395198
rect 30876 388198 30918 388434
rect 31154 388198 31196 388434
rect 30876 381434 31196 388198
rect 30876 381198 30918 381434
rect 31154 381198 31196 381434
rect 30876 374434 31196 381198
rect 30876 374198 30918 374434
rect 31154 374198 31196 374434
rect 30876 367434 31196 374198
rect 30876 367198 30918 367434
rect 31154 367198 31196 367434
rect 30876 360434 31196 367198
rect 30876 360198 30918 360434
rect 31154 360198 31196 360434
rect 30876 353434 31196 360198
rect 30876 353198 30918 353434
rect 31154 353198 31196 353434
rect 30876 346434 31196 353198
rect 30876 346198 30918 346434
rect 31154 346198 31196 346434
rect 30876 339434 31196 346198
rect 30876 339198 30918 339434
rect 31154 339198 31196 339434
rect 30876 332434 31196 339198
rect 30876 332198 30918 332434
rect 31154 332198 31196 332434
rect 30876 325434 31196 332198
rect 30876 325198 30918 325434
rect 31154 325198 31196 325434
rect 30876 318434 31196 325198
rect 30876 318198 30918 318434
rect 31154 318198 31196 318434
rect 30876 311434 31196 318198
rect 30876 311198 30918 311434
rect 31154 311198 31196 311434
rect 30876 304434 31196 311198
rect 30876 304198 30918 304434
rect 31154 304198 31196 304434
rect 30876 297434 31196 304198
rect 30876 297198 30918 297434
rect 31154 297198 31196 297434
rect 30876 290434 31196 297198
rect 30876 290198 30918 290434
rect 31154 290198 31196 290434
rect 30876 283434 31196 290198
rect 30876 283198 30918 283434
rect 31154 283198 31196 283434
rect 30876 276434 31196 283198
rect 30876 276198 30918 276434
rect 31154 276198 31196 276434
rect 30876 269434 31196 276198
rect 30876 269198 30918 269434
rect 31154 269198 31196 269434
rect 30876 262434 31196 269198
rect 30876 262198 30918 262434
rect 31154 262198 31196 262434
rect 30876 255434 31196 262198
rect 30876 255198 30918 255434
rect 31154 255198 31196 255434
rect 30876 248434 31196 255198
rect 30876 248198 30918 248434
rect 31154 248198 31196 248434
rect 30876 241434 31196 248198
rect 30876 241198 30918 241434
rect 31154 241198 31196 241434
rect 30876 234434 31196 241198
rect 30876 234198 30918 234434
rect 31154 234198 31196 234434
rect 30876 227434 31196 234198
rect 30876 227198 30918 227434
rect 31154 227198 31196 227434
rect 30876 220434 31196 227198
rect 30876 220198 30918 220434
rect 31154 220198 31196 220434
rect 30876 213434 31196 220198
rect 30876 213198 30918 213434
rect 31154 213198 31196 213434
rect 30876 206434 31196 213198
rect 30876 206198 30918 206434
rect 31154 206198 31196 206434
rect 30876 199434 31196 206198
rect 30876 199198 30918 199434
rect 31154 199198 31196 199434
rect 30876 192434 31196 199198
rect 30876 192198 30918 192434
rect 31154 192198 31196 192434
rect 30876 185434 31196 192198
rect 30876 185198 30918 185434
rect 31154 185198 31196 185434
rect 30876 178434 31196 185198
rect 30876 178198 30918 178434
rect 31154 178198 31196 178434
rect 30876 171434 31196 178198
rect 30876 171198 30918 171434
rect 31154 171198 31196 171434
rect 30876 164434 31196 171198
rect 30876 164198 30918 164434
rect 31154 164198 31196 164434
rect 30876 157434 31196 164198
rect 30876 157198 30918 157434
rect 31154 157198 31196 157434
rect 30876 150434 31196 157198
rect 30876 150198 30918 150434
rect 31154 150198 31196 150434
rect 30876 143434 31196 150198
rect 30876 143198 30918 143434
rect 31154 143198 31196 143434
rect 30876 136434 31196 143198
rect 30876 136198 30918 136434
rect 31154 136198 31196 136434
rect 30876 129434 31196 136198
rect 30876 129198 30918 129434
rect 31154 129198 31196 129434
rect 30876 122434 31196 129198
rect 30876 122198 30918 122434
rect 31154 122198 31196 122434
rect 30876 115434 31196 122198
rect 30876 115198 30918 115434
rect 31154 115198 31196 115434
rect 30876 108434 31196 115198
rect 30876 108198 30918 108434
rect 31154 108198 31196 108434
rect 30876 101434 31196 108198
rect 30876 101198 30918 101434
rect 31154 101198 31196 101434
rect 30876 94434 31196 101198
rect 30876 94198 30918 94434
rect 31154 94198 31196 94434
rect 30876 87434 31196 94198
rect 30876 87198 30918 87434
rect 31154 87198 31196 87434
rect 30876 80434 31196 87198
rect 30876 80198 30918 80434
rect 31154 80198 31196 80434
rect 30876 73434 31196 80198
rect 30876 73198 30918 73434
rect 31154 73198 31196 73434
rect 30876 66434 31196 73198
rect 30876 66198 30918 66434
rect 31154 66198 31196 66434
rect 30876 59434 31196 66198
rect 30876 59198 30918 59434
rect 31154 59198 31196 59434
rect 30876 52434 31196 59198
rect 30876 52198 30918 52434
rect 31154 52198 31196 52434
rect 30876 45434 31196 52198
rect 30876 45198 30918 45434
rect 31154 45198 31196 45434
rect 30876 38434 31196 45198
rect 30876 38198 30918 38434
rect 31154 38198 31196 38434
rect 30876 31434 31196 38198
rect 30876 31198 30918 31434
rect 31154 31198 31196 31434
rect 30876 24434 31196 31198
rect 30876 24198 30918 24434
rect 31154 24198 31196 24434
rect 30876 17434 31196 24198
rect 30876 17198 30918 17434
rect 31154 17198 31196 17434
rect 30876 10434 31196 17198
rect 30876 10198 30918 10434
rect 31154 10198 31196 10434
rect 30876 3434 31196 10198
rect 30876 3198 30918 3434
rect 31154 3198 31196 3434
rect 30876 -1706 31196 3198
rect 30876 -1942 30918 -1706
rect 31154 -1942 31196 -1706
rect 30876 -2026 31196 -1942
rect 30876 -2262 30918 -2026
rect 31154 -2262 31196 -2026
rect 30876 -2294 31196 -2262
rect 36144 705238 36464 706230
rect 36144 705002 36186 705238
rect 36422 705002 36464 705238
rect 36144 704918 36464 705002
rect 36144 704682 36186 704918
rect 36422 704682 36464 704918
rect 36144 695494 36464 704682
rect 36144 695258 36186 695494
rect 36422 695258 36464 695494
rect 36144 688494 36464 695258
rect 36144 688258 36186 688494
rect 36422 688258 36464 688494
rect 36144 681494 36464 688258
rect 36144 681258 36186 681494
rect 36422 681258 36464 681494
rect 36144 674494 36464 681258
rect 36144 674258 36186 674494
rect 36422 674258 36464 674494
rect 36144 667494 36464 674258
rect 36144 667258 36186 667494
rect 36422 667258 36464 667494
rect 36144 660494 36464 667258
rect 36144 660258 36186 660494
rect 36422 660258 36464 660494
rect 36144 653494 36464 660258
rect 36144 653258 36186 653494
rect 36422 653258 36464 653494
rect 36144 646494 36464 653258
rect 36144 646258 36186 646494
rect 36422 646258 36464 646494
rect 36144 639494 36464 646258
rect 36144 639258 36186 639494
rect 36422 639258 36464 639494
rect 36144 632494 36464 639258
rect 36144 632258 36186 632494
rect 36422 632258 36464 632494
rect 36144 625494 36464 632258
rect 36144 625258 36186 625494
rect 36422 625258 36464 625494
rect 36144 618494 36464 625258
rect 36144 618258 36186 618494
rect 36422 618258 36464 618494
rect 36144 611494 36464 618258
rect 36144 611258 36186 611494
rect 36422 611258 36464 611494
rect 36144 604494 36464 611258
rect 36144 604258 36186 604494
rect 36422 604258 36464 604494
rect 36144 597494 36464 604258
rect 36144 597258 36186 597494
rect 36422 597258 36464 597494
rect 36144 590494 36464 597258
rect 36144 590258 36186 590494
rect 36422 590258 36464 590494
rect 36144 583494 36464 590258
rect 36144 583258 36186 583494
rect 36422 583258 36464 583494
rect 36144 576494 36464 583258
rect 36144 576258 36186 576494
rect 36422 576258 36464 576494
rect 36144 569494 36464 576258
rect 36144 569258 36186 569494
rect 36422 569258 36464 569494
rect 36144 562494 36464 569258
rect 36144 562258 36186 562494
rect 36422 562258 36464 562494
rect 36144 555494 36464 562258
rect 36144 555258 36186 555494
rect 36422 555258 36464 555494
rect 36144 548494 36464 555258
rect 36144 548258 36186 548494
rect 36422 548258 36464 548494
rect 36144 541494 36464 548258
rect 36144 541258 36186 541494
rect 36422 541258 36464 541494
rect 36144 534494 36464 541258
rect 36144 534258 36186 534494
rect 36422 534258 36464 534494
rect 36144 527494 36464 534258
rect 36144 527258 36186 527494
rect 36422 527258 36464 527494
rect 36144 520494 36464 527258
rect 36144 520258 36186 520494
rect 36422 520258 36464 520494
rect 36144 513494 36464 520258
rect 36144 513258 36186 513494
rect 36422 513258 36464 513494
rect 36144 506494 36464 513258
rect 36144 506258 36186 506494
rect 36422 506258 36464 506494
rect 36144 499494 36464 506258
rect 36144 499258 36186 499494
rect 36422 499258 36464 499494
rect 36144 492494 36464 499258
rect 36144 492258 36186 492494
rect 36422 492258 36464 492494
rect 36144 485494 36464 492258
rect 36144 485258 36186 485494
rect 36422 485258 36464 485494
rect 36144 478494 36464 485258
rect 36144 478258 36186 478494
rect 36422 478258 36464 478494
rect 36144 471494 36464 478258
rect 36144 471258 36186 471494
rect 36422 471258 36464 471494
rect 36144 464494 36464 471258
rect 36144 464258 36186 464494
rect 36422 464258 36464 464494
rect 36144 457494 36464 464258
rect 36144 457258 36186 457494
rect 36422 457258 36464 457494
rect 36144 450494 36464 457258
rect 36144 450258 36186 450494
rect 36422 450258 36464 450494
rect 36144 443494 36464 450258
rect 36144 443258 36186 443494
rect 36422 443258 36464 443494
rect 36144 436494 36464 443258
rect 36144 436258 36186 436494
rect 36422 436258 36464 436494
rect 36144 429494 36464 436258
rect 36144 429258 36186 429494
rect 36422 429258 36464 429494
rect 36144 422494 36464 429258
rect 36144 422258 36186 422494
rect 36422 422258 36464 422494
rect 36144 415494 36464 422258
rect 36144 415258 36186 415494
rect 36422 415258 36464 415494
rect 36144 408494 36464 415258
rect 36144 408258 36186 408494
rect 36422 408258 36464 408494
rect 36144 401494 36464 408258
rect 36144 401258 36186 401494
rect 36422 401258 36464 401494
rect 36144 394494 36464 401258
rect 36144 394258 36186 394494
rect 36422 394258 36464 394494
rect 36144 387494 36464 394258
rect 36144 387258 36186 387494
rect 36422 387258 36464 387494
rect 36144 380494 36464 387258
rect 36144 380258 36186 380494
rect 36422 380258 36464 380494
rect 36144 373494 36464 380258
rect 36144 373258 36186 373494
rect 36422 373258 36464 373494
rect 36144 366494 36464 373258
rect 36144 366258 36186 366494
rect 36422 366258 36464 366494
rect 36144 359494 36464 366258
rect 36144 359258 36186 359494
rect 36422 359258 36464 359494
rect 36144 352494 36464 359258
rect 36144 352258 36186 352494
rect 36422 352258 36464 352494
rect 36144 345494 36464 352258
rect 36144 345258 36186 345494
rect 36422 345258 36464 345494
rect 36144 338494 36464 345258
rect 36144 338258 36186 338494
rect 36422 338258 36464 338494
rect 36144 331494 36464 338258
rect 36144 331258 36186 331494
rect 36422 331258 36464 331494
rect 36144 324494 36464 331258
rect 36144 324258 36186 324494
rect 36422 324258 36464 324494
rect 36144 317494 36464 324258
rect 36144 317258 36186 317494
rect 36422 317258 36464 317494
rect 36144 310494 36464 317258
rect 36144 310258 36186 310494
rect 36422 310258 36464 310494
rect 36144 303494 36464 310258
rect 36144 303258 36186 303494
rect 36422 303258 36464 303494
rect 36144 296494 36464 303258
rect 36144 296258 36186 296494
rect 36422 296258 36464 296494
rect 36144 289494 36464 296258
rect 36144 289258 36186 289494
rect 36422 289258 36464 289494
rect 36144 282494 36464 289258
rect 36144 282258 36186 282494
rect 36422 282258 36464 282494
rect 36144 275494 36464 282258
rect 36144 275258 36186 275494
rect 36422 275258 36464 275494
rect 36144 268494 36464 275258
rect 36144 268258 36186 268494
rect 36422 268258 36464 268494
rect 36144 261494 36464 268258
rect 36144 261258 36186 261494
rect 36422 261258 36464 261494
rect 36144 254494 36464 261258
rect 36144 254258 36186 254494
rect 36422 254258 36464 254494
rect 36144 247494 36464 254258
rect 36144 247258 36186 247494
rect 36422 247258 36464 247494
rect 36144 240494 36464 247258
rect 36144 240258 36186 240494
rect 36422 240258 36464 240494
rect 36144 233494 36464 240258
rect 36144 233258 36186 233494
rect 36422 233258 36464 233494
rect 36144 226494 36464 233258
rect 36144 226258 36186 226494
rect 36422 226258 36464 226494
rect 36144 219494 36464 226258
rect 36144 219258 36186 219494
rect 36422 219258 36464 219494
rect 36144 212494 36464 219258
rect 36144 212258 36186 212494
rect 36422 212258 36464 212494
rect 36144 205494 36464 212258
rect 36144 205258 36186 205494
rect 36422 205258 36464 205494
rect 36144 198494 36464 205258
rect 36144 198258 36186 198494
rect 36422 198258 36464 198494
rect 36144 191494 36464 198258
rect 36144 191258 36186 191494
rect 36422 191258 36464 191494
rect 36144 184494 36464 191258
rect 36144 184258 36186 184494
rect 36422 184258 36464 184494
rect 36144 177494 36464 184258
rect 36144 177258 36186 177494
rect 36422 177258 36464 177494
rect 36144 170494 36464 177258
rect 36144 170258 36186 170494
rect 36422 170258 36464 170494
rect 36144 163494 36464 170258
rect 36144 163258 36186 163494
rect 36422 163258 36464 163494
rect 36144 156494 36464 163258
rect 36144 156258 36186 156494
rect 36422 156258 36464 156494
rect 36144 149494 36464 156258
rect 36144 149258 36186 149494
rect 36422 149258 36464 149494
rect 36144 142494 36464 149258
rect 36144 142258 36186 142494
rect 36422 142258 36464 142494
rect 36144 135494 36464 142258
rect 36144 135258 36186 135494
rect 36422 135258 36464 135494
rect 36144 128494 36464 135258
rect 36144 128258 36186 128494
rect 36422 128258 36464 128494
rect 36144 121494 36464 128258
rect 36144 121258 36186 121494
rect 36422 121258 36464 121494
rect 36144 114494 36464 121258
rect 36144 114258 36186 114494
rect 36422 114258 36464 114494
rect 36144 107494 36464 114258
rect 36144 107258 36186 107494
rect 36422 107258 36464 107494
rect 36144 100494 36464 107258
rect 36144 100258 36186 100494
rect 36422 100258 36464 100494
rect 36144 93494 36464 100258
rect 36144 93258 36186 93494
rect 36422 93258 36464 93494
rect 36144 86494 36464 93258
rect 36144 86258 36186 86494
rect 36422 86258 36464 86494
rect 36144 79494 36464 86258
rect 36144 79258 36186 79494
rect 36422 79258 36464 79494
rect 36144 72494 36464 79258
rect 36144 72258 36186 72494
rect 36422 72258 36464 72494
rect 36144 65494 36464 72258
rect 36144 65258 36186 65494
rect 36422 65258 36464 65494
rect 36144 58494 36464 65258
rect 36144 58258 36186 58494
rect 36422 58258 36464 58494
rect 36144 51494 36464 58258
rect 36144 51258 36186 51494
rect 36422 51258 36464 51494
rect 36144 44494 36464 51258
rect 36144 44258 36186 44494
rect 36422 44258 36464 44494
rect 36144 37494 36464 44258
rect 36144 37258 36186 37494
rect 36422 37258 36464 37494
rect 36144 30494 36464 37258
rect 36144 30258 36186 30494
rect 36422 30258 36464 30494
rect 36144 23494 36464 30258
rect 36144 23258 36186 23494
rect 36422 23258 36464 23494
rect 36144 16494 36464 23258
rect 36144 16258 36186 16494
rect 36422 16258 36464 16494
rect 36144 9494 36464 16258
rect 36144 9258 36186 9494
rect 36422 9258 36464 9494
rect 36144 2494 36464 9258
rect 36144 2258 36186 2494
rect 36422 2258 36464 2494
rect 36144 -746 36464 2258
rect 36144 -982 36186 -746
rect 36422 -982 36464 -746
rect 36144 -1066 36464 -982
rect 36144 -1302 36186 -1066
rect 36422 -1302 36464 -1066
rect 36144 -2294 36464 -1302
rect 37876 706198 38196 706230
rect 37876 705962 37918 706198
rect 38154 705962 38196 706198
rect 37876 705878 38196 705962
rect 37876 705642 37918 705878
rect 38154 705642 38196 705878
rect 37876 696434 38196 705642
rect 37876 696198 37918 696434
rect 38154 696198 38196 696434
rect 37876 689434 38196 696198
rect 37876 689198 37918 689434
rect 38154 689198 38196 689434
rect 37876 682434 38196 689198
rect 37876 682198 37918 682434
rect 38154 682198 38196 682434
rect 37876 675434 38196 682198
rect 37876 675198 37918 675434
rect 38154 675198 38196 675434
rect 37876 668434 38196 675198
rect 37876 668198 37918 668434
rect 38154 668198 38196 668434
rect 37876 661434 38196 668198
rect 37876 661198 37918 661434
rect 38154 661198 38196 661434
rect 37876 654434 38196 661198
rect 37876 654198 37918 654434
rect 38154 654198 38196 654434
rect 37876 647434 38196 654198
rect 37876 647198 37918 647434
rect 38154 647198 38196 647434
rect 37876 640434 38196 647198
rect 37876 640198 37918 640434
rect 38154 640198 38196 640434
rect 37876 633434 38196 640198
rect 37876 633198 37918 633434
rect 38154 633198 38196 633434
rect 37876 626434 38196 633198
rect 37876 626198 37918 626434
rect 38154 626198 38196 626434
rect 37876 619434 38196 626198
rect 37876 619198 37918 619434
rect 38154 619198 38196 619434
rect 37876 612434 38196 619198
rect 37876 612198 37918 612434
rect 38154 612198 38196 612434
rect 37876 605434 38196 612198
rect 37876 605198 37918 605434
rect 38154 605198 38196 605434
rect 37876 598434 38196 605198
rect 37876 598198 37918 598434
rect 38154 598198 38196 598434
rect 37876 591434 38196 598198
rect 37876 591198 37918 591434
rect 38154 591198 38196 591434
rect 37876 584434 38196 591198
rect 37876 584198 37918 584434
rect 38154 584198 38196 584434
rect 37876 577434 38196 584198
rect 37876 577198 37918 577434
rect 38154 577198 38196 577434
rect 37876 570434 38196 577198
rect 37876 570198 37918 570434
rect 38154 570198 38196 570434
rect 37876 563434 38196 570198
rect 37876 563198 37918 563434
rect 38154 563198 38196 563434
rect 37876 556434 38196 563198
rect 37876 556198 37918 556434
rect 38154 556198 38196 556434
rect 37876 549434 38196 556198
rect 37876 549198 37918 549434
rect 38154 549198 38196 549434
rect 37876 542434 38196 549198
rect 37876 542198 37918 542434
rect 38154 542198 38196 542434
rect 37876 535434 38196 542198
rect 37876 535198 37918 535434
rect 38154 535198 38196 535434
rect 37876 528434 38196 535198
rect 37876 528198 37918 528434
rect 38154 528198 38196 528434
rect 37876 521434 38196 528198
rect 37876 521198 37918 521434
rect 38154 521198 38196 521434
rect 37876 514434 38196 521198
rect 37876 514198 37918 514434
rect 38154 514198 38196 514434
rect 37876 507434 38196 514198
rect 37876 507198 37918 507434
rect 38154 507198 38196 507434
rect 37876 500434 38196 507198
rect 37876 500198 37918 500434
rect 38154 500198 38196 500434
rect 37876 493434 38196 500198
rect 37876 493198 37918 493434
rect 38154 493198 38196 493434
rect 37876 486434 38196 493198
rect 37876 486198 37918 486434
rect 38154 486198 38196 486434
rect 37876 479434 38196 486198
rect 37876 479198 37918 479434
rect 38154 479198 38196 479434
rect 37876 472434 38196 479198
rect 37876 472198 37918 472434
rect 38154 472198 38196 472434
rect 37876 465434 38196 472198
rect 37876 465198 37918 465434
rect 38154 465198 38196 465434
rect 37876 458434 38196 465198
rect 37876 458198 37918 458434
rect 38154 458198 38196 458434
rect 37876 451434 38196 458198
rect 37876 451198 37918 451434
rect 38154 451198 38196 451434
rect 37876 444434 38196 451198
rect 37876 444198 37918 444434
rect 38154 444198 38196 444434
rect 37876 437434 38196 444198
rect 37876 437198 37918 437434
rect 38154 437198 38196 437434
rect 37876 430434 38196 437198
rect 37876 430198 37918 430434
rect 38154 430198 38196 430434
rect 37876 423434 38196 430198
rect 37876 423198 37918 423434
rect 38154 423198 38196 423434
rect 37876 416434 38196 423198
rect 37876 416198 37918 416434
rect 38154 416198 38196 416434
rect 37876 409434 38196 416198
rect 37876 409198 37918 409434
rect 38154 409198 38196 409434
rect 37876 402434 38196 409198
rect 37876 402198 37918 402434
rect 38154 402198 38196 402434
rect 37876 395434 38196 402198
rect 37876 395198 37918 395434
rect 38154 395198 38196 395434
rect 37876 388434 38196 395198
rect 37876 388198 37918 388434
rect 38154 388198 38196 388434
rect 37876 381434 38196 388198
rect 37876 381198 37918 381434
rect 38154 381198 38196 381434
rect 37876 374434 38196 381198
rect 37876 374198 37918 374434
rect 38154 374198 38196 374434
rect 37876 367434 38196 374198
rect 37876 367198 37918 367434
rect 38154 367198 38196 367434
rect 37876 360434 38196 367198
rect 37876 360198 37918 360434
rect 38154 360198 38196 360434
rect 37876 353434 38196 360198
rect 37876 353198 37918 353434
rect 38154 353198 38196 353434
rect 37876 346434 38196 353198
rect 37876 346198 37918 346434
rect 38154 346198 38196 346434
rect 37876 339434 38196 346198
rect 37876 339198 37918 339434
rect 38154 339198 38196 339434
rect 37876 332434 38196 339198
rect 37876 332198 37918 332434
rect 38154 332198 38196 332434
rect 37876 325434 38196 332198
rect 37876 325198 37918 325434
rect 38154 325198 38196 325434
rect 37876 318434 38196 325198
rect 37876 318198 37918 318434
rect 38154 318198 38196 318434
rect 37876 311434 38196 318198
rect 37876 311198 37918 311434
rect 38154 311198 38196 311434
rect 37876 304434 38196 311198
rect 37876 304198 37918 304434
rect 38154 304198 38196 304434
rect 37876 297434 38196 304198
rect 37876 297198 37918 297434
rect 38154 297198 38196 297434
rect 37876 290434 38196 297198
rect 37876 290198 37918 290434
rect 38154 290198 38196 290434
rect 37876 283434 38196 290198
rect 37876 283198 37918 283434
rect 38154 283198 38196 283434
rect 37876 276434 38196 283198
rect 37876 276198 37918 276434
rect 38154 276198 38196 276434
rect 37876 269434 38196 276198
rect 37876 269198 37918 269434
rect 38154 269198 38196 269434
rect 37876 262434 38196 269198
rect 37876 262198 37918 262434
rect 38154 262198 38196 262434
rect 37876 255434 38196 262198
rect 37876 255198 37918 255434
rect 38154 255198 38196 255434
rect 37876 248434 38196 255198
rect 37876 248198 37918 248434
rect 38154 248198 38196 248434
rect 37876 241434 38196 248198
rect 37876 241198 37918 241434
rect 38154 241198 38196 241434
rect 37876 234434 38196 241198
rect 37876 234198 37918 234434
rect 38154 234198 38196 234434
rect 37876 227434 38196 234198
rect 37876 227198 37918 227434
rect 38154 227198 38196 227434
rect 37876 220434 38196 227198
rect 37876 220198 37918 220434
rect 38154 220198 38196 220434
rect 37876 213434 38196 220198
rect 37876 213198 37918 213434
rect 38154 213198 38196 213434
rect 37876 206434 38196 213198
rect 37876 206198 37918 206434
rect 38154 206198 38196 206434
rect 37876 199434 38196 206198
rect 37876 199198 37918 199434
rect 38154 199198 38196 199434
rect 37876 192434 38196 199198
rect 37876 192198 37918 192434
rect 38154 192198 38196 192434
rect 37876 185434 38196 192198
rect 37876 185198 37918 185434
rect 38154 185198 38196 185434
rect 37876 178434 38196 185198
rect 37876 178198 37918 178434
rect 38154 178198 38196 178434
rect 37876 171434 38196 178198
rect 37876 171198 37918 171434
rect 38154 171198 38196 171434
rect 37876 164434 38196 171198
rect 37876 164198 37918 164434
rect 38154 164198 38196 164434
rect 37876 157434 38196 164198
rect 37876 157198 37918 157434
rect 38154 157198 38196 157434
rect 37876 150434 38196 157198
rect 37876 150198 37918 150434
rect 38154 150198 38196 150434
rect 37876 143434 38196 150198
rect 37876 143198 37918 143434
rect 38154 143198 38196 143434
rect 37876 136434 38196 143198
rect 37876 136198 37918 136434
rect 38154 136198 38196 136434
rect 37876 129434 38196 136198
rect 37876 129198 37918 129434
rect 38154 129198 38196 129434
rect 37876 122434 38196 129198
rect 37876 122198 37918 122434
rect 38154 122198 38196 122434
rect 37876 115434 38196 122198
rect 37876 115198 37918 115434
rect 38154 115198 38196 115434
rect 37876 108434 38196 115198
rect 37876 108198 37918 108434
rect 38154 108198 38196 108434
rect 37876 101434 38196 108198
rect 37876 101198 37918 101434
rect 38154 101198 38196 101434
rect 37876 94434 38196 101198
rect 37876 94198 37918 94434
rect 38154 94198 38196 94434
rect 37876 87434 38196 94198
rect 37876 87198 37918 87434
rect 38154 87198 38196 87434
rect 37876 80434 38196 87198
rect 37876 80198 37918 80434
rect 38154 80198 38196 80434
rect 37876 73434 38196 80198
rect 37876 73198 37918 73434
rect 38154 73198 38196 73434
rect 37876 66434 38196 73198
rect 37876 66198 37918 66434
rect 38154 66198 38196 66434
rect 37876 59434 38196 66198
rect 37876 59198 37918 59434
rect 38154 59198 38196 59434
rect 37876 52434 38196 59198
rect 37876 52198 37918 52434
rect 38154 52198 38196 52434
rect 37876 45434 38196 52198
rect 37876 45198 37918 45434
rect 38154 45198 38196 45434
rect 37876 38434 38196 45198
rect 37876 38198 37918 38434
rect 38154 38198 38196 38434
rect 37876 31434 38196 38198
rect 37876 31198 37918 31434
rect 38154 31198 38196 31434
rect 37876 24434 38196 31198
rect 37876 24198 37918 24434
rect 38154 24198 38196 24434
rect 37876 17434 38196 24198
rect 37876 17198 37918 17434
rect 38154 17198 38196 17434
rect 37876 10434 38196 17198
rect 37876 10198 37918 10434
rect 38154 10198 38196 10434
rect 37876 3434 38196 10198
rect 37876 3198 37918 3434
rect 38154 3198 38196 3434
rect 37876 -1706 38196 3198
rect 37876 -1942 37918 -1706
rect 38154 -1942 38196 -1706
rect 37876 -2026 38196 -1942
rect 37876 -2262 37918 -2026
rect 38154 -2262 38196 -2026
rect 37876 -2294 38196 -2262
rect 43144 705238 43464 706230
rect 43144 705002 43186 705238
rect 43422 705002 43464 705238
rect 43144 704918 43464 705002
rect 43144 704682 43186 704918
rect 43422 704682 43464 704918
rect 43144 695494 43464 704682
rect 43144 695258 43186 695494
rect 43422 695258 43464 695494
rect 43144 688494 43464 695258
rect 43144 688258 43186 688494
rect 43422 688258 43464 688494
rect 43144 681494 43464 688258
rect 43144 681258 43186 681494
rect 43422 681258 43464 681494
rect 43144 674494 43464 681258
rect 43144 674258 43186 674494
rect 43422 674258 43464 674494
rect 43144 667494 43464 674258
rect 43144 667258 43186 667494
rect 43422 667258 43464 667494
rect 43144 660494 43464 667258
rect 43144 660258 43186 660494
rect 43422 660258 43464 660494
rect 43144 653494 43464 660258
rect 43144 653258 43186 653494
rect 43422 653258 43464 653494
rect 43144 646494 43464 653258
rect 43144 646258 43186 646494
rect 43422 646258 43464 646494
rect 43144 639494 43464 646258
rect 43144 639258 43186 639494
rect 43422 639258 43464 639494
rect 43144 632494 43464 639258
rect 43144 632258 43186 632494
rect 43422 632258 43464 632494
rect 43144 625494 43464 632258
rect 43144 625258 43186 625494
rect 43422 625258 43464 625494
rect 43144 618494 43464 625258
rect 43144 618258 43186 618494
rect 43422 618258 43464 618494
rect 43144 611494 43464 618258
rect 43144 611258 43186 611494
rect 43422 611258 43464 611494
rect 43144 604494 43464 611258
rect 43144 604258 43186 604494
rect 43422 604258 43464 604494
rect 43144 597494 43464 604258
rect 43144 597258 43186 597494
rect 43422 597258 43464 597494
rect 43144 590494 43464 597258
rect 43144 590258 43186 590494
rect 43422 590258 43464 590494
rect 43144 583494 43464 590258
rect 43144 583258 43186 583494
rect 43422 583258 43464 583494
rect 43144 576494 43464 583258
rect 43144 576258 43186 576494
rect 43422 576258 43464 576494
rect 43144 569494 43464 576258
rect 43144 569258 43186 569494
rect 43422 569258 43464 569494
rect 43144 562494 43464 569258
rect 43144 562258 43186 562494
rect 43422 562258 43464 562494
rect 43144 555494 43464 562258
rect 43144 555258 43186 555494
rect 43422 555258 43464 555494
rect 43144 548494 43464 555258
rect 43144 548258 43186 548494
rect 43422 548258 43464 548494
rect 43144 541494 43464 548258
rect 43144 541258 43186 541494
rect 43422 541258 43464 541494
rect 43144 534494 43464 541258
rect 43144 534258 43186 534494
rect 43422 534258 43464 534494
rect 43144 527494 43464 534258
rect 43144 527258 43186 527494
rect 43422 527258 43464 527494
rect 43144 520494 43464 527258
rect 43144 520258 43186 520494
rect 43422 520258 43464 520494
rect 43144 513494 43464 520258
rect 43144 513258 43186 513494
rect 43422 513258 43464 513494
rect 43144 506494 43464 513258
rect 43144 506258 43186 506494
rect 43422 506258 43464 506494
rect 43144 499494 43464 506258
rect 43144 499258 43186 499494
rect 43422 499258 43464 499494
rect 43144 492494 43464 499258
rect 43144 492258 43186 492494
rect 43422 492258 43464 492494
rect 43144 485494 43464 492258
rect 43144 485258 43186 485494
rect 43422 485258 43464 485494
rect 43144 478494 43464 485258
rect 43144 478258 43186 478494
rect 43422 478258 43464 478494
rect 43144 471494 43464 478258
rect 43144 471258 43186 471494
rect 43422 471258 43464 471494
rect 43144 464494 43464 471258
rect 43144 464258 43186 464494
rect 43422 464258 43464 464494
rect 43144 457494 43464 464258
rect 43144 457258 43186 457494
rect 43422 457258 43464 457494
rect 43144 450494 43464 457258
rect 43144 450258 43186 450494
rect 43422 450258 43464 450494
rect 43144 443494 43464 450258
rect 43144 443258 43186 443494
rect 43422 443258 43464 443494
rect 43144 436494 43464 443258
rect 43144 436258 43186 436494
rect 43422 436258 43464 436494
rect 43144 429494 43464 436258
rect 43144 429258 43186 429494
rect 43422 429258 43464 429494
rect 43144 422494 43464 429258
rect 43144 422258 43186 422494
rect 43422 422258 43464 422494
rect 43144 415494 43464 422258
rect 43144 415258 43186 415494
rect 43422 415258 43464 415494
rect 43144 408494 43464 415258
rect 43144 408258 43186 408494
rect 43422 408258 43464 408494
rect 43144 401494 43464 408258
rect 43144 401258 43186 401494
rect 43422 401258 43464 401494
rect 43144 394494 43464 401258
rect 43144 394258 43186 394494
rect 43422 394258 43464 394494
rect 43144 387494 43464 394258
rect 43144 387258 43186 387494
rect 43422 387258 43464 387494
rect 43144 380494 43464 387258
rect 43144 380258 43186 380494
rect 43422 380258 43464 380494
rect 43144 373494 43464 380258
rect 43144 373258 43186 373494
rect 43422 373258 43464 373494
rect 43144 366494 43464 373258
rect 43144 366258 43186 366494
rect 43422 366258 43464 366494
rect 43144 359494 43464 366258
rect 43144 359258 43186 359494
rect 43422 359258 43464 359494
rect 43144 352494 43464 359258
rect 43144 352258 43186 352494
rect 43422 352258 43464 352494
rect 43144 345494 43464 352258
rect 43144 345258 43186 345494
rect 43422 345258 43464 345494
rect 43144 338494 43464 345258
rect 43144 338258 43186 338494
rect 43422 338258 43464 338494
rect 43144 331494 43464 338258
rect 43144 331258 43186 331494
rect 43422 331258 43464 331494
rect 43144 324494 43464 331258
rect 43144 324258 43186 324494
rect 43422 324258 43464 324494
rect 43144 317494 43464 324258
rect 43144 317258 43186 317494
rect 43422 317258 43464 317494
rect 43144 310494 43464 317258
rect 43144 310258 43186 310494
rect 43422 310258 43464 310494
rect 43144 303494 43464 310258
rect 43144 303258 43186 303494
rect 43422 303258 43464 303494
rect 43144 296494 43464 303258
rect 43144 296258 43186 296494
rect 43422 296258 43464 296494
rect 43144 289494 43464 296258
rect 43144 289258 43186 289494
rect 43422 289258 43464 289494
rect 43144 282494 43464 289258
rect 43144 282258 43186 282494
rect 43422 282258 43464 282494
rect 43144 275494 43464 282258
rect 43144 275258 43186 275494
rect 43422 275258 43464 275494
rect 43144 268494 43464 275258
rect 43144 268258 43186 268494
rect 43422 268258 43464 268494
rect 43144 261494 43464 268258
rect 43144 261258 43186 261494
rect 43422 261258 43464 261494
rect 43144 254494 43464 261258
rect 43144 254258 43186 254494
rect 43422 254258 43464 254494
rect 43144 247494 43464 254258
rect 43144 247258 43186 247494
rect 43422 247258 43464 247494
rect 43144 240494 43464 247258
rect 43144 240258 43186 240494
rect 43422 240258 43464 240494
rect 43144 233494 43464 240258
rect 43144 233258 43186 233494
rect 43422 233258 43464 233494
rect 43144 226494 43464 233258
rect 43144 226258 43186 226494
rect 43422 226258 43464 226494
rect 43144 219494 43464 226258
rect 43144 219258 43186 219494
rect 43422 219258 43464 219494
rect 43144 212494 43464 219258
rect 43144 212258 43186 212494
rect 43422 212258 43464 212494
rect 43144 205494 43464 212258
rect 43144 205258 43186 205494
rect 43422 205258 43464 205494
rect 43144 198494 43464 205258
rect 43144 198258 43186 198494
rect 43422 198258 43464 198494
rect 43144 191494 43464 198258
rect 43144 191258 43186 191494
rect 43422 191258 43464 191494
rect 43144 184494 43464 191258
rect 43144 184258 43186 184494
rect 43422 184258 43464 184494
rect 43144 177494 43464 184258
rect 43144 177258 43186 177494
rect 43422 177258 43464 177494
rect 43144 170494 43464 177258
rect 43144 170258 43186 170494
rect 43422 170258 43464 170494
rect 43144 163494 43464 170258
rect 43144 163258 43186 163494
rect 43422 163258 43464 163494
rect 43144 156494 43464 163258
rect 43144 156258 43186 156494
rect 43422 156258 43464 156494
rect 43144 149494 43464 156258
rect 43144 149258 43186 149494
rect 43422 149258 43464 149494
rect 43144 142494 43464 149258
rect 43144 142258 43186 142494
rect 43422 142258 43464 142494
rect 43144 135494 43464 142258
rect 43144 135258 43186 135494
rect 43422 135258 43464 135494
rect 43144 128494 43464 135258
rect 43144 128258 43186 128494
rect 43422 128258 43464 128494
rect 43144 121494 43464 128258
rect 43144 121258 43186 121494
rect 43422 121258 43464 121494
rect 43144 114494 43464 121258
rect 43144 114258 43186 114494
rect 43422 114258 43464 114494
rect 43144 107494 43464 114258
rect 43144 107258 43186 107494
rect 43422 107258 43464 107494
rect 43144 100494 43464 107258
rect 43144 100258 43186 100494
rect 43422 100258 43464 100494
rect 43144 93494 43464 100258
rect 43144 93258 43186 93494
rect 43422 93258 43464 93494
rect 43144 86494 43464 93258
rect 43144 86258 43186 86494
rect 43422 86258 43464 86494
rect 43144 79494 43464 86258
rect 43144 79258 43186 79494
rect 43422 79258 43464 79494
rect 43144 72494 43464 79258
rect 43144 72258 43186 72494
rect 43422 72258 43464 72494
rect 43144 65494 43464 72258
rect 43144 65258 43186 65494
rect 43422 65258 43464 65494
rect 43144 58494 43464 65258
rect 43144 58258 43186 58494
rect 43422 58258 43464 58494
rect 43144 51494 43464 58258
rect 43144 51258 43186 51494
rect 43422 51258 43464 51494
rect 43144 44494 43464 51258
rect 43144 44258 43186 44494
rect 43422 44258 43464 44494
rect 43144 37494 43464 44258
rect 43144 37258 43186 37494
rect 43422 37258 43464 37494
rect 43144 30494 43464 37258
rect 43144 30258 43186 30494
rect 43422 30258 43464 30494
rect 43144 23494 43464 30258
rect 43144 23258 43186 23494
rect 43422 23258 43464 23494
rect 43144 16494 43464 23258
rect 43144 16258 43186 16494
rect 43422 16258 43464 16494
rect 43144 9494 43464 16258
rect 43144 9258 43186 9494
rect 43422 9258 43464 9494
rect 43144 2494 43464 9258
rect 43144 2258 43186 2494
rect 43422 2258 43464 2494
rect 43144 -746 43464 2258
rect 43144 -982 43186 -746
rect 43422 -982 43464 -746
rect 43144 -1066 43464 -982
rect 43144 -1302 43186 -1066
rect 43422 -1302 43464 -1066
rect 43144 -2294 43464 -1302
rect 44876 706198 45196 706230
rect 44876 705962 44918 706198
rect 45154 705962 45196 706198
rect 44876 705878 45196 705962
rect 44876 705642 44918 705878
rect 45154 705642 45196 705878
rect 44876 696434 45196 705642
rect 44876 696198 44918 696434
rect 45154 696198 45196 696434
rect 44876 689434 45196 696198
rect 44876 689198 44918 689434
rect 45154 689198 45196 689434
rect 44876 682434 45196 689198
rect 44876 682198 44918 682434
rect 45154 682198 45196 682434
rect 44876 675434 45196 682198
rect 44876 675198 44918 675434
rect 45154 675198 45196 675434
rect 44876 668434 45196 675198
rect 44876 668198 44918 668434
rect 45154 668198 45196 668434
rect 44876 661434 45196 668198
rect 44876 661198 44918 661434
rect 45154 661198 45196 661434
rect 44876 654434 45196 661198
rect 44876 654198 44918 654434
rect 45154 654198 45196 654434
rect 44876 647434 45196 654198
rect 44876 647198 44918 647434
rect 45154 647198 45196 647434
rect 44876 640434 45196 647198
rect 44876 640198 44918 640434
rect 45154 640198 45196 640434
rect 44876 633434 45196 640198
rect 44876 633198 44918 633434
rect 45154 633198 45196 633434
rect 44876 626434 45196 633198
rect 44876 626198 44918 626434
rect 45154 626198 45196 626434
rect 44876 619434 45196 626198
rect 44876 619198 44918 619434
rect 45154 619198 45196 619434
rect 44876 612434 45196 619198
rect 44876 612198 44918 612434
rect 45154 612198 45196 612434
rect 44876 605434 45196 612198
rect 44876 605198 44918 605434
rect 45154 605198 45196 605434
rect 44876 598434 45196 605198
rect 44876 598198 44918 598434
rect 45154 598198 45196 598434
rect 44876 591434 45196 598198
rect 44876 591198 44918 591434
rect 45154 591198 45196 591434
rect 44876 584434 45196 591198
rect 44876 584198 44918 584434
rect 45154 584198 45196 584434
rect 44876 577434 45196 584198
rect 44876 577198 44918 577434
rect 45154 577198 45196 577434
rect 44876 570434 45196 577198
rect 44876 570198 44918 570434
rect 45154 570198 45196 570434
rect 44876 563434 45196 570198
rect 44876 563198 44918 563434
rect 45154 563198 45196 563434
rect 44876 556434 45196 563198
rect 44876 556198 44918 556434
rect 45154 556198 45196 556434
rect 44876 549434 45196 556198
rect 44876 549198 44918 549434
rect 45154 549198 45196 549434
rect 44876 542434 45196 549198
rect 44876 542198 44918 542434
rect 45154 542198 45196 542434
rect 44876 535434 45196 542198
rect 44876 535198 44918 535434
rect 45154 535198 45196 535434
rect 44876 528434 45196 535198
rect 44876 528198 44918 528434
rect 45154 528198 45196 528434
rect 44876 521434 45196 528198
rect 44876 521198 44918 521434
rect 45154 521198 45196 521434
rect 44876 514434 45196 521198
rect 44876 514198 44918 514434
rect 45154 514198 45196 514434
rect 44876 507434 45196 514198
rect 44876 507198 44918 507434
rect 45154 507198 45196 507434
rect 44876 500434 45196 507198
rect 44876 500198 44918 500434
rect 45154 500198 45196 500434
rect 44876 493434 45196 500198
rect 44876 493198 44918 493434
rect 45154 493198 45196 493434
rect 44876 486434 45196 493198
rect 44876 486198 44918 486434
rect 45154 486198 45196 486434
rect 44876 479434 45196 486198
rect 44876 479198 44918 479434
rect 45154 479198 45196 479434
rect 44876 472434 45196 479198
rect 44876 472198 44918 472434
rect 45154 472198 45196 472434
rect 44876 465434 45196 472198
rect 44876 465198 44918 465434
rect 45154 465198 45196 465434
rect 44876 458434 45196 465198
rect 44876 458198 44918 458434
rect 45154 458198 45196 458434
rect 44876 451434 45196 458198
rect 44876 451198 44918 451434
rect 45154 451198 45196 451434
rect 44876 444434 45196 451198
rect 44876 444198 44918 444434
rect 45154 444198 45196 444434
rect 44876 437434 45196 444198
rect 44876 437198 44918 437434
rect 45154 437198 45196 437434
rect 44876 430434 45196 437198
rect 44876 430198 44918 430434
rect 45154 430198 45196 430434
rect 44876 423434 45196 430198
rect 44876 423198 44918 423434
rect 45154 423198 45196 423434
rect 44876 416434 45196 423198
rect 44876 416198 44918 416434
rect 45154 416198 45196 416434
rect 44876 409434 45196 416198
rect 44876 409198 44918 409434
rect 45154 409198 45196 409434
rect 44876 402434 45196 409198
rect 44876 402198 44918 402434
rect 45154 402198 45196 402434
rect 44876 395434 45196 402198
rect 44876 395198 44918 395434
rect 45154 395198 45196 395434
rect 44876 388434 45196 395198
rect 44876 388198 44918 388434
rect 45154 388198 45196 388434
rect 44876 381434 45196 388198
rect 44876 381198 44918 381434
rect 45154 381198 45196 381434
rect 44876 374434 45196 381198
rect 44876 374198 44918 374434
rect 45154 374198 45196 374434
rect 44876 367434 45196 374198
rect 44876 367198 44918 367434
rect 45154 367198 45196 367434
rect 44876 360434 45196 367198
rect 44876 360198 44918 360434
rect 45154 360198 45196 360434
rect 44876 353434 45196 360198
rect 44876 353198 44918 353434
rect 45154 353198 45196 353434
rect 44876 346434 45196 353198
rect 44876 346198 44918 346434
rect 45154 346198 45196 346434
rect 44876 339434 45196 346198
rect 44876 339198 44918 339434
rect 45154 339198 45196 339434
rect 44876 332434 45196 339198
rect 44876 332198 44918 332434
rect 45154 332198 45196 332434
rect 44876 325434 45196 332198
rect 44876 325198 44918 325434
rect 45154 325198 45196 325434
rect 44876 318434 45196 325198
rect 44876 318198 44918 318434
rect 45154 318198 45196 318434
rect 44876 311434 45196 318198
rect 44876 311198 44918 311434
rect 45154 311198 45196 311434
rect 44876 304434 45196 311198
rect 44876 304198 44918 304434
rect 45154 304198 45196 304434
rect 44876 297434 45196 304198
rect 44876 297198 44918 297434
rect 45154 297198 45196 297434
rect 44876 290434 45196 297198
rect 44876 290198 44918 290434
rect 45154 290198 45196 290434
rect 44876 283434 45196 290198
rect 44876 283198 44918 283434
rect 45154 283198 45196 283434
rect 44876 276434 45196 283198
rect 44876 276198 44918 276434
rect 45154 276198 45196 276434
rect 44876 269434 45196 276198
rect 44876 269198 44918 269434
rect 45154 269198 45196 269434
rect 44876 262434 45196 269198
rect 44876 262198 44918 262434
rect 45154 262198 45196 262434
rect 44876 255434 45196 262198
rect 44876 255198 44918 255434
rect 45154 255198 45196 255434
rect 44876 248434 45196 255198
rect 44876 248198 44918 248434
rect 45154 248198 45196 248434
rect 44876 241434 45196 248198
rect 44876 241198 44918 241434
rect 45154 241198 45196 241434
rect 44876 234434 45196 241198
rect 44876 234198 44918 234434
rect 45154 234198 45196 234434
rect 44876 227434 45196 234198
rect 44876 227198 44918 227434
rect 45154 227198 45196 227434
rect 44876 220434 45196 227198
rect 44876 220198 44918 220434
rect 45154 220198 45196 220434
rect 44876 213434 45196 220198
rect 44876 213198 44918 213434
rect 45154 213198 45196 213434
rect 44876 206434 45196 213198
rect 44876 206198 44918 206434
rect 45154 206198 45196 206434
rect 44876 199434 45196 206198
rect 44876 199198 44918 199434
rect 45154 199198 45196 199434
rect 44876 192434 45196 199198
rect 44876 192198 44918 192434
rect 45154 192198 45196 192434
rect 44876 185434 45196 192198
rect 44876 185198 44918 185434
rect 45154 185198 45196 185434
rect 44876 178434 45196 185198
rect 44876 178198 44918 178434
rect 45154 178198 45196 178434
rect 44876 171434 45196 178198
rect 44876 171198 44918 171434
rect 45154 171198 45196 171434
rect 44876 164434 45196 171198
rect 44876 164198 44918 164434
rect 45154 164198 45196 164434
rect 44876 157434 45196 164198
rect 44876 157198 44918 157434
rect 45154 157198 45196 157434
rect 44876 150434 45196 157198
rect 44876 150198 44918 150434
rect 45154 150198 45196 150434
rect 44876 143434 45196 150198
rect 44876 143198 44918 143434
rect 45154 143198 45196 143434
rect 44876 136434 45196 143198
rect 44876 136198 44918 136434
rect 45154 136198 45196 136434
rect 44876 129434 45196 136198
rect 44876 129198 44918 129434
rect 45154 129198 45196 129434
rect 44876 122434 45196 129198
rect 44876 122198 44918 122434
rect 45154 122198 45196 122434
rect 44876 115434 45196 122198
rect 44876 115198 44918 115434
rect 45154 115198 45196 115434
rect 44876 108434 45196 115198
rect 44876 108198 44918 108434
rect 45154 108198 45196 108434
rect 44876 101434 45196 108198
rect 44876 101198 44918 101434
rect 45154 101198 45196 101434
rect 44876 94434 45196 101198
rect 44876 94198 44918 94434
rect 45154 94198 45196 94434
rect 44876 87434 45196 94198
rect 44876 87198 44918 87434
rect 45154 87198 45196 87434
rect 44876 80434 45196 87198
rect 44876 80198 44918 80434
rect 45154 80198 45196 80434
rect 44876 73434 45196 80198
rect 44876 73198 44918 73434
rect 45154 73198 45196 73434
rect 44876 66434 45196 73198
rect 44876 66198 44918 66434
rect 45154 66198 45196 66434
rect 44876 59434 45196 66198
rect 44876 59198 44918 59434
rect 45154 59198 45196 59434
rect 44876 52434 45196 59198
rect 44876 52198 44918 52434
rect 45154 52198 45196 52434
rect 44876 45434 45196 52198
rect 44876 45198 44918 45434
rect 45154 45198 45196 45434
rect 44876 38434 45196 45198
rect 44876 38198 44918 38434
rect 45154 38198 45196 38434
rect 44876 31434 45196 38198
rect 44876 31198 44918 31434
rect 45154 31198 45196 31434
rect 44876 24434 45196 31198
rect 44876 24198 44918 24434
rect 45154 24198 45196 24434
rect 44876 17434 45196 24198
rect 44876 17198 44918 17434
rect 45154 17198 45196 17434
rect 44876 10434 45196 17198
rect 44876 10198 44918 10434
rect 45154 10198 45196 10434
rect 44876 3434 45196 10198
rect 44876 3198 44918 3434
rect 45154 3198 45196 3434
rect 44876 -1706 45196 3198
rect 44876 -1942 44918 -1706
rect 45154 -1942 45196 -1706
rect 44876 -2026 45196 -1942
rect 44876 -2262 44918 -2026
rect 45154 -2262 45196 -2026
rect 44876 -2294 45196 -2262
rect 50144 705238 50464 706230
rect 50144 705002 50186 705238
rect 50422 705002 50464 705238
rect 50144 704918 50464 705002
rect 50144 704682 50186 704918
rect 50422 704682 50464 704918
rect 50144 695494 50464 704682
rect 50144 695258 50186 695494
rect 50422 695258 50464 695494
rect 50144 688494 50464 695258
rect 50144 688258 50186 688494
rect 50422 688258 50464 688494
rect 50144 681494 50464 688258
rect 50144 681258 50186 681494
rect 50422 681258 50464 681494
rect 50144 674494 50464 681258
rect 50144 674258 50186 674494
rect 50422 674258 50464 674494
rect 50144 667494 50464 674258
rect 50144 667258 50186 667494
rect 50422 667258 50464 667494
rect 50144 660494 50464 667258
rect 50144 660258 50186 660494
rect 50422 660258 50464 660494
rect 50144 653494 50464 660258
rect 50144 653258 50186 653494
rect 50422 653258 50464 653494
rect 50144 646494 50464 653258
rect 50144 646258 50186 646494
rect 50422 646258 50464 646494
rect 50144 639494 50464 646258
rect 50144 639258 50186 639494
rect 50422 639258 50464 639494
rect 50144 632494 50464 639258
rect 50144 632258 50186 632494
rect 50422 632258 50464 632494
rect 50144 625494 50464 632258
rect 50144 625258 50186 625494
rect 50422 625258 50464 625494
rect 50144 618494 50464 625258
rect 50144 618258 50186 618494
rect 50422 618258 50464 618494
rect 50144 611494 50464 618258
rect 50144 611258 50186 611494
rect 50422 611258 50464 611494
rect 50144 604494 50464 611258
rect 50144 604258 50186 604494
rect 50422 604258 50464 604494
rect 50144 597494 50464 604258
rect 50144 597258 50186 597494
rect 50422 597258 50464 597494
rect 50144 590494 50464 597258
rect 50144 590258 50186 590494
rect 50422 590258 50464 590494
rect 50144 583494 50464 590258
rect 50144 583258 50186 583494
rect 50422 583258 50464 583494
rect 50144 576494 50464 583258
rect 50144 576258 50186 576494
rect 50422 576258 50464 576494
rect 50144 569494 50464 576258
rect 50144 569258 50186 569494
rect 50422 569258 50464 569494
rect 50144 562494 50464 569258
rect 50144 562258 50186 562494
rect 50422 562258 50464 562494
rect 50144 555494 50464 562258
rect 50144 555258 50186 555494
rect 50422 555258 50464 555494
rect 50144 548494 50464 555258
rect 50144 548258 50186 548494
rect 50422 548258 50464 548494
rect 50144 541494 50464 548258
rect 50144 541258 50186 541494
rect 50422 541258 50464 541494
rect 50144 534494 50464 541258
rect 50144 534258 50186 534494
rect 50422 534258 50464 534494
rect 50144 527494 50464 534258
rect 50144 527258 50186 527494
rect 50422 527258 50464 527494
rect 50144 520494 50464 527258
rect 50144 520258 50186 520494
rect 50422 520258 50464 520494
rect 50144 513494 50464 520258
rect 50144 513258 50186 513494
rect 50422 513258 50464 513494
rect 50144 506494 50464 513258
rect 50144 506258 50186 506494
rect 50422 506258 50464 506494
rect 50144 499494 50464 506258
rect 50144 499258 50186 499494
rect 50422 499258 50464 499494
rect 50144 492494 50464 499258
rect 50144 492258 50186 492494
rect 50422 492258 50464 492494
rect 50144 485494 50464 492258
rect 50144 485258 50186 485494
rect 50422 485258 50464 485494
rect 50144 478494 50464 485258
rect 50144 478258 50186 478494
rect 50422 478258 50464 478494
rect 50144 471494 50464 478258
rect 50144 471258 50186 471494
rect 50422 471258 50464 471494
rect 50144 464494 50464 471258
rect 50144 464258 50186 464494
rect 50422 464258 50464 464494
rect 50144 457494 50464 464258
rect 50144 457258 50186 457494
rect 50422 457258 50464 457494
rect 50144 450494 50464 457258
rect 50144 450258 50186 450494
rect 50422 450258 50464 450494
rect 50144 443494 50464 450258
rect 50144 443258 50186 443494
rect 50422 443258 50464 443494
rect 50144 436494 50464 443258
rect 50144 436258 50186 436494
rect 50422 436258 50464 436494
rect 50144 429494 50464 436258
rect 50144 429258 50186 429494
rect 50422 429258 50464 429494
rect 50144 422494 50464 429258
rect 50144 422258 50186 422494
rect 50422 422258 50464 422494
rect 50144 415494 50464 422258
rect 50144 415258 50186 415494
rect 50422 415258 50464 415494
rect 50144 408494 50464 415258
rect 50144 408258 50186 408494
rect 50422 408258 50464 408494
rect 50144 401494 50464 408258
rect 50144 401258 50186 401494
rect 50422 401258 50464 401494
rect 50144 394494 50464 401258
rect 50144 394258 50186 394494
rect 50422 394258 50464 394494
rect 50144 387494 50464 394258
rect 50144 387258 50186 387494
rect 50422 387258 50464 387494
rect 50144 380494 50464 387258
rect 50144 380258 50186 380494
rect 50422 380258 50464 380494
rect 50144 373494 50464 380258
rect 50144 373258 50186 373494
rect 50422 373258 50464 373494
rect 50144 366494 50464 373258
rect 50144 366258 50186 366494
rect 50422 366258 50464 366494
rect 50144 359494 50464 366258
rect 50144 359258 50186 359494
rect 50422 359258 50464 359494
rect 50144 352494 50464 359258
rect 50144 352258 50186 352494
rect 50422 352258 50464 352494
rect 50144 345494 50464 352258
rect 50144 345258 50186 345494
rect 50422 345258 50464 345494
rect 50144 338494 50464 345258
rect 50144 338258 50186 338494
rect 50422 338258 50464 338494
rect 50144 331494 50464 338258
rect 50144 331258 50186 331494
rect 50422 331258 50464 331494
rect 50144 324494 50464 331258
rect 50144 324258 50186 324494
rect 50422 324258 50464 324494
rect 50144 317494 50464 324258
rect 50144 317258 50186 317494
rect 50422 317258 50464 317494
rect 50144 310494 50464 317258
rect 50144 310258 50186 310494
rect 50422 310258 50464 310494
rect 50144 303494 50464 310258
rect 50144 303258 50186 303494
rect 50422 303258 50464 303494
rect 50144 296494 50464 303258
rect 50144 296258 50186 296494
rect 50422 296258 50464 296494
rect 50144 289494 50464 296258
rect 50144 289258 50186 289494
rect 50422 289258 50464 289494
rect 50144 282494 50464 289258
rect 50144 282258 50186 282494
rect 50422 282258 50464 282494
rect 50144 275494 50464 282258
rect 50144 275258 50186 275494
rect 50422 275258 50464 275494
rect 50144 268494 50464 275258
rect 50144 268258 50186 268494
rect 50422 268258 50464 268494
rect 50144 261494 50464 268258
rect 50144 261258 50186 261494
rect 50422 261258 50464 261494
rect 50144 254494 50464 261258
rect 50144 254258 50186 254494
rect 50422 254258 50464 254494
rect 50144 247494 50464 254258
rect 50144 247258 50186 247494
rect 50422 247258 50464 247494
rect 50144 240494 50464 247258
rect 50144 240258 50186 240494
rect 50422 240258 50464 240494
rect 50144 233494 50464 240258
rect 50144 233258 50186 233494
rect 50422 233258 50464 233494
rect 50144 226494 50464 233258
rect 50144 226258 50186 226494
rect 50422 226258 50464 226494
rect 50144 219494 50464 226258
rect 50144 219258 50186 219494
rect 50422 219258 50464 219494
rect 50144 212494 50464 219258
rect 50144 212258 50186 212494
rect 50422 212258 50464 212494
rect 50144 205494 50464 212258
rect 50144 205258 50186 205494
rect 50422 205258 50464 205494
rect 50144 198494 50464 205258
rect 50144 198258 50186 198494
rect 50422 198258 50464 198494
rect 50144 191494 50464 198258
rect 50144 191258 50186 191494
rect 50422 191258 50464 191494
rect 50144 184494 50464 191258
rect 50144 184258 50186 184494
rect 50422 184258 50464 184494
rect 50144 177494 50464 184258
rect 50144 177258 50186 177494
rect 50422 177258 50464 177494
rect 50144 170494 50464 177258
rect 50144 170258 50186 170494
rect 50422 170258 50464 170494
rect 50144 163494 50464 170258
rect 50144 163258 50186 163494
rect 50422 163258 50464 163494
rect 50144 156494 50464 163258
rect 50144 156258 50186 156494
rect 50422 156258 50464 156494
rect 50144 149494 50464 156258
rect 50144 149258 50186 149494
rect 50422 149258 50464 149494
rect 50144 142494 50464 149258
rect 50144 142258 50186 142494
rect 50422 142258 50464 142494
rect 50144 135494 50464 142258
rect 50144 135258 50186 135494
rect 50422 135258 50464 135494
rect 50144 128494 50464 135258
rect 50144 128258 50186 128494
rect 50422 128258 50464 128494
rect 50144 121494 50464 128258
rect 50144 121258 50186 121494
rect 50422 121258 50464 121494
rect 50144 114494 50464 121258
rect 50144 114258 50186 114494
rect 50422 114258 50464 114494
rect 50144 107494 50464 114258
rect 50144 107258 50186 107494
rect 50422 107258 50464 107494
rect 50144 100494 50464 107258
rect 50144 100258 50186 100494
rect 50422 100258 50464 100494
rect 50144 93494 50464 100258
rect 50144 93258 50186 93494
rect 50422 93258 50464 93494
rect 50144 86494 50464 93258
rect 50144 86258 50186 86494
rect 50422 86258 50464 86494
rect 50144 79494 50464 86258
rect 50144 79258 50186 79494
rect 50422 79258 50464 79494
rect 50144 72494 50464 79258
rect 50144 72258 50186 72494
rect 50422 72258 50464 72494
rect 50144 65494 50464 72258
rect 50144 65258 50186 65494
rect 50422 65258 50464 65494
rect 50144 58494 50464 65258
rect 50144 58258 50186 58494
rect 50422 58258 50464 58494
rect 50144 51494 50464 58258
rect 50144 51258 50186 51494
rect 50422 51258 50464 51494
rect 50144 44494 50464 51258
rect 50144 44258 50186 44494
rect 50422 44258 50464 44494
rect 50144 37494 50464 44258
rect 50144 37258 50186 37494
rect 50422 37258 50464 37494
rect 50144 30494 50464 37258
rect 50144 30258 50186 30494
rect 50422 30258 50464 30494
rect 50144 23494 50464 30258
rect 50144 23258 50186 23494
rect 50422 23258 50464 23494
rect 50144 16494 50464 23258
rect 50144 16258 50186 16494
rect 50422 16258 50464 16494
rect 50144 9494 50464 16258
rect 50144 9258 50186 9494
rect 50422 9258 50464 9494
rect 50144 2494 50464 9258
rect 50144 2258 50186 2494
rect 50422 2258 50464 2494
rect 50144 -746 50464 2258
rect 50144 -982 50186 -746
rect 50422 -982 50464 -746
rect 50144 -1066 50464 -982
rect 50144 -1302 50186 -1066
rect 50422 -1302 50464 -1066
rect 50144 -2294 50464 -1302
rect 51876 706198 52196 706230
rect 51876 705962 51918 706198
rect 52154 705962 52196 706198
rect 51876 705878 52196 705962
rect 51876 705642 51918 705878
rect 52154 705642 52196 705878
rect 51876 696434 52196 705642
rect 51876 696198 51918 696434
rect 52154 696198 52196 696434
rect 51876 689434 52196 696198
rect 51876 689198 51918 689434
rect 52154 689198 52196 689434
rect 51876 682434 52196 689198
rect 51876 682198 51918 682434
rect 52154 682198 52196 682434
rect 51876 675434 52196 682198
rect 51876 675198 51918 675434
rect 52154 675198 52196 675434
rect 51876 668434 52196 675198
rect 51876 668198 51918 668434
rect 52154 668198 52196 668434
rect 51876 661434 52196 668198
rect 51876 661198 51918 661434
rect 52154 661198 52196 661434
rect 51876 654434 52196 661198
rect 51876 654198 51918 654434
rect 52154 654198 52196 654434
rect 51876 647434 52196 654198
rect 51876 647198 51918 647434
rect 52154 647198 52196 647434
rect 51876 640434 52196 647198
rect 51876 640198 51918 640434
rect 52154 640198 52196 640434
rect 51876 633434 52196 640198
rect 51876 633198 51918 633434
rect 52154 633198 52196 633434
rect 51876 626434 52196 633198
rect 51876 626198 51918 626434
rect 52154 626198 52196 626434
rect 51876 619434 52196 626198
rect 51876 619198 51918 619434
rect 52154 619198 52196 619434
rect 51876 612434 52196 619198
rect 51876 612198 51918 612434
rect 52154 612198 52196 612434
rect 51876 605434 52196 612198
rect 51876 605198 51918 605434
rect 52154 605198 52196 605434
rect 51876 598434 52196 605198
rect 51876 598198 51918 598434
rect 52154 598198 52196 598434
rect 51876 591434 52196 598198
rect 51876 591198 51918 591434
rect 52154 591198 52196 591434
rect 51876 584434 52196 591198
rect 51876 584198 51918 584434
rect 52154 584198 52196 584434
rect 51876 577434 52196 584198
rect 51876 577198 51918 577434
rect 52154 577198 52196 577434
rect 51876 570434 52196 577198
rect 51876 570198 51918 570434
rect 52154 570198 52196 570434
rect 51876 563434 52196 570198
rect 51876 563198 51918 563434
rect 52154 563198 52196 563434
rect 51876 556434 52196 563198
rect 51876 556198 51918 556434
rect 52154 556198 52196 556434
rect 51876 549434 52196 556198
rect 51876 549198 51918 549434
rect 52154 549198 52196 549434
rect 51876 542434 52196 549198
rect 51876 542198 51918 542434
rect 52154 542198 52196 542434
rect 51876 535434 52196 542198
rect 51876 535198 51918 535434
rect 52154 535198 52196 535434
rect 51876 528434 52196 535198
rect 51876 528198 51918 528434
rect 52154 528198 52196 528434
rect 51876 521434 52196 528198
rect 51876 521198 51918 521434
rect 52154 521198 52196 521434
rect 51876 514434 52196 521198
rect 51876 514198 51918 514434
rect 52154 514198 52196 514434
rect 51876 507434 52196 514198
rect 51876 507198 51918 507434
rect 52154 507198 52196 507434
rect 51876 500434 52196 507198
rect 51876 500198 51918 500434
rect 52154 500198 52196 500434
rect 51876 493434 52196 500198
rect 51876 493198 51918 493434
rect 52154 493198 52196 493434
rect 51876 486434 52196 493198
rect 51876 486198 51918 486434
rect 52154 486198 52196 486434
rect 51876 479434 52196 486198
rect 51876 479198 51918 479434
rect 52154 479198 52196 479434
rect 51876 472434 52196 479198
rect 51876 472198 51918 472434
rect 52154 472198 52196 472434
rect 51876 465434 52196 472198
rect 51876 465198 51918 465434
rect 52154 465198 52196 465434
rect 51876 458434 52196 465198
rect 51876 458198 51918 458434
rect 52154 458198 52196 458434
rect 51876 451434 52196 458198
rect 51876 451198 51918 451434
rect 52154 451198 52196 451434
rect 51876 444434 52196 451198
rect 51876 444198 51918 444434
rect 52154 444198 52196 444434
rect 51876 437434 52196 444198
rect 51876 437198 51918 437434
rect 52154 437198 52196 437434
rect 51876 430434 52196 437198
rect 51876 430198 51918 430434
rect 52154 430198 52196 430434
rect 51876 423434 52196 430198
rect 51876 423198 51918 423434
rect 52154 423198 52196 423434
rect 51876 416434 52196 423198
rect 51876 416198 51918 416434
rect 52154 416198 52196 416434
rect 51876 409434 52196 416198
rect 51876 409198 51918 409434
rect 52154 409198 52196 409434
rect 51876 402434 52196 409198
rect 51876 402198 51918 402434
rect 52154 402198 52196 402434
rect 51876 395434 52196 402198
rect 51876 395198 51918 395434
rect 52154 395198 52196 395434
rect 51876 388434 52196 395198
rect 51876 388198 51918 388434
rect 52154 388198 52196 388434
rect 51876 381434 52196 388198
rect 51876 381198 51918 381434
rect 52154 381198 52196 381434
rect 51876 374434 52196 381198
rect 51876 374198 51918 374434
rect 52154 374198 52196 374434
rect 51876 367434 52196 374198
rect 51876 367198 51918 367434
rect 52154 367198 52196 367434
rect 51876 360434 52196 367198
rect 51876 360198 51918 360434
rect 52154 360198 52196 360434
rect 51876 353434 52196 360198
rect 51876 353198 51918 353434
rect 52154 353198 52196 353434
rect 51876 346434 52196 353198
rect 51876 346198 51918 346434
rect 52154 346198 52196 346434
rect 51876 339434 52196 346198
rect 51876 339198 51918 339434
rect 52154 339198 52196 339434
rect 51876 332434 52196 339198
rect 51876 332198 51918 332434
rect 52154 332198 52196 332434
rect 51876 325434 52196 332198
rect 51876 325198 51918 325434
rect 52154 325198 52196 325434
rect 51876 318434 52196 325198
rect 51876 318198 51918 318434
rect 52154 318198 52196 318434
rect 51876 311434 52196 318198
rect 51876 311198 51918 311434
rect 52154 311198 52196 311434
rect 51876 304434 52196 311198
rect 51876 304198 51918 304434
rect 52154 304198 52196 304434
rect 51876 297434 52196 304198
rect 51876 297198 51918 297434
rect 52154 297198 52196 297434
rect 51876 290434 52196 297198
rect 51876 290198 51918 290434
rect 52154 290198 52196 290434
rect 51876 283434 52196 290198
rect 51876 283198 51918 283434
rect 52154 283198 52196 283434
rect 51876 276434 52196 283198
rect 51876 276198 51918 276434
rect 52154 276198 52196 276434
rect 51876 269434 52196 276198
rect 51876 269198 51918 269434
rect 52154 269198 52196 269434
rect 51876 262434 52196 269198
rect 51876 262198 51918 262434
rect 52154 262198 52196 262434
rect 51876 255434 52196 262198
rect 51876 255198 51918 255434
rect 52154 255198 52196 255434
rect 51876 248434 52196 255198
rect 51876 248198 51918 248434
rect 52154 248198 52196 248434
rect 51876 241434 52196 248198
rect 51876 241198 51918 241434
rect 52154 241198 52196 241434
rect 51876 234434 52196 241198
rect 51876 234198 51918 234434
rect 52154 234198 52196 234434
rect 51876 227434 52196 234198
rect 51876 227198 51918 227434
rect 52154 227198 52196 227434
rect 51876 220434 52196 227198
rect 51876 220198 51918 220434
rect 52154 220198 52196 220434
rect 51876 213434 52196 220198
rect 51876 213198 51918 213434
rect 52154 213198 52196 213434
rect 51876 206434 52196 213198
rect 51876 206198 51918 206434
rect 52154 206198 52196 206434
rect 51876 199434 52196 206198
rect 51876 199198 51918 199434
rect 52154 199198 52196 199434
rect 51876 192434 52196 199198
rect 51876 192198 51918 192434
rect 52154 192198 52196 192434
rect 51876 185434 52196 192198
rect 51876 185198 51918 185434
rect 52154 185198 52196 185434
rect 51876 178434 52196 185198
rect 51876 178198 51918 178434
rect 52154 178198 52196 178434
rect 51876 171434 52196 178198
rect 51876 171198 51918 171434
rect 52154 171198 52196 171434
rect 51876 164434 52196 171198
rect 51876 164198 51918 164434
rect 52154 164198 52196 164434
rect 51876 157434 52196 164198
rect 51876 157198 51918 157434
rect 52154 157198 52196 157434
rect 51876 150434 52196 157198
rect 51876 150198 51918 150434
rect 52154 150198 52196 150434
rect 51876 143434 52196 150198
rect 51876 143198 51918 143434
rect 52154 143198 52196 143434
rect 51876 136434 52196 143198
rect 51876 136198 51918 136434
rect 52154 136198 52196 136434
rect 51876 129434 52196 136198
rect 51876 129198 51918 129434
rect 52154 129198 52196 129434
rect 51876 122434 52196 129198
rect 51876 122198 51918 122434
rect 52154 122198 52196 122434
rect 51876 115434 52196 122198
rect 51876 115198 51918 115434
rect 52154 115198 52196 115434
rect 51876 108434 52196 115198
rect 51876 108198 51918 108434
rect 52154 108198 52196 108434
rect 51876 101434 52196 108198
rect 51876 101198 51918 101434
rect 52154 101198 52196 101434
rect 51876 94434 52196 101198
rect 51876 94198 51918 94434
rect 52154 94198 52196 94434
rect 51876 87434 52196 94198
rect 51876 87198 51918 87434
rect 52154 87198 52196 87434
rect 51876 80434 52196 87198
rect 51876 80198 51918 80434
rect 52154 80198 52196 80434
rect 51876 73434 52196 80198
rect 51876 73198 51918 73434
rect 52154 73198 52196 73434
rect 51876 66434 52196 73198
rect 51876 66198 51918 66434
rect 52154 66198 52196 66434
rect 51876 59434 52196 66198
rect 51876 59198 51918 59434
rect 52154 59198 52196 59434
rect 51876 52434 52196 59198
rect 51876 52198 51918 52434
rect 52154 52198 52196 52434
rect 51876 45434 52196 52198
rect 51876 45198 51918 45434
rect 52154 45198 52196 45434
rect 51876 38434 52196 45198
rect 51876 38198 51918 38434
rect 52154 38198 52196 38434
rect 51876 31434 52196 38198
rect 51876 31198 51918 31434
rect 52154 31198 52196 31434
rect 51876 24434 52196 31198
rect 51876 24198 51918 24434
rect 52154 24198 52196 24434
rect 51876 17434 52196 24198
rect 51876 17198 51918 17434
rect 52154 17198 52196 17434
rect 51876 10434 52196 17198
rect 51876 10198 51918 10434
rect 52154 10198 52196 10434
rect 51876 3434 52196 10198
rect 51876 3198 51918 3434
rect 52154 3198 52196 3434
rect 51876 -1706 52196 3198
rect 51876 -1942 51918 -1706
rect 52154 -1942 52196 -1706
rect 51876 -2026 52196 -1942
rect 51876 -2262 51918 -2026
rect 52154 -2262 52196 -2026
rect 51876 -2294 52196 -2262
rect 57144 705238 57464 706230
rect 57144 705002 57186 705238
rect 57422 705002 57464 705238
rect 57144 704918 57464 705002
rect 57144 704682 57186 704918
rect 57422 704682 57464 704918
rect 57144 695494 57464 704682
rect 57144 695258 57186 695494
rect 57422 695258 57464 695494
rect 57144 688494 57464 695258
rect 57144 688258 57186 688494
rect 57422 688258 57464 688494
rect 57144 681494 57464 688258
rect 57144 681258 57186 681494
rect 57422 681258 57464 681494
rect 57144 674494 57464 681258
rect 57144 674258 57186 674494
rect 57422 674258 57464 674494
rect 57144 667494 57464 674258
rect 57144 667258 57186 667494
rect 57422 667258 57464 667494
rect 57144 660494 57464 667258
rect 57144 660258 57186 660494
rect 57422 660258 57464 660494
rect 57144 653494 57464 660258
rect 57144 653258 57186 653494
rect 57422 653258 57464 653494
rect 57144 646494 57464 653258
rect 57144 646258 57186 646494
rect 57422 646258 57464 646494
rect 57144 639494 57464 646258
rect 57144 639258 57186 639494
rect 57422 639258 57464 639494
rect 57144 632494 57464 639258
rect 57144 632258 57186 632494
rect 57422 632258 57464 632494
rect 57144 625494 57464 632258
rect 57144 625258 57186 625494
rect 57422 625258 57464 625494
rect 57144 618494 57464 625258
rect 57144 618258 57186 618494
rect 57422 618258 57464 618494
rect 57144 611494 57464 618258
rect 57144 611258 57186 611494
rect 57422 611258 57464 611494
rect 57144 604494 57464 611258
rect 57144 604258 57186 604494
rect 57422 604258 57464 604494
rect 57144 597494 57464 604258
rect 57144 597258 57186 597494
rect 57422 597258 57464 597494
rect 57144 590494 57464 597258
rect 57144 590258 57186 590494
rect 57422 590258 57464 590494
rect 57144 583494 57464 590258
rect 57144 583258 57186 583494
rect 57422 583258 57464 583494
rect 57144 576494 57464 583258
rect 57144 576258 57186 576494
rect 57422 576258 57464 576494
rect 57144 569494 57464 576258
rect 57144 569258 57186 569494
rect 57422 569258 57464 569494
rect 57144 562494 57464 569258
rect 57144 562258 57186 562494
rect 57422 562258 57464 562494
rect 57144 555494 57464 562258
rect 57144 555258 57186 555494
rect 57422 555258 57464 555494
rect 57144 548494 57464 555258
rect 57144 548258 57186 548494
rect 57422 548258 57464 548494
rect 57144 541494 57464 548258
rect 57144 541258 57186 541494
rect 57422 541258 57464 541494
rect 57144 534494 57464 541258
rect 57144 534258 57186 534494
rect 57422 534258 57464 534494
rect 57144 527494 57464 534258
rect 57144 527258 57186 527494
rect 57422 527258 57464 527494
rect 57144 520494 57464 527258
rect 57144 520258 57186 520494
rect 57422 520258 57464 520494
rect 57144 513494 57464 520258
rect 57144 513258 57186 513494
rect 57422 513258 57464 513494
rect 57144 506494 57464 513258
rect 57144 506258 57186 506494
rect 57422 506258 57464 506494
rect 57144 499494 57464 506258
rect 57144 499258 57186 499494
rect 57422 499258 57464 499494
rect 57144 492494 57464 499258
rect 57144 492258 57186 492494
rect 57422 492258 57464 492494
rect 57144 485494 57464 492258
rect 57144 485258 57186 485494
rect 57422 485258 57464 485494
rect 57144 478494 57464 485258
rect 57144 478258 57186 478494
rect 57422 478258 57464 478494
rect 57144 471494 57464 478258
rect 57144 471258 57186 471494
rect 57422 471258 57464 471494
rect 57144 464494 57464 471258
rect 57144 464258 57186 464494
rect 57422 464258 57464 464494
rect 57144 457494 57464 464258
rect 57144 457258 57186 457494
rect 57422 457258 57464 457494
rect 57144 450494 57464 457258
rect 57144 450258 57186 450494
rect 57422 450258 57464 450494
rect 57144 443494 57464 450258
rect 57144 443258 57186 443494
rect 57422 443258 57464 443494
rect 57144 436494 57464 443258
rect 57144 436258 57186 436494
rect 57422 436258 57464 436494
rect 57144 429494 57464 436258
rect 57144 429258 57186 429494
rect 57422 429258 57464 429494
rect 57144 422494 57464 429258
rect 57144 422258 57186 422494
rect 57422 422258 57464 422494
rect 57144 415494 57464 422258
rect 57144 415258 57186 415494
rect 57422 415258 57464 415494
rect 57144 408494 57464 415258
rect 57144 408258 57186 408494
rect 57422 408258 57464 408494
rect 57144 401494 57464 408258
rect 57144 401258 57186 401494
rect 57422 401258 57464 401494
rect 57144 394494 57464 401258
rect 57144 394258 57186 394494
rect 57422 394258 57464 394494
rect 57144 387494 57464 394258
rect 57144 387258 57186 387494
rect 57422 387258 57464 387494
rect 57144 380494 57464 387258
rect 57144 380258 57186 380494
rect 57422 380258 57464 380494
rect 57144 373494 57464 380258
rect 57144 373258 57186 373494
rect 57422 373258 57464 373494
rect 57144 366494 57464 373258
rect 57144 366258 57186 366494
rect 57422 366258 57464 366494
rect 57144 359494 57464 366258
rect 57144 359258 57186 359494
rect 57422 359258 57464 359494
rect 57144 352494 57464 359258
rect 57144 352258 57186 352494
rect 57422 352258 57464 352494
rect 57144 345494 57464 352258
rect 57144 345258 57186 345494
rect 57422 345258 57464 345494
rect 57144 338494 57464 345258
rect 57144 338258 57186 338494
rect 57422 338258 57464 338494
rect 57144 331494 57464 338258
rect 57144 331258 57186 331494
rect 57422 331258 57464 331494
rect 57144 324494 57464 331258
rect 57144 324258 57186 324494
rect 57422 324258 57464 324494
rect 57144 317494 57464 324258
rect 57144 317258 57186 317494
rect 57422 317258 57464 317494
rect 57144 310494 57464 317258
rect 57144 310258 57186 310494
rect 57422 310258 57464 310494
rect 57144 303494 57464 310258
rect 57144 303258 57186 303494
rect 57422 303258 57464 303494
rect 57144 296494 57464 303258
rect 57144 296258 57186 296494
rect 57422 296258 57464 296494
rect 57144 289494 57464 296258
rect 57144 289258 57186 289494
rect 57422 289258 57464 289494
rect 57144 282494 57464 289258
rect 57144 282258 57186 282494
rect 57422 282258 57464 282494
rect 57144 275494 57464 282258
rect 57144 275258 57186 275494
rect 57422 275258 57464 275494
rect 57144 268494 57464 275258
rect 57144 268258 57186 268494
rect 57422 268258 57464 268494
rect 57144 261494 57464 268258
rect 57144 261258 57186 261494
rect 57422 261258 57464 261494
rect 57144 254494 57464 261258
rect 57144 254258 57186 254494
rect 57422 254258 57464 254494
rect 57144 247494 57464 254258
rect 57144 247258 57186 247494
rect 57422 247258 57464 247494
rect 57144 240494 57464 247258
rect 57144 240258 57186 240494
rect 57422 240258 57464 240494
rect 57144 233494 57464 240258
rect 57144 233258 57186 233494
rect 57422 233258 57464 233494
rect 57144 226494 57464 233258
rect 57144 226258 57186 226494
rect 57422 226258 57464 226494
rect 57144 219494 57464 226258
rect 57144 219258 57186 219494
rect 57422 219258 57464 219494
rect 57144 212494 57464 219258
rect 57144 212258 57186 212494
rect 57422 212258 57464 212494
rect 57144 205494 57464 212258
rect 57144 205258 57186 205494
rect 57422 205258 57464 205494
rect 57144 198494 57464 205258
rect 57144 198258 57186 198494
rect 57422 198258 57464 198494
rect 57144 191494 57464 198258
rect 57144 191258 57186 191494
rect 57422 191258 57464 191494
rect 57144 184494 57464 191258
rect 57144 184258 57186 184494
rect 57422 184258 57464 184494
rect 57144 177494 57464 184258
rect 57144 177258 57186 177494
rect 57422 177258 57464 177494
rect 57144 170494 57464 177258
rect 57144 170258 57186 170494
rect 57422 170258 57464 170494
rect 57144 163494 57464 170258
rect 57144 163258 57186 163494
rect 57422 163258 57464 163494
rect 57144 156494 57464 163258
rect 57144 156258 57186 156494
rect 57422 156258 57464 156494
rect 57144 149494 57464 156258
rect 57144 149258 57186 149494
rect 57422 149258 57464 149494
rect 57144 142494 57464 149258
rect 57144 142258 57186 142494
rect 57422 142258 57464 142494
rect 57144 135494 57464 142258
rect 57144 135258 57186 135494
rect 57422 135258 57464 135494
rect 57144 128494 57464 135258
rect 57144 128258 57186 128494
rect 57422 128258 57464 128494
rect 57144 121494 57464 128258
rect 57144 121258 57186 121494
rect 57422 121258 57464 121494
rect 57144 114494 57464 121258
rect 57144 114258 57186 114494
rect 57422 114258 57464 114494
rect 57144 107494 57464 114258
rect 57144 107258 57186 107494
rect 57422 107258 57464 107494
rect 57144 100494 57464 107258
rect 57144 100258 57186 100494
rect 57422 100258 57464 100494
rect 57144 93494 57464 100258
rect 57144 93258 57186 93494
rect 57422 93258 57464 93494
rect 57144 86494 57464 93258
rect 57144 86258 57186 86494
rect 57422 86258 57464 86494
rect 57144 79494 57464 86258
rect 57144 79258 57186 79494
rect 57422 79258 57464 79494
rect 57144 72494 57464 79258
rect 57144 72258 57186 72494
rect 57422 72258 57464 72494
rect 57144 65494 57464 72258
rect 57144 65258 57186 65494
rect 57422 65258 57464 65494
rect 57144 58494 57464 65258
rect 57144 58258 57186 58494
rect 57422 58258 57464 58494
rect 57144 51494 57464 58258
rect 57144 51258 57186 51494
rect 57422 51258 57464 51494
rect 57144 44494 57464 51258
rect 57144 44258 57186 44494
rect 57422 44258 57464 44494
rect 57144 37494 57464 44258
rect 57144 37258 57186 37494
rect 57422 37258 57464 37494
rect 57144 30494 57464 37258
rect 57144 30258 57186 30494
rect 57422 30258 57464 30494
rect 57144 23494 57464 30258
rect 57144 23258 57186 23494
rect 57422 23258 57464 23494
rect 57144 16494 57464 23258
rect 57144 16258 57186 16494
rect 57422 16258 57464 16494
rect 57144 9494 57464 16258
rect 57144 9258 57186 9494
rect 57422 9258 57464 9494
rect 57144 2494 57464 9258
rect 57144 2258 57186 2494
rect 57422 2258 57464 2494
rect 57144 -746 57464 2258
rect 57144 -982 57186 -746
rect 57422 -982 57464 -746
rect 57144 -1066 57464 -982
rect 57144 -1302 57186 -1066
rect 57422 -1302 57464 -1066
rect 57144 -2294 57464 -1302
rect 58876 706198 59196 706230
rect 58876 705962 58918 706198
rect 59154 705962 59196 706198
rect 58876 705878 59196 705962
rect 58876 705642 58918 705878
rect 59154 705642 59196 705878
rect 58876 696434 59196 705642
rect 58876 696198 58918 696434
rect 59154 696198 59196 696434
rect 58876 689434 59196 696198
rect 58876 689198 58918 689434
rect 59154 689198 59196 689434
rect 58876 682434 59196 689198
rect 58876 682198 58918 682434
rect 59154 682198 59196 682434
rect 58876 675434 59196 682198
rect 58876 675198 58918 675434
rect 59154 675198 59196 675434
rect 58876 668434 59196 675198
rect 58876 668198 58918 668434
rect 59154 668198 59196 668434
rect 58876 661434 59196 668198
rect 58876 661198 58918 661434
rect 59154 661198 59196 661434
rect 58876 654434 59196 661198
rect 58876 654198 58918 654434
rect 59154 654198 59196 654434
rect 58876 647434 59196 654198
rect 58876 647198 58918 647434
rect 59154 647198 59196 647434
rect 58876 640434 59196 647198
rect 58876 640198 58918 640434
rect 59154 640198 59196 640434
rect 58876 633434 59196 640198
rect 58876 633198 58918 633434
rect 59154 633198 59196 633434
rect 58876 626434 59196 633198
rect 58876 626198 58918 626434
rect 59154 626198 59196 626434
rect 58876 619434 59196 626198
rect 58876 619198 58918 619434
rect 59154 619198 59196 619434
rect 58876 612434 59196 619198
rect 58876 612198 58918 612434
rect 59154 612198 59196 612434
rect 58876 605434 59196 612198
rect 58876 605198 58918 605434
rect 59154 605198 59196 605434
rect 58876 598434 59196 605198
rect 58876 598198 58918 598434
rect 59154 598198 59196 598434
rect 58876 591434 59196 598198
rect 58876 591198 58918 591434
rect 59154 591198 59196 591434
rect 58876 584434 59196 591198
rect 58876 584198 58918 584434
rect 59154 584198 59196 584434
rect 58876 577434 59196 584198
rect 58876 577198 58918 577434
rect 59154 577198 59196 577434
rect 58876 570434 59196 577198
rect 58876 570198 58918 570434
rect 59154 570198 59196 570434
rect 58876 563434 59196 570198
rect 58876 563198 58918 563434
rect 59154 563198 59196 563434
rect 58876 556434 59196 563198
rect 58876 556198 58918 556434
rect 59154 556198 59196 556434
rect 58876 549434 59196 556198
rect 58876 549198 58918 549434
rect 59154 549198 59196 549434
rect 58876 542434 59196 549198
rect 58876 542198 58918 542434
rect 59154 542198 59196 542434
rect 58876 535434 59196 542198
rect 58876 535198 58918 535434
rect 59154 535198 59196 535434
rect 58876 528434 59196 535198
rect 58876 528198 58918 528434
rect 59154 528198 59196 528434
rect 58876 521434 59196 528198
rect 58876 521198 58918 521434
rect 59154 521198 59196 521434
rect 58876 514434 59196 521198
rect 58876 514198 58918 514434
rect 59154 514198 59196 514434
rect 58876 507434 59196 514198
rect 58876 507198 58918 507434
rect 59154 507198 59196 507434
rect 58876 500434 59196 507198
rect 58876 500198 58918 500434
rect 59154 500198 59196 500434
rect 58876 493434 59196 500198
rect 58876 493198 58918 493434
rect 59154 493198 59196 493434
rect 58876 486434 59196 493198
rect 58876 486198 58918 486434
rect 59154 486198 59196 486434
rect 58876 479434 59196 486198
rect 58876 479198 58918 479434
rect 59154 479198 59196 479434
rect 58876 472434 59196 479198
rect 58876 472198 58918 472434
rect 59154 472198 59196 472434
rect 58876 465434 59196 472198
rect 58876 465198 58918 465434
rect 59154 465198 59196 465434
rect 58876 458434 59196 465198
rect 58876 458198 58918 458434
rect 59154 458198 59196 458434
rect 58876 451434 59196 458198
rect 58876 451198 58918 451434
rect 59154 451198 59196 451434
rect 58876 444434 59196 451198
rect 58876 444198 58918 444434
rect 59154 444198 59196 444434
rect 58876 437434 59196 444198
rect 58876 437198 58918 437434
rect 59154 437198 59196 437434
rect 58876 430434 59196 437198
rect 58876 430198 58918 430434
rect 59154 430198 59196 430434
rect 58876 423434 59196 430198
rect 58876 423198 58918 423434
rect 59154 423198 59196 423434
rect 58876 416434 59196 423198
rect 58876 416198 58918 416434
rect 59154 416198 59196 416434
rect 58876 409434 59196 416198
rect 58876 409198 58918 409434
rect 59154 409198 59196 409434
rect 58876 402434 59196 409198
rect 58876 402198 58918 402434
rect 59154 402198 59196 402434
rect 58876 395434 59196 402198
rect 58876 395198 58918 395434
rect 59154 395198 59196 395434
rect 58876 388434 59196 395198
rect 58876 388198 58918 388434
rect 59154 388198 59196 388434
rect 58876 381434 59196 388198
rect 58876 381198 58918 381434
rect 59154 381198 59196 381434
rect 58876 374434 59196 381198
rect 58876 374198 58918 374434
rect 59154 374198 59196 374434
rect 58876 367434 59196 374198
rect 58876 367198 58918 367434
rect 59154 367198 59196 367434
rect 58876 360434 59196 367198
rect 58876 360198 58918 360434
rect 59154 360198 59196 360434
rect 58876 353434 59196 360198
rect 58876 353198 58918 353434
rect 59154 353198 59196 353434
rect 58876 346434 59196 353198
rect 58876 346198 58918 346434
rect 59154 346198 59196 346434
rect 58876 339434 59196 346198
rect 58876 339198 58918 339434
rect 59154 339198 59196 339434
rect 58876 332434 59196 339198
rect 58876 332198 58918 332434
rect 59154 332198 59196 332434
rect 58876 325434 59196 332198
rect 58876 325198 58918 325434
rect 59154 325198 59196 325434
rect 58876 318434 59196 325198
rect 58876 318198 58918 318434
rect 59154 318198 59196 318434
rect 58876 311434 59196 318198
rect 58876 311198 58918 311434
rect 59154 311198 59196 311434
rect 58876 304434 59196 311198
rect 58876 304198 58918 304434
rect 59154 304198 59196 304434
rect 58876 297434 59196 304198
rect 58876 297198 58918 297434
rect 59154 297198 59196 297434
rect 58876 290434 59196 297198
rect 58876 290198 58918 290434
rect 59154 290198 59196 290434
rect 58876 283434 59196 290198
rect 58876 283198 58918 283434
rect 59154 283198 59196 283434
rect 58876 276434 59196 283198
rect 58876 276198 58918 276434
rect 59154 276198 59196 276434
rect 58876 269434 59196 276198
rect 58876 269198 58918 269434
rect 59154 269198 59196 269434
rect 58876 262434 59196 269198
rect 58876 262198 58918 262434
rect 59154 262198 59196 262434
rect 58876 255434 59196 262198
rect 58876 255198 58918 255434
rect 59154 255198 59196 255434
rect 58876 248434 59196 255198
rect 58876 248198 58918 248434
rect 59154 248198 59196 248434
rect 58876 241434 59196 248198
rect 58876 241198 58918 241434
rect 59154 241198 59196 241434
rect 58876 234434 59196 241198
rect 58876 234198 58918 234434
rect 59154 234198 59196 234434
rect 58876 227434 59196 234198
rect 58876 227198 58918 227434
rect 59154 227198 59196 227434
rect 58876 220434 59196 227198
rect 58876 220198 58918 220434
rect 59154 220198 59196 220434
rect 58876 213434 59196 220198
rect 58876 213198 58918 213434
rect 59154 213198 59196 213434
rect 58876 206434 59196 213198
rect 58876 206198 58918 206434
rect 59154 206198 59196 206434
rect 58876 199434 59196 206198
rect 58876 199198 58918 199434
rect 59154 199198 59196 199434
rect 58876 192434 59196 199198
rect 58876 192198 58918 192434
rect 59154 192198 59196 192434
rect 58876 185434 59196 192198
rect 58876 185198 58918 185434
rect 59154 185198 59196 185434
rect 58876 178434 59196 185198
rect 58876 178198 58918 178434
rect 59154 178198 59196 178434
rect 58876 171434 59196 178198
rect 58876 171198 58918 171434
rect 59154 171198 59196 171434
rect 58876 164434 59196 171198
rect 58876 164198 58918 164434
rect 59154 164198 59196 164434
rect 58876 157434 59196 164198
rect 58876 157198 58918 157434
rect 59154 157198 59196 157434
rect 58876 150434 59196 157198
rect 58876 150198 58918 150434
rect 59154 150198 59196 150434
rect 58876 143434 59196 150198
rect 58876 143198 58918 143434
rect 59154 143198 59196 143434
rect 58876 136434 59196 143198
rect 58876 136198 58918 136434
rect 59154 136198 59196 136434
rect 58876 129434 59196 136198
rect 58876 129198 58918 129434
rect 59154 129198 59196 129434
rect 58876 122434 59196 129198
rect 58876 122198 58918 122434
rect 59154 122198 59196 122434
rect 58876 115434 59196 122198
rect 58876 115198 58918 115434
rect 59154 115198 59196 115434
rect 58876 108434 59196 115198
rect 58876 108198 58918 108434
rect 59154 108198 59196 108434
rect 58876 101434 59196 108198
rect 58876 101198 58918 101434
rect 59154 101198 59196 101434
rect 58876 94434 59196 101198
rect 58876 94198 58918 94434
rect 59154 94198 59196 94434
rect 58876 87434 59196 94198
rect 58876 87198 58918 87434
rect 59154 87198 59196 87434
rect 58876 80434 59196 87198
rect 58876 80198 58918 80434
rect 59154 80198 59196 80434
rect 58876 73434 59196 80198
rect 58876 73198 58918 73434
rect 59154 73198 59196 73434
rect 58876 66434 59196 73198
rect 58876 66198 58918 66434
rect 59154 66198 59196 66434
rect 58876 59434 59196 66198
rect 58876 59198 58918 59434
rect 59154 59198 59196 59434
rect 58876 52434 59196 59198
rect 58876 52198 58918 52434
rect 59154 52198 59196 52434
rect 58876 45434 59196 52198
rect 58876 45198 58918 45434
rect 59154 45198 59196 45434
rect 58876 38434 59196 45198
rect 58876 38198 58918 38434
rect 59154 38198 59196 38434
rect 58876 31434 59196 38198
rect 58876 31198 58918 31434
rect 59154 31198 59196 31434
rect 58876 24434 59196 31198
rect 58876 24198 58918 24434
rect 59154 24198 59196 24434
rect 58876 17434 59196 24198
rect 58876 17198 58918 17434
rect 59154 17198 59196 17434
rect 58876 10434 59196 17198
rect 58876 10198 58918 10434
rect 59154 10198 59196 10434
rect 58876 3434 59196 10198
rect 58876 3198 58918 3434
rect 59154 3198 59196 3434
rect 58876 -1706 59196 3198
rect 58876 -1942 58918 -1706
rect 59154 -1942 59196 -1706
rect 58876 -2026 59196 -1942
rect 58876 -2262 58918 -2026
rect 59154 -2262 59196 -2026
rect 58876 -2294 59196 -2262
rect 64144 705238 64464 706230
rect 64144 705002 64186 705238
rect 64422 705002 64464 705238
rect 64144 704918 64464 705002
rect 64144 704682 64186 704918
rect 64422 704682 64464 704918
rect 64144 695494 64464 704682
rect 64144 695258 64186 695494
rect 64422 695258 64464 695494
rect 64144 688494 64464 695258
rect 64144 688258 64186 688494
rect 64422 688258 64464 688494
rect 64144 681494 64464 688258
rect 64144 681258 64186 681494
rect 64422 681258 64464 681494
rect 64144 674494 64464 681258
rect 64144 674258 64186 674494
rect 64422 674258 64464 674494
rect 64144 667494 64464 674258
rect 64144 667258 64186 667494
rect 64422 667258 64464 667494
rect 64144 660494 64464 667258
rect 64144 660258 64186 660494
rect 64422 660258 64464 660494
rect 64144 653494 64464 660258
rect 64144 653258 64186 653494
rect 64422 653258 64464 653494
rect 64144 646494 64464 653258
rect 64144 646258 64186 646494
rect 64422 646258 64464 646494
rect 64144 639494 64464 646258
rect 64144 639258 64186 639494
rect 64422 639258 64464 639494
rect 64144 632494 64464 639258
rect 64144 632258 64186 632494
rect 64422 632258 64464 632494
rect 64144 625494 64464 632258
rect 64144 625258 64186 625494
rect 64422 625258 64464 625494
rect 64144 618494 64464 625258
rect 64144 618258 64186 618494
rect 64422 618258 64464 618494
rect 64144 611494 64464 618258
rect 64144 611258 64186 611494
rect 64422 611258 64464 611494
rect 64144 604494 64464 611258
rect 64144 604258 64186 604494
rect 64422 604258 64464 604494
rect 64144 597494 64464 604258
rect 64144 597258 64186 597494
rect 64422 597258 64464 597494
rect 64144 590494 64464 597258
rect 64144 590258 64186 590494
rect 64422 590258 64464 590494
rect 64144 583494 64464 590258
rect 64144 583258 64186 583494
rect 64422 583258 64464 583494
rect 64144 576494 64464 583258
rect 64144 576258 64186 576494
rect 64422 576258 64464 576494
rect 64144 569494 64464 576258
rect 64144 569258 64186 569494
rect 64422 569258 64464 569494
rect 64144 562494 64464 569258
rect 64144 562258 64186 562494
rect 64422 562258 64464 562494
rect 64144 555494 64464 562258
rect 64144 555258 64186 555494
rect 64422 555258 64464 555494
rect 64144 548494 64464 555258
rect 64144 548258 64186 548494
rect 64422 548258 64464 548494
rect 64144 541494 64464 548258
rect 64144 541258 64186 541494
rect 64422 541258 64464 541494
rect 64144 534494 64464 541258
rect 64144 534258 64186 534494
rect 64422 534258 64464 534494
rect 64144 527494 64464 534258
rect 64144 527258 64186 527494
rect 64422 527258 64464 527494
rect 64144 520494 64464 527258
rect 64144 520258 64186 520494
rect 64422 520258 64464 520494
rect 64144 513494 64464 520258
rect 64144 513258 64186 513494
rect 64422 513258 64464 513494
rect 64144 506494 64464 513258
rect 64144 506258 64186 506494
rect 64422 506258 64464 506494
rect 64144 499494 64464 506258
rect 64144 499258 64186 499494
rect 64422 499258 64464 499494
rect 64144 492494 64464 499258
rect 64144 492258 64186 492494
rect 64422 492258 64464 492494
rect 64144 485494 64464 492258
rect 64144 485258 64186 485494
rect 64422 485258 64464 485494
rect 64144 478494 64464 485258
rect 64144 478258 64186 478494
rect 64422 478258 64464 478494
rect 64144 471494 64464 478258
rect 64144 471258 64186 471494
rect 64422 471258 64464 471494
rect 64144 464494 64464 471258
rect 64144 464258 64186 464494
rect 64422 464258 64464 464494
rect 64144 457494 64464 464258
rect 64144 457258 64186 457494
rect 64422 457258 64464 457494
rect 64144 450494 64464 457258
rect 64144 450258 64186 450494
rect 64422 450258 64464 450494
rect 64144 443494 64464 450258
rect 64144 443258 64186 443494
rect 64422 443258 64464 443494
rect 64144 436494 64464 443258
rect 64144 436258 64186 436494
rect 64422 436258 64464 436494
rect 64144 429494 64464 436258
rect 64144 429258 64186 429494
rect 64422 429258 64464 429494
rect 64144 422494 64464 429258
rect 64144 422258 64186 422494
rect 64422 422258 64464 422494
rect 64144 415494 64464 422258
rect 64144 415258 64186 415494
rect 64422 415258 64464 415494
rect 64144 408494 64464 415258
rect 64144 408258 64186 408494
rect 64422 408258 64464 408494
rect 64144 401494 64464 408258
rect 64144 401258 64186 401494
rect 64422 401258 64464 401494
rect 64144 394494 64464 401258
rect 64144 394258 64186 394494
rect 64422 394258 64464 394494
rect 64144 387494 64464 394258
rect 64144 387258 64186 387494
rect 64422 387258 64464 387494
rect 64144 380494 64464 387258
rect 64144 380258 64186 380494
rect 64422 380258 64464 380494
rect 64144 373494 64464 380258
rect 64144 373258 64186 373494
rect 64422 373258 64464 373494
rect 64144 366494 64464 373258
rect 64144 366258 64186 366494
rect 64422 366258 64464 366494
rect 64144 359494 64464 366258
rect 64144 359258 64186 359494
rect 64422 359258 64464 359494
rect 64144 352494 64464 359258
rect 64144 352258 64186 352494
rect 64422 352258 64464 352494
rect 64144 345494 64464 352258
rect 64144 345258 64186 345494
rect 64422 345258 64464 345494
rect 64144 338494 64464 345258
rect 64144 338258 64186 338494
rect 64422 338258 64464 338494
rect 64144 331494 64464 338258
rect 64144 331258 64186 331494
rect 64422 331258 64464 331494
rect 64144 324494 64464 331258
rect 64144 324258 64186 324494
rect 64422 324258 64464 324494
rect 64144 317494 64464 324258
rect 64144 317258 64186 317494
rect 64422 317258 64464 317494
rect 64144 310494 64464 317258
rect 64144 310258 64186 310494
rect 64422 310258 64464 310494
rect 64144 303494 64464 310258
rect 64144 303258 64186 303494
rect 64422 303258 64464 303494
rect 64144 296494 64464 303258
rect 64144 296258 64186 296494
rect 64422 296258 64464 296494
rect 64144 289494 64464 296258
rect 64144 289258 64186 289494
rect 64422 289258 64464 289494
rect 64144 282494 64464 289258
rect 64144 282258 64186 282494
rect 64422 282258 64464 282494
rect 64144 275494 64464 282258
rect 64144 275258 64186 275494
rect 64422 275258 64464 275494
rect 64144 268494 64464 275258
rect 64144 268258 64186 268494
rect 64422 268258 64464 268494
rect 64144 261494 64464 268258
rect 64144 261258 64186 261494
rect 64422 261258 64464 261494
rect 64144 254494 64464 261258
rect 64144 254258 64186 254494
rect 64422 254258 64464 254494
rect 64144 247494 64464 254258
rect 64144 247258 64186 247494
rect 64422 247258 64464 247494
rect 64144 240494 64464 247258
rect 64144 240258 64186 240494
rect 64422 240258 64464 240494
rect 64144 233494 64464 240258
rect 64144 233258 64186 233494
rect 64422 233258 64464 233494
rect 64144 226494 64464 233258
rect 64144 226258 64186 226494
rect 64422 226258 64464 226494
rect 64144 219494 64464 226258
rect 64144 219258 64186 219494
rect 64422 219258 64464 219494
rect 64144 212494 64464 219258
rect 64144 212258 64186 212494
rect 64422 212258 64464 212494
rect 64144 205494 64464 212258
rect 64144 205258 64186 205494
rect 64422 205258 64464 205494
rect 64144 198494 64464 205258
rect 64144 198258 64186 198494
rect 64422 198258 64464 198494
rect 64144 191494 64464 198258
rect 64144 191258 64186 191494
rect 64422 191258 64464 191494
rect 64144 184494 64464 191258
rect 64144 184258 64186 184494
rect 64422 184258 64464 184494
rect 64144 177494 64464 184258
rect 64144 177258 64186 177494
rect 64422 177258 64464 177494
rect 64144 170494 64464 177258
rect 64144 170258 64186 170494
rect 64422 170258 64464 170494
rect 64144 163494 64464 170258
rect 64144 163258 64186 163494
rect 64422 163258 64464 163494
rect 64144 156494 64464 163258
rect 64144 156258 64186 156494
rect 64422 156258 64464 156494
rect 64144 149494 64464 156258
rect 64144 149258 64186 149494
rect 64422 149258 64464 149494
rect 64144 142494 64464 149258
rect 64144 142258 64186 142494
rect 64422 142258 64464 142494
rect 64144 135494 64464 142258
rect 64144 135258 64186 135494
rect 64422 135258 64464 135494
rect 64144 128494 64464 135258
rect 64144 128258 64186 128494
rect 64422 128258 64464 128494
rect 64144 121494 64464 128258
rect 64144 121258 64186 121494
rect 64422 121258 64464 121494
rect 64144 114494 64464 121258
rect 64144 114258 64186 114494
rect 64422 114258 64464 114494
rect 64144 107494 64464 114258
rect 64144 107258 64186 107494
rect 64422 107258 64464 107494
rect 64144 100494 64464 107258
rect 64144 100258 64186 100494
rect 64422 100258 64464 100494
rect 64144 93494 64464 100258
rect 64144 93258 64186 93494
rect 64422 93258 64464 93494
rect 64144 86494 64464 93258
rect 64144 86258 64186 86494
rect 64422 86258 64464 86494
rect 64144 79494 64464 86258
rect 64144 79258 64186 79494
rect 64422 79258 64464 79494
rect 64144 72494 64464 79258
rect 64144 72258 64186 72494
rect 64422 72258 64464 72494
rect 64144 65494 64464 72258
rect 64144 65258 64186 65494
rect 64422 65258 64464 65494
rect 64144 58494 64464 65258
rect 64144 58258 64186 58494
rect 64422 58258 64464 58494
rect 64144 51494 64464 58258
rect 64144 51258 64186 51494
rect 64422 51258 64464 51494
rect 64144 44494 64464 51258
rect 64144 44258 64186 44494
rect 64422 44258 64464 44494
rect 64144 37494 64464 44258
rect 64144 37258 64186 37494
rect 64422 37258 64464 37494
rect 64144 30494 64464 37258
rect 64144 30258 64186 30494
rect 64422 30258 64464 30494
rect 64144 23494 64464 30258
rect 64144 23258 64186 23494
rect 64422 23258 64464 23494
rect 64144 16494 64464 23258
rect 64144 16258 64186 16494
rect 64422 16258 64464 16494
rect 64144 9494 64464 16258
rect 64144 9258 64186 9494
rect 64422 9258 64464 9494
rect 64144 2494 64464 9258
rect 64144 2258 64186 2494
rect 64422 2258 64464 2494
rect 64144 -746 64464 2258
rect 64144 -982 64186 -746
rect 64422 -982 64464 -746
rect 64144 -1066 64464 -982
rect 64144 -1302 64186 -1066
rect 64422 -1302 64464 -1066
rect 64144 -2294 64464 -1302
rect 65876 706198 66196 706230
rect 65876 705962 65918 706198
rect 66154 705962 66196 706198
rect 65876 705878 66196 705962
rect 65876 705642 65918 705878
rect 66154 705642 66196 705878
rect 65876 696434 66196 705642
rect 65876 696198 65918 696434
rect 66154 696198 66196 696434
rect 65876 689434 66196 696198
rect 65876 689198 65918 689434
rect 66154 689198 66196 689434
rect 65876 682434 66196 689198
rect 65876 682198 65918 682434
rect 66154 682198 66196 682434
rect 65876 675434 66196 682198
rect 65876 675198 65918 675434
rect 66154 675198 66196 675434
rect 65876 668434 66196 675198
rect 65876 668198 65918 668434
rect 66154 668198 66196 668434
rect 65876 661434 66196 668198
rect 65876 661198 65918 661434
rect 66154 661198 66196 661434
rect 65876 654434 66196 661198
rect 65876 654198 65918 654434
rect 66154 654198 66196 654434
rect 65876 647434 66196 654198
rect 65876 647198 65918 647434
rect 66154 647198 66196 647434
rect 65876 640434 66196 647198
rect 65876 640198 65918 640434
rect 66154 640198 66196 640434
rect 65876 633434 66196 640198
rect 65876 633198 65918 633434
rect 66154 633198 66196 633434
rect 65876 626434 66196 633198
rect 65876 626198 65918 626434
rect 66154 626198 66196 626434
rect 65876 619434 66196 626198
rect 65876 619198 65918 619434
rect 66154 619198 66196 619434
rect 65876 612434 66196 619198
rect 65876 612198 65918 612434
rect 66154 612198 66196 612434
rect 65876 605434 66196 612198
rect 65876 605198 65918 605434
rect 66154 605198 66196 605434
rect 65876 598434 66196 605198
rect 65876 598198 65918 598434
rect 66154 598198 66196 598434
rect 65876 591434 66196 598198
rect 65876 591198 65918 591434
rect 66154 591198 66196 591434
rect 65876 584434 66196 591198
rect 65876 584198 65918 584434
rect 66154 584198 66196 584434
rect 65876 577434 66196 584198
rect 65876 577198 65918 577434
rect 66154 577198 66196 577434
rect 65876 570434 66196 577198
rect 65876 570198 65918 570434
rect 66154 570198 66196 570434
rect 65876 563434 66196 570198
rect 65876 563198 65918 563434
rect 66154 563198 66196 563434
rect 65876 556434 66196 563198
rect 65876 556198 65918 556434
rect 66154 556198 66196 556434
rect 65876 549434 66196 556198
rect 65876 549198 65918 549434
rect 66154 549198 66196 549434
rect 65876 542434 66196 549198
rect 65876 542198 65918 542434
rect 66154 542198 66196 542434
rect 65876 535434 66196 542198
rect 65876 535198 65918 535434
rect 66154 535198 66196 535434
rect 65876 528434 66196 535198
rect 65876 528198 65918 528434
rect 66154 528198 66196 528434
rect 65876 521434 66196 528198
rect 65876 521198 65918 521434
rect 66154 521198 66196 521434
rect 65876 514434 66196 521198
rect 65876 514198 65918 514434
rect 66154 514198 66196 514434
rect 65876 507434 66196 514198
rect 65876 507198 65918 507434
rect 66154 507198 66196 507434
rect 65876 500434 66196 507198
rect 65876 500198 65918 500434
rect 66154 500198 66196 500434
rect 65876 493434 66196 500198
rect 65876 493198 65918 493434
rect 66154 493198 66196 493434
rect 65876 486434 66196 493198
rect 65876 486198 65918 486434
rect 66154 486198 66196 486434
rect 65876 479434 66196 486198
rect 65876 479198 65918 479434
rect 66154 479198 66196 479434
rect 65876 472434 66196 479198
rect 65876 472198 65918 472434
rect 66154 472198 66196 472434
rect 65876 465434 66196 472198
rect 65876 465198 65918 465434
rect 66154 465198 66196 465434
rect 65876 458434 66196 465198
rect 65876 458198 65918 458434
rect 66154 458198 66196 458434
rect 65876 451434 66196 458198
rect 65876 451198 65918 451434
rect 66154 451198 66196 451434
rect 65876 444434 66196 451198
rect 65876 444198 65918 444434
rect 66154 444198 66196 444434
rect 65876 437434 66196 444198
rect 65876 437198 65918 437434
rect 66154 437198 66196 437434
rect 65876 430434 66196 437198
rect 65876 430198 65918 430434
rect 66154 430198 66196 430434
rect 65876 423434 66196 430198
rect 65876 423198 65918 423434
rect 66154 423198 66196 423434
rect 65876 416434 66196 423198
rect 65876 416198 65918 416434
rect 66154 416198 66196 416434
rect 65876 409434 66196 416198
rect 65876 409198 65918 409434
rect 66154 409198 66196 409434
rect 65876 402434 66196 409198
rect 65876 402198 65918 402434
rect 66154 402198 66196 402434
rect 65876 395434 66196 402198
rect 65876 395198 65918 395434
rect 66154 395198 66196 395434
rect 65876 388434 66196 395198
rect 65876 388198 65918 388434
rect 66154 388198 66196 388434
rect 65876 381434 66196 388198
rect 65876 381198 65918 381434
rect 66154 381198 66196 381434
rect 65876 374434 66196 381198
rect 65876 374198 65918 374434
rect 66154 374198 66196 374434
rect 65876 367434 66196 374198
rect 65876 367198 65918 367434
rect 66154 367198 66196 367434
rect 65876 360434 66196 367198
rect 65876 360198 65918 360434
rect 66154 360198 66196 360434
rect 65876 353434 66196 360198
rect 65876 353198 65918 353434
rect 66154 353198 66196 353434
rect 65876 346434 66196 353198
rect 65876 346198 65918 346434
rect 66154 346198 66196 346434
rect 65876 339434 66196 346198
rect 65876 339198 65918 339434
rect 66154 339198 66196 339434
rect 65876 332434 66196 339198
rect 65876 332198 65918 332434
rect 66154 332198 66196 332434
rect 65876 325434 66196 332198
rect 65876 325198 65918 325434
rect 66154 325198 66196 325434
rect 65876 318434 66196 325198
rect 65876 318198 65918 318434
rect 66154 318198 66196 318434
rect 65876 311434 66196 318198
rect 65876 311198 65918 311434
rect 66154 311198 66196 311434
rect 65876 304434 66196 311198
rect 65876 304198 65918 304434
rect 66154 304198 66196 304434
rect 65876 297434 66196 304198
rect 65876 297198 65918 297434
rect 66154 297198 66196 297434
rect 65876 290434 66196 297198
rect 65876 290198 65918 290434
rect 66154 290198 66196 290434
rect 65876 283434 66196 290198
rect 65876 283198 65918 283434
rect 66154 283198 66196 283434
rect 65876 276434 66196 283198
rect 65876 276198 65918 276434
rect 66154 276198 66196 276434
rect 65876 269434 66196 276198
rect 65876 269198 65918 269434
rect 66154 269198 66196 269434
rect 65876 262434 66196 269198
rect 65876 262198 65918 262434
rect 66154 262198 66196 262434
rect 65876 255434 66196 262198
rect 65876 255198 65918 255434
rect 66154 255198 66196 255434
rect 65876 248434 66196 255198
rect 65876 248198 65918 248434
rect 66154 248198 66196 248434
rect 65876 241434 66196 248198
rect 65876 241198 65918 241434
rect 66154 241198 66196 241434
rect 65876 234434 66196 241198
rect 65876 234198 65918 234434
rect 66154 234198 66196 234434
rect 65876 227434 66196 234198
rect 65876 227198 65918 227434
rect 66154 227198 66196 227434
rect 65876 220434 66196 227198
rect 65876 220198 65918 220434
rect 66154 220198 66196 220434
rect 65876 213434 66196 220198
rect 65876 213198 65918 213434
rect 66154 213198 66196 213434
rect 65876 206434 66196 213198
rect 65876 206198 65918 206434
rect 66154 206198 66196 206434
rect 65876 199434 66196 206198
rect 65876 199198 65918 199434
rect 66154 199198 66196 199434
rect 65876 192434 66196 199198
rect 65876 192198 65918 192434
rect 66154 192198 66196 192434
rect 65876 185434 66196 192198
rect 65876 185198 65918 185434
rect 66154 185198 66196 185434
rect 65876 178434 66196 185198
rect 65876 178198 65918 178434
rect 66154 178198 66196 178434
rect 65876 171434 66196 178198
rect 65876 171198 65918 171434
rect 66154 171198 66196 171434
rect 65876 164434 66196 171198
rect 65876 164198 65918 164434
rect 66154 164198 66196 164434
rect 65876 157434 66196 164198
rect 65876 157198 65918 157434
rect 66154 157198 66196 157434
rect 65876 150434 66196 157198
rect 65876 150198 65918 150434
rect 66154 150198 66196 150434
rect 65876 143434 66196 150198
rect 65876 143198 65918 143434
rect 66154 143198 66196 143434
rect 65876 136434 66196 143198
rect 65876 136198 65918 136434
rect 66154 136198 66196 136434
rect 65876 129434 66196 136198
rect 65876 129198 65918 129434
rect 66154 129198 66196 129434
rect 65876 122434 66196 129198
rect 65876 122198 65918 122434
rect 66154 122198 66196 122434
rect 65876 115434 66196 122198
rect 65876 115198 65918 115434
rect 66154 115198 66196 115434
rect 65876 108434 66196 115198
rect 65876 108198 65918 108434
rect 66154 108198 66196 108434
rect 65876 101434 66196 108198
rect 65876 101198 65918 101434
rect 66154 101198 66196 101434
rect 65876 94434 66196 101198
rect 65876 94198 65918 94434
rect 66154 94198 66196 94434
rect 65876 87434 66196 94198
rect 65876 87198 65918 87434
rect 66154 87198 66196 87434
rect 65876 80434 66196 87198
rect 65876 80198 65918 80434
rect 66154 80198 66196 80434
rect 65876 73434 66196 80198
rect 65876 73198 65918 73434
rect 66154 73198 66196 73434
rect 65876 66434 66196 73198
rect 65876 66198 65918 66434
rect 66154 66198 66196 66434
rect 65876 59434 66196 66198
rect 65876 59198 65918 59434
rect 66154 59198 66196 59434
rect 65876 52434 66196 59198
rect 65876 52198 65918 52434
rect 66154 52198 66196 52434
rect 65876 45434 66196 52198
rect 65876 45198 65918 45434
rect 66154 45198 66196 45434
rect 65876 38434 66196 45198
rect 65876 38198 65918 38434
rect 66154 38198 66196 38434
rect 65876 31434 66196 38198
rect 65876 31198 65918 31434
rect 66154 31198 66196 31434
rect 65876 24434 66196 31198
rect 65876 24198 65918 24434
rect 66154 24198 66196 24434
rect 65876 17434 66196 24198
rect 65876 17198 65918 17434
rect 66154 17198 66196 17434
rect 65876 10434 66196 17198
rect 65876 10198 65918 10434
rect 66154 10198 66196 10434
rect 65876 3434 66196 10198
rect 65876 3198 65918 3434
rect 66154 3198 66196 3434
rect 65876 -1706 66196 3198
rect 65876 -1942 65918 -1706
rect 66154 -1942 66196 -1706
rect 65876 -2026 66196 -1942
rect 65876 -2262 65918 -2026
rect 66154 -2262 66196 -2026
rect 65876 -2294 66196 -2262
rect 71144 705238 71464 706230
rect 71144 705002 71186 705238
rect 71422 705002 71464 705238
rect 71144 704918 71464 705002
rect 71144 704682 71186 704918
rect 71422 704682 71464 704918
rect 71144 695494 71464 704682
rect 71144 695258 71186 695494
rect 71422 695258 71464 695494
rect 71144 688494 71464 695258
rect 71144 688258 71186 688494
rect 71422 688258 71464 688494
rect 71144 681494 71464 688258
rect 71144 681258 71186 681494
rect 71422 681258 71464 681494
rect 71144 674494 71464 681258
rect 71144 674258 71186 674494
rect 71422 674258 71464 674494
rect 71144 667494 71464 674258
rect 71144 667258 71186 667494
rect 71422 667258 71464 667494
rect 71144 660494 71464 667258
rect 71144 660258 71186 660494
rect 71422 660258 71464 660494
rect 71144 653494 71464 660258
rect 71144 653258 71186 653494
rect 71422 653258 71464 653494
rect 71144 646494 71464 653258
rect 71144 646258 71186 646494
rect 71422 646258 71464 646494
rect 71144 639494 71464 646258
rect 71144 639258 71186 639494
rect 71422 639258 71464 639494
rect 71144 632494 71464 639258
rect 71144 632258 71186 632494
rect 71422 632258 71464 632494
rect 71144 625494 71464 632258
rect 71144 625258 71186 625494
rect 71422 625258 71464 625494
rect 71144 618494 71464 625258
rect 71144 618258 71186 618494
rect 71422 618258 71464 618494
rect 71144 611494 71464 618258
rect 71144 611258 71186 611494
rect 71422 611258 71464 611494
rect 71144 604494 71464 611258
rect 71144 604258 71186 604494
rect 71422 604258 71464 604494
rect 71144 597494 71464 604258
rect 71144 597258 71186 597494
rect 71422 597258 71464 597494
rect 71144 590494 71464 597258
rect 71144 590258 71186 590494
rect 71422 590258 71464 590494
rect 71144 583494 71464 590258
rect 71144 583258 71186 583494
rect 71422 583258 71464 583494
rect 71144 576494 71464 583258
rect 71144 576258 71186 576494
rect 71422 576258 71464 576494
rect 71144 569494 71464 576258
rect 71144 569258 71186 569494
rect 71422 569258 71464 569494
rect 71144 562494 71464 569258
rect 71144 562258 71186 562494
rect 71422 562258 71464 562494
rect 71144 555494 71464 562258
rect 71144 555258 71186 555494
rect 71422 555258 71464 555494
rect 71144 548494 71464 555258
rect 71144 548258 71186 548494
rect 71422 548258 71464 548494
rect 71144 541494 71464 548258
rect 71144 541258 71186 541494
rect 71422 541258 71464 541494
rect 71144 534494 71464 541258
rect 71144 534258 71186 534494
rect 71422 534258 71464 534494
rect 71144 527494 71464 534258
rect 71144 527258 71186 527494
rect 71422 527258 71464 527494
rect 71144 520494 71464 527258
rect 71144 520258 71186 520494
rect 71422 520258 71464 520494
rect 71144 513494 71464 520258
rect 71144 513258 71186 513494
rect 71422 513258 71464 513494
rect 71144 506494 71464 513258
rect 71144 506258 71186 506494
rect 71422 506258 71464 506494
rect 71144 499494 71464 506258
rect 71144 499258 71186 499494
rect 71422 499258 71464 499494
rect 71144 492494 71464 499258
rect 71144 492258 71186 492494
rect 71422 492258 71464 492494
rect 71144 485494 71464 492258
rect 71144 485258 71186 485494
rect 71422 485258 71464 485494
rect 71144 478494 71464 485258
rect 71144 478258 71186 478494
rect 71422 478258 71464 478494
rect 71144 471494 71464 478258
rect 71144 471258 71186 471494
rect 71422 471258 71464 471494
rect 71144 464494 71464 471258
rect 71144 464258 71186 464494
rect 71422 464258 71464 464494
rect 71144 457494 71464 464258
rect 71144 457258 71186 457494
rect 71422 457258 71464 457494
rect 71144 450494 71464 457258
rect 71144 450258 71186 450494
rect 71422 450258 71464 450494
rect 71144 443494 71464 450258
rect 71144 443258 71186 443494
rect 71422 443258 71464 443494
rect 71144 436494 71464 443258
rect 71144 436258 71186 436494
rect 71422 436258 71464 436494
rect 71144 429494 71464 436258
rect 71144 429258 71186 429494
rect 71422 429258 71464 429494
rect 71144 422494 71464 429258
rect 71144 422258 71186 422494
rect 71422 422258 71464 422494
rect 71144 415494 71464 422258
rect 71144 415258 71186 415494
rect 71422 415258 71464 415494
rect 71144 408494 71464 415258
rect 71144 408258 71186 408494
rect 71422 408258 71464 408494
rect 71144 401494 71464 408258
rect 71144 401258 71186 401494
rect 71422 401258 71464 401494
rect 71144 394494 71464 401258
rect 71144 394258 71186 394494
rect 71422 394258 71464 394494
rect 71144 387494 71464 394258
rect 71144 387258 71186 387494
rect 71422 387258 71464 387494
rect 71144 380494 71464 387258
rect 71144 380258 71186 380494
rect 71422 380258 71464 380494
rect 71144 373494 71464 380258
rect 71144 373258 71186 373494
rect 71422 373258 71464 373494
rect 71144 366494 71464 373258
rect 71144 366258 71186 366494
rect 71422 366258 71464 366494
rect 71144 359494 71464 366258
rect 71144 359258 71186 359494
rect 71422 359258 71464 359494
rect 71144 352494 71464 359258
rect 71144 352258 71186 352494
rect 71422 352258 71464 352494
rect 71144 345494 71464 352258
rect 71144 345258 71186 345494
rect 71422 345258 71464 345494
rect 71144 338494 71464 345258
rect 71144 338258 71186 338494
rect 71422 338258 71464 338494
rect 71144 331494 71464 338258
rect 71144 331258 71186 331494
rect 71422 331258 71464 331494
rect 71144 324494 71464 331258
rect 71144 324258 71186 324494
rect 71422 324258 71464 324494
rect 71144 317494 71464 324258
rect 71144 317258 71186 317494
rect 71422 317258 71464 317494
rect 71144 310494 71464 317258
rect 71144 310258 71186 310494
rect 71422 310258 71464 310494
rect 71144 303494 71464 310258
rect 71144 303258 71186 303494
rect 71422 303258 71464 303494
rect 71144 296494 71464 303258
rect 71144 296258 71186 296494
rect 71422 296258 71464 296494
rect 71144 289494 71464 296258
rect 71144 289258 71186 289494
rect 71422 289258 71464 289494
rect 71144 282494 71464 289258
rect 71144 282258 71186 282494
rect 71422 282258 71464 282494
rect 71144 275494 71464 282258
rect 71144 275258 71186 275494
rect 71422 275258 71464 275494
rect 71144 268494 71464 275258
rect 71144 268258 71186 268494
rect 71422 268258 71464 268494
rect 71144 261494 71464 268258
rect 71144 261258 71186 261494
rect 71422 261258 71464 261494
rect 71144 254494 71464 261258
rect 71144 254258 71186 254494
rect 71422 254258 71464 254494
rect 71144 247494 71464 254258
rect 71144 247258 71186 247494
rect 71422 247258 71464 247494
rect 71144 240494 71464 247258
rect 71144 240258 71186 240494
rect 71422 240258 71464 240494
rect 71144 233494 71464 240258
rect 71144 233258 71186 233494
rect 71422 233258 71464 233494
rect 71144 226494 71464 233258
rect 71144 226258 71186 226494
rect 71422 226258 71464 226494
rect 71144 219494 71464 226258
rect 71144 219258 71186 219494
rect 71422 219258 71464 219494
rect 71144 212494 71464 219258
rect 71144 212258 71186 212494
rect 71422 212258 71464 212494
rect 71144 205494 71464 212258
rect 71144 205258 71186 205494
rect 71422 205258 71464 205494
rect 71144 198494 71464 205258
rect 71144 198258 71186 198494
rect 71422 198258 71464 198494
rect 71144 191494 71464 198258
rect 71144 191258 71186 191494
rect 71422 191258 71464 191494
rect 71144 184494 71464 191258
rect 71144 184258 71186 184494
rect 71422 184258 71464 184494
rect 71144 177494 71464 184258
rect 71144 177258 71186 177494
rect 71422 177258 71464 177494
rect 71144 170494 71464 177258
rect 71144 170258 71186 170494
rect 71422 170258 71464 170494
rect 71144 163494 71464 170258
rect 71144 163258 71186 163494
rect 71422 163258 71464 163494
rect 71144 156494 71464 163258
rect 71144 156258 71186 156494
rect 71422 156258 71464 156494
rect 71144 149494 71464 156258
rect 71144 149258 71186 149494
rect 71422 149258 71464 149494
rect 71144 142494 71464 149258
rect 71144 142258 71186 142494
rect 71422 142258 71464 142494
rect 71144 135494 71464 142258
rect 71144 135258 71186 135494
rect 71422 135258 71464 135494
rect 71144 128494 71464 135258
rect 71144 128258 71186 128494
rect 71422 128258 71464 128494
rect 71144 121494 71464 128258
rect 71144 121258 71186 121494
rect 71422 121258 71464 121494
rect 71144 114494 71464 121258
rect 71144 114258 71186 114494
rect 71422 114258 71464 114494
rect 71144 107494 71464 114258
rect 71144 107258 71186 107494
rect 71422 107258 71464 107494
rect 71144 100494 71464 107258
rect 71144 100258 71186 100494
rect 71422 100258 71464 100494
rect 71144 93494 71464 100258
rect 71144 93258 71186 93494
rect 71422 93258 71464 93494
rect 71144 86494 71464 93258
rect 71144 86258 71186 86494
rect 71422 86258 71464 86494
rect 71144 79494 71464 86258
rect 71144 79258 71186 79494
rect 71422 79258 71464 79494
rect 71144 72494 71464 79258
rect 71144 72258 71186 72494
rect 71422 72258 71464 72494
rect 71144 65494 71464 72258
rect 71144 65258 71186 65494
rect 71422 65258 71464 65494
rect 71144 58494 71464 65258
rect 71144 58258 71186 58494
rect 71422 58258 71464 58494
rect 71144 51494 71464 58258
rect 71144 51258 71186 51494
rect 71422 51258 71464 51494
rect 71144 44494 71464 51258
rect 71144 44258 71186 44494
rect 71422 44258 71464 44494
rect 71144 37494 71464 44258
rect 71144 37258 71186 37494
rect 71422 37258 71464 37494
rect 71144 30494 71464 37258
rect 71144 30258 71186 30494
rect 71422 30258 71464 30494
rect 71144 23494 71464 30258
rect 71144 23258 71186 23494
rect 71422 23258 71464 23494
rect 71144 16494 71464 23258
rect 71144 16258 71186 16494
rect 71422 16258 71464 16494
rect 71144 9494 71464 16258
rect 71144 9258 71186 9494
rect 71422 9258 71464 9494
rect 71144 2494 71464 9258
rect 71144 2258 71186 2494
rect 71422 2258 71464 2494
rect 71144 -746 71464 2258
rect 71144 -982 71186 -746
rect 71422 -982 71464 -746
rect 71144 -1066 71464 -982
rect 71144 -1302 71186 -1066
rect 71422 -1302 71464 -1066
rect 71144 -2294 71464 -1302
rect 72876 706198 73196 706230
rect 72876 705962 72918 706198
rect 73154 705962 73196 706198
rect 72876 705878 73196 705962
rect 72876 705642 72918 705878
rect 73154 705642 73196 705878
rect 72876 696434 73196 705642
rect 72876 696198 72918 696434
rect 73154 696198 73196 696434
rect 72876 689434 73196 696198
rect 72876 689198 72918 689434
rect 73154 689198 73196 689434
rect 72876 682434 73196 689198
rect 72876 682198 72918 682434
rect 73154 682198 73196 682434
rect 72876 675434 73196 682198
rect 72876 675198 72918 675434
rect 73154 675198 73196 675434
rect 72876 668434 73196 675198
rect 72876 668198 72918 668434
rect 73154 668198 73196 668434
rect 72876 661434 73196 668198
rect 72876 661198 72918 661434
rect 73154 661198 73196 661434
rect 72876 654434 73196 661198
rect 72876 654198 72918 654434
rect 73154 654198 73196 654434
rect 72876 647434 73196 654198
rect 72876 647198 72918 647434
rect 73154 647198 73196 647434
rect 72876 640434 73196 647198
rect 72876 640198 72918 640434
rect 73154 640198 73196 640434
rect 72876 633434 73196 640198
rect 72876 633198 72918 633434
rect 73154 633198 73196 633434
rect 72876 626434 73196 633198
rect 72876 626198 72918 626434
rect 73154 626198 73196 626434
rect 72876 619434 73196 626198
rect 72876 619198 72918 619434
rect 73154 619198 73196 619434
rect 72876 612434 73196 619198
rect 72876 612198 72918 612434
rect 73154 612198 73196 612434
rect 72876 605434 73196 612198
rect 72876 605198 72918 605434
rect 73154 605198 73196 605434
rect 72876 598434 73196 605198
rect 72876 598198 72918 598434
rect 73154 598198 73196 598434
rect 72876 591434 73196 598198
rect 72876 591198 72918 591434
rect 73154 591198 73196 591434
rect 72876 584434 73196 591198
rect 72876 584198 72918 584434
rect 73154 584198 73196 584434
rect 72876 577434 73196 584198
rect 72876 577198 72918 577434
rect 73154 577198 73196 577434
rect 72876 570434 73196 577198
rect 72876 570198 72918 570434
rect 73154 570198 73196 570434
rect 72876 563434 73196 570198
rect 72876 563198 72918 563434
rect 73154 563198 73196 563434
rect 72876 556434 73196 563198
rect 72876 556198 72918 556434
rect 73154 556198 73196 556434
rect 72876 549434 73196 556198
rect 72876 549198 72918 549434
rect 73154 549198 73196 549434
rect 72876 542434 73196 549198
rect 72876 542198 72918 542434
rect 73154 542198 73196 542434
rect 72876 535434 73196 542198
rect 72876 535198 72918 535434
rect 73154 535198 73196 535434
rect 72876 528434 73196 535198
rect 72876 528198 72918 528434
rect 73154 528198 73196 528434
rect 72876 521434 73196 528198
rect 72876 521198 72918 521434
rect 73154 521198 73196 521434
rect 72876 514434 73196 521198
rect 72876 514198 72918 514434
rect 73154 514198 73196 514434
rect 72876 507434 73196 514198
rect 72876 507198 72918 507434
rect 73154 507198 73196 507434
rect 72876 500434 73196 507198
rect 72876 500198 72918 500434
rect 73154 500198 73196 500434
rect 72876 493434 73196 500198
rect 72876 493198 72918 493434
rect 73154 493198 73196 493434
rect 72876 486434 73196 493198
rect 72876 486198 72918 486434
rect 73154 486198 73196 486434
rect 72876 479434 73196 486198
rect 72876 479198 72918 479434
rect 73154 479198 73196 479434
rect 72876 472434 73196 479198
rect 72876 472198 72918 472434
rect 73154 472198 73196 472434
rect 72876 465434 73196 472198
rect 72876 465198 72918 465434
rect 73154 465198 73196 465434
rect 72876 458434 73196 465198
rect 72876 458198 72918 458434
rect 73154 458198 73196 458434
rect 72876 451434 73196 458198
rect 72876 451198 72918 451434
rect 73154 451198 73196 451434
rect 72876 444434 73196 451198
rect 72876 444198 72918 444434
rect 73154 444198 73196 444434
rect 72876 437434 73196 444198
rect 72876 437198 72918 437434
rect 73154 437198 73196 437434
rect 72876 430434 73196 437198
rect 72876 430198 72918 430434
rect 73154 430198 73196 430434
rect 72876 423434 73196 430198
rect 72876 423198 72918 423434
rect 73154 423198 73196 423434
rect 72876 416434 73196 423198
rect 72876 416198 72918 416434
rect 73154 416198 73196 416434
rect 72876 409434 73196 416198
rect 72876 409198 72918 409434
rect 73154 409198 73196 409434
rect 72876 402434 73196 409198
rect 72876 402198 72918 402434
rect 73154 402198 73196 402434
rect 72876 395434 73196 402198
rect 72876 395198 72918 395434
rect 73154 395198 73196 395434
rect 72876 388434 73196 395198
rect 72876 388198 72918 388434
rect 73154 388198 73196 388434
rect 72876 381434 73196 388198
rect 72876 381198 72918 381434
rect 73154 381198 73196 381434
rect 72876 374434 73196 381198
rect 72876 374198 72918 374434
rect 73154 374198 73196 374434
rect 72876 367434 73196 374198
rect 72876 367198 72918 367434
rect 73154 367198 73196 367434
rect 72876 360434 73196 367198
rect 72876 360198 72918 360434
rect 73154 360198 73196 360434
rect 72876 353434 73196 360198
rect 72876 353198 72918 353434
rect 73154 353198 73196 353434
rect 72876 346434 73196 353198
rect 72876 346198 72918 346434
rect 73154 346198 73196 346434
rect 72876 339434 73196 346198
rect 72876 339198 72918 339434
rect 73154 339198 73196 339434
rect 72876 332434 73196 339198
rect 72876 332198 72918 332434
rect 73154 332198 73196 332434
rect 72876 325434 73196 332198
rect 72876 325198 72918 325434
rect 73154 325198 73196 325434
rect 72876 318434 73196 325198
rect 72876 318198 72918 318434
rect 73154 318198 73196 318434
rect 72876 311434 73196 318198
rect 72876 311198 72918 311434
rect 73154 311198 73196 311434
rect 72876 304434 73196 311198
rect 72876 304198 72918 304434
rect 73154 304198 73196 304434
rect 72876 297434 73196 304198
rect 72876 297198 72918 297434
rect 73154 297198 73196 297434
rect 72876 290434 73196 297198
rect 72876 290198 72918 290434
rect 73154 290198 73196 290434
rect 72876 283434 73196 290198
rect 72876 283198 72918 283434
rect 73154 283198 73196 283434
rect 72876 276434 73196 283198
rect 72876 276198 72918 276434
rect 73154 276198 73196 276434
rect 72876 269434 73196 276198
rect 72876 269198 72918 269434
rect 73154 269198 73196 269434
rect 72876 262434 73196 269198
rect 72876 262198 72918 262434
rect 73154 262198 73196 262434
rect 72876 255434 73196 262198
rect 72876 255198 72918 255434
rect 73154 255198 73196 255434
rect 72876 248434 73196 255198
rect 72876 248198 72918 248434
rect 73154 248198 73196 248434
rect 72876 241434 73196 248198
rect 72876 241198 72918 241434
rect 73154 241198 73196 241434
rect 72876 234434 73196 241198
rect 72876 234198 72918 234434
rect 73154 234198 73196 234434
rect 72876 227434 73196 234198
rect 72876 227198 72918 227434
rect 73154 227198 73196 227434
rect 72876 220434 73196 227198
rect 72876 220198 72918 220434
rect 73154 220198 73196 220434
rect 72876 213434 73196 220198
rect 72876 213198 72918 213434
rect 73154 213198 73196 213434
rect 72876 206434 73196 213198
rect 72876 206198 72918 206434
rect 73154 206198 73196 206434
rect 72876 199434 73196 206198
rect 72876 199198 72918 199434
rect 73154 199198 73196 199434
rect 72876 192434 73196 199198
rect 72876 192198 72918 192434
rect 73154 192198 73196 192434
rect 72876 185434 73196 192198
rect 72876 185198 72918 185434
rect 73154 185198 73196 185434
rect 72876 178434 73196 185198
rect 72876 178198 72918 178434
rect 73154 178198 73196 178434
rect 72876 171434 73196 178198
rect 72876 171198 72918 171434
rect 73154 171198 73196 171434
rect 72876 164434 73196 171198
rect 72876 164198 72918 164434
rect 73154 164198 73196 164434
rect 72876 157434 73196 164198
rect 72876 157198 72918 157434
rect 73154 157198 73196 157434
rect 72876 150434 73196 157198
rect 72876 150198 72918 150434
rect 73154 150198 73196 150434
rect 72876 143434 73196 150198
rect 72876 143198 72918 143434
rect 73154 143198 73196 143434
rect 72876 136434 73196 143198
rect 72876 136198 72918 136434
rect 73154 136198 73196 136434
rect 72876 129434 73196 136198
rect 72876 129198 72918 129434
rect 73154 129198 73196 129434
rect 72876 122434 73196 129198
rect 72876 122198 72918 122434
rect 73154 122198 73196 122434
rect 72876 115434 73196 122198
rect 72876 115198 72918 115434
rect 73154 115198 73196 115434
rect 72876 108434 73196 115198
rect 72876 108198 72918 108434
rect 73154 108198 73196 108434
rect 72876 101434 73196 108198
rect 72876 101198 72918 101434
rect 73154 101198 73196 101434
rect 72876 94434 73196 101198
rect 72876 94198 72918 94434
rect 73154 94198 73196 94434
rect 72876 87434 73196 94198
rect 72876 87198 72918 87434
rect 73154 87198 73196 87434
rect 72876 80434 73196 87198
rect 72876 80198 72918 80434
rect 73154 80198 73196 80434
rect 72876 73434 73196 80198
rect 72876 73198 72918 73434
rect 73154 73198 73196 73434
rect 72876 66434 73196 73198
rect 72876 66198 72918 66434
rect 73154 66198 73196 66434
rect 72876 59434 73196 66198
rect 72876 59198 72918 59434
rect 73154 59198 73196 59434
rect 72876 52434 73196 59198
rect 72876 52198 72918 52434
rect 73154 52198 73196 52434
rect 72876 45434 73196 52198
rect 72876 45198 72918 45434
rect 73154 45198 73196 45434
rect 72876 38434 73196 45198
rect 72876 38198 72918 38434
rect 73154 38198 73196 38434
rect 72876 31434 73196 38198
rect 72876 31198 72918 31434
rect 73154 31198 73196 31434
rect 72876 24434 73196 31198
rect 72876 24198 72918 24434
rect 73154 24198 73196 24434
rect 72876 17434 73196 24198
rect 72876 17198 72918 17434
rect 73154 17198 73196 17434
rect 72876 10434 73196 17198
rect 72876 10198 72918 10434
rect 73154 10198 73196 10434
rect 72876 3434 73196 10198
rect 72876 3198 72918 3434
rect 73154 3198 73196 3434
rect 72876 -1706 73196 3198
rect 72876 -1942 72918 -1706
rect 73154 -1942 73196 -1706
rect 72876 -2026 73196 -1942
rect 72876 -2262 72918 -2026
rect 73154 -2262 73196 -2026
rect 72876 -2294 73196 -2262
rect 78144 705238 78464 706230
rect 78144 705002 78186 705238
rect 78422 705002 78464 705238
rect 78144 704918 78464 705002
rect 78144 704682 78186 704918
rect 78422 704682 78464 704918
rect 78144 695494 78464 704682
rect 78144 695258 78186 695494
rect 78422 695258 78464 695494
rect 78144 688494 78464 695258
rect 78144 688258 78186 688494
rect 78422 688258 78464 688494
rect 78144 681494 78464 688258
rect 78144 681258 78186 681494
rect 78422 681258 78464 681494
rect 78144 674494 78464 681258
rect 78144 674258 78186 674494
rect 78422 674258 78464 674494
rect 78144 667494 78464 674258
rect 78144 667258 78186 667494
rect 78422 667258 78464 667494
rect 78144 660494 78464 667258
rect 78144 660258 78186 660494
rect 78422 660258 78464 660494
rect 78144 653494 78464 660258
rect 78144 653258 78186 653494
rect 78422 653258 78464 653494
rect 78144 646494 78464 653258
rect 78144 646258 78186 646494
rect 78422 646258 78464 646494
rect 78144 639494 78464 646258
rect 78144 639258 78186 639494
rect 78422 639258 78464 639494
rect 78144 632494 78464 639258
rect 78144 632258 78186 632494
rect 78422 632258 78464 632494
rect 78144 625494 78464 632258
rect 78144 625258 78186 625494
rect 78422 625258 78464 625494
rect 78144 618494 78464 625258
rect 78144 618258 78186 618494
rect 78422 618258 78464 618494
rect 78144 611494 78464 618258
rect 78144 611258 78186 611494
rect 78422 611258 78464 611494
rect 78144 604494 78464 611258
rect 78144 604258 78186 604494
rect 78422 604258 78464 604494
rect 78144 597494 78464 604258
rect 78144 597258 78186 597494
rect 78422 597258 78464 597494
rect 78144 590494 78464 597258
rect 78144 590258 78186 590494
rect 78422 590258 78464 590494
rect 78144 583494 78464 590258
rect 78144 583258 78186 583494
rect 78422 583258 78464 583494
rect 78144 576494 78464 583258
rect 78144 576258 78186 576494
rect 78422 576258 78464 576494
rect 78144 569494 78464 576258
rect 78144 569258 78186 569494
rect 78422 569258 78464 569494
rect 78144 562494 78464 569258
rect 78144 562258 78186 562494
rect 78422 562258 78464 562494
rect 78144 555494 78464 562258
rect 78144 555258 78186 555494
rect 78422 555258 78464 555494
rect 78144 548494 78464 555258
rect 78144 548258 78186 548494
rect 78422 548258 78464 548494
rect 78144 541494 78464 548258
rect 78144 541258 78186 541494
rect 78422 541258 78464 541494
rect 78144 534494 78464 541258
rect 78144 534258 78186 534494
rect 78422 534258 78464 534494
rect 78144 527494 78464 534258
rect 78144 527258 78186 527494
rect 78422 527258 78464 527494
rect 78144 520494 78464 527258
rect 78144 520258 78186 520494
rect 78422 520258 78464 520494
rect 78144 513494 78464 520258
rect 78144 513258 78186 513494
rect 78422 513258 78464 513494
rect 78144 506494 78464 513258
rect 78144 506258 78186 506494
rect 78422 506258 78464 506494
rect 78144 499494 78464 506258
rect 78144 499258 78186 499494
rect 78422 499258 78464 499494
rect 78144 492494 78464 499258
rect 78144 492258 78186 492494
rect 78422 492258 78464 492494
rect 78144 485494 78464 492258
rect 78144 485258 78186 485494
rect 78422 485258 78464 485494
rect 78144 478494 78464 485258
rect 78144 478258 78186 478494
rect 78422 478258 78464 478494
rect 78144 471494 78464 478258
rect 78144 471258 78186 471494
rect 78422 471258 78464 471494
rect 78144 464494 78464 471258
rect 78144 464258 78186 464494
rect 78422 464258 78464 464494
rect 78144 457494 78464 464258
rect 78144 457258 78186 457494
rect 78422 457258 78464 457494
rect 78144 450494 78464 457258
rect 78144 450258 78186 450494
rect 78422 450258 78464 450494
rect 78144 443494 78464 450258
rect 78144 443258 78186 443494
rect 78422 443258 78464 443494
rect 78144 436494 78464 443258
rect 78144 436258 78186 436494
rect 78422 436258 78464 436494
rect 78144 429494 78464 436258
rect 78144 429258 78186 429494
rect 78422 429258 78464 429494
rect 78144 422494 78464 429258
rect 78144 422258 78186 422494
rect 78422 422258 78464 422494
rect 78144 415494 78464 422258
rect 78144 415258 78186 415494
rect 78422 415258 78464 415494
rect 78144 408494 78464 415258
rect 78144 408258 78186 408494
rect 78422 408258 78464 408494
rect 78144 401494 78464 408258
rect 78144 401258 78186 401494
rect 78422 401258 78464 401494
rect 78144 394494 78464 401258
rect 78144 394258 78186 394494
rect 78422 394258 78464 394494
rect 78144 387494 78464 394258
rect 78144 387258 78186 387494
rect 78422 387258 78464 387494
rect 78144 380494 78464 387258
rect 78144 380258 78186 380494
rect 78422 380258 78464 380494
rect 78144 373494 78464 380258
rect 78144 373258 78186 373494
rect 78422 373258 78464 373494
rect 78144 366494 78464 373258
rect 78144 366258 78186 366494
rect 78422 366258 78464 366494
rect 78144 359494 78464 366258
rect 78144 359258 78186 359494
rect 78422 359258 78464 359494
rect 78144 352494 78464 359258
rect 78144 352258 78186 352494
rect 78422 352258 78464 352494
rect 78144 345494 78464 352258
rect 78144 345258 78186 345494
rect 78422 345258 78464 345494
rect 78144 338494 78464 345258
rect 78144 338258 78186 338494
rect 78422 338258 78464 338494
rect 78144 331494 78464 338258
rect 78144 331258 78186 331494
rect 78422 331258 78464 331494
rect 78144 324494 78464 331258
rect 78144 324258 78186 324494
rect 78422 324258 78464 324494
rect 78144 317494 78464 324258
rect 78144 317258 78186 317494
rect 78422 317258 78464 317494
rect 78144 310494 78464 317258
rect 78144 310258 78186 310494
rect 78422 310258 78464 310494
rect 78144 303494 78464 310258
rect 78144 303258 78186 303494
rect 78422 303258 78464 303494
rect 78144 296494 78464 303258
rect 78144 296258 78186 296494
rect 78422 296258 78464 296494
rect 78144 289494 78464 296258
rect 78144 289258 78186 289494
rect 78422 289258 78464 289494
rect 78144 282494 78464 289258
rect 78144 282258 78186 282494
rect 78422 282258 78464 282494
rect 78144 275494 78464 282258
rect 78144 275258 78186 275494
rect 78422 275258 78464 275494
rect 78144 268494 78464 275258
rect 78144 268258 78186 268494
rect 78422 268258 78464 268494
rect 78144 261494 78464 268258
rect 78144 261258 78186 261494
rect 78422 261258 78464 261494
rect 78144 254494 78464 261258
rect 78144 254258 78186 254494
rect 78422 254258 78464 254494
rect 78144 247494 78464 254258
rect 78144 247258 78186 247494
rect 78422 247258 78464 247494
rect 78144 240494 78464 247258
rect 78144 240258 78186 240494
rect 78422 240258 78464 240494
rect 78144 233494 78464 240258
rect 78144 233258 78186 233494
rect 78422 233258 78464 233494
rect 78144 226494 78464 233258
rect 78144 226258 78186 226494
rect 78422 226258 78464 226494
rect 78144 219494 78464 226258
rect 78144 219258 78186 219494
rect 78422 219258 78464 219494
rect 78144 212494 78464 219258
rect 78144 212258 78186 212494
rect 78422 212258 78464 212494
rect 78144 205494 78464 212258
rect 78144 205258 78186 205494
rect 78422 205258 78464 205494
rect 78144 198494 78464 205258
rect 78144 198258 78186 198494
rect 78422 198258 78464 198494
rect 78144 191494 78464 198258
rect 78144 191258 78186 191494
rect 78422 191258 78464 191494
rect 78144 184494 78464 191258
rect 78144 184258 78186 184494
rect 78422 184258 78464 184494
rect 78144 177494 78464 184258
rect 78144 177258 78186 177494
rect 78422 177258 78464 177494
rect 78144 170494 78464 177258
rect 78144 170258 78186 170494
rect 78422 170258 78464 170494
rect 78144 163494 78464 170258
rect 78144 163258 78186 163494
rect 78422 163258 78464 163494
rect 78144 156494 78464 163258
rect 78144 156258 78186 156494
rect 78422 156258 78464 156494
rect 78144 149494 78464 156258
rect 78144 149258 78186 149494
rect 78422 149258 78464 149494
rect 78144 142494 78464 149258
rect 78144 142258 78186 142494
rect 78422 142258 78464 142494
rect 78144 135494 78464 142258
rect 78144 135258 78186 135494
rect 78422 135258 78464 135494
rect 78144 128494 78464 135258
rect 78144 128258 78186 128494
rect 78422 128258 78464 128494
rect 78144 121494 78464 128258
rect 78144 121258 78186 121494
rect 78422 121258 78464 121494
rect 78144 114494 78464 121258
rect 78144 114258 78186 114494
rect 78422 114258 78464 114494
rect 78144 107494 78464 114258
rect 78144 107258 78186 107494
rect 78422 107258 78464 107494
rect 78144 100494 78464 107258
rect 78144 100258 78186 100494
rect 78422 100258 78464 100494
rect 78144 93494 78464 100258
rect 78144 93258 78186 93494
rect 78422 93258 78464 93494
rect 78144 86494 78464 93258
rect 78144 86258 78186 86494
rect 78422 86258 78464 86494
rect 78144 79494 78464 86258
rect 78144 79258 78186 79494
rect 78422 79258 78464 79494
rect 78144 72494 78464 79258
rect 78144 72258 78186 72494
rect 78422 72258 78464 72494
rect 78144 65494 78464 72258
rect 78144 65258 78186 65494
rect 78422 65258 78464 65494
rect 78144 58494 78464 65258
rect 78144 58258 78186 58494
rect 78422 58258 78464 58494
rect 78144 51494 78464 58258
rect 78144 51258 78186 51494
rect 78422 51258 78464 51494
rect 78144 44494 78464 51258
rect 78144 44258 78186 44494
rect 78422 44258 78464 44494
rect 78144 37494 78464 44258
rect 78144 37258 78186 37494
rect 78422 37258 78464 37494
rect 78144 30494 78464 37258
rect 78144 30258 78186 30494
rect 78422 30258 78464 30494
rect 78144 23494 78464 30258
rect 78144 23258 78186 23494
rect 78422 23258 78464 23494
rect 78144 16494 78464 23258
rect 78144 16258 78186 16494
rect 78422 16258 78464 16494
rect 78144 9494 78464 16258
rect 78144 9258 78186 9494
rect 78422 9258 78464 9494
rect 78144 2494 78464 9258
rect 78144 2258 78186 2494
rect 78422 2258 78464 2494
rect 78144 -746 78464 2258
rect 78144 -982 78186 -746
rect 78422 -982 78464 -746
rect 78144 -1066 78464 -982
rect 78144 -1302 78186 -1066
rect 78422 -1302 78464 -1066
rect 78144 -2294 78464 -1302
rect 79876 706198 80196 706230
rect 79876 705962 79918 706198
rect 80154 705962 80196 706198
rect 79876 705878 80196 705962
rect 79876 705642 79918 705878
rect 80154 705642 80196 705878
rect 79876 696434 80196 705642
rect 79876 696198 79918 696434
rect 80154 696198 80196 696434
rect 79876 689434 80196 696198
rect 79876 689198 79918 689434
rect 80154 689198 80196 689434
rect 79876 682434 80196 689198
rect 79876 682198 79918 682434
rect 80154 682198 80196 682434
rect 79876 675434 80196 682198
rect 79876 675198 79918 675434
rect 80154 675198 80196 675434
rect 79876 668434 80196 675198
rect 79876 668198 79918 668434
rect 80154 668198 80196 668434
rect 79876 661434 80196 668198
rect 79876 661198 79918 661434
rect 80154 661198 80196 661434
rect 79876 654434 80196 661198
rect 79876 654198 79918 654434
rect 80154 654198 80196 654434
rect 79876 647434 80196 654198
rect 79876 647198 79918 647434
rect 80154 647198 80196 647434
rect 79876 640434 80196 647198
rect 79876 640198 79918 640434
rect 80154 640198 80196 640434
rect 79876 633434 80196 640198
rect 79876 633198 79918 633434
rect 80154 633198 80196 633434
rect 79876 626434 80196 633198
rect 79876 626198 79918 626434
rect 80154 626198 80196 626434
rect 79876 619434 80196 626198
rect 79876 619198 79918 619434
rect 80154 619198 80196 619434
rect 79876 612434 80196 619198
rect 79876 612198 79918 612434
rect 80154 612198 80196 612434
rect 79876 605434 80196 612198
rect 79876 605198 79918 605434
rect 80154 605198 80196 605434
rect 79876 598434 80196 605198
rect 79876 598198 79918 598434
rect 80154 598198 80196 598434
rect 79876 591434 80196 598198
rect 79876 591198 79918 591434
rect 80154 591198 80196 591434
rect 79876 584434 80196 591198
rect 79876 584198 79918 584434
rect 80154 584198 80196 584434
rect 79876 577434 80196 584198
rect 79876 577198 79918 577434
rect 80154 577198 80196 577434
rect 79876 570434 80196 577198
rect 79876 570198 79918 570434
rect 80154 570198 80196 570434
rect 79876 563434 80196 570198
rect 79876 563198 79918 563434
rect 80154 563198 80196 563434
rect 79876 556434 80196 563198
rect 79876 556198 79918 556434
rect 80154 556198 80196 556434
rect 79876 549434 80196 556198
rect 79876 549198 79918 549434
rect 80154 549198 80196 549434
rect 79876 542434 80196 549198
rect 79876 542198 79918 542434
rect 80154 542198 80196 542434
rect 79876 535434 80196 542198
rect 79876 535198 79918 535434
rect 80154 535198 80196 535434
rect 79876 528434 80196 535198
rect 79876 528198 79918 528434
rect 80154 528198 80196 528434
rect 79876 521434 80196 528198
rect 79876 521198 79918 521434
rect 80154 521198 80196 521434
rect 79876 514434 80196 521198
rect 79876 514198 79918 514434
rect 80154 514198 80196 514434
rect 79876 507434 80196 514198
rect 79876 507198 79918 507434
rect 80154 507198 80196 507434
rect 79876 500434 80196 507198
rect 79876 500198 79918 500434
rect 80154 500198 80196 500434
rect 79876 493434 80196 500198
rect 79876 493198 79918 493434
rect 80154 493198 80196 493434
rect 79876 486434 80196 493198
rect 79876 486198 79918 486434
rect 80154 486198 80196 486434
rect 79876 479434 80196 486198
rect 79876 479198 79918 479434
rect 80154 479198 80196 479434
rect 79876 472434 80196 479198
rect 79876 472198 79918 472434
rect 80154 472198 80196 472434
rect 79876 465434 80196 472198
rect 79876 465198 79918 465434
rect 80154 465198 80196 465434
rect 79876 458434 80196 465198
rect 79876 458198 79918 458434
rect 80154 458198 80196 458434
rect 79876 451434 80196 458198
rect 79876 451198 79918 451434
rect 80154 451198 80196 451434
rect 79876 444434 80196 451198
rect 79876 444198 79918 444434
rect 80154 444198 80196 444434
rect 79876 437434 80196 444198
rect 79876 437198 79918 437434
rect 80154 437198 80196 437434
rect 79876 430434 80196 437198
rect 79876 430198 79918 430434
rect 80154 430198 80196 430434
rect 79876 423434 80196 430198
rect 79876 423198 79918 423434
rect 80154 423198 80196 423434
rect 79876 416434 80196 423198
rect 79876 416198 79918 416434
rect 80154 416198 80196 416434
rect 79876 409434 80196 416198
rect 79876 409198 79918 409434
rect 80154 409198 80196 409434
rect 79876 402434 80196 409198
rect 79876 402198 79918 402434
rect 80154 402198 80196 402434
rect 79876 395434 80196 402198
rect 79876 395198 79918 395434
rect 80154 395198 80196 395434
rect 79876 388434 80196 395198
rect 79876 388198 79918 388434
rect 80154 388198 80196 388434
rect 79876 381434 80196 388198
rect 79876 381198 79918 381434
rect 80154 381198 80196 381434
rect 79876 374434 80196 381198
rect 79876 374198 79918 374434
rect 80154 374198 80196 374434
rect 79876 367434 80196 374198
rect 79876 367198 79918 367434
rect 80154 367198 80196 367434
rect 79876 360434 80196 367198
rect 79876 360198 79918 360434
rect 80154 360198 80196 360434
rect 79876 353434 80196 360198
rect 79876 353198 79918 353434
rect 80154 353198 80196 353434
rect 79876 346434 80196 353198
rect 79876 346198 79918 346434
rect 80154 346198 80196 346434
rect 79876 339434 80196 346198
rect 79876 339198 79918 339434
rect 80154 339198 80196 339434
rect 79876 332434 80196 339198
rect 79876 332198 79918 332434
rect 80154 332198 80196 332434
rect 79876 325434 80196 332198
rect 79876 325198 79918 325434
rect 80154 325198 80196 325434
rect 79876 318434 80196 325198
rect 79876 318198 79918 318434
rect 80154 318198 80196 318434
rect 79876 311434 80196 318198
rect 79876 311198 79918 311434
rect 80154 311198 80196 311434
rect 79876 304434 80196 311198
rect 79876 304198 79918 304434
rect 80154 304198 80196 304434
rect 79876 297434 80196 304198
rect 79876 297198 79918 297434
rect 80154 297198 80196 297434
rect 79876 290434 80196 297198
rect 79876 290198 79918 290434
rect 80154 290198 80196 290434
rect 79876 283434 80196 290198
rect 79876 283198 79918 283434
rect 80154 283198 80196 283434
rect 79876 276434 80196 283198
rect 79876 276198 79918 276434
rect 80154 276198 80196 276434
rect 79876 269434 80196 276198
rect 79876 269198 79918 269434
rect 80154 269198 80196 269434
rect 79876 262434 80196 269198
rect 79876 262198 79918 262434
rect 80154 262198 80196 262434
rect 79876 255434 80196 262198
rect 79876 255198 79918 255434
rect 80154 255198 80196 255434
rect 79876 248434 80196 255198
rect 79876 248198 79918 248434
rect 80154 248198 80196 248434
rect 79876 241434 80196 248198
rect 79876 241198 79918 241434
rect 80154 241198 80196 241434
rect 79876 234434 80196 241198
rect 79876 234198 79918 234434
rect 80154 234198 80196 234434
rect 79876 227434 80196 234198
rect 79876 227198 79918 227434
rect 80154 227198 80196 227434
rect 79876 220434 80196 227198
rect 79876 220198 79918 220434
rect 80154 220198 80196 220434
rect 79876 213434 80196 220198
rect 79876 213198 79918 213434
rect 80154 213198 80196 213434
rect 79876 206434 80196 213198
rect 79876 206198 79918 206434
rect 80154 206198 80196 206434
rect 79876 199434 80196 206198
rect 79876 199198 79918 199434
rect 80154 199198 80196 199434
rect 79876 192434 80196 199198
rect 79876 192198 79918 192434
rect 80154 192198 80196 192434
rect 79876 185434 80196 192198
rect 79876 185198 79918 185434
rect 80154 185198 80196 185434
rect 79876 178434 80196 185198
rect 79876 178198 79918 178434
rect 80154 178198 80196 178434
rect 79876 171434 80196 178198
rect 79876 171198 79918 171434
rect 80154 171198 80196 171434
rect 79876 164434 80196 171198
rect 79876 164198 79918 164434
rect 80154 164198 80196 164434
rect 79876 157434 80196 164198
rect 79876 157198 79918 157434
rect 80154 157198 80196 157434
rect 79876 150434 80196 157198
rect 79876 150198 79918 150434
rect 80154 150198 80196 150434
rect 79876 143434 80196 150198
rect 79876 143198 79918 143434
rect 80154 143198 80196 143434
rect 79876 136434 80196 143198
rect 79876 136198 79918 136434
rect 80154 136198 80196 136434
rect 79876 129434 80196 136198
rect 79876 129198 79918 129434
rect 80154 129198 80196 129434
rect 79876 122434 80196 129198
rect 79876 122198 79918 122434
rect 80154 122198 80196 122434
rect 79876 115434 80196 122198
rect 79876 115198 79918 115434
rect 80154 115198 80196 115434
rect 79876 108434 80196 115198
rect 79876 108198 79918 108434
rect 80154 108198 80196 108434
rect 79876 101434 80196 108198
rect 79876 101198 79918 101434
rect 80154 101198 80196 101434
rect 79876 94434 80196 101198
rect 79876 94198 79918 94434
rect 80154 94198 80196 94434
rect 79876 87434 80196 94198
rect 79876 87198 79918 87434
rect 80154 87198 80196 87434
rect 79876 80434 80196 87198
rect 79876 80198 79918 80434
rect 80154 80198 80196 80434
rect 79876 73434 80196 80198
rect 79876 73198 79918 73434
rect 80154 73198 80196 73434
rect 79876 66434 80196 73198
rect 79876 66198 79918 66434
rect 80154 66198 80196 66434
rect 79876 59434 80196 66198
rect 79876 59198 79918 59434
rect 80154 59198 80196 59434
rect 79876 52434 80196 59198
rect 79876 52198 79918 52434
rect 80154 52198 80196 52434
rect 79876 45434 80196 52198
rect 79876 45198 79918 45434
rect 80154 45198 80196 45434
rect 79876 38434 80196 45198
rect 79876 38198 79918 38434
rect 80154 38198 80196 38434
rect 79876 31434 80196 38198
rect 79876 31198 79918 31434
rect 80154 31198 80196 31434
rect 79876 24434 80196 31198
rect 79876 24198 79918 24434
rect 80154 24198 80196 24434
rect 79876 17434 80196 24198
rect 79876 17198 79918 17434
rect 80154 17198 80196 17434
rect 79876 10434 80196 17198
rect 79876 10198 79918 10434
rect 80154 10198 80196 10434
rect 79876 3434 80196 10198
rect 79876 3198 79918 3434
rect 80154 3198 80196 3434
rect 79876 -1706 80196 3198
rect 79876 -1942 79918 -1706
rect 80154 -1942 80196 -1706
rect 79876 -2026 80196 -1942
rect 79876 -2262 79918 -2026
rect 80154 -2262 80196 -2026
rect 79876 -2294 80196 -2262
rect 85144 705238 85464 706230
rect 85144 705002 85186 705238
rect 85422 705002 85464 705238
rect 85144 704918 85464 705002
rect 85144 704682 85186 704918
rect 85422 704682 85464 704918
rect 85144 695494 85464 704682
rect 85144 695258 85186 695494
rect 85422 695258 85464 695494
rect 85144 688494 85464 695258
rect 85144 688258 85186 688494
rect 85422 688258 85464 688494
rect 85144 681494 85464 688258
rect 85144 681258 85186 681494
rect 85422 681258 85464 681494
rect 85144 674494 85464 681258
rect 85144 674258 85186 674494
rect 85422 674258 85464 674494
rect 85144 667494 85464 674258
rect 85144 667258 85186 667494
rect 85422 667258 85464 667494
rect 85144 660494 85464 667258
rect 85144 660258 85186 660494
rect 85422 660258 85464 660494
rect 85144 653494 85464 660258
rect 85144 653258 85186 653494
rect 85422 653258 85464 653494
rect 85144 646494 85464 653258
rect 85144 646258 85186 646494
rect 85422 646258 85464 646494
rect 85144 639494 85464 646258
rect 85144 639258 85186 639494
rect 85422 639258 85464 639494
rect 85144 632494 85464 639258
rect 85144 632258 85186 632494
rect 85422 632258 85464 632494
rect 85144 625494 85464 632258
rect 85144 625258 85186 625494
rect 85422 625258 85464 625494
rect 85144 618494 85464 625258
rect 85144 618258 85186 618494
rect 85422 618258 85464 618494
rect 85144 611494 85464 618258
rect 85144 611258 85186 611494
rect 85422 611258 85464 611494
rect 85144 604494 85464 611258
rect 85144 604258 85186 604494
rect 85422 604258 85464 604494
rect 85144 597494 85464 604258
rect 85144 597258 85186 597494
rect 85422 597258 85464 597494
rect 85144 590494 85464 597258
rect 85144 590258 85186 590494
rect 85422 590258 85464 590494
rect 85144 583494 85464 590258
rect 85144 583258 85186 583494
rect 85422 583258 85464 583494
rect 85144 576494 85464 583258
rect 85144 576258 85186 576494
rect 85422 576258 85464 576494
rect 85144 569494 85464 576258
rect 85144 569258 85186 569494
rect 85422 569258 85464 569494
rect 85144 562494 85464 569258
rect 85144 562258 85186 562494
rect 85422 562258 85464 562494
rect 85144 555494 85464 562258
rect 85144 555258 85186 555494
rect 85422 555258 85464 555494
rect 85144 548494 85464 555258
rect 85144 548258 85186 548494
rect 85422 548258 85464 548494
rect 85144 541494 85464 548258
rect 85144 541258 85186 541494
rect 85422 541258 85464 541494
rect 85144 534494 85464 541258
rect 85144 534258 85186 534494
rect 85422 534258 85464 534494
rect 85144 527494 85464 534258
rect 85144 527258 85186 527494
rect 85422 527258 85464 527494
rect 85144 520494 85464 527258
rect 85144 520258 85186 520494
rect 85422 520258 85464 520494
rect 85144 513494 85464 520258
rect 85144 513258 85186 513494
rect 85422 513258 85464 513494
rect 85144 506494 85464 513258
rect 85144 506258 85186 506494
rect 85422 506258 85464 506494
rect 85144 499494 85464 506258
rect 85144 499258 85186 499494
rect 85422 499258 85464 499494
rect 85144 492494 85464 499258
rect 85144 492258 85186 492494
rect 85422 492258 85464 492494
rect 85144 485494 85464 492258
rect 85144 485258 85186 485494
rect 85422 485258 85464 485494
rect 85144 478494 85464 485258
rect 85144 478258 85186 478494
rect 85422 478258 85464 478494
rect 85144 471494 85464 478258
rect 85144 471258 85186 471494
rect 85422 471258 85464 471494
rect 85144 464494 85464 471258
rect 85144 464258 85186 464494
rect 85422 464258 85464 464494
rect 85144 457494 85464 464258
rect 85144 457258 85186 457494
rect 85422 457258 85464 457494
rect 85144 450494 85464 457258
rect 85144 450258 85186 450494
rect 85422 450258 85464 450494
rect 85144 443494 85464 450258
rect 85144 443258 85186 443494
rect 85422 443258 85464 443494
rect 85144 436494 85464 443258
rect 85144 436258 85186 436494
rect 85422 436258 85464 436494
rect 85144 429494 85464 436258
rect 85144 429258 85186 429494
rect 85422 429258 85464 429494
rect 85144 422494 85464 429258
rect 85144 422258 85186 422494
rect 85422 422258 85464 422494
rect 85144 415494 85464 422258
rect 85144 415258 85186 415494
rect 85422 415258 85464 415494
rect 85144 408494 85464 415258
rect 85144 408258 85186 408494
rect 85422 408258 85464 408494
rect 85144 401494 85464 408258
rect 85144 401258 85186 401494
rect 85422 401258 85464 401494
rect 85144 394494 85464 401258
rect 85144 394258 85186 394494
rect 85422 394258 85464 394494
rect 85144 387494 85464 394258
rect 85144 387258 85186 387494
rect 85422 387258 85464 387494
rect 85144 380494 85464 387258
rect 85144 380258 85186 380494
rect 85422 380258 85464 380494
rect 85144 373494 85464 380258
rect 85144 373258 85186 373494
rect 85422 373258 85464 373494
rect 85144 366494 85464 373258
rect 85144 366258 85186 366494
rect 85422 366258 85464 366494
rect 85144 359494 85464 366258
rect 85144 359258 85186 359494
rect 85422 359258 85464 359494
rect 85144 352494 85464 359258
rect 85144 352258 85186 352494
rect 85422 352258 85464 352494
rect 85144 345494 85464 352258
rect 85144 345258 85186 345494
rect 85422 345258 85464 345494
rect 85144 338494 85464 345258
rect 85144 338258 85186 338494
rect 85422 338258 85464 338494
rect 85144 331494 85464 338258
rect 85144 331258 85186 331494
rect 85422 331258 85464 331494
rect 85144 324494 85464 331258
rect 85144 324258 85186 324494
rect 85422 324258 85464 324494
rect 85144 317494 85464 324258
rect 85144 317258 85186 317494
rect 85422 317258 85464 317494
rect 85144 310494 85464 317258
rect 85144 310258 85186 310494
rect 85422 310258 85464 310494
rect 85144 303494 85464 310258
rect 85144 303258 85186 303494
rect 85422 303258 85464 303494
rect 85144 296494 85464 303258
rect 85144 296258 85186 296494
rect 85422 296258 85464 296494
rect 85144 289494 85464 296258
rect 85144 289258 85186 289494
rect 85422 289258 85464 289494
rect 85144 282494 85464 289258
rect 85144 282258 85186 282494
rect 85422 282258 85464 282494
rect 85144 275494 85464 282258
rect 85144 275258 85186 275494
rect 85422 275258 85464 275494
rect 85144 268494 85464 275258
rect 85144 268258 85186 268494
rect 85422 268258 85464 268494
rect 85144 261494 85464 268258
rect 85144 261258 85186 261494
rect 85422 261258 85464 261494
rect 85144 254494 85464 261258
rect 85144 254258 85186 254494
rect 85422 254258 85464 254494
rect 85144 247494 85464 254258
rect 85144 247258 85186 247494
rect 85422 247258 85464 247494
rect 85144 240494 85464 247258
rect 85144 240258 85186 240494
rect 85422 240258 85464 240494
rect 85144 233494 85464 240258
rect 85144 233258 85186 233494
rect 85422 233258 85464 233494
rect 85144 226494 85464 233258
rect 85144 226258 85186 226494
rect 85422 226258 85464 226494
rect 85144 219494 85464 226258
rect 85144 219258 85186 219494
rect 85422 219258 85464 219494
rect 85144 212494 85464 219258
rect 85144 212258 85186 212494
rect 85422 212258 85464 212494
rect 85144 205494 85464 212258
rect 85144 205258 85186 205494
rect 85422 205258 85464 205494
rect 85144 198494 85464 205258
rect 85144 198258 85186 198494
rect 85422 198258 85464 198494
rect 85144 191494 85464 198258
rect 85144 191258 85186 191494
rect 85422 191258 85464 191494
rect 85144 184494 85464 191258
rect 85144 184258 85186 184494
rect 85422 184258 85464 184494
rect 85144 177494 85464 184258
rect 85144 177258 85186 177494
rect 85422 177258 85464 177494
rect 85144 170494 85464 177258
rect 85144 170258 85186 170494
rect 85422 170258 85464 170494
rect 85144 163494 85464 170258
rect 85144 163258 85186 163494
rect 85422 163258 85464 163494
rect 85144 156494 85464 163258
rect 85144 156258 85186 156494
rect 85422 156258 85464 156494
rect 85144 149494 85464 156258
rect 85144 149258 85186 149494
rect 85422 149258 85464 149494
rect 85144 142494 85464 149258
rect 85144 142258 85186 142494
rect 85422 142258 85464 142494
rect 85144 135494 85464 142258
rect 85144 135258 85186 135494
rect 85422 135258 85464 135494
rect 85144 128494 85464 135258
rect 85144 128258 85186 128494
rect 85422 128258 85464 128494
rect 85144 121494 85464 128258
rect 85144 121258 85186 121494
rect 85422 121258 85464 121494
rect 85144 114494 85464 121258
rect 85144 114258 85186 114494
rect 85422 114258 85464 114494
rect 85144 107494 85464 114258
rect 85144 107258 85186 107494
rect 85422 107258 85464 107494
rect 85144 100494 85464 107258
rect 85144 100258 85186 100494
rect 85422 100258 85464 100494
rect 85144 93494 85464 100258
rect 85144 93258 85186 93494
rect 85422 93258 85464 93494
rect 85144 86494 85464 93258
rect 85144 86258 85186 86494
rect 85422 86258 85464 86494
rect 85144 79494 85464 86258
rect 85144 79258 85186 79494
rect 85422 79258 85464 79494
rect 85144 72494 85464 79258
rect 85144 72258 85186 72494
rect 85422 72258 85464 72494
rect 85144 65494 85464 72258
rect 85144 65258 85186 65494
rect 85422 65258 85464 65494
rect 85144 58494 85464 65258
rect 85144 58258 85186 58494
rect 85422 58258 85464 58494
rect 85144 51494 85464 58258
rect 85144 51258 85186 51494
rect 85422 51258 85464 51494
rect 85144 44494 85464 51258
rect 85144 44258 85186 44494
rect 85422 44258 85464 44494
rect 85144 37494 85464 44258
rect 85144 37258 85186 37494
rect 85422 37258 85464 37494
rect 85144 30494 85464 37258
rect 85144 30258 85186 30494
rect 85422 30258 85464 30494
rect 85144 23494 85464 30258
rect 85144 23258 85186 23494
rect 85422 23258 85464 23494
rect 85144 16494 85464 23258
rect 85144 16258 85186 16494
rect 85422 16258 85464 16494
rect 85144 9494 85464 16258
rect 85144 9258 85186 9494
rect 85422 9258 85464 9494
rect 85144 2494 85464 9258
rect 85144 2258 85186 2494
rect 85422 2258 85464 2494
rect 85144 -746 85464 2258
rect 85144 -982 85186 -746
rect 85422 -982 85464 -746
rect 85144 -1066 85464 -982
rect 85144 -1302 85186 -1066
rect 85422 -1302 85464 -1066
rect 85144 -2294 85464 -1302
rect 86876 706198 87196 706230
rect 86876 705962 86918 706198
rect 87154 705962 87196 706198
rect 86876 705878 87196 705962
rect 86876 705642 86918 705878
rect 87154 705642 87196 705878
rect 86876 696434 87196 705642
rect 86876 696198 86918 696434
rect 87154 696198 87196 696434
rect 86876 689434 87196 696198
rect 86876 689198 86918 689434
rect 87154 689198 87196 689434
rect 86876 682434 87196 689198
rect 86876 682198 86918 682434
rect 87154 682198 87196 682434
rect 86876 675434 87196 682198
rect 86876 675198 86918 675434
rect 87154 675198 87196 675434
rect 86876 668434 87196 675198
rect 86876 668198 86918 668434
rect 87154 668198 87196 668434
rect 86876 661434 87196 668198
rect 86876 661198 86918 661434
rect 87154 661198 87196 661434
rect 86876 654434 87196 661198
rect 86876 654198 86918 654434
rect 87154 654198 87196 654434
rect 86876 647434 87196 654198
rect 86876 647198 86918 647434
rect 87154 647198 87196 647434
rect 86876 640434 87196 647198
rect 86876 640198 86918 640434
rect 87154 640198 87196 640434
rect 86876 633434 87196 640198
rect 86876 633198 86918 633434
rect 87154 633198 87196 633434
rect 86876 626434 87196 633198
rect 86876 626198 86918 626434
rect 87154 626198 87196 626434
rect 86876 619434 87196 626198
rect 86876 619198 86918 619434
rect 87154 619198 87196 619434
rect 86876 612434 87196 619198
rect 86876 612198 86918 612434
rect 87154 612198 87196 612434
rect 86876 605434 87196 612198
rect 86876 605198 86918 605434
rect 87154 605198 87196 605434
rect 86876 598434 87196 605198
rect 86876 598198 86918 598434
rect 87154 598198 87196 598434
rect 86876 591434 87196 598198
rect 86876 591198 86918 591434
rect 87154 591198 87196 591434
rect 86876 584434 87196 591198
rect 86876 584198 86918 584434
rect 87154 584198 87196 584434
rect 86876 577434 87196 584198
rect 86876 577198 86918 577434
rect 87154 577198 87196 577434
rect 86876 570434 87196 577198
rect 86876 570198 86918 570434
rect 87154 570198 87196 570434
rect 86876 563434 87196 570198
rect 86876 563198 86918 563434
rect 87154 563198 87196 563434
rect 86876 556434 87196 563198
rect 86876 556198 86918 556434
rect 87154 556198 87196 556434
rect 86876 549434 87196 556198
rect 86876 549198 86918 549434
rect 87154 549198 87196 549434
rect 86876 542434 87196 549198
rect 86876 542198 86918 542434
rect 87154 542198 87196 542434
rect 86876 535434 87196 542198
rect 86876 535198 86918 535434
rect 87154 535198 87196 535434
rect 86876 528434 87196 535198
rect 86876 528198 86918 528434
rect 87154 528198 87196 528434
rect 86876 521434 87196 528198
rect 86876 521198 86918 521434
rect 87154 521198 87196 521434
rect 86876 514434 87196 521198
rect 86876 514198 86918 514434
rect 87154 514198 87196 514434
rect 86876 507434 87196 514198
rect 86876 507198 86918 507434
rect 87154 507198 87196 507434
rect 86876 500434 87196 507198
rect 86876 500198 86918 500434
rect 87154 500198 87196 500434
rect 86876 493434 87196 500198
rect 86876 493198 86918 493434
rect 87154 493198 87196 493434
rect 86876 486434 87196 493198
rect 86876 486198 86918 486434
rect 87154 486198 87196 486434
rect 86876 479434 87196 486198
rect 86876 479198 86918 479434
rect 87154 479198 87196 479434
rect 86876 472434 87196 479198
rect 86876 472198 86918 472434
rect 87154 472198 87196 472434
rect 86876 465434 87196 472198
rect 86876 465198 86918 465434
rect 87154 465198 87196 465434
rect 86876 458434 87196 465198
rect 86876 458198 86918 458434
rect 87154 458198 87196 458434
rect 86876 451434 87196 458198
rect 86876 451198 86918 451434
rect 87154 451198 87196 451434
rect 86876 444434 87196 451198
rect 86876 444198 86918 444434
rect 87154 444198 87196 444434
rect 86876 437434 87196 444198
rect 86876 437198 86918 437434
rect 87154 437198 87196 437434
rect 86876 430434 87196 437198
rect 86876 430198 86918 430434
rect 87154 430198 87196 430434
rect 86876 423434 87196 430198
rect 86876 423198 86918 423434
rect 87154 423198 87196 423434
rect 86876 416434 87196 423198
rect 86876 416198 86918 416434
rect 87154 416198 87196 416434
rect 86876 409434 87196 416198
rect 86876 409198 86918 409434
rect 87154 409198 87196 409434
rect 86876 402434 87196 409198
rect 86876 402198 86918 402434
rect 87154 402198 87196 402434
rect 86876 395434 87196 402198
rect 86876 395198 86918 395434
rect 87154 395198 87196 395434
rect 86876 388434 87196 395198
rect 86876 388198 86918 388434
rect 87154 388198 87196 388434
rect 86876 381434 87196 388198
rect 86876 381198 86918 381434
rect 87154 381198 87196 381434
rect 86876 374434 87196 381198
rect 86876 374198 86918 374434
rect 87154 374198 87196 374434
rect 86876 367434 87196 374198
rect 86876 367198 86918 367434
rect 87154 367198 87196 367434
rect 86876 360434 87196 367198
rect 86876 360198 86918 360434
rect 87154 360198 87196 360434
rect 86876 353434 87196 360198
rect 86876 353198 86918 353434
rect 87154 353198 87196 353434
rect 86876 346434 87196 353198
rect 86876 346198 86918 346434
rect 87154 346198 87196 346434
rect 86876 339434 87196 346198
rect 86876 339198 86918 339434
rect 87154 339198 87196 339434
rect 86876 332434 87196 339198
rect 86876 332198 86918 332434
rect 87154 332198 87196 332434
rect 86876 325434 87196 332198
rect 86876 325198 86918 325434
rect 87154 325198 87196 325434
rect 86876 318434 87196 325198
rect 86876 318198 86918 318434
rect 87154 318198 87196 318434
rect 86876 311434 87196 318198
rect 86876 311198 86918 311434
rect 87154 311198 87196 311434
rect 86876 304434 87196 311198
rect 86876 304198 86918 304434
rect 87154 304198 87196 304434
rect 86876 297434 87196 304198
rect 86876 297198 86918 297434
rect 87154 297198 87196 297434
rect 86876 290434 87196 297198
rect 86876 290198 86918 290434
rect 87154 290198 87196 290434
rect 86876 283434 87196 290198
rect 86876 283198 86918 283434
rect 87154 283198 87196 283434
rect 86876 276434 87196 283198
rect 86876 276198 86918 276434
rect 87154 276198 87196 276434
rect 86876 269434 87196 276198
rect 86876 269198 86918 269434
rect 87154 269198 87196 269434
rect 86876 262434 87196 269198
rect 86876 262198 86918 262434
rect 87154 262198 87196 262434
rect 86876 255434 87196 262198
rect 86876 255198 86918 255434
rect 87154 255198 87196 255434
rect 86876 248434 87196 255198
rect 86876 248198 86918 248434
rect 87154 248198 87196 248434
rect 86876 241434 87196 248198
rect 86876 241198 86918 241434
rect 87154 241198 87196 241434
rect 86876 234434 87196 241198
rect 86876 234198 86918 234434
rect 87154 234198 87196 234434
rect 86876 227434 87196 234198
rect 86876 227198 86918 227434
rect 87154 227198 87196 227434
rect 86876 220434 87196 227198
rect 86876 220198 86918 220434
rect 87154 220198 87196 220434
rect 86876 213434 87196 220198
rect 86876 213198 86918 213434
rect 87154 213198 87196 213434
rect 86876 206434 87196 213198
rect 86876 206198 86918 206434
rect 87154 206198 87196 206434
rect 86876 199434 87196 206198
rect 86876 199198 86918 199434
rect 87154 199198 87196 199434
rect 86876 192434 87196 199198
rect 86876 192198 86918 192434
rect 87154 192198 87196 192434
rect 86876 185434 87196 192198
rect 86876 185198 86918 185434
rect 87154 185198 87196 185434
rect 86876 178434 87196 185198
rect 86876 178198 86918 178434
rect 87154 178198 87196 178434
rect 86876 171434 87196 178198
rect 86876 171198 86918 171434
rect 87154 171198 87196 171434
rect 86876 164434 87196 171198
rect 86876 164198 86918 164434
rect 87154 164198 87196 164434
rect 86876 157434 87196 164198
rect 86876 157198 86918 157434
rect 87154 157198 87196 157434
rect 86876 150434 87196 157198
rect 86876 150198 86918 150434
rect 87154 150198 87196 150434
rect 86876 143434 87196 150198
rect 86876 143198 86918 143434
rect 87154 143198 87196 143434
rect 86876 136434 87196 143198
rect 86876 136198 86918 136434
rect 87154 136198 87196 136434
rect 86876 129434 87196 136198
rect 86876 129198 86918 129434
rect 87154 129198 87196 129434
rect 86876 122434 87196 129198
rect 86876 122198 86918 122434
rect 87154 122198 87196 122434
rect 86876 115434 87196 122198
rect 86876 115198 86918 115434
rect 87154 115198 87196 115434
rect 86876 108434 87196 115198
rect 86876 108198 86918 108434
rect 87154 108198 87196 108434
rect 86876 101434 87196 108198
rect 86876 101198 86918 101434
rect 87154 101198 87196 101434
rect 86876 94434 87196 101198
rect 86876 94198 86918 94434
rect 87154 94198 87196 94434
rect 86876 87434 87196 94198
rect 86876 87198 86918 87434
rect 87154 87198 87196 87434
rect 86876 80434 87196 87198
rect 86876 80198 86918 80434
rect 87154 80198 87196 80434
rect 86876 73434 87196 80198
rect 86876 73198 86918 73434
rect 87154 73198 87196 73434
rect 86876 66434 87196 73198
rect 86876 66198 86918 66434
rect 87154 66198 87196 66434
rect 86876 59434 87196 66198
rect 86876 59198 86918 59434
rect 87154 59198 87196 59434
rect 86876 52434 87196 59198
rect 86876 52198 86918 52434
rect 87154 52198 87196 52434
rect 86876 45434 87196 52198
rect 86876 45198 86918 45434
rect 87154 45198 87196 45434
rect 86876 38434 87196 45198
rect 86876 38198 86918 38434
rect 87154 38198 87196 38434
rect 86876 31434 87196 38198
rect 86876 31198 86918 31434
rect 87154 31198 87196 31434
rect 86876 24434 87196 31198
rect 86876 24198 86918 24434
rect 87154 24198 87196 24434
rect 86876 17434 87196 24198
rect 86876 17198 86918 17434
rect 87154 17198 87196 17434
rect 86876 10434 87196 17198
rect 86876 10198 86918 10434
rect 87154 10198 87196 10434
rect 86876 3434 87196 10198
rect 86876 3198 86918 3434
rect 87154 3198 87196 3434
rect 86876 -1706 87196 3198
rect 86876 -1942 86918 -1706
rect 87154 -1942 87196 -1706
rect 86876 -2026 87196 -1942
rect 86876 -2262 86918 -2026
rect 87154 -2262 87196 -2026
rect 86876 -2294 87196 -2262
rect 92144 705238 92464 706230
rect 92144 705002 92186 705238
rect 92422 705002 92464 705238
rect 92144 704918 92464 705002
rect 92144 704682 92186 704918
rect 92422 704682 92464 704918
rect 92144 695494 92464 704682
rect 92144 695258 92186 695494
rect 92422 695258 92464 695494
rect 92144 688494 92464 695258
rect 92144 688258 92186 688494
rect 92422 688258 92464 688494
rect 92144 681494 92464 688258
rect 92144 681258 92186 681494
rect 92422 681258 92464 681494
rect 92144 674494 92464 681258
rect 92144 674258 92186 674494
rect 92422 674258 92464 674494
rect 92144 667494 92464 674258
rect 92144 667258 92186 667494
rect 92422 667258 92464 667494
rect 92144 660494 92464 667258
rect 92144 660258 92186 660494
rect 92422 660258 92464 660494
rect 92144 653494 92464 660258
rect 92144 653258 92186 653494
rect 92422 653258 92464 653494
rect 92144 646494 92464 653258
rect 92144 646258 92186 646494
rect 92422 646258 92464 646494
rect 92144 639494 92464 646258
rect 92144 639258 92186 639494
rect 92422 639258 92464 639494
rect 92144 632494 92464 639258
rect 92144 632258 92186 632494
rect 92422 632258 92464 632494
rect 92144 625494 92464 632258
rect 92144 625258 92186 625494
rect 92422 625258 92464 625494
rect 92144 618494 92464 625258
rect 92144 618258 92186 618494
rect 92422 618258 92464 618494
rect 92144 611494 92464 618258
rect 92144 611258 92186 611494
rect 92422 611258 92464 611494
rect 92144 604494 92464 611258
rect 92144 604258 92186 604494
rect 92422 604258 92464 604494
rect 92144 597494 92464 604258
rect 92144 597258 92186 597494
rect 92422 597258 92464 597494
rect 92144 590494 92464 597258
rect 92144 590258 92186 590494
rect 92422 590258 92464 590494
rect 92144 583494 92464 590258
rect 92144 583258 92186 583494
rect 92422 583258 92464 583494
rect 92144 576494 92464 583258
rect 92144 576258 92186 576494
rect 92422 576258 92464 576494
rect 92144 569494 92464 576258
rect 92144 569258 92186 569494
rect 92422 569258 92464 569494
rect 92144 562494 92464 569258
rect 92144 562258 92186 562494
rect 92422 562258 92464 562494
rect 92144 555494 92464 562258
rect 92144 555258 92186 555494
rect 92422 555258 92464 555494
rect 92144 548494 92464 555258
rect 92144 548258 92186 548494
rect 92422 548258 92464 548494
rect 92144 541494 92464 548258
rect 92144 541258 92186 541494
rect 92422 541258 92464 541494
rect 92144 534494 92464 541258
rect 92144 534258 92186 534494
rect 92422 534258 92464 534494
rect 92144 527494 92464 534258
rect 92144 527258 92186 527494
rect 92422 527258 92464 527494
rect 92144 520494 92464 527258
rect 92144 520258 92186 520494
rect 92422 520258 92464 520494
rect 92144 513494 92464 520258
rect 92144 513258 92186 513494
rect 92422 513258 92464 513494
rect 92144 506494 92464 513258
rect 92144 506258 92186 506494
rect 92422 506258 92464 506494
rect 92144 499494 92464 506258
rect 92144 499258 92186 499494
rect 92422 499258 92464 499494
rect 92144 492494 92464 499258
rect 92144 492258 92186 492494
rect 92422 492258 92464 492494
rect 92144 485494 92464 492258
rect 92144 485258 92186 485494
rect 92422 485258 92464 485494
rect 92144 478494 92464 485258
rect 92144 478258 92186 478494
rect 92422 478258 92464 478494
rect 92144 471494 92464 478258
rect 92144 471258 92186 471494
rect 92422 471258 92464 471494
rect 92144 464494 92464 471258
rect 92144 464258 92186 464494
rect 92422 464258 92464 464494
rect 92144 457494 92464 464258
rect 92144 457258 92186 457494
rect 92422 457258 92464 457494
rect 92144 450494 92464 457258
rect 92144 450258 92186 450494
rect 92422 450258 92464 450494
rect 92144 443494 92464 450258
rect 92144 443258 92186 443494
rect 92422 443258 92464 443494
rect 92144 436494 92464 443258
rect 92144 436258 92186 436494
rect 92422 436258 92464 436494
rect 92144 429494 92464 436258
rect 92144 429258 92186 429494
rect 92422 429258 92464 429494
rect 92144 422494 92464 429258
rect 92144 422258 92186 422494
rect 92422 422258 92464 422494
rect 92144 415494 92464 422258
rect 92144 415258 92186 415494
rect 92422 415258 92464 415494
rect 92144 408494 92464 415258
rect 92144 408258 92186 408494
rect 92422 408258 92464 408494
rect 92144 401494 92464 408258
rect 92144 401258 92186 401494
rect 92422 401258 92464 401494
rect 92144 394494 92464 401258
rect 92144 394258 92186 394494
rect 92422 394258 92464 394494
rect 92144 387494 92464 394258
rect 92144 387258 92186 387494
rect 92422 387258 92464 387494
rect 92144 380494 92464 387258
rect 92144 380258 92186 380494
rect 92422 380258 92464 380494
rect 92144 373494 92464 380258
rect 92144 373258 92186 373494
rect 92422 373258 92464 373494
rect 92144 366494 92464 373258
rect 92144 366258 92186 366494
rect 92422 366258 92464 366494
rect 92144 359494 92464 366258
rect 92144 359258 92186 359494
rect 92422 359258 92464 359494
rect 92144 352494 92464 359258
rect 92144 352258 92186 352494
rect 92422 352258 92464 352494
rect 92144 345494 92464 352258
rect 92144 345258 92186 345494
rect 92422 345258 92464 345494
rect 92144 338494 92464 345258
rect 92144 338258 92186 338494
rect 92422 338258 92464 338494
rect 92144 331494 92464 338258
rect 92144 331258 92186 331494
rect 92422 331258 92464 331494
rect 92144 324494 92464 331258
rect 92144 324258 92186 324494
rect 92422 324258 92464 324494
rect 92144 317494 92464 324258
rect 92144 317258 92186 317494
rect 92422 317258 92464 317494
rect 92144 310494 92464 317258
rect 92144 310258 92186 310494
rect 92422 310258 92464 310494
rect 92144 303494 92464 310258
rect 92144 303258 92186 303494
rect 92422 303258 92464 303494
rect 92144 296494 92464 303258
rect 92144 296258 92186 296494
rect 92422 296258 92464 296494
rect 92144 289494 92464 296258
rect 92144 289258 92186 289494
rect 92422 289258 92464 289494
rect 92144 282494 92464 289258
rect 92144 282258 92186 282494
rect 92422 282258 92464 282494
rect 92144 275494 92464 282258
rect 92144 275258 92186 275494
rect 92422 275258 92464 275494
rect 92144 268494 92464 275258
rect 92144 268258 92186 268494
rect 92422 268258 92464 268494
rect 92144 261494 92464 268258
rect 92144 261258 92186 261494
rect 92422 261258 92464 261494
rect 92144 254494 92464 261258
rect 92144 254258 92186 254494
rect 92422 254258 92464 254494
rect 92144 247494 92464 254258
rect 92144 247258 92186 247494
rect 92422 247258 92464 247494
rect 92144 240494 92464 247258
rect 92144 240258 92186 240494
rect 92422 240258 92464 240494
rect 92144 233494 92464 240258
rect 92144 233258 92186 233494
rect 92422 233258 92464 233494
rect 92144 226494 92464 233258
rect 92144 226258 92186 226494
rect 92422 226258 92464 226494
rect 92144 219494 92464 226258
rect 92144 219258 92186 219494
rect 92422 219258 92464 219494
rect 92144 212494 92464 219258
rect 92144 212258 92186 212494
rect 92422 212258 92464 212494
rect 92144 205494 92464 212258
rect 92144 205258 92186 205494
rect 92422 205258 92464 205494
rect 92144 198494 92464 205258
rect 92144 198258 92186 198494
rect 92422 198258 92464 198494
rect 92144 191494 92464 198258
rect 92144 191258 92186 191494
rect 92422 191258 92464 191494
rect 92144 184494 92464 191258
rect 92144 184258 92186 184494
rect 92422 184258 92464 184494
rect 92144 177494 92464 184258
rect 92144 177258 92186 177494
rect 92422 177258 92464 177494
rect 92144 170494 92464 177258
rect 92144 170258 92186 170494
rect 92422 170258 92464 170494
rect 92144 163494 92464 170258
rect 92144 163258 92186 163494
rect 92422 163258 92464 163494
rect 92144 156494 92464 163258
rect 92144 156258 92186 156494
rect 92422 156258 92464 156494
rect 92144 149494 92464 156258
rect 92144 149258 92186 149494
rect 92422 149258 92464 149494
rect 92144 142494 92464 149258
rect 92144 142258 92186 142494
rect 92422 142258 92464 142494
rect 92144 135494 92464 142258
rect 92144 135258 92186 135494
rect 92422 135258 92464 135494
rect 92144 128494 92464 135258
rect 92144 128258 92186 128494
rect 92422 128258 92464 128494
rect 92144 121494 92464 128258
rect 92144 121258 92186 121494
rect 92422 121258 92464 121494
rect 92144 114494 92464 121258
rect 92144 114258 92186 114494
rect 92422 114258 92464 114494
rect 92144 107494 92464 114258
rect 92144 107258 92186 107494
rect 92422 107258 92464 107494
rect 92144 100494 92464 107258
rect 92144 100258 92186 100494
rect 92422 100258 92464 100494
rect 92144 93494 92464 100258
rect 92144 93258 92186 93494
rect 92422 93258 92464 93494
rect 92144 86494 92464 93258
rect 92144 86258 92186 86494
rect 92422 86258 92464 86494
rect 92144 79494 92464 86258
rect 92144 79258 92186 79494
rect 92422 79258 92464 79494
rect 92144 72494 92464 79258
rect 92144 72258 92186 72494
rect 92422 72258 92464 72494
rect 92144 65494 92464 72258
rect 92144 65258 92186 65494
rect 92422 65258 92464 65494
rect 92144 58494 92464 65258
rect 92144 58258 92186 58494
rect 92422 58258 92464 58494
rect 92144 51494 92464 58258
rect 92144 51258 92186 51494
rect 92422 51258 92464 51494
rect 92144 44494 92464 51258
rect 92144 44258 92186 44494
rect 92422 44258 92464 44494
rect 92144 37494 92464 44258
rect 92144 37258 92186 37494
rect 92422 37258 92464 37494
rect 92144 30494 92464 37258
rect 92144 30258 92186 30494
rect 92422 30258 92464 30494
rect 92144 23494 92464 30258
rect 92144 23258 92186 23494
rect 92422 23258 92464 23494
rect 92144 16494 92464 23258
rect 92144 16258 92186 16494
rect 92422 16258 92464 16494
rect 92144 9494 92464 16258
rect 92144 9258 92186 9494
rect 92422 9258 92464 9494
rect 92144 2494 92464 9258
rect 92144 2258 92186 2494
rect 92422 2258 92464 2494
rect 92144 -746 92464 2258
rect 92144 -982 92186 -746
rect 92422 -982 92464 -746
rect 92144 -1066 92464 -982
rect 92144 -1302 92186 -1066
rect 92422 -1302 92464 -1066
rect 92144 -2294 92464 -1302
rect 93876 706198 94196 706230
rect 93876 705962 93918 706198
rect 94154 705962 94196 706198
rect 93876 705878 94196 705962
rect 93876 705642 93918 705878
rect 94154 705642 94196 705878
rect 93876 696434 94196 705642
rect 93876 696198 93918 696434
rect 94154 696198 94196 696434
rect 93876 689434 94196 696198
rect 93876 689198 93918 689434
rect 94154 689198 94196 689434
rect 93876 682434 94196 689198
rect 93876 682198 93918 682434
rect 94154 682198 94196 682434
rect 93876 675434 94196 682198
rect 93876 675198 93918 675434
rect 94154 675198 94196 675434
rect 93876 668434 94196 675198
rect 93876 668198 93918 668434
rect 94154 668198 94196 668434
rect 93876 661434 94196 668198
rect 93876 661198 93918 661434
rect 94154 661198 94196 661434
rect 93876 654434 94196 661198
rect 93876 654198 93918 654434
rect 94154 654198 94196 654434
rect 93876 647434 94196 654198
rect 93876 647198 93918 647434
rect 94154 647198 94196 647434
rect 93876 640434 94196 647198
rect 93876 640198 93918 640434
rect 94154 640198 94196 640434
rect 93876 633434 94196 640198
rect 93876 633198 93918 633434
rect 94154 633198 94196 633434
rect 93876 626434 94196 633198
rect 93876 626198 93918 626434
rect 94154 626198 94196 626434
rect 93876 619434 94196 626198
rect 93876 619198 93918 619434
rect 94154 619198 94196 619434
rect 93876 612434 94196 619198
rect 93876 612198 93918 612434
rect 94154 612198 94196 612434
rect 93876 605434 94196 612198
rect 93876 605198 93918 605434
rect 94154 605198 94196 605434
rect 93876 598434 94196 605198
rect 93876 598198 93918 598434
rect 94154 598198 94196 598434
rect 93876 591434 94196 598198
rect 93876 591198 93918 591434
rect 94154 591198 94196 591434
rect 93876 584434 94196 591198
rect 93876 584198 93918 584434
rect 94154 584198 94196 584434
rect 93876 577434 94196 584198
rect 93876 577198 93918 577434
rect 94154 577198 94196 577434
rect 93876 570434 94196 577198
rect 93876 570198 93918 570434
rect 94154 570198 94196 570434
rect 93876 563434 94196 570198
rect 93876 563198 93918 563434
rect 94154 563198 94196 563434
rect 93876 556434 94196 563198
rect 93876 556198 93918 556434
rect 94154 556198 94196 556434
rect 93876 549434 94196 556198
rect 93876 549198 93918 549434
rect 94154 549198 94196 549434
rect 93876 542434 94196 549198
rect 93876 542198 93918 542434
rect 94154 542198 94196 542434
rect 93876 535434 94196 542198
rect 93876 535198 93918 535434
rect 94154 535198 94196 535434
rect 93876 528434 94196 535198
rect 93876 528198 93918 528434
rect 94154 528198 94196 528434
rect 93876 521434 94196 528198
rect 93876 521198 93918 521434
rect 94154 521198 94196 521434
rect 93876 514434 94196 521198
rect 93876 514198 93918 514434
rect 94154 514198 94196 514434
rect 93876 507434 94196 514198
rect 93876 507198 93918 507434
rect 94154 507198 94196 507434
rect 93876 500434 94196 507198
rect 93876 500198 93918 500434
rect 94154 500198 94196 500434
rect 93876 493434 94196 500198
rect 93876 493198 93918 493434
rect 94154 493198 94196 493434
rect 93876 486434 94196 493198
rect 93876 486198 93918 486434
rect 94154 486198 94196 486434
rect 93876 479434 94196 486198
rect 93876 479198 93918 479434
rect 94154 479198 94196 479434
rect 93876 472434 94196 479198
rect 93876 472198 93918 472434
rect 94154 472198 94196 472434
rect 93876 465434 94196 472198
rect 93876 465198 93918 465434
rect 94154 465198 94196 465434
rect 93876 458434 94196 465198
rect 93876 458198 93918 458434
rect 94154 458198 94196 458434
rect 93876 451434 94196 458198
rect 93876 451198 93918 451434
rect 94154 451198 94196 451434
rect 93876 444434 94196 451198
rect 93876 444198 93918 444434
rect 94154 444198 94196 444434
rect 93876 437434 94196 444198
rect 93876 437198 93918 437434
rect 94154 437198 94196 437434
rect 93876 430434 94196 437198
rect 93876 430198 93918 430434
rect 94154 430198 94196 430434
rect 93876 423434 94196 430198
rect 93876 423198 93918 423434
rect 94154 423198 94196 423434
rect 93876 416434 94196 423198
rect 93876 416198 93918 416434
rect 94154 416198 94196 416434
rect 93876 409434 94196 416198
rect 93876 409198 93918 409434
rect 94154 409198 94196 409434
rect 93876 402434 94196 409198
rect 93876 402198 93918 402434
rect 94154 402198 94196 402434
rect 93876 395434 94196 402198
rect 93876 395198 93918 395434
rect 94154 395198 94196 395434
rect 93876 388434 94196 395198
rect 93876 388198 93918 388434
rect 94154 388198 94196 388434
rect 93876 381434 94196 388198
rect 93876 381198 93918 381434
rect 94154 381198 94196 381434
rect 93876 374434 94196 381198
rect 93876 374198 93918 374434
rect 94154 374198 94196 374434
rect 93876 367434 94196 374198
rect 93876 367198 93918 367434
rect 94154 367198 94196 367434
rect 93876 360434 94196 367198
rect 93876 360198 93918 360434
rect 94154 360198 94196 360434
rect 93876 353434 94196 360198
rect 93876 353198 93918 353434
rect 94154 353198 94196 353434
rect 93876 346434 94196 353198
rect 93876 346198 93918 346434
rect 94154 346198 94196 346434
rect 93876 339434 94196 346198
rect 93876 339198 93918 339434
rect 94154 339198 94196 339434
rect 93876 332434 94196 339198
rect 93876 332198 93918 332434
rect 94154 332198 94196 332434
rect 93876 325434 94196 332198
rect 93876 325198 93918 325434
rect 94154 325198 94196 325434
rect 93876 318434 94196 325198
rect 93876 318198 93918 318434
rect 94154 318198 94196 318434
rect 93876 311434 94196 318198
rect 93876 311198 93918 311434
rect 94154 311198 94196 311434
rect 93876 304434 94196 311198
rect 93876 304198 93918 304434
rect 94154 304198 94196 304434
rect 93876 297434 94196 304198
rect 93876 297198 93918 297434
rect 94154 297198 94196 297434
rect 93876 290434 94196 297198
rect 93876 290198 93918 290434
rect 94154 290198 94196 290434
rect 93876 283434 94196 290198
rect 93876 283198 93918 283434
rect 94154 283198 94196 283434
rect 93876 276434 94196 283198
rect 93876 276198 93918 276434
rect 94154 276198 94196 276434
rect 93876 269434 94196 276198
rect 93876 269198 93918 269434
rect 94154 269198 94196 269434
rect 93876 262434 94196 269198
rect 93876 262198 93918 262434
rect 94154 262198 94196 262434
rect 93876 255434 94196 262198
rect 93876 255198 93918 255434
rect 94154 255198 94196 255434
rect 93876 248434 94196 255198
rect 93876 248198 93918 248434
rect 94154 248198 94196 248434
rect 93876 241434 94196 248198
rect 93876 241198 93918 241434
rect 94154 241198 94196 241434
rect 93876 234434 94196 241198
rect 93876 234198 93918 234434
rect 94154 234198 94196 234434
rect 93876 227434 94196 234198
rect 93876 227198 93918 227434
rect 94154 227198 94196 227434
rect 93876 220434 94196 227198
rect 93876 220198 93918 220434
rect 94154 220198 94196 220434
rect 93876 213434 94196 220198
rect 93876 213198 93918 213434
rect 94154 213198 94196 213434
rect 93876 206434 94196 213198
rect 93876 206198 93918 206434
rect 94154 206198 94196 206434
rect 93876 199434 94196 206198
rect 93876 199198 93918 199434
rect 94154 199198 94196 199434
rect 93876 192434 94196 199198
rect 93876 192198 93918 192434
rect 94154 192198 94196 192434
rect 93876 185434 94196 192198
rect 93876 185198 93918 185434
rect 94154 185198 94196 185434
rect 93876 178434 94196 185198
rect 93876 178198 93918 178434
rect 94154 178198 94196 178434
rect 93876 171434 94196 178198
rect 93876 171198 93918 171434
rect 94154 171198 94196 171434
rect 93876 164434 94196 171198
rect 93876 164198 93918 164434
rect 94154 164198 94196 164434
rect 93876 157434 94196 164198
rect 93876 157198 93918 157434
rect 94154 157198 94196 157434
rect 93876 150434 94196 157198
rect 93876 150198 93918 150434
rect 94154 150198 94196 150434
rect 93876 143434 94196 150198
rect 93876 143198 93918 143434
rect 94154 143198 94196 143434
rect 93876 136434 94196 143198
rect 93876 136198 93918 136434
rect 94154 136198 94196 136434
rect 93876 129434 94196 136198
rect 93876 129198 93918 129434
rect 94154 129198 94196 129434
rect 93876 122434 94196 129198
rect 93876 122198 93918 122434
rect 94154 122198 94196 122434
rect 93876 115434 94196 122198
rect 93876 115198 93918 115434
rect 94154 115198 94196 115434
rect 93876 108434 94196 115198
rect 93876 108198 93918 108434
rect 94154 108198 94196 108434
rect 93876 101434 94196 108198
rect 93876 101198 93918 101434
rect 94154 101198 94196 101434
rect 93876 94434 94196 101198
rect 93876 94198 93918 94434
rect 94154 94198 94196 94434
rect 93876 87434 94196 94198
rect 93876 87198 93918 87434
rect 94154 87198 94196 87434
rect 93876 80434 94196 87198
rect 93876 80198 93918 80434
rect 94154 80198 94196 80434
rect 93876 73434 94196 80198
rect 93876 73198 93918 73434
rect 94154 73198 94196 73434
rect 93876 66434 94196 73198
rect 93876 66198 93918 66434
rect 94154 66198 94196 66434
rect 93876 59434 94196 66198
rect 93876 59198 93918 59434
rect 94154 59198 94196 59434
rect 93876 52434 94196 59198
rect 93876 52198 93918 52434
rect 94154 52198 94196 52434
rect 93876 45434 94196 52198
rect 93876 45198 93918 45434
rect 94154 45198 94196 45434
rect 93876 38434 94196 45198
rect 93876 38198 93918 38434
rect 94154 38198 94196 38434
rect 93876 31434 94196 38198
rect 93876 31198 93918 31434
rect 94154 31198 94196 31434
rect 93876 24434 94196 31198
rect 93876 24198 93918 24434
rect 94154 24198 94196 24434
rect 93876 17434 94196 24198
rect 93876 17198 93918 17434
rect 94154 17198 94196 17434
rect 93876 10434 94196 17198
rect 93876 10198 93918 10434
rect 94154 10198 94196 10434
rect 93876 3434 94196 10198
rect 93876 3198 93918 3434
rect 94154 3198 94196 3434
rect 93876 -1706 94196 3198
rect 93876 -1942 93918 -1706
rect 94154 -1942 94196 -1706
rect 93876 -2026 94196 -1942
rect 93876 -2262 93918 -2026
rect 94154 -2262 94196 -2026
rect 93876 -2294 94196 -2262
rect 99144 705238 99464 706230
rect 99144 705002 99186 705238
rect 99422 705002 99464 705238
rect 99144 704918 99464 705002
rect 99144 704682 99186 704918
rect 99422 704682 99464 704918
rect 99144 695494 99464 704682
rect 99144 695258 99186 695494
rect 99422 695258 99464 695494
rect 99144 688494 99464 695258
rect 99144 688258 99186 688494
rect 99422 688258 99464 688494
rect 99144 681494 99464 688258
rect 99144 681258 99186 681494
rect 99422 681258 99464 681494
rect 99144 674494 99464 681258
rect 99144 674258 99186 674494
rect 99422 674258 99464 674494
rect 99144 667494 99464 674258
rect 99144 667258 99186 667494
rect 99422 667258 99464 667494
rect 99144 660494 99464 667258
rect 99144 660258 99186 660494
rect 99422 660258 99464 660494
rect 99144 653494 99464 660258
rect 99144 653258 99186 653494
rect 99422 653258 99464 653494
rect 99144 646494 99464 653258
rect 99144 646258 99186 646494
rect 99422 646258 99464 646494
rect 99144 639494 99464 646258
rect 99144 639258 99186 639494
rect 99422 639258 99464 639494
rect 99144 632494 99464 639258
rect 99144 632258 99186 632494
rect 99422 632258 99464 632494
rect 99144 625494 99464 632258
rect 99144 625258 99186 625494
rect 99422 625258 99464 625494
rect 99144 618494 99464 625258
rect 99144 618258 99186 618494
rect 99422 618258 99464 618494
rect 99144 611494 99464 618258
rect 99144 611258 99186 611494
rect 99422 611258 99464 611494
rect 99144 604494 99464 611258
rect 99144 604258 99186 604494
rect 99422 604258 99464 604494
rect 99144 597494 99464 604258
rect 99144 597258 99186 597494
rect 99422 597258 99464 597494
rect 99144 590494 99464 597258
rect 99144 590258 99186 590494
rect 99422 590258 99464 590494
rect 99144 583494 99464 590258
rect 99144 583258 99186 583494
rect 99422 583258 99464 583494
rect 99144 576494 99464 583258
rect 99144 576258 99186 576494
rect 99422 576258 99464 576494
rect 99144 569494 99464 576258
rect 99144 569258 99186 569494
rect 99422 569258 99464 569494
rect 99144 562494 99464 569258
rect 99144 562258 99186 562494
rect 99422 562258 99464 562494
rect 99144 555494 99464 562258
rect 99144 555258 99186 555494
rect 99422 555258 99464 555494
rect 99144 548494 99464 555258
rect 99144 548258 99186 548494
rect 99422 548258 99464 548494
rect 99144 541494 99464 548258
rect 99144 541258 99186 541494
rect 99422 541258 99464 541494
rect 99144 534494 99464 541258
rect 99144 534258 99186 534494
rect 99422 534258 99464 534494
rect 99144 527494 99464 534258
rect 99144 527258 99186 527494
rect 99422 527258 99464 527494
rect 99144 520494 99464 527258
rect 99144 520258 99186 520494
rect 99422 520258 99464 520494
rect 99144 513494 99464 520258
rect 99144 513258 99186 513494
rect 99422 513258 99464 513494
rect 99144 506494 99464 513258
rect 99144 506258 99186 506494
rect 99422 506258 99464 506494
rect 99144 499494 99464 506258
rect 99144 499258 99186 499494
rect 99422 499258 99464 499494
rect 99144 492494 99464 499258
rect 99144 492258 99186 492494
rect 99422 492258 99464 492494
rect 99144 485494 99464 492258
rect 99144 485258 99186 485494
rect 99422 485258 99464 485494
rect 99144 478494 99464 485258
rect 99144 478258 99186 478494
rect 99422 478258 99464 478494
rect 99144 471494 99464 478258
rect 99144 471258 99186 471494
rect 99422 471258 99464 471494
rect 99144 464494 99464 471258
rect 99144 464258 99186 464494
rect 99422 464258 99464 464494
rect 99144 457494 99464 464258
rect 99144 457258 99186 457494
rect 99422 457258 99464 457494
rect 99144 450494 99464 457258
rect 99144 450258 99186 450494
rect 99422 450258 99464 450494
rect 99144 443494 99464 450258
rect 99144 443258 99186 443494
rect 99422 443258 99464 443494
rect 99144 436494 99464 443258
rect 99144 436258 99186 436494
rect 99422 436258 99464 436494
rect 99144 429494 99464 436258
rect 99144 429258 99186 429494
rect 99422 429258 99464 429494
rect 99144 422494 99464 429258
rect 99144 422258 99186 422494
rect 99422 422258 99464 422494
rect 99144 415494 99464 422258
rect 99144 415258 99186 415494
rect 99422 415258 99464 415494
rect 99144 408494 99464 415258
rect 99144 408258 99186 408494
rect 99422 408258 99464 408494
rect 99144 401494 99464 408258
rect 99144 401258 99186 401494
rect 99422 401258 99464 401494
rect 99144 394494 99464 401258
rect 99144 394258 99186 394494
rect 99422 394258 99464 394494
rect 99144 387494 99464 394258
rect 99144 387258 99186 387494
rect 99422 387258 99464 387494
rect 99144 380494 99464 387258
rect 99144 380258 99186 380494
rect 99422 380258 99464 380494
rect 99144 373494 99464 380258
rect 99144 373258 99186 373494
rect 99422 373258 99464 373494
rect 99144 366494 99464 373258
rect 99144 366258 99186 366494
rect 99422 366258 99464 366494
rect 99144 359494 99464 366258
rect 99144 359258 99186 359494
rect 99422 359258 99464 359494
rect 99144 352494 99464 359258
rect 99144 352258 99186 352494
rect 99422 352258 99464 352494
rect 99144 345494 99464 352258
rect 99144 345258 99186 345494
rect 99422 345258 99464 345494
rect 99144 338494 99464 345258
rect 99144 338258 99186 338494
rect 99422 338258 99464 338494
rect 99144 331494 99464 338258
rect 99144 331258 99186 331494
rect 99422 331258 99464 331494
rect 99144 324494 99464 331258
rect 99144 324258 99186 324494
rect 99422 324258 99464 324494
rect 99144 317494 99464 324258
rect 99144 317258 99186 317494
rect 99422 317258 99464 317494
rect 99144 310494 99464 317258
rect 99144 310258 99186 310494
rect 99422 310258 99464 310494
rect 99144 303494 99464 310258
rect 99144 303258 99186 303494
rect 99422 303258 99464 303494
rect 99144 296494 99464 303258
rect 99144 296258 99186 296494
rect 99422 296258 99464 296494
rect 99144 289494 99464 296258
rect 99144 289258 99186 289494
rect 99422 289258 99464 289494
rect 99144 282494 99464 289258
rect 99144 282258 99186 282494
rect 99422 282258 99464 282494
rect 99144 275494 99464 282258
rect 99144 275258 99186 275494
rect 99422 275258 99464 275494
rect 99144 268494 99464 275258
rect 99144 268258 99186 268494
rect 99422 268258 99464 268494
rect 99144 261494 99464 268258
rect 99144 261258 99186 261494
rect 99422 261258 99464 261494
rect 99144 254494 99464 261258
rect 99144 254258 99186 254494
rect 99422 254258 99464 254494
rect 99144 247494 99464 254258
rect 99144 247258 99186 247494
rect 99422 247258 99464 247494
rect 99144 240494 99464 247258
rect 99144 240258 99186 240494
rect 99422 240258 99464 240494
rect 99144 233494 99464 240258
rect 99144 233258 99186 233494
rect 99422 233258 99464 233494
rect 99144 226494 99464 233258
rect 99144 226258 99186 226494
rect 99422 226258 99464 226494
rect 99144 219494 99464 226258
rect 99144 219258 99186 219494
rect 99422 219258 99464 219494
rect 99144 212494 99464 219258
rect 99144 212258 99186 212494
rect 99422 212258 99464 212494
rect 99144 205494 99464 212258
rect 99144 205258 99186 205494
rect 99422 205258 99464 205494
rect 99144 198494 99464 205258
rect 99144 198258 99186 198494
rect 99422 198258 99464 198494
rect 99144 191494 99464 198258
rect 99144 191258 99186 191494
rect 99422 191258 99464 191494
rect 99144 184494 99464 191258
rect 99144 184258 99186 184494
rect 99422 184258 99464 184494
rect 99144 177494 99464 184258
rect 99144 177258 99186 177494
rect 99422 177258 99464 177494
rect 99144 170494 99464 177258
rect 99144 170258 99186 170494
rect 99422 170258 99464 170494
rect 99144 163494 99464 170258
rect 99144 163258 99186 163494
rect 99422 163258 99464 163494
rect 99144 156494 99464 163258
rect 99144 156258 99186 156494
rect 99422 156258 99464 156494
rect 99144 149494 99464 156258
rect 99144 149258 99186 149494
rect 99422 149258 99464 149494
rect 99144 142494 99464 149258
rect 99144 142258 99186 142494
rect 99422 142258 99464 142494
rect 99144 135494 99464 142258
rect 99144 135258 99186 135494
rect 99422 135258 99464 135494
rect 99144 128494 99464 135258
rect 99144 128258 99186 128494
rect 99422 128258 99464 128494
rect 99144 121494 99464 128258
rect 99144 121258 99186 121494
rect 99422 121258 99464 121494
rect 99144 114494 99464 121258
rect 99144 114258 99186 114494
rect 99422 114258 99464 114494
rect 99144 107494 99464 114258
rect 99144 107258 99186 107494
rect 99422 107258 99464 107494
rect 99144 100494 99464 107258
rect 99144 100258 99186 100494
rect 99422 100258 99464 100494
rect 99144 93494 99464 100258
rect 99144 93258 99186 93494
rect 99422 93258 99464 93494
rect 99144 86494 99464 93258
rect 99144 86258 99186 86494
rect 99422 86258 99464 86494
rect 99144 79494 99464 86258
rect 99144 79258 99186 79494
rect 99422 79258 99464 79494
rect 99144 72494 99464 79258
rect 99144 72258 99186 72494
rect 99422 72258 99464 72494
rect 99144 65494 99464 72258
rect 99144 65258 99186 65494
rect 99422 65258 99464 65494
rect 99144 58494 99464 65258
rect 99144 58258 99186 58494
rect 99422 58258 99464 58494
rect 99144 51494 99464 58258
rect 99144 51258 99186 51494
rect 99422 51258 99464 51494
rect 99144 44494 99464 51258
rect 99144 44258 99186 44494
rect 99422 44258 99464 44494
rect 99144 37494 99464 44258
rect 99144 37258 99186 37494
rect 99422 37258 99464 37494
rect 99144 30494 99464 37258
rect 99144 30258 99186 30494
rect 99422 30258 99464 30494
rect 99144 23494 99464 30258
rect 99144 23258 99186 23494
rect 99422 23258 99464 23494
rect 99144 16494 99464 23258
rect 99144 16258 99186 16494
rect 99422 16258 99464 16494
rect 99144 9494 99464 16258
rect 99144 9258 99186 9494
rect 99422 9258 99464 9494
rect 99144 2494 99464 9258
rect 99144 2258 99186 2494
rect 99422 2258 99464 2494
rect 99144 -746 99464 2258
rect 99144 -982 99186 -746
rect 99422 -982 99464 -746
rect 99144 -1066 99464 -982
rect 99144 -1302 99186 -1066
rect 99422 -1302 99464 -1066
rect 99144 -2294 99464 -1302
rect 100876 706198 101196 706230
rect 100876 705962 100918 706198
rect 101154 705962 101196 706198
rect 100876 705878 101196 705962
rect 100876 705642 100918 705878
rect 101154 705642 101196 705878
rect 100876 696434 101196 705642
rect 100876 696198 100918 696434
rect 101154 696198 101196 696434
rect 100876 689434 101196 696198
rect 100876 689198 100918 689434
rect 101154 689198 101196 689434
rect 100876 682434 101196 689198
rect 100876 682198 100918 682434
rect 101154 682198 101196 682434
rect 100876 675434 101196 682198
rect 100876 675198 100918 675434
rect 101154 675198 101196 675434
rect 100876 668434 101196 675198
rect 100876 668198 100918 668434
rect 101154 668198 101196 668434
rect 100876 661434 101196 668198
rect 100876 661198 100918 661434
rect 101154 661198 101196 661434
rect 100876 654434 101196 661198
rect 100876 654198 100918 654434
rect 101154 654198 101196 654434
rect 100876 647434 101196 654198
rect 100876 647198 100918 647434
rect 101154 647198 101196 647434
rect 100876 640434 101196 647198
rect 100876 640198 100918 640434
rect 101154 640198 101196 640434
rect 100876 633434 101196 640198
rect 100876 633198 100918 633434
rect 101154 633198 101196 633434
rect 100876 626434 101196 633198
rect 100876 626198 100918 626434
rect 101154 626198 101196 626434
rect 100876 619434 101196 626198
rect 100876 619198 100918 619434
rect 101154 619198 101196 619434
rect 100876 612434 101196 619198
rect 100876 612198 100918 612434
rect 101154 612198 101196 612434
rect 100876 605434 101196 612198
rect 100876 605198 100918 605434
rect 101154 605198 101196 605434
rect 100876 598434 101196 605198
rect 100876 598198 100918 598434
rect 101154 598198 101196 598434
rect 100876 591434 101196 598198
rect 100876 591198 100918 591434
rect 101154 591198 101196 591434
rect 100876 584434 101196 591198
rect 100876 584198 100918 584434
rect 101154 584198 101196 584434
rect 100876 577434 101196 584198
rect 100876 577198 100918 577434
rect 101154 577198 101196 577434
rect 100876 570434 101196 577198
rect 100876 570198 100918 570434
rect 101154 570198 101196 570434
rect 100876 563434 101196 570198
rect 100876 563198 100918 563434
rect 101154 563198 101196 563434
rect 100876 556434 101196 563198
rect 100876 556198 100918 556434
rect 101154 556198 101196 556434
rect 100876 549434 101196 556198
rect 100876 549198 100918 549434
rect 101154 549198 101196 549434
rect 100876 542434 101196 549198
rect 100876 542198 100918 542434
rect 101154 542198 101196 542434
rect 100876 535434 101196 542198
rect 100876 535198 100918 535434
rect 101154 535198 101196 535434
rect 100876 528434 101196 535198
rect 100876 528198 100918 528434
rect 101154 528198 101196 528434
rect 100876 521434 101196 528198
rect 100876 521198 100918 521434
rect 101154 521198 101196 521434
rect 100876 514434 101196 521198
rect 100876 514198 100918 514434
rect 101154 514198 101196 514434
rect 100876 507434 101196 514198
rect 100876 507198 100918 507434
rect 101154 507198 101196 507434
rect 100876 500434 101196 507198
rect 100876 500198 100918 500434
rect 101154 500198 101196 500434
rect 100876 493434 101196 500198
rect 100876 493198 100918 493434
rect 101154 493198 101196 493434
rect 100876 486434 101196 493198
rect 100876 486198 100918 486434
rect 101154 486198 101196 486434
rect 100876 479434 101196 486198
rect 100876 479198 100918 479434
rect 101154 479198 101196 479434
rect 100876 472434 101196 479198
rect 100876 472198 100918 472434
rect 101154 472198 101196 472434
rect 100876 465434 101196 472198
rect 100876 465198 100918 465434
rect 101154 465198 101196 465434
rect 100876 458434 101196 465198
rect 100876 458198 100918 458434
rect 101154 458198 101196 458434
rect 100876 451434 101196 458198
rect 100876 451198 100918 451434
rect 101154 451198 101196 451434
rect 100876 444434 101196 451198
rect 100876 444198 100918 444434
rect 101154 444198 101196 444434
rect 100876 437434 101196 444198
rect 100876 437198 100918 437434
rect 101154 437198 101196 437434
rect 100876 430434 101196 437198
rect 100876 430198 100918 430434
rect 101154 430198 101196 430434
rect 100876 423434 101196 430198
rect 100876 423198 100918 423434
rect 101154 423198 101196 423434
rect 100876 416434 101196 423198
rect 100876 416198 100918 416434
rect 101154 416198 101196 416434
rect 100876 409434 101196 416198
rect 100876 409198 100918 409434
rect 101154 409198 101196 409434
rect 100876 402434 101196 409198
rect 100876 402198 100918 402434
rect 101154 402198 101196 402434
rect 100876 395434 101196 402198
rect 100876 395198 100918 395434
rect 101154 395198 101196 395434
rect 100876 388434 101196 395198
rect 100876 388198 100918 388434
rect 101154 388198 101196 388434
rect 100876 381434 101196 388198
rect 100876 381198 100918 381434
rect 101154 381198 101196 381434
rect 100876 374434 101196 381198
rect 100876 374198 100918 374434
rect 101154 374198 101196 374434
rect 100876 367434 101196 374198
rect 100876 367198 100918 367434
rect 101154 367198 101196 367434
rect 100876 360434 101196 367198
rect 100876 360198 100918 360434
rect 101154 360198 101196 360434
rect 100876 353434 101196 360198
rect 100876 353198 100918 353434
rect 101154 353198 101196 353434
rect 100876 346434 101196 353198
rect 100876 346198 100918 346434
rect 101154 346198 101196 346434
rect 100876 339434 101196 346198
rect 100876 339198 100918 339434
rect 101154 339198 101196 339434
rect 100876 332434 101196 339198
rect 100876 332198 100918 332434
rect 101154 332198 101196 332434
rect 100876 325434 101196 332198
rect 100876 325198 100918 325434
rect 101154 325198 101196 325434
rect 100876 318434 101196 325198
rect 100876 318198 100918 318434
rect 101154 318198 101196 318434
rect 100876 311434 101196 318198
rect 100876 311198 100918 311434
rect 101154 311198 101196 311434
rect 100876 304434 101196 311198
rect 100876 304198 100918 304434
rect 101154 304198 101196 304434
rect 100876 297434 101196 304198
rect 100876 297198 100918 297434
rect 101154 297198 101196 297434
rect 100876 290434 101196 297198
rect 100876 290198 100918 290434
rect 101154 290198 101196 290434
rect 100876 283434 101196 290198
rect 100876 283198 100918 283434
rect 101154 283198 101196 283434
rect 100876 276434 101196 283198
rect 100876 276198 100918 276434
rect 101154 276198 101196 276434
rect 100876 269434 101196 276198
rect 100876 269198 100918 269434
rect 101154 269198 101196 269434
rect 100876 262434 101196 269198
rect 100876 262198 100918 262434
rect 101154 262198 101196 262434
rect 100876 255434 101196 262198
rect 100876 255198 100918 255434
rect 101154 255198 101196 255434
rect 100876 248434 101196 255198
rect 100876 248198 100918 248434
rect 101154 248198 101196 248434
rect 100876 241434 101196 248198
rect 100876 241198 100918 241434
rect 101154 241198 101196 241434
rect 100876 234434 101196 241198
rect 100876 234198 100918 234434
rect 101154 234198 101196 234434
rect 100876 227434 101196 234198
rect 100876 227198 100918 227434
rect 101154 227198 101196 227434
rect 100876 220434 101196 227198
rect 100876 220198 100918 220434
rect 101154 220198 101196 220434
rect 100876 213434 101196 220198
rect 100876 213198 100918 213434
rect 101154 213198 101196 213434
rect 100876 206434 101196 213198
rect 100876 206198 100918 206434
rect 101154 206198 101196 206434
rect 100876 199434 101196 206198
rect 100876 199198 100918 199434
rect 101154 199198 101196 199434
rect 100876 192434 101196 199198
rect 100876 192198 100918 192434
rect 101154 192198 101196 192434
rect 100876 185434 101196 192198
rect 100876 185198 100918 185434
rect 101154 185198 101196 185434
rect 100876 178434 101196 185198
rect 100876 178198 100918 178434
rect 101154 178198 101196 178434
rect 100876 171434 101196 178198
rect 100876 171198 100918 171434
rect 101154 171198 101196 171434
rect 100876 164434 101196 171198
rect 100876 164198 100918 164434
rect 101154 164198 101196 164434
rect 100876 157434 101196 164198
rect 100876 157198 100918 157434
rect 101154 157198 101196 157434
rect 100876 150434 101196 157198
rect 100876 150198 100918 150434
rect 101154 150198 101196 150434
rect 100876 143434 101196 150198
rect 100876 143198 100918 143434
rect 101154 143198 101196 143434
rect 100876 136434 101196 143198
rect 100876 136198 100918 136434
rect 101154 136198 101196 136434
rect 100876 129434 101196 136198
rect 100876 129198 100918 129434
rect 101154 129198 101196 129434
rect 100876 122434 101196 129198
rect 100876 122198 100918 122434
rect 101154 122198 101196 122434
rect 100876 115434 101196 122198
rect 100876 115198 100918 115434
rect 101154 115198 101196 115434
rect 100876 108434 101196 115198
rect 100876 108198 100918 108434
rect 101154 108198 101196 108434
rect 100876 101434 101196 108198
rect 100876 101198 100918 101434
rect 101154 101198 101196 101434
rect 100876 94434 101196 101198
rect 100876 94198 100918 94434
rect 101154 94198 101196 94434
rect 100876 87434 101196 94198
rect 100876 87198 100918 87434
rect 101154 87198 101196 87434
rect 100876 80434 101196 87198
rect 100876 80198 100918 80434
rect 101154 80198 101196 80434
rect 100876 73434 101196 80198
rect 100876 73198 100918 73434
rect 101154 73198 101196 73434
rect 100876 66434 101196 73198
rect 100876 66198 100918 66434
rect 101154 66198 101196 66434
rect 100876 59434 101196 66198
rect 100876 59198 100918 59434
rect 101154 59198 101196 59434
rect 100876 52434 101196 59198
rect 100876 52198 100918 52434
rect 101154 52198 101196 52434
rect 100876 45434 101196 52198
rect 100876 45198 100918 45434
rect 101154 45198 101196 45434
rect 100876 38434 101196 45198
rect 100876 38198 100918 38434
rect 101154 38198 101196 38434
rect 100876 31434 101196 38198
rect 100876 31198 100918 31434
rect 101154 31198 101196 31434
rect 100876 24434 101196 31198
rect 100876 24198 100918 24434
rect 101154 24198 101196 24434
rect 100876 17434 101196 24198
rect 100876 17198 100918 17434
rect 101154 17198 101196 17434
rect 100876 10434 101196 17198
rect 100876 10198 100918 10434
rect 101154 10198 101196 10434
rect 100876 3434 101196 10198
rect 100876 3198 100918 3434
rect 101154 3198 101196 3434
rect 100876 -1706 101196 3198
rect 100876 -1942 100918 -1706
rect 101154 -1942 101196 -1706
rect 100876 -2026 101196 -1942
rect 100876 -2262 100918 -2026
rect 101154 -2262 101196 -2026
rect 100876 -2294 101196 -2262
rect 106144 705238 106464 706230
rect 106144 705002 106186 705238
rect 106422 705002 106464 705238
rect 106144 704918 106464 705002
rect 106144 704682 106186 704918
rect 106422 704682 106464 704918
rect 106144 695494 106464 704682
rect 106144 695258 106186 695494
rect 106422 695258 106464 695494
rect 106144 688494 106464 695258
rect 106144 688258 106186 688494
rect 106422 688258 106464 688494
rect 106144 681494 106464 688258
rect 106144 681258 106186 681494
rect 106422 681258 106464 681494
rect 106144 674494 106464 681258
rect 106144 674258 106186 674494
rect 106422 674258 106464 674494
rect 106144 667494 106464 674258
rect 106144 667258 106186 667494
rect 106422 667258 106464 667494
rect 106144 660494 106464 667258
rect 106144 660258 106186 660494
rect 106422 660258 106464 660494
rect 106144 653494 106464 660258
rect 106144 653258 106186 653494
rect 106422 653258 106464 653494
rect 106144 646494 106464 653258
rect 106144 646258 106186 646494
rect 106422 646258 106464 646494
rect 106144 639494 106464 646258
rect 106144 639258 106186 639494
rect 106422 639258 106464 639494
rect 106144 632494 106464 639258
rect 106144 632258 106186 632494
rect 106422 632258 106464 632494
rect 106144 625494 106464 632258
rect 106144 625258 106186 625494
rect 106422 625258 106464 625494
rect 106144 618494 106464 625258
rect 106144 618258 106186 618494
rect 106422 618258 106464 618494
rect 106144 611494 106464 618258
rect 106144 611258 106186 611494
rect 106422 611258 106464 611494
rect 106144 604494 106464 611258
rect 106144 604258 106186 604494
rect 106422 604258 106464 604494
rect 106144 597494 106464 604258
rect 106144 597258 106186 597494
rect 106422 597258 106464 597494
rect 106144 590494 106464 597258
rect 106144 590258 106186 590494
rect 106422 590258 106464 590494
rect 106144 583494 106464 590258
rect 106144 583258 106186 583494
rect 106422 583258 106464 583494
rect 106144 576494 106464 583258
rect 106144 576258 106186 576494
rect 106422 576258 106464 576494
rect 106144 569494 106464 576258
rect 106144 569258 106186 569494
rect 106422 569258 106464 569494
rect 106144 562494 106464 569258
rect 106144 562258 106186 562494
rect 106422 562258 106464 562494
rect 106144 555494 106464 562258
rect 106144 555258 106186 555494
rect 106422 555258 106464 555494
rect 106144 548494 106464 555258
rect 106144 548258 106186 548494
rect 106422 548258 106464 548494
rect 106144 541494 106464 548258
rect 106144 541258 106186 541494
rect 106422 541258 106464 541494
rect 106144 534494 106464 541258
rect 106144 534258 106186 534494
rect 106422 534258 106464 534494
rect 106144 527494 106464 534258
rect 106144 527258 106186 527494
rect 106422 527258 106464 527494
rect 106144 520494 106464 527258
rect 106144 520258 106186 520494
rect 106422 520258 106464 520494
rect 106144 513494 106464 520258
rect 106144 513258 106186 513494
rect 106422 513258 106464 513494
rect 106144 506494 106464 513258
rect 106144 506258 106186 506494
rect 106422 506258 106464 506494
rect 106144 499494 106464 506258
rect 106144 499258 106186 499494
rect 106422 499258 106464 499494
rect 106144 492494 106464 499258
rect 106144 492258 106186 492494
rect 106422 492258 106464 492494
rect 106144 485494 106464 492258
rect 106144 485258 106186 485494
rect 106422 485258 106464 485494
rect 106144 478494 106464 485258
rect 106144 478258 106186 478494
rect 106422 478258 106464 478494
rect 106144 471494 106464 478258
rect 106144 471258 106186 471494
rect 106422 471258 106464 471494
rect 106144 464494 106464 471258
rect 106144 464258 106186 464494
rect 106422 464258 106464 464494
rect 106144 457494 106464 464258
rect 106144 457258 106186 457494
rect 106422 457258 106464 457494
rect 106144 450494 106464 457258
rect 106144 450258 106186 450494
rect 106422 450258 106464 450494
rect 106144 443494 106464 450258
rect 106144 443258 106186 443494
rect 106422 443258 106464 443494
rect 106144 436494 106464 443258
rect 106144 436258 106186 436494
rect 106422 436258 106464 436494
rect 106144 429494 106464 436258
rect 106144 429258 106186 429494
rect 106422 429258 106464 429494
rect 106144 422494 106464 429258
rect 106144 422258 106186 422494
rect 106422 422258 106464 422494
rect 106144 415494 106464 422258
rect 106144 415258 106186 415494
rect 106422 415258 106464 415494
rect 106144 408494 106464 415258
rect 106144 408258 106186 408494
rect 106422 408258 106464 408494
rect 106144 401494 106464 408258
rect 106144 401258 106186 401494
rect 106422 401258 106464 401494
rect 106144 394494 106464 401258
rect 106144 394258 106186 394494
rect 106422 394258 106464 394494
rect 106144 387494 106464 394258
rect 106144 387258 106186 387494
rect 106422 387258 106464 387494
rect 106144 380494 106464 387258
rect 106144 380258 106186 380494
rect 106422 380258 106464 380494
rect 106144 373494 106464 380258
rect 106144 373258 106186 373494
rect 106422 373258 106464 373494
rect 106144 366494 106464 373258
rect 106144 366258 106186 366494
rect 106422 366258 106464 366494
rect 106144 359494 106464 366258
rect 106144 359258 106186 359494
rect 106422 359258 106464 359494
rect 106144 352494 106464 359258
rect 106144 352258 106186 352494
rect 106422 352258 106464 352494
rect 106144 345494 106464 352258
rect 106144 345258 106186 345494
rect 106422 345258 106464 345494
rect 106144 338494 106464 345258
rect 106144 338258 106186 338494
rect 106422 338258 106464 338494
rect 106144 331494 106464 338258
rect 106144 331258 106186 331494
rect 106422 331258 106464 331494
rect 106144 324494 106464 331258
rect 106144 324258 106186 324494
rect 106422 324258 106464 324494
rect 106144 317494 106464 324258
rect 106144 317258 106186 317494
rect 106422 317258 106464 317494
rect 106144 310494 106464 317258
rect 106144 310258 106186 310494
rect 106422 310258 106464 310494
rect 106144 303494 106464 310258
rect 106144 303258 106186 303494
rect 106422 303258 106464 303494
rect 106144 296494 106464 303258
rect 106144 296258 106186 296494
rect 106422 296258 106464 296494
rect 106144 289494 106464 296258
rect 106144 289258 106186 289494
rect 106422 289258 106464 289494
rect 106144 282494 106464 289258
rect 106144 282258 106186 282494
rect 106422 282258 106464 282494
rect 106144 275494 106464 282258
rect 106144 275258 106186 275494
rect 106422 275258 106464 275494
rect 106144 268494 106464 275258
rect 106144 268258 106186 268494
rect 106422 268258 106464 268494
rect 106144 261494 106464 268258
rect 106144 261258 106186 261494
rect 106422 261258 106464 261494
rect 106144 254494 106464 261258
rect 106144 254258 106186 254494
rect 106422 254258 106464 254494
rect 106144 247494 106464 254258
rect 106144 247258 106186 247494
rect 106422 247258 106464 247494
rect 106144 240494 106464 247258
rect 106144 240258 106186 240494
rect 106422 240258 106464 240494
rect 106144 233494 106464 240258
rect 106144 233258 106186 233494
rect 106422 233258 106464 233494
rect 106144 226494 106464 233258
rect 106144 226258 106186 226494
rect 106422 226258 106464 226494
rect 106144 219494 106464 226258
rect 106144 219258 106186 219494
rect 106422 219258 106464 219494
rect 106144 212494 106464 219258
rect 106144 212258 106186 212494
rect 106422 212258 106464 212494
rect 106144 205494 106464 212258
rect 106144 205258 106186 205494
rect 106422 205258 106464 205494
rect 106144 198494 106464 205258
rect 106144 198258 106186 198494
rect 106422 198258 106464 198494
rect 106144 191494 106464 198258
rect 106144 191258 106186 191494
rect 106422 191258 106464 191494
rect 106144 184494 106464 191258
rect 106144 184258 106186 184494
rect 106422 184258 106464 184494
rect 106144 177494 106464 184258
rect 106144 177258 106186 177494
rect 106422 177258 106464 177494
rect 106144 170494 106464 177258
rect 106144 170258 106186 170494
rect 106422 170258 106464 170494
rect 106144 163494 106464 170258
rect 106144 163258 106186 163494
rect 106422 163258 106464 163494
rect 106144 156494 106464 163258
rect 106144 156258 106186 156494
rect 106422 156258 106464 156494
rect 106144 149494 106464 156258
rect 106144 149258 106186 149494
rect 106422 149258 106464 149494
rect 106144 142494 106464 149258
rect 106144 142258 106186 142494
rect 106422 142258 106464 142494
rect 106144 135494 106464 142258
rect 106144 135258 106186 135494
rect 106422 135258 106464 135494
rect 106144 128494 106464 135258
rect 106144 128258 106186 128494
rect 106422 128258 106464 128494
rect 106144 121494 106464 128258
rect 106144 121258 106186 121494
rect 106422 121258 106464 121494
rect 106144 114494 106464 121258
rect 106144 114258 106186 114494
rect 106422 114258 106464 114494
rect 106144 107494 106464 114258
rect 106144 107258 106186 107494
rect 106422 107258 106464 107494
rect 106144 100494 106464 107258
rect 106144 100258 106186 100494
rect 106422 100258 106464 100494
rect 106144 93494 106464 100258
rect 106144 93258 106186 93494
rect 106422 93258 106464 93494
rect 106144 86494 106464 93258
rect 106144 86258 106186 86494
rect 106422 86258 106464 86494
rect 106144 79494 106464 86258
rect 106144 79258 106186 79494
rect 106422 79258 106464 79494
rect 106144 72494 106464 79258
rect 106144 72258 106186 72494
rect 106422 72258 106464 72494
rect 106144 65494 106464 72258
rect 106144 65258 106186 65494
rect 106422 65258 106464 65494
rect 106144 58494 106464 65258
rect 106144 58258 106186 58494
rect 106422 58258 106464 58494
rect 106144 51494 106464 58258
rect 106144 51258 106186 51494
rect 106422 51258 106464 51494
rect 106144 44494 106464 51258
rect 106144 44258 106186 44494
rect 106422 44258 106464 44494
rect 106144 37494 106464 44258
rect 106144 37258 106186 37494
rect 106422 37258 106464 37494
rect 106144 30494 106464 37258
rect 106144 30258 106186 30494
rect 106422 30258 106464 30494
rect 106144 23494 106464 30258
rect 106144 23258 106186 23494
rect 106422 23258 106464 23494
rect 106144 16494 106464 23258
rect 106144 16258 106186 16494
rect 106422 16258 106464 16494
rect 106144 9494 106464 16258
rect 106144 9258 106186 9494
rect 106422 9258 106464 9494
rect 106144 2494 106464 9258
rect 106144 2258 106186 2494
rect 106422 2258 106464 2494
rect 106144 -746 106464 2258
rect 106144 -982 106186 -746
rect 106422 -982 106464 -746
rect 106144 -1066 106464 -982
rect 106144 -1302 106186 -1066
rect 106422 -1302 106464 -1066
rect 106144 -2294 106464 -1302
rect 107876 706198 108196 706230
rect 107876 705962 107918 706198
rect 108154 705962 108196 706198
rect 107876 705878 108196 705962
rect 107876 705642 107918 705878
rect 108154 705642 108196 705878
rect 107876 696434 108196 705642
rect 107876 696198 107918 696434
rect 108154 696198 108196 696434
rect 107876 689434 108196 696198
rect 107876 689198 107918 689434
rect 108154 689198 108196 689434
rect 107876 682434 108196 689198
rect 107876 682198 107918 682434
rect 108154 682198 108196 682434
rect 107876 675434 108196 682198
rect 107876 675198 107918 675434
rect 108154 675198 108196 675434
rect 107876 668434 108196 675198
rect 107876 668198 107918 668434
rect 108154 668198 108196 668434
rect 107876 661434 108196 668198
rect 107876 661198 107918 661434
rect 108154 661198 108196 661434
rect 107876 654434 108196 661198
rect 107876 654198 107918 654434
rect 108154 654198 108196 654434
rect 107876 647434 108196 654198
rect 107876 647198 107918 647434
rect 108154 647198 108196 647434
rect 107876 640434 108196 647198
rect 107876 640198 107918 640434
rect 108154 640198 108196 640434
rect 107876 633434 108196 640198
rect 107876 633198 107918 633434
rect 108154 633198 108196 633434
rect 107876 626434 108196 633198
rect 107876 626198 107918 626434
rect 108154 626198 108196 626434
rect 107876 619434 108196 626198
rect 107876 619198 107918 619434
rect 108154 619198 108196 619434
rect 107876 612434 108196 619198
rect 107876 612198 107918 612434
rect 108154 612198 108196 612434
rect 107876 605434 108196 612198
rect 107876 605198 107918 605434
rect 108154 605198 108196 605434
rect 107876 598434 108196 605198
rect 107876 598198 107918 598434
rect 108154 598198 108196 598434
rect 107876 591434 108196 598198
rect 107876 591198 107918 591434
rect 108154 591198 108196 591434
rect 107876 584434 108196 591198
rect 107876 584198 107918 584434
rect 108154 584198 108196 584434
rect 107876 577434 108196 584198
rect 107876 577198 107918 577434
rect 108154 577198 108196 577434
rect 107876 570434 108196 577198
rect 107876 570198 107918 570434
rect 108154 570198 108196 570434
rect 107876 563434 108196 570198
rect 107876 563198 107918 563434
rect 108154 563198 108196 563434
rect 107876 556434 108196 563198
rect 107876 556198 107918 556434
rect 108154 556198 108196 556434
rect 107876 549434 108196 556198
rect 107876 549198 107918 549434
rect 108154 549198 108196 549434
rect 107876 542434 108196 549198
rect 107876 542198 107918 542434
rect 108154 542198 108196 542434
rect 107876 535434 108196 542198
rect 107876 535198 107918 535434
rect 108154 535198 108196 535434
rect 107876 528434 108196 535198
rect 107876 528198 107918 528434
rect 108154 528198 108196 528434
rect 107876 521434 108196 528198
rect 107876 521198 107918 521434
rect 108154 521198 108196 521434
rect 107876 514434 108196 521198
rect 107876 514198 107918 514434
rect 108154 514198 108196 514434
rect 107876 507434 108196 514198
rect 107876 507198 107918 507434
rect 108154 507198 108196 507434
rect 107876 500434 108196 507198
rect 107876 500198 107918 500434
rect 108154 500198 108196 500434
rect 107876 493434 108196 500198
rect 107876 493198 107918 493434
rect 108154 493198 108196 493434
rect 107876 486434 108196 493198
rect 107876 486198 107918 486434
rect 108154 486198 108196 486434
rect 107876 479434 108196 486198
rect 107876 479198 107918 479434
rect 108154 479198 108196 479434
rect 107876 472434 108196 479198
rect 107876 472198 107918 472434
rect 108154 472198 108196 472434
rect 107876 465434 108196 472198
rect 107876 465198 107918 465434
rect 108154 465198 108196 465434
rect 107876 458434 108196 465198
rect 107876 458198 107918 458434
rect 108154 458198 108196 458434
rect 107876 451434 108196 458198
rect 107876 451198 107918 451434
rect 108154 451198 108196 451434
rect 107876 444434 108196 451198
rect 107876 444198 107918 444434
rect 108154 444198 108196 444434
rect 107876 437434 108196 444198
rect 107876 437198 107918 437434
rect 108154 437198 108196 437434
rect 107876 430434 108196 437198
rect 107876 430198 107918 430434
rect 108154 430198 108196 430434
rect 107876 423434 108196 430198
rect 107876 423198 107918 423434
rect 108154 423198 108196 423434
rect 107876 416434 108196 423198
rect 107876 416198 107918 416434
rect 108154 416198 108196 416434
rect 107876 409434 108196 416198
rect 107876 409198 107918 409434
rect 108154 409198 108196 409434
rect 107876 402434 108196 409198
rect 107876 402198 107918 402434
rect 108154 402198 108196 402434
rect 107876 395434 108196 402198
rect 107876 395198 107918 395434
rect 108154 395198 108196 395434
rect 107876 388434 108196 395198
rect 107876 388198 107918 388434
rect 108154 388198 108196 388434
rect 107876 381434 108196 388198
rect 107876 381198 107918 381434
rect 108154 381198 108196 381434
rect 107876 374434 108196 381198
rect 107876 374198 107918 374434
rect 108154 374198 108196 374434
rect 107876 367434 108196 374198
rect 107876 367198 107918 367434
rect 108154 367198 108196 367434
rect 107876 360434 108196 367198
rect 107876 360198 107918 360434
rect 108154 360198 108196 360434
rect 107876 353434 108196 360198
rect 107876 353198 107918 353434
rect 108154 353198 108196 353434
rect 107876 346434 108196 353198
rect 107876 346198 107918 346434
rect 108154 346198 108196 346434
rect 107876 339434 108196 346198
rect 107876 339198 107918 339434
rect 108154 339198 108196 339434
rect 107876 332434 108196 339198
rect 107876 332198 107918 332434
rect 108154 332198 108196 332434
rect 107876 325434 108196 332198
rect 107876 325198 107918 325434
rect 108154 325198 108196 325434
rect 107876 318434 108196 325198
rect 107876 318198 107918 318434
rect 108154 318198 108196 318434
rect 107876 311434 108196 318198
rect 107876 311198 107918 311434
rect 108154 311198 108196 311434
rect 107876 304434 108196 311198
rect 107876 304198 107918 304434
rect 108154 304198 108196 304434
rect 107876 297434 108196 304198
rect 107876 297198 107918 297434
rect 108154 297198 108196 297434
rect 107876 290434 108196 297198
rect 107876 290198 107918 290434
rect 108154 290198 108196 290434
rect 107876 283434 108196 290198
rect 107876 283198 107918 283434
rect 108154 283198 108196 283434
rect 107876 276434 108196 283198
rect 107876 276198 107918 276434
rect 108154 276198 108196 276434
rect 107876 269434 108196 276198
rect 107876 269198 107918 269434
rect 108154 269198 108196 269434
rect 107876 262434 108196 269198
rect 107876 262198 107918 262434
rect 108154 262198 108196 262434
rect 107876 255434 108196 262198
rect 107876 255198 107918 255434
rect 108154 255198 108196 255434
rect 107876 248434 108196 255198
rect 107876 248198 107918 248434
rect 108154 248198 108196 248434
rect 107876 241434 108196 248198
rect 107876 241198 107918 241434
rect 108154 241198 108196 241434
rect 107876 234434 108196 241198
rect 107876 234198 107918 234434
rect 108154 234198 108196 234434
rect 107876 227434 108196 234198
rect 107876 227198 107918 227434
rect 108154 227198 108196 227434
rect 107876 220434 108196 227198
rect 107876 220198 107918 220434
rect 108154 220198 108196 220434
rect 107876 213434 108196 220198
rect 107876 213198 107918 213434
rect 108154 213198 108196 213434
rect 107876 206434 108196 213198
rect 107876 206198 107918 206434
rect 108154 206198 108196 206434
rect 107876 199434 108196 206198
rect 107876 199198 107918 199434
rect 108154 199198 108196 199434
rect 107876 192434 108196 199198
rect 107876 192198 107918 192434
rect 108154 192198 108196 192434
rect 107876 185434 108196 192198
rect 107876 185198 107918 185434
rect 108154 185198 108196 185434
rect 107876 178434 108196 185198
rect 107876 178198 107918 178434
rect 108154 178198 108196 178434
rect 107876 171434 108196 178198
rect 107876 171198 107918 171434
rect 108154 171198 108196 171434
rect 107876 164434 108196 171198
rect 107876 164198 107918 164434
rect 108154 164198 108196 164434
rect 107876 157434 108196 164198
rect 107876 157198 107918 157434
rect 108154 157198 108196 157434
rect 107876 150434 108196 157198
rect 107876 150198 107918 150434
rect 108154 150198 108196 150434
rect 107876 143434 108196 150198
rect 107876 143198 107918 143434
rect 108154 143198 108196 143434
rect 107876 136434 108196 143198
rect 107876 136198 107918 136434
rect 108154 136198 108196 136434
rect 107876 129434 108196 136198
rect 107876 129198 107918 129434
rect 108154 129198 108196 129434
rect 107876 122434 108196 129198
rect 107876 122198 107918 122434
rect 108154 122198 108196 122434
rect 107876 115434 108196 122198
rect 107876 115198 107918 115434
rect 108154 115198 108196 115434
rect 107876 108434 108196 115198
rect 107876 108198 107918 108434
rect 108154 108198 108196 108434
rect 107876 101434 108196 108198
rect 107876 101198 107918 101434
rect 108154 101198 108196 101434
rect 107876 94434 108196 101198
rect 107876 94198 107918 94434
rect 108154 94198 108196 94434
rect 107876 87434 108196 94198
rect 107876 87198 107918 87434
rect 108154 87198 108196 87434
rect 107876 80434 108196 87198
rect 107876 80198 107918 80434
rect 108154 80198 108196 80434
rect 107876 73434 108196 80198
rect 107876 73198 107918 73434
rect 108154 73198 108196 73434
rect 107876 66434 108196 73198
rect 107876 66198 107918 66434
rect 108154 66198 108196 66434
rect 107876 59434 108196 66198
rect 107876 59198 107918 59434
rect 108154 59198 108196 59434
rect 107876 52434 108196 59198
rect 107876 52198 107918 52434
rect 108154 52198 108196 52434
rect 107876 45434 108196 52198
rect 107876 45198 107918 45434
rect 108154 45198 108196 45434
rect 107876 38434 108196 45198
rect 107876 38198 107918 38434
rect 108154 38198 108196 38434
rect 107876 31434 108196 38198
rect 107876 31198 107918 31434
rect 108154 31198 108196 31434
rect 107876 24434 108196 31198
rect 107876 24198 107918 24434
rect 108154 24198 108196 24434
rect 107876 17434 108196 24198
rect 107876 17198 107918 17434
rect 108154 17198 108196 17434
rect 107876 10434 108196 17198
rect 107876 10198 107918 10434
rect 108154 10198 108196 10434
rect 107876 3434 108196 10198
rect 107876 3198 107918 3434
rect 108154 3198 108196 3434
rect 107876 -1706 108196 3198
rect 107876 -1942 107918 -1706
rect 108154 -1942 108196 -1706
rect 107876 -2026 108196 -1942
rect 107876 -2262 107918 -2026
rect 108154 -2262 108196 -2026
rect 107876 -2294 108196 -2262
rect 113144 705238 113464 706230
rect 113144 705002 113186 705238
rect 113422 705002 113464 705238
rect 113144 704918 113464 705002
rect 113144 704682 113186 704918
rect 113422 704682 113464 704918
rect 113144 695494 113464 704682
rect 113144 695258 113186 695494
rect 113422 695258 113464 695494
rect 113144 688494 113464 695258
rect 113144 688258 113186 688494
rect 113422 688258 113464 688494
rect 113144 681494 113464 688258
rect 113144 681258 113186 681494
rect 113422 681258 113464 681494
rect 113144 674494 113464 681258
rect 113144 674258 113186 674494
rect 113422 674258 113464 674494
rect 113144 667494 113464 674258
rect 113144 667258 113186 667494
rect 113422 667258 113464 667494
rect 113144 660494 113464 667258
rect 113144 660258 113186 660494
rect 113422 660258 113464 660494
rect 113144 653494 113464 660258
rect 113144 653258 113186 653494
rect 113422 653258 113464 653494
rect 113144 646494 113464 653258
rect 113144 646258 113186 646494
rect 113422 646258 113464 646494
rect 113144 639494 113464 646258
rect 113144 639258 113186 639494
rect 113422 639258 113464 639494
rect 113144 632494 113464 639258
rect 113144 632258 113186 632494
rect 113422 632258 113464 632494
rect 113144 625494 113464 632258
rect 113144 625258 113186 625494
rect 113422 625258 113464 625494
rect 113144 618494 113464 625258
rect 113144 618258 113186 618494
rect 113422 618258 113464 618494
rect 113144 611494 113464 618258
rect 113144 611258 113186 611494
rect 113422 611258 113464 611494
rect 113144 604494 113464 611258
rect 113144 604258 113186 604494
rect 113422 604258 113464 604494
rect 113144 597494 113464 604258
rect 113144 597258 113186 597494
rect 113422 597258 113464 597494
rect 113144 590494 113464 597258
rect 113144 590258 113186 590494
rect 113422 590258 113464 590494
rect 113144 583494 113464 590258
rect 113144 583258 113186 583494
rect 113422 583258 113464 583494
rect 113144 576494 113464 583258
rect 113144 576258 113186 576494
rect 113422 576258 113464 576494
rect 113144 569494 113464 576258
rect 113144 569258 113186 569494
rect 113422 569258 113464 569494
rect 113144 562494 113464 569258
rect 113144 562258 113186 562494
rect 113422 562258 113464 562494
rect 113144 555494 113464 562258
rect 113144 555258 113186 555494
rect 113422 555258 113464 555494
rect 113144 548494 113464 555258
rect 113144 548258 113186 548494
rect 113422 548258 113464 548494
rect 113144 541494 113464 548258
rect 113144 541258 113186 541494
rect 113422 541258 113464 541494
rect 113144 534494 113464 541258
rect 113144 534258 113186 534494
rect 113422 534258 113464 534494
rect 113144 527494 113464 534258
rect 113144 527258 113186 527494
rect 113422 527258 113464 527494
rect 113144 520494 113464 527258
rect 113144 520258 113186 520494
rect 113422 520258 113464 520494
rect 113144 513494 113464 520258
rect 113144 513258 113186 513494
rect 113422 513258 113464 513494
rect 113144 506494 113464 513258
rect 113144 506258 113186 506494
rect 113422 506258 113464 506494
rect 113144 499494 113464 506258
rect 113144 499258 113186 499494
rect 113422 499258 113464 499494
rect 113144 492494 113464 499258
rect 113144 492258 113186 492494
rect 113422 492258 113464 492494
rect 113144 485494 113464 492258
rect 113144 485258 113186 485494
rect 113422 485258 113464 485494
rect 113144 478494 113464 485258
rect 113144 478258 113186 478494
rect 113422 478258 113464 478494
rect 113144 471494 113464 478258
rect 113144 471258 113186 471494
rect 113422 471258 113464 471494
rect 113144 464494 113464 471258
rect 113144 464258 113186 464494
rect 113422 464258 113464 464494
rect 113144 457494 113464 464258
rect 113144 457258 113186 457494
rect 113422 457258 113464 457494
rect 113144 450494 113464 457258
rect 113144 450258 113186 450494
rect 113422 450258 113464 450494
rect 113144 443494 113464 450258
rect 113144 443258 113186 443494
rect 113422 443258 113464 443494
rect 113144 436494 113464 443258
rect 113144 436258 113186 436494
rect 113422 436258 113464 436494
rect 113144 429494 113464 436258
rect 113144 429258 113186 429494
rect 113422 429258 113464 429494
rect 113144 422494 113464 429258
rect 113144 422258 113186 422494
rect 113422 422258 113464 422494
rect 113144 415494 113464 422258
rect 113144 415258 113186 415494
rect 113422 415258 113464 415494
rect 113144 408494 113464 415258
rect 113144 408258 113186 408494
rect 113422 408258 113464 408494
rect 113144 401494 113464 408258
rect 113144 401258 113186 401494
rect 113422 401258 113464 401494
rect 113144 394494 113464 401258
rect 113144 394258 113186 394494
rect 113422 394258 113464 394494
rect 113144 387494 113464 394258
rect 113144 387258 113186 387494
rect 113422 387258 113464 387494
rect 113144 380494 113464 387258
rect 113144 380258 113186 380494
rect 113422 380258 113464 380494
rect 113144 373494 113464 380258
rect 113144 373258 113186 373494
rect 113422 373258 113464 373494
rect 113144 366494 113464 373258
rect 113144 366258 113186 366494
rect 113422 366258 113464 366494
rect 113144 359494 113464 366258
rect 113144 359258 113186 359494
rect 113422 359258 113464 359494
rect 113144 352494 113464 359258
rect 113144 352258 113186 352494
rect 113422 352258 113464 352494
rect 113144 345494 113464 352258
rect 113144 345258 113186 345494
rect 113422 345258 113464 345494
rect 113144 338494 113464 345258
rect 113144 338258 113186 338494
rect 113422 338258 113464 338494
rect 113144 331494 113464 338258
rect 113144 331258 113186 331494
rect 113422 331258 113464 331494
rect 113144 324494 113464 331258
rect 113144 324258 113186 324494
rect 113422 324258 113464 324494
rect 113144 317494 113464 324258
rect 113144 317258 113186 317494
rect 113422 317258 113464 317494
rect 113144 310494 113464 317258
rect 113144 310258 113186 310494
rect 113422 310258 113464 310494
rect 113144 303494 113464 310258
rect 113144 303258 113186 303494
rect 113422 303258 113464 303494
rect 113144 296494 113464 303258
rect 113144 296258 113186 296494
rect 113422 296258 113464 296494
rect 113144 289494 113464 296258
rect 113144 289258 113186 289494
rect 113422 289258 113464 289494
rect 113144 282494 113464 289258
rect 113144 282258 113186 282494
rect 113422 282258 113464 282494
rect 113144 275494 113464 282258
rect 113144 275258 113186 275494
rect 113422 275258 113464 275494
rect 113144 268494 113464 275258
rect 113144 268258 113186 268494
rect 113422 268258 113464 268494
rect 113144 261494 113464 268258
rect 113144 261258 113186 261494
rect 113422 261258 113464 261494
rect 113144 254494 113464 261258
rect 113144 254258 113186 254494
rect 113422 254258 113464 254494
rect 113144 247494 113464 254258
rect 113144 247258 113186 247494
rect 113422 247258 113464 247494
rect 113144 240494 113464 247258
rect 113144 240258 113186 240494
rect 113422 240258 113464 240494
rect 113144 233494 113464 240258
rect 113144 233258 113186 233494
rect 113422 233258 113464 233494
rect 113144 226494 113464 233258
rect 113144 226258 113186 226494
rect 113422 226258 113464 226494
rect 113144 219494 113464 226258
rect 113144 219258 113186 219494
rect 113422 219258 113464 219494
rect 113144 212494 113464 219258
rect 113144 212258 113186 212494
rect 113422 212258 113464 212494
rect 113144 205494 113464 212258
rect 113144 205258 113186 205494
rect 113422 205258 113464 205494
rect 113144 198494 113464 205258
rect 113144 198258 113186 198494
rect 113422 198258 113464 198494
rect 113144 191494 113464 198258
rect 113144 191258 113186 191494
rect 113422 191258 113464 191494
rect 113144 184494 113464 191258
rect 113144 184258 113186 184494
rect 113422 184258 113464 184494
rect 113144 177494 113464 184258
rect 113144 177258 113186 177494
rect 113422 177258 113464 177494
rect 113144 170494 113464 177258
rect 113144 170258 113186 170494
rect 113422 170258 113464 170494
rect 113144 163494 113464 170258
rect 113144 163258 113186 163494
rect 113422 163258 113464 163494
rect 113144 156494 113464 163258
rect 113144 156258 113186 156494
rect 113422 156258 113464 156494
rect 113144 149494 113464 156258
rect 113144 149258 113186 149494
rect 113422 149258 113464 149494
rect 113144 142494 113464 149258
rect 113144 142258 113186 142494
rect 113422 142258 113464 142494
rect 113144 135494 113464 142258
rect 113144 135258 113186 135494
rect 113422 135258 113464 135494
rect 113144 128494 113464 135258
rect 113144 128258 113186 128494
rect 113422 128258 113464 128494
rect 113144 121494 113464 128258
rect 113144 121258 113186 121494
rect 113422 121258 113464 121494
rect 113144 114494 113464 121258
rect 113144 114258 113186 114494
rect 113422 114258 113464 114494
rect 113144 107494 113464 114258
rect 113144 107258 113186 107494
rect 113422 107258 113464 107494
rect 113144 100494 113464 107258
rect 113144 100258 113186 100494
rect 113422 100258 113464 100494
rect 113144 93494 113464 100258
rect 113144 93258 113186 93494
rect 113422 93258 113464 93494
rect 113144 86494 113464 93258
rect 113144 86258 113186 86494
rect 113422 86258 113464 86494
rect 113144 79494 113464 86258
rect 113144 79258 113186 79494
rect 113422 79258 113464 79494
rect 113144 72494 113464 79258
rect 113144 72258 113186 72494
rect 113422 72258 113464 72494
rect 113144 65494 113464 72258
rect 113144 65258 113186 65494
rect 113422 65258 113464 65494
rect 113144 58494 113464 65258
rect 113144 58258 113186 58494
rect 113422 58258 113464 58494
rect 113144 51494 113464 58258
rect 113144 51258 113186 51494
rect 113422 51258 113464 51494
rect 113144 44494 113464 51258
rect 113144 44258 113186 44494
rect 113422 44258 113464 44494
rect 113144 37494 113464 44258
rect 113144 37258 113186 37494
rect 113422 37258 113464 37494
rect 113144 30494 113464 37258
rect 113144 30258 113186 30494
rect 113422 30258 113464 30494
rect 113144 23494 113464 30258
rect 113144 23258 113186 23494
rect 113422 23258 113464 23494
rect 113144 16494 113464 23258
rect 113144 16258 113186 16494
rect 113422 16258 113464 16494
rect 113144 9494 113464 16258
rect 113144 9258 113186 9494
rect 113422 9258 113464 9494
rect 113144 2494 113464 9258
rect 113144 2258 113186 2494
rect 113422 2258 113464 2494
rect 113144 -746 113464 2258
rect 113144 -982 113186 -746
rect 113422 -982 113464 -746
rect 113144 -1066 113464 -982
rect 113144 -1302 113186 -1066
rect 113422 -1302 113464 -1066
rect 113144 -2294 113464 -1302
rect 114876 706198 115196 706230
rect 114876 705962 114918 706198
rect 115154 705962 115196 706198
rect 114876 705878 115196 705962
rect 114876 705642 114918 705878
rect 115154 705642 115196 705878
rect 114876 696434 115196 705642
rect 114876 696198 114918 696434
rect 115154 696198 115196 696434
rect 114876 689434 115196 696198
rect 114876 689198 114918 689434
rect 115154 689198 115196 689434
rect 114876 682434 115196 689198
rect 114876 682198 114918 682434
rect 115154 682198 115196 682434
rect 114876 675434 115196 682198
rect 114876 675198 114918 675434
rect 115154 675198 115196 675434
rect 114876 668434 115196 675198
rect 114876 668198 114918 668434
rect 115154 668198 115196 668434
rect 114876 661434 115196 668198
rect 114876 661198 114918 661434
rect 115154 661198 115196 661434
rect 114876 654434 115196 661198
rect 114876 654198 114918 654434
rect 115154 654198 115196 654434
rect 114876 647434 115196 654198
rect 114876 647198 114918 647434
rect 115154 647198 115196 647434
rect 114876 640434 115196 647198
rect 114876 640198 114918 640434
rect 115154 640198 115196 640434
rect 114876 633434 115196 640198
rect 114876 633198 114918 633434
rect 115154 633198 115196 633434
rect 114876 626434 115196 633198
rect 114876 626198 114918 626434
rect 115154 626198 115196 626434
rect 114876 619434 115196 626198
rect 114876 619198 114918 619434
rect 115154 619198 115196 619434
rect 114876 612434 115196 619198
rect 114876 612198 114918 612434
rect 115154 612198 115196 612434
rect 114876 605434 115196 612198
rect 114876 605198 114918 605434
rect 115154 605198 115196 605434
rect 114876 598434 115196 605198
rect 114876 598198 114918 598434
rect 115154 598198 115196 598434
rect 114876 591434 115196 598198
rect 114876 591198 114918 591434
rect 115154 591198 115196 591434
rect 114876 584434 115196 591198
rect 114876 584198 114918 584434
rect 115154 584198 115196 584434
rect 114876 577434 115196 584198
rect 114876 577198 114918 577434
rect 115154 577198 115196 577434
rect 114876 570434 115196 577198
rect 114876 570198 114918 570434
rect 115154 570198 115196 570434
rect 114876 563434 115196 570198
rect 114876 563198 114918 563434
rect 115154 563198 115196 563434
rect 114876 556434 115196 563198
rect 114876 556198 114918 556434
rect 115154 556198 115196 556434
rect 114876 549434 115196 556198
rect 114876 549198 114918 549434
rect 115154 549198 115196 549434
rect 114876 542434 115196 549198
rect 114876 542198 114918 542434
rect 115154 542198 115196 542434
rect 114876 535434 115196 542198
rect 114876 535198 114918 535434
rect 115154 535198 115196 535434
rect 114876 528434 115196 535198
rect 114876 528198 114918 528434
rect 115154 528198 115196 528434
rect 114876 521434 115196 528198
rect 114876 521198 114918 521434
rect 115154 521198 115196 521434
rect 114876 514434 115196 521198
rect 114876 514198 114918 514434
rect 115154 514198 115196 514434
rect 114876 507434 115196 514198
rect 114876 507198 114918 507434
rect 115154 507198 115196 507434
rect 114876 500434 115196 507198
rect 114876 500198 114918 500434
rect 115154 500198 115196 500434
rect 114876 493434 115196 500198
rect 114876 493198 114918 493434
rect 115154 493198 115196 493434
rect 114876 486434 115196 493198
rect 114876 486198 114918 486434
rect 115154 486198 115196 486434
rect 114876 479434 115196 486198
rect 114876 479198 114918 479434
rect 115154 479198 115196 479434
rect 114876 472434 115196 479198
rect 114876 472198 114918 472434
rect 115154 472198 115196 472434
rect 114876 465434 115196 472198
rect 114876 465198 114918 465434
rect 115154 465198 115196 465434
rect 114876 458434 115196 465198
rect 114876 458198 114918 458434
rect 115154 458198 115196 458434
rect 114876 451434 115196 458198
rect 114876 451198 114918 451434
rect 115154 451198 115196 451434
rect 114876 444434 115196 451198
rect 114876 444198 114918 444434
rect 115154 444198 115196 444434
rect 114876 437434 115196 444198
rect 114876 437198 114918 437434
rect 115154 437198 115196 437434
rect 114876 430434 115196 437198
rect 114876 430198 114918 430434
rect 115154 430198 115196 430434
rect 114876 423434 115196 430198
rect 114876 423198 114918 423434
rect 115154 423198 115196 423434
rect 114876 416434 115196 423198
rect 114876 416198 114918 416434
rect 115154 416198 115196 416434
rect 114876 409434 115196 416198
rect 114876 409198 114918 409434
rect 115154 409198 115196 409434
rect 114876 402434 115196 409198
rect 114876 402198 114918 402434
rect 115154 402198 115196 402434
rect 114876 395434 115196 402198
rect 114876 395198 114918 395434
rect 115154 395198 115196 395434
rect 114876 388434 115196 395198
rect 114876 388198 114918 388434
rect 115154 388198 115196 388434
rect 114876 381434 115196 388198
rect 114876 381198 114918 381434
rect 115154 381198 115196 381434
rect 114876 374434 115196 381198
rect 114876 374198 114918 374434
rect 115154 374198 115196 374434
rect 114876 367434 115196 374198
rect 114876 367198 114918 367434
rect 115154 367198 115196 367434
rect 114876 360434 115196 367198
rect 114876 360198 114918 360434
rect 115154 360198 115196 360434
rect 114876 353434 115196 360198
rect 114876 353198 114918 353434
rect 115154 353198 115196 353434
rect 114876 346434 115196 353198
rect 114876 346198 114918 346434
rect 115154 346198 115196 346434
rect 114876 339434 115196 346198
rect 114876 339198 114918 339434
rect 115154 339198 115196 339434
rect 114876 332434 115196 339198
rect 114876 332198 114918 332434
rect 115154 332198 115196 332434
rect 114876 325434 115196 332198
rect 114876 325198 114918 325434
rect 115154 325198 115196 325434
rect 114876 318434 115196 325198
rect 114876 318198 114918 318434
rect 115154 318198 115196 318434
rect 114876 311434 115196 318198
rect 114876 311198 114918 311434
rect 115154 311198 115196 311434
rect 114876 304434 115196 311198
rect 114876 304198 114918 304434
rect 115154 304198 115196 304434
rect 114876 297434 115196 304198
rect 114876 297198 114918 297434
rect 115154 297198 115196 297434
rect 114876 290434 115196 297198
rect 114876 290198 114918 290434
rect 115154 290198 115196 290434
rect 114876 283434 115196 290198
rect 114876 283198 114918 283434
rect 115154 283198 115196 283434
rect 114876 276434 115196 283198
rect 114876 276198 114918 276434
rect 115154 276198 115196 276434
rect 114876 269434 115196 276198
rect 114876 269198 114918 269434
rect 115154 269198 115196 269434
rect 114876 262434 115196 269198
rect 114876 262198 114918 262434
rect 115154 262198 115196 262434
rect 114876 255434 115196 262198
rect 114876 255198 114918 255434
rect 115154 255198 115196 255434
rect 114876 248434 115196 255198
rect 114876 248198 114918 248434
rect 115154 248198 115196 248434
rect 114876 241434 115196 248198
rect 114876 241198 114918 241434
rect 115154 241198 115196 241434
rect 114876 234434 115196 241198
rect 114876 234198 114918 234434
rect 115154 234198 115196 234434
rect 114876 227434 115196 234198
rect 114876 227198 114918 227434
rect 115154 227198 115196 227434
rect 114876 220434 115196 227198
rect 114876 220198 114918 220434
rect 115154 220198 115196 220434
rect 114876 213434 115196 220198
rect 114876 213198 114918 213434
rect 115154 213198 115196 213434
rect 114876 206434 115196 213198
rect 114876 206198 114918 206434
rect 115154 206198 115196 206434
rect 114876 199434 115196 206198
rect 114876 199198 114918 199434
rect 115154 199198 115196 199434
rect 114876 192434 115196 199198
rect 114876 192198 114918 192434
rect 115154 192198 115196 192434
rect 114876 185434 115196 192198
rect 114876 185198 114918 185434
rect 115154 185198 115196 185434
rect 114876 178434 115196 185198
rect 114876 178198 114918 178434
rect 115154 178198 115196 178434
rect 114876 171434 115196 178198
rect 114876 171198 114918 171434
rect 115154 171198 115196 171434
rect 114876 164434 115196 171198
rect 114876 164198 114918 164434
rect 115154 164198 115196 164434
rect 114876 157434 115196 164198
rect 114876 157198 114918 157434
rect 115154 157198 115196 157434
rect 114876 150434 115196 157198
rect 114876 150198 114918 150434
rect 115154 150198 115196 150434
rect 114876 143434 115196 150198
rect 114876 143198 114918 143434
rect 115154 143198 115196 143434
rect 114876 136434 115196 143198
rect 114876 136198 114918 136434
rect 115154 136198 115196 136434
rect 114876 129434 115196 136198
rect 114876 129198 114918 129434
rect 115154 129198 115196 129434
rect 114876 122434 115196 129198
rect 114876 122198 114918 122434
rect 115154 122198 115196 122434
rect 114876 115434 115196 122198
rect 114876 115198 114918 115434
rect 115154 115198 115196 115434
rect 114876 108434 115196 115198
rect 114876 108198 114918 108434
rect 115154 108198 115196 108434
rect 114876 101434 115196 108198
rect 114876 101198 114918 101434
rect 115154 101198 115196 101434
rect 114876 94434 115196 101198
rect 114876 94198 114918 94434
rect 115154 94198 115196 94434
rect 114876 87434 115196 94198
rect 114876 87198 114918 87434
rect 115154 87198 115196 87434
rect 114876 80434 115196 87198
rect 114876 80198 114918 80434
rect 115154 80198 115196 80434
rect 114876 73434 115196 80198
rect 114876 73198 114918 73434
rect 115154 73198 115196 73434
rect 114876 66434 115196 73198
rect 114876 66198 114918 66434
rect 115154 66198 115196 66434
rect 114876 59434 115196 66198
rect 114876 59198 114918 59434
rect 115154 59198 115196 59434
rect 114876 52434 115196 59198
rect 114876 52198 114918 52434
rect 115154 52198 115196 52434
rect 114876 45434 115196 52198
rect 114876 45198 114918 45434
rect 115154 45198 115196 45434
rect 114876 38434 115196 45198
rect 114876 38198 114918 38434
rect 115154 38198 115196 38434
rect 114876 31434 115196 38198
rect 114876 31198 114918 31434
rect 115154 31198 115196 31434
rect 114876 24434 115196 31198
rect 114876 24198 114918 24434
rect 115154 24198 115196 24434
rect 114876 17434 115196 24198
rect 114876 17198 114918 17434
rect 115154 17198 115196 17434
rect 114876 10434 115196 17198
rect 114876 10198 114918 10434
rect 115154 10198 115196 10434
rect 114876 3434 115196 10198
rect 114876 3198 114918 3434
rect 115154 3198 115196 3434
rect 114876 -1706 115196 3198
rect 114876 -1942 114918 -1706
rect 115154 -1942 115196 -1706
rect 114876 -2026 115196 -1942
rect 114876 -2262 114918 -2026
rect 115154 -2262 115196 -2026
rect 114876 -2294 115196 -2262
rect 120144 705238 120464 706230
rect 120144 705002 120186 705238
rect 120422 705002 120464 705238
rect 120144 704918 120464 705002
rect 120144 704682 120186 704918
rect 120422 704682 120464 704918
rect 120144 695494 120464 704682
rect 120144 695258 120186 695494
rect 120422 695258 120464 695494
rect 120144 688494 120464 695258
rect 120144 688258 120186 688494
rect 120422 688258 120464 688494
rect 120144 681494 120464 688258
rect 120144 681258 120186 681494
rect 120422 681258 120464 681494
rect 120144 674494 120464 681258
rect 120144 674258 120186 674494
rect 120422 674258 120464 674494
rect 120144 667494 120464 674258
rect 120144 667258 120186 667494
rect 120422 667258 120464 667494
rect 120144 660494 120464 667258
rect 120144 660258 120186 660494
rect 120422 660258 120464 660494
rect 120144 653494 120464 660258
rect 120144 653258 120186 653494
rect 120422 653258 120464 653494
rect 120144 646494 120464 653258
rect 120144 646258 120186 646494
rect 120422 646258 120464 646494
rect 120144 639494 120464 646258
rect 120144 639258 120186 639494
rect 120422 639258 120464 639494
rect 120144 632494 120464 639258
rect 120144 632258 120186 632494
rect 120422 632258 120464 632494
rect 120144 625494 120464 632258
rect 120144 625258 120186 625494
rect 120422 625258 120464 625494
rect 120144 618494 120464 625258
rect 120144 618258 120186 618494
rect 120422 618258 120464 618494
rect 120144 611494 120464 618258
rect 120144 611258 120186 611494
rect 120422 611258 120464 611494
rect 120144 604494 120464 611258
rect 120144 604258 120186 604494
rect 120422 604258 120464 604494
rect 120144 597494 120464 604258
rect 120144 597258 120186 597494
rect 120422 597258 120464 597494
rect 120144 590494 120464 597258
rect 120144 590258 120186 590494
rect 120422 590258 120464 590494
rect 120144 583494 120464 590258
rect 120144 583258 120186 583494
rect 120422 583258 120464 583494
rect 120144 576494 120464 583258
rect 120144 576258 120186 576494
rect 120422 576258 120464 576494
rect 120144 569494 120464 576258
rect 120144 569258 120186 569494
rect 120422 569258 120464 569494
rect 120144 562494 120464 569258
rect 120144 562258 120186 562494
rect 120422 562258 120464 562494
rect 120144 555494 120464 562258
rect 120144 555258 120186 555494
rect 120422 555258 120464 555494
rect 120144 548494 120464 555258
rect 120144 548258 120186 548494
rect 120422 548258 120464 548494
rect 120144 541494 120464 548258
rect 120144 541258 120186 541494
rect 120422 541258 120464 541494
rect 120144 534494 120464 541258
rect 120144 534258 120186 534494
rect 120422 534258 120464 534494
rect 120144 527494 120464 534258
rect 120144 527258 120186 527494
rect 120422 527258 120464 527494
rect 120144 520494 120464 527258
rect 120144 520258 120186 520494
rect 120422 520258 120464 520494
rect 120144 513494 120464 520258
rect 120144 513258 120186 513494
rect 120422 513258 120464 513494
rect 120144 506494 120464 513258
rect 120144 506258 120186 506494
rect 120422 506258 120464 506494
rect 120144 499494 120464 506258
rect 120144 499258 120186 499494
rect 120422 499258 120464 499494
rect 120144 492494 120464 499258
rect 120144 492258 120186 492494
rect 120422 492258 120464 492494
rect 120144 485494 120464 492258
rect 120144 485258 120186 485494
rect 120422 485258 120464 485494
rect 120144 478494 120464 485258
rect 120144 478258 120186 478494
rect 120422 478258 120464 478494
rect 120144 471494 120464 478258
rect 120144 471258 120186 471494
rect 120422 471258 120464 471494
rect 120144 464494 120464 471258
rect 120144 464258 120186 464494
rect 120422 464258 120464 464494
rect 120144 457494 120464 464258
rect 120144 457258 120186 457494
rect 120422 457258 120464 457494
rect 120144 450494 120464 457258
rect 120144 450258 120186 450494
rect 120422 450258 120464 450494
rect 120144 443494 120464 450258
rect 120144 443258 120186 443494
rect 120422 443258 120464 443494
rect 120144 436494 120464 443258
rect 120144 436258 120186 436494
rect 120422 436258 120464 436494
rect 120144 429494 120464 436258
rect 120144 429258 120186 429494
rect 120422 429258 120464 429494
rect 120144 422494 120464 429258
rect 120144 422258 120186 422494
rect 120422 422258 120464 422494
rect 120144 415494 120464 422258
rect 120144 415258 120186 415494
rect 120422 415258 120464 415494
rect 120144 408494 120464 415258
rect 120144 408258 120186 408494
rect 120422 408258 120464 408494
rect 120144 401494 120464 408258
rect 120144 401258 120186 401494
rect 120422 401258 120464 401494
rect 120144 394494 120464 401258
rect 120144 394258 120186 394494
rect 120422 394258 120464 394494
rect 120144 387494 120464 394258
rect 120144 387258 120186 387494
rect 120422 387258 120464 387494
rect 120144 380494 120464 387258
rect 120144 380258 120186 380494
rect 120422 380258 120464 380494
rect 120144 373494 120464 380258
rect 120144 373258 120186 373494
rect 120422 373258 120464 373494
rect 120144 366494 120464 373258
rect 120144 366258 120186 366494
rect 120422 366258 120464 366494
rect 120144 359494 120464 366258
rect 120144 359258 120186 359494
rect 120422 359258 120464 359494
rect 120144 352494 120464 359258
rect 120144 352258 120186 352494
rect 120422 352258 120464 352494
rect 120144 345494 120464 352258
rect 120144 345258 120186 345494
rect 120422 345258 120464 345494
rect 120144 338494 120464 345258
rect 120144 338258 120186 338494
rect 120422 338258 120464 338494
rect 120144 331494 120464 338258
rect 120144 331258 120186 331494
rect 120422 331258 120464 331494
rect 120144 324494 120464 331258
rect 120144 324258 120186 324494
rect 120422 324258 120464 324494
rect 120144 317494 120464 324258
rect 120144 317258 120186 317494
rect 120422 317258 120464 317494
rect 120144 310494 120464 317258
rect 120144 310258 120186 310494
rect 120422 310258 120464 310494
rect 120144 303494 120464 310258
rect 120144 303258 120186 303494
rect 120422 303258 120464 303494
rect 120144 296494 120464 303258
rect 120144 296258 120186 296494
rect 120422 296258 120464 296494
rect 120144 289494 120464 296258
rect 120144 289258 120186 289494
rect 120422 289258 120464 289494
rect 120144 282494 120464 289258
rect 120144 282258 120186 282494
rect 120422 282258 120464 282494
rect 120144 275494 120464 282258
rect 120144 275258 120186 275494
rect 120422 275258 120464 275494
rect 120144 268494 120464 275258
rect 120144 268258 120186 268494
rect 120422 268258 120464 268494
rect 120144 261494 120464 268258
rect 120144 261258 120186 261494
rect 120422 261258 120464 261494
rect 120144 254494 120464 261258
rect 120144 254258 120186 254494
rect 120422 254258 120464 254494
rect 120144 247494 120464 254258
rect 120144 247258 120186 247494
rect 120422 247258 120464 247494
rect 120144 240494 120464 247258
rect 120144 240258 120186 240494
rect 120422 240258 120464 240494
rect 120144 233494 120464 240258
rect 120144 233258 120186 233494
rect 120422 233258 120464 233494
rect 120144 226494 120464 233258
rect 120144 226258 120186 226494
rect 120422 226258 120464 226494
rect 120144 219494 120464 226258
rect 120144 219258 120186 219494
rect 120422 219258 120464 219494
rect 120144 212494 120464 219258
rect 120144 212258 120186 212494
rect 120422 212258 120464 212494
rect 120144 205494 120464 212258
rect 120144 205258 120186 205494
rect 120422 205258 120464 205494
rect 120144 198494 120464 205258
rect 120144 198258 120186 198494
rect 120422 198258 120464 198494
rect 120144 191494 120464 198258
rect 120144 191258 120186 191494
rect 120422 191258 120464 191494
rect 120144 184494 120464 191258
rect 120144 184258 120186 184494
rect 120422 184258 120464 184494
rect 120144 177494 120464 184258
rect 120144 177258 120186 177494
rect 120422 177258 120464 177494
rect 120144 170494 120464 177258
rect 120144 170258 120186 170494
rect 120422 170258 120464 170494
rect 120144 163494 120464 170258
rect 120144 163258 120186 163494
rect 120422 163258 120464 163494
rect 120144 156494 120464 163258
rect 120144 156258 120186 156494
rect 120422 156258 120464 156494
rect 120144 149494 120464 156258
rect 120144 149258 120186 149494
rect 120422 149258 120464 149494
rect 120144 142494 120464 149258
rect 120144 142258 120186 142494
rect 120422 142258 120464 142494
rect 120144 135494 120464 142258
rect 120144 135258 120186 135494
rect 120422 135258 120464 135494
rect 120144 128494 120464 135258
rect 120144 128258 120186 128494
rect 120422 128258 120464 128494
rect 120144 121494 120464 128258
rect 120144 121258 120186 121494
rect 120422 121258 120464 121494
rect 120144 114494 120464 121258
rect 120144 114258 120186 114494
rect 120422 114258 120464 114494
rect 120144 107494 120464 114258
rect 120144 107258 120186 107494
rect 120422 107258 120464 107494
rect 120144 100494 120464 107258
rect 120144 100258 120186 100494
rect 120422 100258 120464 100494
rect 120144 93494 120464 100258
rect 120144 93258 120186 93494
rect 120422 93258 120464 93494
rect 120144 86494 120464 93258
rect 120144 86258 120186 86494
rect 120422 86258 120464 86494
rect 120144 79494 120464 86258
rect 120144 79258 120186 79494
rect 120422 79258 120464 79494
rect 120144 72494 120464 79258
rect 120144 72258 120186 72494
rect 120422 72258 120464 72494
rect 120144 65494 120464 72258
rect 120144 65258 120186 65494
rect 120422 65258 120464 65494
rect 120144 58494 120464 65258
rect 120144 58258 120186 58494
rect 120422 58258 120464 58494
rect 120144 51494 120464 58258
rect 120144 51258 120186 51494
rect 120422 51258 120464 51494
rect 120144 44494 120464 51258
rect 120144 44258 120186 44494
rect 120422 44258 120464 44494
rect 120144 37494 120464 44258
rect 120144 37258 120186 37494
rect 120422 37258 120464 37494
rect 120144 30494 120464 37258
rect 120144 30258 120186 30494
rect 120422 30258 120464 30494
rect 120144 23494 120464 30258
rect 120144 23258 120186 23494
rect 120422 23258 120464 23494
rect 120144 16494 120464 23258
rect 120144 16258 120186 16494
rect 120422 16258 120464 16494
rect 120144 9494 120464 16258
rect 120144 9258 120186 9494
rect 120422 9258 120464 9494
rect 120144 2494 120464 9258
rect 120144 2258 120186 2494
rect 120422 2258 120464 2494
rect 120144 -746 120464 2258
rect 120144 -982 120186 -746
rect 120422 -982 120464 -746
rect 120144 -1066 120464 -982
rect 120144 -1302 120186 -1066
rect 120422 -1302 120464 -1066
rect 120144 -2294 120464 -1302
rect 121876 706198 122196 706230
rect 121876 705962 121918 706198
rect 122154 705962 122196 706198
rect 121876 705878 122196 705962
rect 121876 705642 121918 705878
rect 122154 705642 122196 705878
rect 121876 696434 122196 705642
rect 121876 696198 121918 696434
rect 122154 696198 122196 696434
rect 121876 689434 122196 696198
rect 121876 689198 121918 689434
rect 122154 689198 122196 689434
rect 121876 682434 122196 689198
rect 121876 682198 121918 682434
rect 122154 682198 122196 682434
rect 121876 675434 122196 682198
rect 121876 675198 121918 675434
rect 122154 675198 122196 675434
rect 121876 668434 122196 675198
rect 121876 668198 121918 668434
rect 122154 668198 122196 668434
rect 121876 661434 122196 668198
rect 121876 661198 121918 661434
rect 122154 661198 122196 661434
rect 121876 654434 122196 661198
rect 121876 654198 121918 654434
rect 122154 654198 122196 654434
rect 121876 647434 122196 654198
rect 121876 647198 121918 647434
rect 122154 647198 122196 647434
rect 121876 640434 122196 647198
rect 121876 640198 121918 640434
rect 122154 640198 122196 640434
rect 121876 633434 122196 640198
rect 121876 633198 121918 633434
rect 122154 633198 122196 633434
rect 121876 626434 122196 633198
rect 121876 626198 121918 626434
rect 122154 626198 122196 626434
rect 121876 619434 122196 626198
rect 121876 619198 121918 619434
rect 122154 619198 122196 619434
rect 121876 612434 122196 619198
rect 121876 612198 121918 612434
rect 122154 612198 122196 612434
rect 121876 605434 122196 612198
rect 121876 605198 121918 605434
rect 122154 605198 122196 605434
rect 121876 598434 122196 605198
rect 121876 598198 121918 598434
rect 122154 598198 122196 598434
rect 121876 591434 122196 598198
rect 121876 591198 121918 591434
rect 122154 591198 122196 591434
rect 121876 584434 122196 591198
rect 121876 584198 121918 584434
rect 122154 584198 122196 584434
rect 121876 577434 122196 584198
rect 121876 577198 121918 577434
rect 122154 577198 122196 577434
rect 121876 570434 122196 577198
rect 121876 570198 121918 570434
rect 122154 570198 122196 570434
rect 121876 563434 122196 570198
rect 121876 563198 121918 563434
rect 122154 563198 122196 563434
rect 121876 556434 122196 563198
rect 121876 556198 121918 556434
rect 122154 556198 122196 556434
rect 121876 549434 122196 556198
rect 121876 549198 121918 549434
rect 122154 549198 122196 549434
rect 121876 542434 122196 549198
rect 121876 542198 121918 542434
rect 122154 542198 122196 542434
rect 121876 535434 122196 542198
rect 121876 535198 121918 535434
rect 122154 535198 122196 535434
rect 121876 528434 122196 535198
rect 121876 528198 121918 528434
rect 122154 528198 122196 528434
rect 121876 521434 122196 528198
rect 121876 521198 121918 521434
rect 122154 521198 122196 521434
rect 121876 514434 122196 521198
rect 121876 514198 121918 514434
rect 122154 514198 122196 514434
rect 121876 507434 122196 514198
rect 121876 507198 121918 507434
rect 122154 507198 122196 507434
rect 121876 500434 122196 507198
rect 121876 500198 121918 500434
rect 122154 500198 122196 500434
rect 121876 493434 122196 500198
rect 121876 493198 121918 493434
rect 122154 493198 122196 493434
rect 121876 486434 122196 493198
rect 121876 486198 121918 486434
rect 122154 486198 122196 486434
rect 121876 479434 122196 486198
rect 121876 479198 121918 479434
rect 122154 479198 122196 479434
rect 121876 472434 122196 479198
rect 121876 472198 121918 472434
rect 122154 472198 122196 472434
rect 121876 465434 122196 472198
rect 121876 465198 121918 465434
rect 122154 465198 122196 465434
rect 121876 458434 122196 465198
rect 121876 458198 121918 458434
rect 122154 458198 122196 458434
rect 121876 451434 122196 458198
rect 121876 451198 121918 451434
rect 122154 451198 122196 451434
rect 121876 444434 122196 451198
rect 121876 444198 121918 444434
rect 122154 444198 122196 444434
rect 121876 437434 122196 444198
rect 121876 437198 121918 437434
rect 122154 437198 122196 437434
rect 121876 430434 122196 437198
rect 121876 430198 121918 430434
rect 122154 430198 122196 430434
rect 121876 423434 122196 430198
rect 121876 423198 121918 423434
rect 122154 423198 122196 423434
rect 121876 416434 122196 423198
rect 121876 416198 121918 416434
rect 122154 416198 122196 416434
rect 121876 409434 122196 416198
rect 121876 409198 121918 409434
rect 122154 409198 122196 409434
rect 121876 402434 122196 409198
rect 121876 402198 121918 402434
rect 122154 402198 122196 402434
rect 121876 395434 122196 402198
rect 121876 395198 121918 395434
rect 122154 395198 122196 395434
rect 121876 388434 122196 395198
rect 121876 388198 121918 388434
rect 122154 388198 122196 388434
rect 121876 381434 122196 388198
rect 121876 381198 121918 381434
rect 122154 381198 122196 381434
rect 121876 374434 122196 381198
rect 121876 374198 121918 374434
rect 122154 374198 122196 374434
rect 121876 367434 122196 374198
rect 121876 367198 121918 367434
rect 122154 367198 122196 367434
rect 121876 360434 122196 367198
rect 121876 360198 121918 360434
rect 122154 360198 122196 360434
rect 121876 353434 122196 360198
rect 121876 353198 121918 353434
rect 122154 353198 122196 353434
rect 121876 346434 122196 353198
rect 121876 346198 121918 346434
rect 122154 346198 122196 346434
rect 121876 339434 122196 346198
rect 121876 339198 121918 339434
rect 122154 339198 122196 339434
rect 121876 332434 122196 339198
rect 121876 332198 121918 332434
rect 122154 332198 122196 332434
rect 121876 325434 122196 332198
rect 121876 325198 121918 325434
rect 122154 325198 122196 325434
rect 121876 318434 122196 325198
rect 121876 318198 121918 318434
rect 122154 318198 122196 318434
rect 121876 311434 122196 318198
rect 121876 311198 121918 311434
rect 122154 311198 122196 311434
rect 121876 304434 122196 311198
rect 121876 304198 121918 304434
rect 122154 304198 122196 304434
rect 121876 297434 122196 304198
rect 121876 297198 121918 297434
rect 122154 297198 122196 297434
rect 121876 290434 122196 297198
rect 121876 290198 121918 290434
rect 122154 290198 122196 290434
rect 121876 283434 122196 290198
rect 121876 283198 121918 283434
rect 122154 283198 122196 283434
rect 121876 276434 122196 283198
rect 121876 276198 121918 276434
rect 122154 276198 122196 276434
rect 121876 269434 122196 276198
rect 121876 269198 121918 269434
rect 122154 269198 122196 269434
rect 121876 262434 122196 269198
rect 121876 262198 121918 262434
rect 122154 262198 122196 262434
rect 121876 255434 122196 262198
rect 121876 255198 121918 255434
rect 122154 255198 122196 255434
rect 121876 248434 122196 255198
rect 121876 248198 121918 248434
rect 122154 248198 122196 248434
rect 121876 241434 122196 248198
rect 121876 241198 121918 241434
rect 122154 241198 122196 241434
rect 121876 234434 122196 241198
rect 121876 234198 121918 234434
rect 122154 234198 122196 234434
rect 121876 227434 122196 234198
rect 121876 227198 121918 227434
rect 122154 227198 122196 227434
rect 121876 220434 122196 227198
rect 121876 220198 121918 220434
rect 122154 220198 122196 220434
rect 121876 213434 122196 220198
rect 121876 213198 121918 213434
rect 122154 213198 122196 213434
rect 121876 206434 122196 213198
rect 121876 206198 121918 206434
rect 122154 206198 122196 206434
rect 121876 199434 122196 206198
rect 121876 199198 121918 199434
rect 122154 199198 122196 199434
rect 121876 192434 122196 199198
rect 121876 192198 121918 192434
rect 122154 192198 122196 192434
rect 121876 185434 122196 192198
rect 121876 185198 121918 185434
rect 122154 185198 122196 185434
rect 121876 178434 122196 185198
rect 121876 178198 121918 178434
rect 122154 178198 122196 178434
rect 121876 171434 122196 178198
rect 121876 171198 121918 171434
rect 122154 171198 122196 171434
rect 121876 164434 122196 171198
rect 121876 164198 121918 164434
rect 122154 164198 122196 164434
rect 121876 157434 122196 164198
rect 121876 157198 121918 157434
rect 122154 157198 122196 157434
rect 121876 150434 122196 157198
rect 121876 150198 121918 150434
rect 122154 150198 122196 150434
rect 121876 143434 122196 150198
rect 121876 143198 121918 143434
rect 122154 143198 122196 143434
rect 121876 136434 122196 143198
rect 121876 136198 121918 136434
rect 122154 136198 122196 136434
rect 121876 129434 122196 136198
rect 121876 129198 121918 129434
rect 122154 129198 122196 129434
rect 121876 122434 122196 129198
rect 121876 122198 121918 122434
rect 122154 122198 122196 122434
rect 121876 115434 122196 122198
rect 121876 115198 121918 115434
rect 122154 115198 122196 115434
rect 121876 108434 122196 115198
rect 121876 108198 121918 108434
rect 122154 108198 122196 108434
rect 121876 101434 122196 108198
rect 121876 101198 121918 101434
rect 122154 101198 122196 101434
rect 121876 94434 122196 101198
rect 121876 94198 121918 94434
rect 122154 94198 122196 94434
rect 121876 87434 122196 94198
rect 121876 87198 121918 87434
rect 122154 87198 122196 87434
rect 121876 80434 122196 87198
rect 121876 80198 121918 80434
rect 122154 80198 122196 80434
rect 121876 73434 122196 80198
rect 121876 73198 121918 73434
rect 122154 73198 122196 73434
rect 121876 66434 122196 73198
rect 121876 66198 121918 66434
rect 122154 66198 122196 66434
rect 121876 59434 122196 66198
rect 121876 59198 121918 59434
rect 122154 59198 122196 59434
rect 121876 52434 122196 59198
rect 121876 52198 121918 52434
rect 122154 52198 122196 52434
rect 121876 45434 122196 52198
rect 121876 45198 121918 45434
rect 122154 45198 122196 45434
rect 121876 38434 122196 45198
rect 121876 38198 121918 38434
rect 122154 38198 122196 38434
rect 121876 31434 122196 38198
rect 121876 31198 121918 31434
rect 122154 31198 122196 31434
rect 121876 24434 122196 31198
rect 121876 24198 121918 24434
rect 122154 24198 122196 24434
rect 121876 17434 122196 24198
rect 121876 17198 121918 17434
rect 122154 17198 122196 17434
rect 121876 10434 122196 17198
rect 121876 10198 121918 10434
rect 122154 10198 122196 10434
rect 121876 3434 122196 10198
rect 121876 3198 121918 3434
rect 122154 3198 122196 3434
rect 121876 -1706 122196 3198
rect 121876 -1942 121918 -1706
rect 122154 -1942 122196 -1706
rect 121876 -2026 122196 -1942
rect 121876 -2262 121918 -2026
rect 122154 -2262 122196 -2026
rect 121876 -2294 122196 -2262
rect 127144 705238 127464 706230
rect 127144 705002 127186 705238
rect 127422 705002 127464 705238
rect 127144 704918 127464 705002
rect 127144 704682 127186 704918
rect 127422 704682 127464 704918
rect 127144 695494 127464 704682
rect 127144 695258 127186 695494
rect 127422 695258 127464 695494
rect 127144 688494 127464 695258
rect 127144 688258 127186 688494
rect 127422 688258 127464 688494
rect 127144 681494 127464 688258
rect 127144 681258 127186 681494
rect 127422 681258 127464 681494
rect 127144 674494 127464 681258
rect 127144 674258 127186 674494
rect 127422 674258 127464 674494
rect 127144 667494 127464 674258
rect 127144 667258 127186 667494
rect 127422 667258 127464 667494
rect 127144 660494 127464 667258
rect 127144 660258 127186 660494
rect 127422 660258 127464 660494
rect 127144 653494 127464 660258
rect 127144 653258 127186 653494
rect 127422 653258 127464 653494
rect 127144 646494 127464 653258
rect 127144 646258 127186 646494
rect 127422 646258 127464 646494
rect 127144 639494 127464 646258
rect 127144 639258 127186 639494
rect 127422 639258 127464 639494
rect 127144 632494 127464 639258
rect 127144 632258 127186 632494
rect 127422 632258 127464 632494
rect 127144 625494 127464 632258
rect 127144 625258 127186 625494
rect 127422 625258 127464 625494
rect 127144 618494 127464 625258
rect 127144 618258 127186 618494
rect 127422 618258 127464 618494
rect 127144 611494 127464 618258
rect 127144 611258 127186 611494
rect 127422 611258 127464 611494
rect 127144 604494 127464 611258
rect 127144 604258 127186 604494
rect 127422 604258 127464 604494
rect 127144 597494 127464 604258
rect 127144 597258 127186 597494
rect 127422 597258 127464 597494
rect 127144 590494 127464 597258
rect 127144 590258 127186 590494
rect 127422 590258 127464 590494
rect 127144 583494 127464 590258
rect 127144 583258 127186 583494
rect 127422 583258 127464 583494
rect 127144 576494 127464 583258
rect 127144 576258 127186 576494
rect 127422 576258 127464 576494
rect 127144 569494 127464 576258
rect 127144 569258 127186 569494
rect 127422 569258 127464 569494
rect 127144 562494 127464 569258
rect 127144 562258 127186 562494
rect 127422 562258 127464 562494
rect 127144 555494 127464 562258
rect 127144 555258 127186 555494
rect 127422 555258 127464 555494
rect 127144 548494 127464 555258
rect 127144 548258 127186 548494
rect 127422 548258 127464 548494
rect 127144 541494 127464 548258
rect 127144 541258 127186 541494
rect 127422 541258 127464 541494
rect 127144 534494 127464 541258
rect 127144 534258 127186 534494
rect 127422 534258 127464 534494
rect 127144 527494 127464 534258
rect 127144 527258 127186 527494
rect 127422 527258 127464 527494
rect 127144 520494 127464 527258
rect 127144 520258 127186 520494
rect 127422 520258 127464 520494
rect 127144 513494 127464 520258
rect 127144 513258 127186 513494
rect 127422 513258 127464 513494
rect 127144 506494 127464 513258
rect 127144 506258 127186 506494
rect 127422 506258 127464 506494
rect 127144 499494 127464 506258
rect 127144 499258 127186 499494
rect 127422 499258 127464 499494
rect 127144 492494 127464 499258
rect 127144 492258 127186 492494
rect 127422 492258 127464 492494
rect 127144 485494 127464 492258
rect 127144 485258 127186 485494
rect 127422 485258 127464 485494
rect 127144 478494 127464 485258
rect 127144 478258 127186 478494
rect 127422 478258 127464 478494
rect 127144 471494 127464 478258
rect 127144 471258 127186 471494
rect 127422 471258 127464 471494
rect 127144 464494 127464 471258
rect 127144 464258 127186 464494
rect 127422 464258 127464 464494
rect 127144 457494 127464 464258
rect 127144 457258 127186 457494
rect 127422 457258 127464 457494
rect 127144 450494 127464 457258
rect 127144 450258 127186 450494
rect 127422 450258 127464 450494
rect 127144 443494 127464 450258
rect 127144 443258 127186 443494
rect 127422 443258 127464 443494
rect 127144 436494 127464 443258
rect 127144 436258 127186 436494
rect 127422 436258 127464 436494
rect 127144 429494 127464 436258
rect 127144 429258 127186 429494
rect 127422 429258 127464 429494
rect 127144 422494 127464 429258
rect 127144 422258 127186 422494
rect 127422 422258 127464 422494
rect 127144 415494 127464 422258
rect 127144 415258 127186 415494
rect 127422 415258 127464 415494
rect 127144 408494 127464 415258
rect 127144 408258 127186 408494
rect 127422 408258 127464 408494
rect 127144 401494 127464 408258
rect 127144 401258 127186 401494
rect 127422 401258 127464 401494
rect 127144 394494 127464 401258
rect 127144 394258 127186 394494
rect 127422 394258 127464 394494
rect 127144 387494 127464 394258
rect 127144 387258 127186 387494
rect 127422 387258 127464 387494
rect 127144 380494 127464 387258
rect 127144 380258 127186 380494
rect 127422 380258 127464 380494
rect 127144 373494 127464 380258
rect 127144 373258 127186 373494
rect 127422 373258 127464 373494
rect 127144 366494 127464 373258
rect 127144 366258 127186 366494
rect 127422 366258 127464 366494
rect 127144 359494 127464 366258
rect 127144 359258 127186 359494
rect 127422 359258 127464 359494
rect 127144 352494 127464 359258
rect 127144 352258 127186 352494
rect 127422 352258 127464 352494
rect 127144 345494 127464 352258
rect 127144 345258 127186 345494
rect 127422 345258 127464 345494
rect 127144 338494 127464 345258
rect 127144 338258 127186 338494
rect 127422 338258 127464 338494
rect 127144 331494 127464 338258
rect 127144 331258 127186 331494
rect 127422 331258 127464 331494
rect 127144 324494 127464 331258
rect 127144 324258 127186 324494
rect 127422 324258 127464 324494
rect 127144 317494 127464 324258
rect 127144 317258 127186 317494
rect 127422 317258 127464 317494
rect 127144 310494 127464 317258
rect 127144 310258 127186 310494
rect 127422 310258 127464 310494
rect 127144 303494 127464 310258
rect 127144 303258 127186 303494
rect 127422 303258 127464 303494
rect 127144 296494 127464 303258
rect 127144 296258 127186 296494
rect 127422 296258 127464 296494
rect 127144 289494 127464 296258
rect 127144 289258 127186 289494
rect 127422 289258 127464 289494
rect 127144 282494 127464 289258
rect 127144 282258 127186 282494
rect 127422 282258 127464 282494
rect 127144 275494 127464 282258
rect 127144 275258 127186 275494
rect 127422 275258 127464 275494
rect 127144 268494 127464 275258
rect 127144 268258 127186 268494
rect 127422 268258 127464 268494
rect 127144 261494 127464 268258
rect 127144 261258 127186 261494
rect 127422 261258 127464 261494
rect 127144 254494 127464 261258
rect 127144 254258 127186 254494
rect 127422 254258 127464 254494
rect 127144 247494 127464 254258
rect 127144 247258 127186 247494
rect 127422 247258 127464 247494
rect 127144 240494 127464 247258
rect 127144 240258 127186 240494
rect 127422 240258 127464 240494
rect 127144 233494 127464 240258
rect 127144 233258 127186 233494
rect 127422 233258 127464 233494
rect 127144 226494 127464 233258
rect 127144 226258 127186 226494
rect 127422 226258 127464 226494
rect 127144 219494 127464 226258
rect 127144 219258 127186 219494
rect 127422 219258 127464 219494
rect 127144 212494 127464 219258
rect 127144 212258 127186 212494
rect 127422 212258 127464 212494
rect 127144 205494 127464 212258
rect 127144 205258 127186 205494
rect 127422 205258 127464 205494
rect 127144 198494 127464 205258
rect 127144 198258 127186 198494
rect 127422 198258 127464 198494
rect 127144 191494 127464 198258
rect 127144 191258 127186 191494
rect 127422 191258 127464 191494
rect 127144 184494 127464 191258
rect 127144 184258 127186 184494
rect 127422 184258 127464 184494
rect 127144 177494 127464 184258
rect 127144 177258 127186 177494
rect 127422 177258 127464 177494
rect 127144 170494 127464 177258
rect 127144 170258 127186 170494
rect 127422 170258 127464 170494
rect 127144 163494 127464 170258
rect 127144 163258 127186 163494
rect 127422 163258 127464 163494
rect 127144 156494 127464 163258
rect 127144 156258 127186 156494
rect 127422 156258 127464 156494
rect 127144 149494 127464 156258
rect 127144 149258 127186 149494
rect 127422 149258 127464 149494
rect 127144 142494 127464 149258
rect 127144 142258 127186 142494
rect 127422 142258 127464 142494
rect 127144 135494 127464 142258
rect 127144 135258 127186 135494
rect 127422 135258 127464 135494
rect 127144 128494 127464 135258
rect 127144 128258 127186 128494
rect 127422 128258 127464 128494
rect 127144 121494 127464 128258
rect 127144 121258 127186 121494
rect 127422 121258 127464 121494
rect 127144 114494 127464 121258
rect 127144 114258 127186 114494
rect 127422 114258 127464 114494
rect 127144 107494 127464 114258
rect 127144 107258 127186 107494
rect 127422 107258 127464 107494
rect 127144 100494 127464 107258
rect 127144 100258 127186 100494
rect 127422 100258 127464 100494
rect 127144 93494 127464 100258
rect 127144 93258 127186 93494
rect 127422 93258 127464 93494
rect 127144 86494 127464 93258
rect 127144 86258 127186 86494
rect 127422 86258 127464 86494
rect 127144 79494 127464 86258
rect 127144 79258 127186 79494
rect 127422 79258 127464 79494
rect 127144 72494 127464 79258
rect 127144 72258 127186 72494
rect 127422 72258 127464 72494
rect 127144 65494 127464 72258
rect 127144 65258 127186 65494
rect 127422 65258 127464 65494
rect 127144 58494 127464 65258
rect 127144 58258 127186 58494
rect 127422 58258 127464 58494
rect 127144 51494 127464 58258
rect 127144 51258 127186 51494
rect 127422 51258 127464 51494
rect 127144 44494 127464 51258
rect 127144 44258 127186 44494
rect 127422 44258 127464 44494
rect 127144 37494 127464 44258
rect 127144 37258 127186 37494
rect 127422 37258 127464 37494
rect 127144 30494 127464 37258
rect 127144 30258 127186 30494
rect 127422 30258 127464 30494
rect 127144 23494 127464 30258
rect 127144 23258 127186 23494
rect 127422 23258 127464 23494
rect 127144 16494 127464 23258
rect 127144 16258 127186 16494
rect 127422 16258 127464 16494
rect 127144 9494 127464 16258
rect 127144 9258 127186 9494
rect 127422 9258 127464 9494
rect 127144 2494 127464 9258
rect 127144 2258 127186 2494
rect 127422 2258 127464 2494
rect 127144 -746 127464 2258
rect 127144 -982 127186 -746
rect 127422 -982 127464 -746
rect 127144 -1066 127464 -982
rect 127144 -1302 127186 -1066
rect 127422 -1302 127464 -1066
rect 127144 -2294 127464 -1302
rect 128876 706198 129196 706230
rect 128876 705962 128918 706198
rect 129154 705962 129196 706198
rect 128876 705878 129196 705962
rect 128876 705642 128918 705878
rect 129154 705642 129196 705878
rect 128876 696434 129196 705642
rect 128876 696198 128918 696434
rect 129154 696198 129196 696434
rect 128876 689434 129196 696198
rect 128876 689198 128918 689434
rect 129154 689198 129196 689434
rect 128876 682434 129196 689198
rect 128876 682198 128918 682434
rect 129154 682198 129196 682434
rect 128876 675434 129196 682198
rect 128876 675198 128918 675434
rect 129154 675198 129196 675434
rect 128876 668434 129196 675198
rect 128876 668198 128918 668434
rect 129154 668198 129196 668434
rect 128876 661434 129196 668198
rect 128876 661198 128918 661434
rect 129154 661198 129196 661434
rect 128876 654434 129196 661198
rect 128876 654198 128918 654434
rect 129154 654198 129196 654434
rect 128876 647434 129196 654198
rect 128876 647198 128918 647434
rect 129154 647198 129196 647434
rect 128876 640434 129196 647198
rect 128876 640198 128918 640434
rect 129154 640198 129196 640434
rect 128876 633434 129196 640198
rect 128876 633198 128918 633434
rect 129154 633198 129196 633434
rect 128876 626434 129196 633198
rect 128876 626198 128918 626434
rect 129154 626198 129196 626434
rect 128876 619434 129196 626198
rect 128876 619198 128918 619434
rect 129154 619198 129196 619434
rect 128876 612434 129196 619198
rect 128876 612198 128918 612434
rect 129154 612198 129196 612434
rect 128876 605434 129196 612198
rect 128876 605198 128918 605434
rect 129154 605198 129196 605434
rect 128876 598434 129196 605198
rect 128876 598198 128918 598434
rect 129154 598198 129196 598434
rect 128876 591434 129196 598198
rect 128876 591198 128918 591434
rect 129154 591198 129196 591434
rect 128876 584434 129196 591198
rect 128876 584198 128918 584434
rect 129154 584198 129196 584434
rect 128876 577434 129196 584198
rect 128876 577198 128918 577434
rect 129154 577198 129196 577434
rect 128876 570434 129196 577198
rect 128876 570198 128918 570434
rect 129154 570198 129196 570434
rect 128876 563434 129196 570198
rect 128876 563198 128918 563434
rect 129154 563198 129196 563434
rect 128876 556434 129196 563198
rect 128876 556198 128918 556434
rect 129154 556198 129196 556434
rect 128876 549434 129196 556198
rect 128876 549198 128918 549434
rect 129154 549198 129196 549434
rect 128876 542434 129196 549198
rect 128876 542198 128918 542434
rect 129154 542198 129196 542434
rect 128876 535434 129196 542198
rect 128876 535198 128918 535434
rect 129154 535198 129196 535434
rect 128876 528434 129196 535198
rect 128876 528198 128918 528434
rect 129154 528198 129196 528434
rect 128876 521434 129196 528198
rect 128876 521198 128918 521434
rect 129154 521198 129196 521434
rect 128876 514434 129196 521198
rect 128876 514198 128918 514434
rect 129154 514198 129196 514434
rect 128876 507434 129196 514198
rect 128876 507198 128918 507434
rect 129154 507198 129196 507434
rect 128876 500434 129196 507198
rect 128876 500198 128918 500434
rect 129154 500198 129196 500434
rect 128876 493434 129196 500198
rect 128876 493198 128918 493434
rect 129154 493198 129196 493434
rect 128876 486434 129196 493198
rect 128876 486198 128918 486434
rect 129154 486198 129196 486434
rect 128876 479434 129196 486198
rect 128876 479198 128918 479434
rect 129154 479198 129196 479434
rect 128876 472434 129196 479198
rect 128876 472198 128918 472434
rect 129154 472198 129196 472434
rect 128876 465434 129196 472198
rect 128876 465198 128918 465434
rect 129154 465198 129196 465434
rect 128876 458434 129196 465198
rect 128876 458198 128918 458434
rect 129154 458198 129196 458434
rect 128876 451434 129196 458198
rect 128876 451198 128918 451434
rect 129154 451198 129196 451434
rect 128876 444434 129196 451198
rect 128876 444198 128918 444434
rect 129154 444198 129196 444434
rect 128876 437434 129196 444198
rect 128876 437198 128918 437434
rect 129154 437198 129196 437434
rect 128876 430434 129196 437198
rect 128876 430198 128918 430434
rect 129154 430198 129196 430434
rect 128876 423434 129196 430198
rect 128876 423198 128918 423434
rect 129154 423198 129196 423434
rect 128876 416434 129196 423198
rect 128876 416198 128918 416434
rect 129154 416198 129196 416434
rect 128876 409434 129196 416198
rect 128876 409198 128918 409434
rect 129154 409198 129196 409434
rect 128876 402434 129196 409198
rect 128876 402198 128918 402434
rect 129154 402198 129196 402434
rect 128876 395434 129196 402198
rect 128876 395198 128918 395434
rect 129154 395198 129196 395434
rect 128876 388434 129196 395198
rect 128876 388198 128918 388434
rect 129154 388198 129196 388434
rect 128876 381434 129196 388198
rect 128876 381198 128918 381434
rect 129154 381198 129196 381434
rect 128876 374434 129196 381198
rect 128876 374198 128918 374434
rect 129154 374198 129196 374434
rect 128876 367434 129196 374198
rect 128876 367198 128918 367434
rect 129154 367198 129196 367434
rect 128876 360434 129196 367198
rect 128876 360198 128918 360434
rect 129154 360198 129196 360434
rect 128876 353434 129196 360198
rect 128876 353198 128918 353434
rect 129154 353198 129196 353434
rect 128876 346434 129196 353198
rect 128876 346198 128918 346434
rect 129154 346198 129196 346434
rect 128876 339434 129196 346198
rect 128876 339198 128918 339434
rect 129154 339198 129196 339434
rect 128876 332434 129196 339198
rect 128876 332198 128918 332434
rect 129154 332198 129196 332434
rect 128876 325434 129196 332198
rect 128876 325198 128918 325434
rect 129154 325198 129196 325434
rect 128876 318434 129196 325198
rect 128876 318198 128918 318434
rect 129154 318198 129196 318434
rect 128876 311434 129196 318198
rect 128876 311198 128918 311434
rect 129154 311198 129196 311434
rect 128876 304434 129196 311198
rect 128876 304198 128918 304434
rect 129154 304198 129196 304434
rect 128876 297434 129196 304198
rect 128876 297198 128918 297434
rect 129154 297198 129196 297434
rect 128876 290434 129196 297198
rect 128876 290198 128918 290434
rect 129154 290198 129196 290434
rect 128876 283434 129196 290198
rect 128876 283198 128918 283434
rect 129154 283198 129196 283434
rect 128876 276434 129196 283198
rect 128876 276198 128918 276434
rect 129154 276198 129196 276434
rect 128876 269434 129196 276198
rect 128876 269198 128918 269434
rect 129154 269198 129196 269434
rect 128876 262434 129196 269198
rect 128876 262198 128918 262434
rect 129154 262198 129196 262434
rect 128876 255434 129196 262198
rect 128876 255198 128918 255434
rect 129154 255198 129196 255434
rect 128876 248434 129196 255198
rect 128876 248198 128918 248434
rect 129154 248198 129196 248434
rect 128876 241434 129196 248198
rect 128876 241198 128918 241434
rect 129154 241198 129196 241434
rect 128876 234434 129196 241198
rect 128876 234198 128918 234434
rect 129154 234198 129196 234434
rect 128876 227434 129196 234198
rect 128876 227198 128918 227434
rect 129154 227198 129196 227434
rect 128876 220434 129196 227198
rect 128876 220198 128918 220434
rect 129154 220198 129196 220434
rect 128876 213434 129196 220198
rect 128876 213198 128918 213434
rect 129154 213198 129196 213434
rect 128876 206434 129196 213198
rect 128876 206198 128918 206434
rect 129154 206198 129196 206434
rect 128876 199434 129196 206198
rect 128876 199198 128918 199434
rect 129154 199198 129196 199434
rect 128876 192434 129196 199198
rect 128876 192198 128918 192434
rect 129154 192198 129196 192434
rect 128876 185434 129196 192198
rect 128876 185198 128918 185434
rect 129154 185198 129196 185434
rect 128876 178434 129196 185198
rect 128876 178198 128918 178434
rect 129154 178198 129196 178434
rect 128876 171434 129196 178198
rect 128876 171198 128918 171434
rect 129154 171198 129196 171434
rect 128876 164434 129196 171198
rect 128876 164198 128918 164434
rect 129154 164198 129196 164434
rect 128876 157434 129196 164198
rect 128876 157198 128918 157434
rect 129154 157198 129196 157434
rect 128876 150434 129196 157198
rect 128876 150198 128918 150434
rect 129154 150198 129196 150434
rect 128876 143434 129196 150198
rect 128876 143198 128918 143434
rect 129154 143198 129196 143434
rect 128876 136434 129196 143198
rect 128876 136198 128918 136434
rect 129154 136198 129196 136434
rect 128876 129434 129196 136198
rect 128876 129198 128918 129434
rect 129154 129198 129196 129434
rect 128876 122434 129196 129198
rect 128876 122198 128918 122434
rect 129154 122198 129196 122434
rect 128876 115434 129196 122198
rect 128876 115198 128918 115434
rect 129154 115198 129196 115434
rect 128876 108434 129196 115198
rect 128876 108198 128918 108434
rect 129154 108198 129196 108434
rect 128876 101434 129196 108198
rect 128876 101198 128918 101434
rect 129154 101198 129196 101434
rect 128876 94434 129196 101198
rect 128876 94198 128918 94434
rect 129154 94198 129196 94434
rect 128876 87434 129196 94198
rect 128876 87198 128918 87434
rect 129154 87198 129196 87434
rect 128876 80434 129196 87198
rect 128876 80198 128918 80434
rect 129154 80198 129196 80434
rect 128876 73434 129196 80198
rect 128876 73198 128918 73434
rect 129154 73198 129196 73434
rect 128876 66434 129196 73198
rect 128876 66198 128918 66434
rect 129154 66198 129196 66434
rect 128876 59434 129196 66198
rect 128876 59198 128918 59434
rect 129154 59198 129196 59434
rect 128876 52434 129196 59198
rect 128876 52198 128918 52434
rect 129154 52198 129196 52434
rect 128876 45434 129196 52198
rect 128876 45198 128918 45434
rect 129154 45198 129196 45434
rect 128876 38434 129196 45198
rect 128876 38198 128918 38434
rect 129154 38198 129196 38434
rect 128876 31434 129196 38198
rect 128876 31198 128918 31434
rect 129154 31198 129196 31434
rect 128876 24434 129196 31198
rect 128876 24198 128918 24434
rect 129154 24198 129196 24434
rect 128876 17434 129196 24198
rect 128876 17198 128918 17434
rect 129154 17198 129196 17434
rect 128876 10434 129196 17198
rect 128876 10198 128918 10434
rect 129154 10198 129196 10434
rect 128876 3434 129196 10198
rect 128876 3198 128918 3434
rect 129154 3198 129196 3434
rect 128876 -1706 129196 3198
rect 128876 -1942 128918 -1706
rect 129154 -1942 129196 -1706
rect 128876 -2026 129196 -1942
rect 128876 -2262 128918 -2026
rect 129154 -2262 129196 -2026
rect 128876 -2294 129196 -2262
rect 134144 705238 134464 706230
rect 134144 705002 134186 705238
rect 134422 705002 134464 705238
rect 134144 704918 134464 705002
rect 134144 704682 134186 704918
rect 134422 704682 134464 704918
rect 134144 695494 134464 704682
rect 134144 695258 134186 695494
rect 134422 695258 134464 695494
rect 134144 688494 134464 695258
rect 134144 688258 134186 688494
rect 134422 688258 134464 688494
rect 134144 681494 134464 688258
rect 134144 681258 134186 681494
rect 134422 681258 134464 681494
rect 134144 674494 134464 681258
rect 134144 674258 134186 674494
rect 134422 674258 134464 674494
rect 134144 667494 134464 674258
rect 134144 667258 134186 667494
rect 134422 667258 134464 667494
rect 134144 660494 134464 667258
rect 134144 660258 134186 660494
rect 134422 660258 134464 660494
rect 134144 653494 134464 660258
rect 134144 653258 134186 653494
rect 134422 653258 134464 653494
rect 134144 646494 134464 653258
rect 134144 646258 134186 646494
rect 134422 646258 134464 646494
rect 134144 639494 134464 646258
rect 134144 639258 134186 639494
rect 134422 639258 134464 639494
rect 134144 632494 134464 639258
rect 134144 632258 134186 632494
rect 134422 632258 134464 632494
rect 134144 625494 134464 632258
rect 134144 625258 134186 625494
rect 134422 625258 134464 625494
rect 134144 618494 134464 625258
rect 134144 618258 134186 618494
rect 134422 618258 134464 618494
rect 134144 611494 134464 618258
rect 134144 611258 134186 611494
rect 134422 611258 134464 611494
rect 134144 604494 134464 611258
rect 134144 604258 134186 604494
rect 134422 604258 134464 604494
rect 134144 597494 134464 604258
rect 134144 597258 134186 597494
rect 134422 597258 134464 597494
rect 134144 590494 134464 597258
rect 134144 590258 134186 590494
rect 134422 590258 134464 590494
rect 134144 583494 134464 590258
rect 134144 583258 134186 583494
rect 134422 583258 134464 583494
rect 134144 576494 134464 583258
rect 134144 576258 134186 576494
rect 134422 576258 134464 576494
rect 134144 569494 134464 576258
rect 134144 569258 134186 569494
rect 134422 569258 134464 569494
rect 134144 562494 134464 569258
rect 134144 562258 134186 562494
rect 134422 562258 134464 562494
rect 134144 555494 134464 562258
rect 134144 555258 134186 555494
rect 134422 555258 134464 555494
rect 134144 548494 134464 555258
rect 134144 548258 134186 548494
rect 134422 548258 134464 548494
rect 134144 541494 134464 548258
rect 134144 541258 134186 541494
rect 134422 541258 134464 541494
rect 134144 534494 134464 541258
rect 134144 534258 134186 534494
rect 134422 534258 134464 534494
rect 134144 527494 134464 534258
rect 134144 527258 134186 527494
rect 134422 527258 134464 527494
rect 134144 520494 134464 527258
rect 134144 520258 134186 520494
rect 134422 520258 134464 520494
rect 134144 513494 134464 520258
rect 134144 513258 134186 513494
rect 134422 513258 134464 513494
rect 134144 506494 134464 513258
rect 134144 506258 134186 506494
rect 134422 506258 134464 506494
rect 134144 499494 134464 506258
rect 134144 499258 134186 499494
rect 134422 499258 134464 499494
rect 134144 492494 134464 499258
rect 134144 492258 134186 492494
rect 134422 492258 134464 492494
rect 134144 485494 134464 492258
rect 134144 485258 134186 485494
rect 134422 485258 134464 485494
rect 134144 478494 134464 485258
rect 134144 478258 134186 478494
rect 134422 478258 134464 478494
rect 134144 471494 134464 478258
rect 134144 471258 134186 471494
rect 134422 471258 134464 471494
rect 134144 464494 134464 471258
rect 134144 464258 134186 464494
rect 134422 464258 134464 464494
rect 134144 457494 134464 464258
rect 134144 457258 134186 457494
rect 134422 457258 134464 457494
rect 134144 450494 134464 457258
rect 134144 450258 134186 450494
rect 134422 450258 134464 450494
rect 134144 443494 134464 450258
rect 134144 443258 134186 443494
rect 134422 443258 134464 443494
rect 134144 436494 134464 443258
rect 134144 436258 134186 436494
rect 134422 436258 134464 436494
rect 134144 429494 134464 436258
rect 134144 429258 134186 429494
rect 134422 429258 134464 429494
rect 134144 422494 134464 429258
rect 134144 422258 134186 422494
rect 134422 422258 134464 422494
rect 134144 415494 134464 422258
rect 134144 415258 134186 415494
rect 134422 415258 134464 415494
rect 134144 408494 134464 415258
rect 134144 408258 134186 408494
rect 134422 408258 134464 408494
rect 134144 401494 134464 408258
rect 134144 401258 134186 401494
rect 134422 401258 134464 401494
rect 134144 394494 134464 401258
rect 134144 394258 134186 394494
rect 134422 394258 134464 394494
rect 134144 387494 134464 394258
rect 134144 387258 134186 387494
rect 134422 387258 134464 387494
rect 134144 380494 134464 387258
rect 134144 380258 134186 380494
rect 134422 380258 134464 380494
rect 134144 373494 134464 380258
rect 134144 373258 134186 373494
rect 134422 373258 134464 373494
rect 134144 366494 134464 373258
rect 134144 366258 134186 366494
rect 134422 366258 134464 366494
rect 134144 359494 134464 366258
rect 134144 359258 134186 359494
rect 134422 359258 134464 359494
rect 134144 352494 134464 359258
rect 134144 352258 134186 352494
rect 134422 352258 134464 352494
rect 134144 345494 134464 352258
rect 134144 345258 134186 345494
rect 134422 345258 134464 345494
rect 134144 338494 134464 345258
rect 134144 338258 134186 338494
rect 134422 338258 134464 338494
rect 134144 331494 134464 338258
rect 134144 331258 134186 331494
rect 134422 331258 134464 331494
rect 134144 324494 134464 331258
rect 134144 324258 134186 324494
rect 134422 324258 134464 324494
rect 134144 317494 134464 324258
rect 134144 317258 134186 317494
rect 134422 317258 134464 317494
rect 134144 310494 134464 317258
rect 134144 310258 134186 310494
rect 134422 310258 134464 310494
rect 134144 303494 134464 310258
rect 134144 303258 134186 303494
rect 134422 303258 134464 303494
rect 134144 296494 134464 303258
rect 134144 296258 134186 296494
rect 134422 296258 134464 296494
rect 134144 289494 134464 296258
rect 134144 289258 134186 289494
rect 134422 289258 134464 289494
rect 134144 282494 134464 289258
rect 134144 282258 134186 282494
rect 134422 282258 134464 282494
rect 134144 275494 134464 282258
rect 134144 275258 134186 275494
rect 134422 275258 134464 275494
rect 134144 268494 134464 275258
rect 134144 268258 134186 268494
rect 134422 268258 134464 268494
rect 134144 261494 134464 268258
rect 134144 261258 134186 261494
rect 134422 261258 134464 261494
rect 134144 254494 134464 261258
rect 134144 254258 134186 254494
rect 134422 254258 134464 254494
rect 134144 247494 134464 254258
rect 134144 247258 134186 247494
rect 134422 247258 134464 247494
rect 134144 240494 134464 247258
rect 134144 240258 134186 240494
rect 134422 240258 134464 240494
rect 134144 233494 134464 240258
rect 134144 233258 134186 233494
rect 134422 233258 134464 233494
rect 134144 226494 134464 233258
rect 134144 226258 134186 226494
rect 134422 226258 134464 226494
rect 134144 219494 134464 226258
rect 134144 219258 134186 219494
rect 134422 219258 134464 219494
rect 134144 212494 134464 219258
rect 134144 212258 134186 212494
rect 134422 212258 134464 212494
rect 134144 205494 134464 212258
rect 134144 205258 134186 205494
rect 134422 205258 134464 205494
rect 134144 198494 134464 205258
rect 134144 198258 134186 198494
rect 134422 198258 134464 198494
rect 134144 191494 134464 198258
rect 134144 191258 134186 191494
rect 134422 191258 134464 191494
rect 134144 184494 134464 191258
rect 134144 184258 134186 184494
rect 134422 184258 134464 184494
rect 134144 177494 134464 184258
rect 134144 177258 134186 177494
rect 134422 177258 134464 177494
rect 134144 170494 134464 177258
rect 134144 170258 134186 170494
rect 134422 170258 134464 170494
rect 134144 163494 134464 170258
rect 134144 163258 134186 163494
rect 134422 163258 134464 163494
rect 134144 156494 134464 163258
rect 134144 156258 134186 156494
rect 134422 156258 134464 156494
rect 134144 149494 134464 156258
rect 134144 149258 134186 149494
rect 134422 149258 134464 149494
rect 134144 142494 134464 149258
rect 134144 142258 134186 142494
rect 134422 142258 134464 142494
rect 134144 135494 134464 142258
rect 134144 135258 134186 135494
rect 134422 135258 134464 135494
rect 134144 128494 134464 135258
rect 134144 128258 134186 128494
rect 134422 128258 134464 128494
rect 134144 121494 134464 128258
rect 134144 121258 134186 121494
rect 134422 121258 134464 121494
rect 134144 114494 134464 121258
rect 134144 114258 134186 114494
rect 134422 114258 134464 114494
rect 134144 107494 134464 114258
rect 134144 107258 134186 107494
rect 134422 107258 134464 107494
rect 134144 100494 134464 107258
rect 134144 100258 134186 100494
rect 134422 100258 134464 100494
rect 134144 93494 134464 100258
rect 134144 93258 134186 93494
rect 134422 93258 134464 93494
rect 134144 86494 134464 93258
rect 134144 86258 134186 86494
rect 134422 86258 134464 86494
rect 134144 79494 134464 86258
rect 134144 79258 134186 79494
rect 134422 79258 134464 79494
rect 134144 72494 134464 79258
rect 134144 72258 134186 72494
rect 134422 72258 134464 72494
rect 134144 65494 134464 72258
rect 134144 65258 134186 65494
rect 134422 65258 134464 65494
rect 134144 58494 134464 65258
rect 134144 58258 134186 58494
rect 134422 58258 134464 58494
rect 134144 51494 134464 58258
rect 134144 51258 134186 51494
rect 134422 51258 134464 51494
rect 134144 44494 134464 51258
rect 134144 44258 134186 44494
rect 134422 44258 134464 44494
rect 134144 37494 134464 44258
rect 134144 37258 134186 37494
rect 134422 37258 134464 37494
rect 134144 30494 134464 37258
rect 134144 30258 134186 30494
rect 134422 30258 134464 30494
rect 134144 23494 134464 30258
rect 134144 23258 134186 23494
rect 134422 23258 134464 23494
rect 134144 16494 134464 23258
rect 134144 16258 134186 16494
rect 134422 16258 134464 16494
rect 134144 9494 134464 16258
rect 134144 9258 134186 9494
rect 134422 9258 134464 9494
rect 134144 2494 134464 9258
rect 134144 2258 134186 2494
rect 134422 2258 134464 2494
rect 134144 -746 134464 2258
rect 134144 -982 134186 -746
rect 134422 -982 134464 -746
rect 134144 -1066 134464 -982
rect 134144 -1302 134186 -1066
rect 134422 -1302 134464 -1066
rect 134144 -2294 134464 -1302
rect 135876 706198 136196 706230
rect 135876 705962 135918 706198
rect 136154 705962 136196 706198
rect 135876 705878 136196 705962
rect 135876 705642 135918 705878
rect 136154 705642 136196 705878
rect 135876 696434 136196 705642
rect 135876 696198 135918 696434
rect 136154 696198 136196 696434
rect 135876 689434 136196 696198
rect 135876 689198 135918 689434
rect 136154 689198 136196 689434
rect 135876 682434 136196 689198
rect 135876 682198 135918 682434
rect 136154 682198 136196 682434
rect 135876 675434 136196 682198
rect 135876 675198 135918 675434
rect 136154 675198 136196 675434
rect 135876 668434 136196 675198
rect 135876 668198 135918 668434
rect 136154 668198 136196 668434
rect 135876 661434 136196 668198
rect 135876 661198 135918 661434
rect 136154 661198 136196 661434
rect 135876 654434 136196 661198
rect 135876 654198 135918 654434
rect 136154 654198 136196 654434
rect 135876 647434 136196 654198
rect 135876 647198 135918 647434
rect 136154 647198 136196 647434
rect 135876 640434 136196 647198
rect 135876 640198 135918 640434
rect 136154 640198 136196 640434
rect 135876 633434 136196 640198
rect 135876 633198 135918 633434
rect 136154 633198 136196 633434
rect 135876 626434 136196 633198
rect 135876 626198 135918 626434
rect 136154 626198 136196 626434
rect 135876 619434 136196 626198
rect 135876 619198 135918 619434
rect 136154 619198 136196 619434
rect 135876 612434 136196 619198
rect 135876 612198 135918 612434
rect 136154 612198 136196 612434
rect 135876 605434 136196 612198
rect 135876 605198 135918 605434
rect 136154 605198 136196 605434
rect 135876 598434 136196 605198
rect 135876 598198 135918 598434
rect 136154 598198 136196 598434
rect 135876 591434 136196 598198
rect 135876 591198 135918 591434
rect 136154 591198 136196 591434
rect 135876 584434 136196 591198
rect 135876 584198 135918 584434
rect 136154 584198 136196 584434
rect 135876 577434 136196 584198
rect 135876 577198 135918 577434
rect 136154 577198 136196 577434
rect 135876 570434 136196 577198
rect 135876 570198 135918 570434
rect 136154 570198 136196 570434
rect 135876 563434 136196 570198
rect 135876 563198 135918 563434
rect 136154 563198 136196 563434
rect 135876 556434 136196 563198
rect 135876 556198 135918 556434
rect 136154 556198 136196 556434
rect 135876 549434 136196 556198
rect 135876 549198 135918 549434
rect 136154 549198 136196 549434
rect 135876 542434 136196 549198
rect 135876 542198 135918 542434
rect 136154 542198 136196 542434
rect 135876 535434 136196 542198
rect 135876 535198 135918 535434
rect 136154 535198 136196 535434
rect 135876 528434 136196 535198
rect 135876 528198 135918 528434
rect 136154 528198 136196 528434
rect 135876 521434 136196 528198
rect 135876 521198 135918 521434
rect 136154 521198 136196 521434
rect 135876 514434 136196 521198
rect 135876 514198 135918 514434
rect 136154 514198 136196 514434
rect 135876 507434 136196 514198
rect 135876 507198 135918 507434
rect 136154 507198 136196 507434
rect 135876 500434 136196 507198
rect 135876 500198 135918 500434
rect 136154 500198 136196 500434
rect 135876 493434 136196 500198
rect 135876 493198 135918 493434
rect 136154 493198 136196 493434
rect 135876 486434 136196 493198
rect 135876 486198 135918 486434
rect 136154 486198 136196 486434
rect 135876 479434 136196 486198
rect 135876 479198 135918 479434
rect 136154 479198 136196 479434
rect 135876 472434 136196 479198
rect 135876 472198 135918 472434
rect 136154 472198 136196 472434
rect 135876 465434 136196 472198
rect 135876 465198 135918 465434
rect 136154 465198 136196 465434
rect 135876 458434 136196 465198
rect 135876 458198 135918 458434
rect 136154 458198 136196 458434
rect 135876 451434 136196 458198
rect 135876 451198 135918 451434
rect 136154 451198 136196 451434
rect 135876 444434 136196 451198
rect 135876 444198 135918 444434
rect 136154 444198 136196 444434
rect 135876 437434 136196 444198
rect 135876 437198 135918 437434
rect 136154 437198 136196 437434
rect 135876 430434 136196 437198
rect 135876 430198 135918 430434
rect 136154 430198 136196 430434
rect 135876 423434 136196 430198
rect 135876 423198 135918 423434
rect 136154 423198 136196 423434
rect 135876 416434 136196 423198
rect 135876 416198 135918 416434
rect 136154 416198 136196 416434
rect 135876 409434 136196 416198
rect 135876 409198 135918 409434
rect 136154 409198 136196 409434
rect 135876 402434 136196 409198
rect 135876 402198 135918 402434
rect 136154 402198 136196 402434
rect 135876 395434 136196 402198
rect 135876 395198 135918 395434
rect 136154 395198 136196 395434
rect 135876 388434 136196 395198
rect 135876 388198 135918 388434
rect 136154 388198 136196 388434
rect 135876 381434 136196 388198
rect 135876 381198 135918 381434
rect 136154 381198 136196 381434
rect 135876 374434 136196 381198
rect 135876 374198 135918 374434
rect 136154 374198 136196 374434
rect 135876 367434 136196 374198
rect 135876 367198 135918 367434
rect 136154 367198 136196 367434
rect 135876 360434 136196 367198
rect 135876 360198 135918 360434
rect 136154 360198 136196 360434
rect 135876 353434 136196 360198
rect 135876 353198 135918 353434
rect 136154 353198 136196 353434
rect 135876 346434 136196 353198
rect 135876 346198 135918 346434
rect 136154 346198 136196 346434
rect 135876 339434 136196 346198
rect 135876 339198 135918 339434
rect 136154 339198 136196 339434
rect 135876 332434 136196 339198
rect 135876 332198 135918 332434
rect 136154 332198 136196 332434
rect 135876 325434 136196 332198
rect 135876 325198 135918 325434
rect 136154 325198 136196 325434
rect 135876 318434 136196 325198
rect 135876 318198 135918 318434
rect 136154 318198 136196 318434
rect 135876 311434 136196 318198
rect 135876 311198 135918 311434
rect 136154 311198 136196 311434
rect 135876 304434 136196 311198
rect 135876 304198 135918 304434
rect 136154 304198 136196 304434
rect 135876 297434 136196 304198
rect 135876 297198 135918 297434
rect 136154 297198 136196 297434
rect 135876 290434 136196 297198
rect 135876 290198 135918 290434
rect 136154 290198 136196 290434
rect 135876 283434 136196 290198
rect 135876 283198 135918 283434
rect 136154 283198 136196 283434
rect 135876 276434 136196 283198
rect 135876 276198 135918 276434
rect 136154 276198 136196 276434
rect 135876 269434 136196 276198
rect 135876 269198 135918 269434
rect 136154 269198 136196 269434
rect 135876 262434 136196 269198
rect 135876 262198 135918 262434
rect 136154 262198 136196 262434
rect 135876 255434 136196 262198
rect 135876 255198 135918 255434
rect 136154 255198 136196 255434
rect 135876 248434 136196 255198
rect 135876 248198 135918 248434
rect 136154 248198 136196 248434
rect 135876 241434 136196 248198
rect 135876 241198 135918 241434
rect 136154 241198 136196 241434
rect 135876 234434 136196 241198
rect 135876 234198 135918 234434
rect 136154 234198 136196 234434
rect 135876 227434 136196 234198
rect 135876 227198 135918 227434
rect 136154 227198 136196 227434
rect 135876 220434 136196 227198
rect 135876 220198 135918 220434
rect 136154 220198 136196 220434
rect 135876 213434 136196 220198
rect 135876 213198 135918 213434
rect 136154 213198 136196 213434
rect 135876 206434 136196 213198
rect 135876 206198 135918 206434
rect 136154 206198 136196 206434
rect 135876 199434 136196 206198
rect 135876 199198 135918 199434
rect 136154 199198 136196 199434
rect 135876 192434 136196 199198
rect 135876 192198 135918 192434
rect 136154 192198 136196 192434
rect 135876 185434 136196 192198
rect 135876 185198 135918 185434
rect 136154 185198 136196 185434
rect 135876 178434 136196 185198
rect 135876 178198 135918 178434
rect 136154 178198 136196 178434
rect 135876 171434 136196 178198
rect 135876 171198 135918 171434
rect 136154 171198 136196 171434
rect 135876 164434 136196 171198
rect 135876 164198 135918 164434
rect 136154 164198 136196 164434
rect 135876 157434 136196 164198
rect 135876 157198 135918 157434
rect 136154 157198 136196 157434
rect 135876 150434 136196 157198
rect 135876 150198 135918 150434
rect 136154 150198 136196 150434
rect 135876 143434 136196 150198
rect 135876 143198 135918 143434
rect 136154 143198 136196 143434
rect 135876 136434 136196 143198
rect 135876 136198 135918 136434
rect 136154 136198 136196 136434
rect 135876 129434 136196 136198
rect 135876 129198 135918 129434
rect 136154 129198 136196 129434
rect 135876 122434 136196 129198
rect 135876 122198 135918 122434
rect 136154 122198 136196 122434
rect 135876 115434 136196 122198
rect 135876 115198 135918 115434
rect 136154 115198 136196 115434
rect 135876 108434 136196 115198
rect 135876 108198 135918 108434
rect 136154 108198 136196 108434
rect 135876 101434 136196 108198
rect 135876 101198 135918 101434
rect 136154 101198 136196 101434
rect 135876 94434 136196 101198
rect 135876 94198 135918 94434
rect 136154 94198 136196 94434
rect 135876 87434 136196 94198
rect 135876 87198 135918 87434
rect 136154 87198 136196 87434
rect 135876 80434 136196 87198
rect 135876 80198 135918 80434
rect 136154 80198 136196 80434
rect 135876 73434 136196 80198
rect 135876 73198 135918 73434
rect 136154 73198 136196 73434
rect 135876 66434 136196 73198
rect 135876 66198 135918 66434
rect 136154 66198 136196 66434
rect 135876 59434 136196 66198
rect 135876 59198 135918 59434
rect 136154 59198 136196 59434
rect 135876 52434 136196 59198
rect 135876 52198 135918 52434
rect 136154 52198 136196 52434
rect 135876 45434 136196 52198
rect 135876 45198 135918 45434
rect 136154 45198 136196 45434
rect 135876 38434 136196 45198
rect 135876 38198 135918 38434
rect 136154 38198 136196 38434
rect 135876 31434 136196 38198
rect 135876 31198 135918 31434
rect 136154 31198 136196 31434
rect 135876 24434 136196 31198
rect 135876 24198 135918 24434
rect 136154 24198 136196 24434
rect 135876 17434 136196 24198
rect 135876 17198 135918 17434
rect 136154 17198 136196 17434
rect 135876 10434 136196 17198
rect 135876 10198 135918 10434
rect 136154 10198 136196 10434
rect 135876 3434 136196 10198
rect 135876 3198 135918 3434
rect 136154 3198 136196 3434
rect 135876 -1706 136196 3198
rect 135876 -1942 135918 -1706
rect 136154 -1942 136196 -1706
rect 135876 -2026 136196 -1942
rect 135876 -2262 135918 -2026
rect 136154 -2262 136196 -2026
rect 135876 -2294 136196 -2262
rect 141144 705238 141464 706230
rect 141144 705002 141186 705238
rect 141422 705002 141464 705238
rect 141144 704918 141464 705002
rect 141144 704682 141186 704918
rect 141422 704682 141464 704918
rect 141144 695494 141464 704682
rect 141144 695258 141186 695494
rect 141422 695258 141464 695494
rect 141144 688494 141464 695258
rect 141144 688258 141186 688494
rect 141422 688258 141464 688494
rect 141144 681494 141464 688258
rect 141144 681258 141186 681494
rect 141422 681258 141464 681494
rect 141144 674494 141464 681258
rect 141144 674258 141186 674494
rect 141422 674258 141464 674494
rect 141144 667494 141464 674258
rect 141144 667258 141186 667494
rect 141422 667258 141464 667494
rect 141144 660494 141464 667258
rect 141144 660258 141186 660494
rect 141422 660258 141464 660494
rect 141144 653494 141464 660258
rect 141144 653258 141186 653494
rect 141422 653258 141464 653494
rect 141144 646494 141464 653258
rect 141144 646258 141186 646494
rect 141422 646258 141464 646494
rect 141144 639494 141464 646258
rect 141144 639258 141186 639494
rect 141422 639258 141464 639494
rect 141144 632494 141464 639258
rect 141144 632258 141186 632494
rect 141422 632258 141464 632494
rect 141144 625494 141464 632258
rect 141144 625258 141186 625494
rect 141422 625258 141464 625494
rect 141144 618494 141464 625258
rect 141144 618258 141186 618494
rect 141422 618258 141464 618494
rect 141144 611494 141464 618258
rect 141144 611258 141186 611494
rect 141422 611258 141464 611494
rect 141144 604494 141464 611258
rect 141144 604258 141186 604494
rect 141422 604258 141464 604494
rect 141144 597494 141464 604258
rect 141144 597258 141186 597494
rect 141422 597258 141464 597494
rect 141144 590494 141464 597258
rect 141144 590258 141186 590494
rect 141422 590258 141464 590494
rect 141144 583494 141464 590258
rect 141144 583258 141186 583494
rect 141422 583258 141464 583494
rect 141144 576494 141464 583258
rect 141144 576258 141186 576494
rect 141422 576258 141464 576494
rect 141144 569494 141464 576258
rect 141144 569258 141186 569494
rect 141422 569258 141464 569494
rect 141144 562494 141464 569258
rect 141144 562258 141186 562494
rect 141422 562258 141464 562494
rect 141144 555494 141464 562258
rect 141144 555258 141186 555494
rect 141422 555258 141464 555494
rect 141144 548494 141464 555258
rect 141144 548258 141186 548494
rect 141422 548258 141464 548494
rect 141144 541494 141464 548258
rect 141144 541258 141186 541494
rect 141422 541258 141464 541494
rect 141144 534494 141464 541258
rect 141144 534258 141186 534494
rect 141422 534258 141464 534494
rect 141144 527494 141464 534258
rect 141144 527258 141186 527494
rect 141422 527258 141464 527494
rect 141144 520494 141464 527258
rect 141144 520258 141186 520494
rect 141422 520258 141464 520494
rect 141144 513494 141464 520258
rect 141144 513258 141186 513494
rect 141422 513258 141464 513494
rect 141144 506494 141464 513258
rect 141144 506258 141186 506494
rect 141422 506258 141464 506494
rect 141144 499494 141464 506258
rect 141144 499258 141186 499494
rect 141422 499258 141464 499494
rect 141144 492494 141464 499258
rect 141144 492258 141186 492494
rect 141422 492258 141464 492494
rect 141144 485494 141464 492258
rect 141144 485258 141186 485494
rect 141422 485258 141464 485494
rect 141144 478494 141464 485258
rect 141144 478258 141186 478494
rect 141422 478258 141464 478494
rect 141144 471494 141464 478258
rect 141144 471258 141186 471494
rect 141422 471258 141464 471494
rect 141144 464494 141464 471258
rect 141144 464258 141186 464494
rect 141422 464258 141464 464494
rect 141144 457494 141464 464258
rect 141144 457258 141186 457494
rect 141422 457258 141464 457494
rect 141144 450494 141464 457258
rect 141144 450258 141186 450494
rect 141422 450258 141464 450494
rect 141144 443494 141464 450258
rect 141144 443258 141186 443494
rect 141422 443258 141464 443494
rect 141144 436494 141464 443258
rect 141144 436258 141186 436494
rect 141422 436258 141464 436494
rect 141144 429494 141464 436258
rect 141144 429258 141186 429494
rect 141422 429258 141464 429494
rect 141144 422494 141464 429258
rect 141144 422258 141186 422494
rect 141422 422258 141464 422494
rect 141144 415494 141464 422258
rect 141144 415258 141186 415494
rect 141422 415258 141464 415494
rect 141144 408494 141464 415258
rect 141144 408258 141186 408494
rect 141422 408258 141464 408494
rect 141144 401494 141464 408258
rect 141144 401258 141186 401494
rect 141422 401258 141464 401494
rect 141144 394494 141464 401258
rect 141144 394258 141186 394494
rect 141422 394258 141464 394494
rect 141144 387494 141464 394258
rect 141144 387258 141186 387494
rect 141422 387258 141464 387494
rect 141144 380494 141464 387258
rect 141144 380258 141186 380494
rect 141422 380258 141464 380494
rect 141144 373494 141464 380258
rect 141144 373258 141186 373494
rect 141422 373258 141464 373494
rect 141144 366494 141464 373258
rect 141144 366258 141186 366494
rect 141422 366258 141464 366494
rect 141144 359494 141464 366258
rect 141144 359258 141186 359494
rect 141422 359258 141464 359494
rect 141144 352494 141464 359258
rect 141144 352258 141186 352494
rect 141422 352258 141464 352494
rect 141144 345494 141464 352258
rect 141144 345258 141186 345494
rect 141422 345258 141464 345494
rect 141144 338494 141464 345258
rect 141144 338258 141186 338494
rect 141422 338258 141464 338494
rect 141144 331494 141464 338258
rect 141144 331258 141186 331494
rect 141422 331258 141464 331494
rect 141144 324494 141464 331258
rect 141144 324258 141186 324494
rect 141422 324258 141464 324494
rect 141144 317494 141464 324258
rect 141144 317258 141186 317494
rect 141422 317258 141464 317494
rect 141144 310494 141464 317258
rect 141144 310258 141186 310494
rect 141422 310258 141464 310494
rect 141144 303494 141464 310258
rect 141144 303258 141186 303494
rect 141422 303258 141464 303494
rect 141144 296494 141464 303258
rect 141144 296258 141186 296494
rect 141422 296258 141464 296494
rect 141144 289494 141464 296258
rect 141144 289258 141186 289494
rect 141422 289258 141464 289494
rect 141144 282494 141464 289258
rect 141144 282258 141186 282494
rect 141422 282258 141464 282494
rect 141144 275494 141464 282258
rect 141144 275258 141186 275494
rect 141422 275258 141464 275494
rect 141144 268494 141464 275258
rect 141144 268258 141186 268494
rect 141422 268258 141464 268494
rect 141144 261494 141464 268258
rect 141144 261258 141186 261494
rect 141422 261258 141464 261494
rect 141144 254494 141464 261258
rect 141144 254258 141186 254494
rect 141422 254258 141464 254494
rect 141144 247494 141464 254258
rect 141144 247258 141186 247494
rect 141422 247258 141464 247494
rect 141144 240494 141464 247258
rect 141144 240258 141186 240494
rect 141422 240258 141464 240494
rect 141144 233494 141464 240258
rect 141144 233258 141186 233494
rect 141422 233258 141464 233494
rect 141144 226494 141464 233258
rect 141144 226258 141186 226494
rect 141422 226258 141464 226494
rect 141144 219494 141464 226258
rect 141144 219258 141186 219494
rect 141422 219258 141464 219494
rect 141144 212494 141464 219258
rect 141144 212258 141186 212494
rect 141422 212258 141464 212494
rect 141144 205494 141464 212258
rect 141144 205258 141186 205494
rect 141422 205258 141464 205494
rect 141144 198494 141464 205258
rect 141144 198258 141186 198494
rect 141422 198258 141464 198494
rect 141144 191494 141464 198258
rect 141144 191258 141186 191494
rect 141422 191258 141464 191494
rect 141144 184494 141464 191258
rect 141144 184258 141186 184494
rect 141422 184258 141464 184494
rect 141144 177494 141464 184258
rect 141144 177258 141186 177494
rect 141422 177258 141464 177494
rect 141144 170494 141464 177258
rect 141144 170258 141186 170494
rect 141422 170258 141464 170494
rect 141144 163494 141464 170258
rect 141144 163258 141186 163494
rect 141422 163258 141464 163494
rect 141144 156494 141464 163258
rect 141144 156258 141186 156494
rect 141422 156258 141464 156494
rect 141144 149494 141464 156258
rect 141144 149258 141186 149494
rect 141422 149258 141464 149494
rect 141144 142494 141464 149258
rect 141144 142258 141186 142494
rect 141422 142258 141464 142494
rect 141144 135494 141464 142258
rect 141144 135258 141186 135494
rect 141422 135258 141464 135494
rect 141144 128494 141464 135258
rect 141144 128258 141186 128494
rect 141422 128258 141464 128494
rect 141144 121494 141464 128258
rect 141144 121258 141186 121494
rect 141422 121258 141464 121494
rect 141144 114494 141464 121258
rect 141144 114258 141186 114494
rect 141422 114258 141464 114494
rect 141144 107494 141464 114258
rect 141144 107258 141186 107494
rect 141422 107258 141464 107494
rect 141144 100494 141464 107258
rect 141144 100258 141186 100494
rect 141422 100258 141464 100494
rect 141144 93494 141464 100258
rect 141144 93258 141186 93494
rect 141422 93258 141464 93494
rect 141144 86494 141464 93258
rect 141144 86258 141186 86494
rect 141422 86258 141464 86494
rect 141144 79494 141464 86258
rect 141144 79258 141186 79494
rect 141422 79258 141464 79494
rect 141144 72494 141464 79258
rect 141144 72258 141186 72494
rect 141422 72258 141464 72494
rect 141144 65494 141464 72258
rect 141144 65258 141186 65494
rect 141422 65258 141464 65494
rect 141144 58494 141464 65258
rect 141144 58258 141186 58494
rect 141422 58258 141464 58494
rect 141144 51494 141464 58258
rect 141144 51258 141186 51494
rect 141422 51258 141464 51494
rect 141144 44494 141464 51258
rect 141144 44258 141186 44494
rect 141422 44258 141464 44494
rect 141144 37494 141464 44258
rect 141144 37258 141186 37494
rect 141422 37258 141464 37494
rect 141144 30494 141464 37258
rect 141144 30258 141186 30494
rect 141422 30258 141464 30494
rect 141144 23494 141464 30258
rect 141144 23258 141186 23494
rect 141422 23258 141464 23494
rect 141144 16494 141464 23258
rect 141144 16258 141186 16494
rect 141422 16258 141464 16494
rect 141144 9494 141464 16258
rect 141144 9258 141186 9494
rect 141422 9258 141464 9494
rect 141144 2494 141464 9258
rect 141144 2258 141186 2494
rect 141422 2258 141464 2494
rect 141144 -746 141464 2258
rect 141144 -982 141186 -746
rect 141422 -982 141464 -746
rect 141144 -1066 141464 -982
rect 141144 -1302 141186 -1066
rect 141422 -1302 141464 -1066
rect 141144 -2294 141464 -1302
rect 142876 706198 143196 706230
rect 142876 705962 142918 706198
rect 143154 705962 143196 706198
rect 142876 705878 143196 705962
rect 142876 705642 142918 705878
rect 143154 705642 143196 705878
rect 142876 696434 143196 705642
rect 142876 696198 142918 696434
rect 143154 696198 143196 696434
rect 142876 689434 143196 696198
rect 142876 689198 142918 689434
rect 143154 689198 143196 689434
rect 142876 682434 143196 689198
rect 142876 682198 142918 682434
rect 143154 682198 143196 682434
rect 142876 675434 143196 682198
rect 142876 675198 142918 675434
rect 143154 675198 143196 675434
rect 142876 668434 143196 675198
rect 142876 668198 142918 668434
rect 143154 668198 143196 668434
rect 142876 661434 143196 668198
rect 142876 661198 142918 661434
rect 143154 661198 143196 661434
rect 142876 654434 143196 661198
rect 142876 654198 142918 654434
rect 143154 654198 143196 654434
rect 142876 647434 143196 654198
rect 142876 647198 142918 647434
rect 143154 647198 143196 647434
rect 142876 640434 143196 647198
rect 142876 640198 142918 640434
rect 143154 640198 143196 640434
rect 142876 633434 143196 640198
rect 142876 633198 142918 633434
rect 143154 633198 143196 633434
rect 142876 626434 143196 633198
rect 142876 626198 142918 626434
rect 143154 626198 143196 626434
rect 142876 619434 143196 626198
rect 142876 619198 142918 619434
rect 143154 619198 143196 619434
rect 142876 612434 143196 619198
rect 142876 612198 142918 612434
rect 143154 612198 143196 612434
rect 142876 605434 143196 612198
rect 142876 605198 142918 605434
rect 143154 605198 143196 605434
rect 142876 598434 143196 605198
rect 142876 598198 142918 598434
rect 143154 598198 143196 598434
rect 142876 591434 143196 598198
rect 142876 591198 142918 591434
rect 143154 591198 143196 591434
rect 142876 584434 143196 591198
rect 142876 584198 142918 584434
rect 143154 584198 143196 584434
rect 142876 577434 143196 584198
rect 142876 577198 142918 577434
rect 143154 577198 143196 577434
rect 142876 570434 143196 577198
rect 142876 570198 142918 570434
rect 143154 570198 143196 570434
rect 142876 563434 143196 570198
rect 142876 563198 142918 563434
rect 143154 563198 143196 563434
rect 142876 556434 143196 563198
rect 142876 556198 142918 556434
rect 143154 556198 143196 556434
rect 142876 549434 143196 556198
rect 142876 549198 142918 549434
rect 143154 549198 143196 549434
rect 142876 542434 143196 549198
rect 142876 542198 142918 542434
rect 143154 542198 143196 542434
rect 142876 535434 143196 542198
rect 142876 535198 142918 535434
rect 143154 535198 143196 535434
rect 142876 528434 143196 535198
rect 142876 528198 142918 528434
rect 143154 528198 143196 528434
rect 142876 521434 143196 528198
rect 142876 521198 142918 521434
rect 143154 521198 143196 521434
rect 142876 514434 143196 521198
rect 142876 514198 142918 514434
rect 143154 514198 143196 514434
rect 142876 507434 143196 514198
rect 142876 507198 142918 507434
rect 143154 507198 143196 507434
rect 142876 500434 143196 507198
rect 142876 500198 142918 500434
rect 143154 500198 143196 500434
rect 142876 493434 143196 500198
rect 142876 493198 142918 493434
rect 143154 493198 143196 493434
rect 142876 486434 143196 493198
rect 142876 486198 142918 486434
rect 143154 486198 143196 486434
rect 142876 479434 143196 486198
rect 142876 479198 142918 479434
rect 143154 479198 143196 479434
rect 142876 472434 143196 479198
rect 142876 472198 142918 472434
rect 143154 472198 143196 472434
rect 142876 465434 143196 472198
rect 142876 465198 142918 465434
rect 143154 465198 143196 465434
rect 142876 458434 143196 465198
rect 142876 458198 142918 458434
rect 143154 458198 143196 458434
rect 142876 451434 143196 458198
rect 142876 451198 142918 451434
rect 143154 451198 143196 451434
rect 142876 444434 143196 451198
rect 142876 444198 142918 444434
rect 143154 444198 143196 444434
rect 142876 437434 143196 444198
rect 142876 437198 142918 437434
rect 143154 437198 143196 437434
rect 142876 430434 143196 437198
rect 142876 430198 142918 430434
rect 143154 430198 143196 430434
rect 142876 423434 143196 430198
rect 142876 423198 142918 423434
rect 143154 423198 143196 423434
rect 142876 416434 143196 423198
rect 142876 416198 142918 416434
rect 143154 416198 143196 416434
rect 142876 409434 143196 416198
rect 142876 409198 142918 409434
rect 143154 409198 143196 409434
rect 142876 402434 143196 409198
rect 142876 402198 142918 402434
rect 143154 402198 143196 402434
rect 142876 395434 143196 402198
rect 142876 395198 142918 395434
rect 143154 395198 143196 395434
rect 142876 388434 143196 395198
rect 142876 388198 142918 388434
rect 143154 388198 143196 388434
rect 142876 381434 143196 388198
rect 142876 381198 142918 381434
rect 143154 381198 143196 381434
rect 142876 374434 143196 381198
rect 142876 374198 142918 374434
rect 143154 374198 143196 374434
rect 142876 367434 143196 374198
rect 142876 367198 142918 367434
rect 143154 367198 143196 367434
rect 142876 360434 143196 367198
rect 142876 360198 142918 360434
rect 143154 360198 143196 360434
rect 142876 353434 143196 360198
rect 142876 353198 142918 353434
rect 143154 353198 143196 353434
rect 142876 346434 143196 353198
rect 142876 346198 142918 346434
rect 143154 346198 143196 346434
rect 142876 339434 143196 346198
rect 142876 339198 142918 339434
rect 143154 339198 143196 339434
rect 142876 332434 143196 339198
rect 142876 332198 142918 332434
rect 143154 332198 143196 332434
rect 142876 325434 143196 332198
rect 142876 325198 142918 325434
rect 143154 325198 143196 325434
rect 142876 318434 143196 325198
rect 142876 318198 142918 318434
rect 143154 318198 143196 318434
rect 142876 311434 143196 318198
rect 142876 311198 142918 311434
rect 143154 311198 143196 311434
rect 142876 304434 143196 311198
rect 142876 304198 142918 304434
rect 143154 304198 143196 304434
rect 142876 297434 143196 304198
rect 142876 297198 142918 297434
rect 143154 297198 143196 297434
rect 142876 290434 143196 297198
rect 142876 290198 142918 290434
rect 143154 290198 143196 290434
rect 142876 283434 143196 290198
rect 142876 283198 142918 283434
rect 143154 283198 143196 283434
rect 142876 276434 143196 283198
rect 142876 276198 142918 276434
rect 143154 276198 143196 276434
rect 142876 269434 143196 276198
rect 142876 269198 142918 269434
rect 143154 269198 143196 269434
rect 142876 262434 143196 269198
rect 142876 262198 142918 262434
rect 143154 262198 143196 262434
rect 142876 255434 143196 262198
rect 142876 255198 142918 255434
rect 143154 255198 143196 255434
rect 142876 248434 143196 255198
rect 142876 248198 142918 248434
rect 143154 248198 143196 248434
rect 142876 241434 143196 248198
rect 142876 241198 142918 241434
rect 143154 241198 143196 241434
rect 142876 234434 143196 241198
rect 142876 234198 142918 234434
rect 143154 234198 143196 234434
rect 142876 227434 143196 234198
rect 142876 227198 142918 227434
rect 143154 227198 143196 227434
rect 142876 220434 143196 227198
rect 142876 220198 142918 220434
rect 143154 220198 143196 220434
rect 142876 213434 143196 220198
rect 142876 213198 142918 213434
rect 143154 213198 143196 213434
rect 142876 206434 143196 213198
rect 142876 206198 142918 206434
rect 143154 206198 143196 206434
rect 142876 199434 143196 206198
rect 142876 199198 142918 199434
rect 143154 199198 143196 199434
rect 142876 192434 143196 199198
rect 142876 192198 142918 192434
rect 143154 192198 143196 192434
rect 142876 185434 143196 192198
rect 142876 185198 142918 185434
rect 143154 185198 143196 185434
rect 142876 178434 143196 185198
rect 142876 178198 142918 178434
rect 143154 178198 143196 178434
rect 142876 171434 143196 178198
rect 142876 171198 142918 171434
rect 143154 171198 143196 171434
rect 142876 164434 143196 171198
rect 142876 164198 142918 164434
rect 143154 164198 143196 164434
rect 142876 157434 143196 164198
rect 142876 157198 142918 157434
rect 143154 157198 143196 157434
rect 142876 150434 143196 157198
rect 142876 150198 142918 150434
rect 143154 150198 143196 150434
rect 142876 143434 143196 150198
rect 142876 143198 142918 143434
rect 143154 143198 143196 143434
rect 142876 136434 143196 143198
rect 142876 136198 142918 136434
rect 143154 136198 143196 136434
rect 142876 129434 143196 136198
rect 142876 129198 142918 129434
rect 143154 129198 143196 129434
rect 142876 122434 143196 129198
rect 142876 122198 142918 122434
rect 143154 122198 143196 122434
rect 142876 115434 143196 122198
rect 142876 115198 142918 115434
rect 143154 115198 143196 115434
rect 142876 108434 143196 115198
rect 142876 108198 142918 108434
rect 143154 108198 143196 108434
rect 142876 101434 143196 108198
rect 142876 101198 142918 101434
rect 143154 101198 143196 101434
rect 142876 94434 143196 101198
rect 142876 94198 142918 94434
rect 143154 94198 143196 94434
rect 142876 87434 143196 94198
rect 142876 87198 142918 87434
rect 143154 87198 143196 87434
rect 142876 80434 143196 87198
rect 142876 80198 142918 80434
rect 143154 80198 143196 80434
rect 142876 73434 143196 80198
rect 142876 73198 142918 73434
rect 143154 73198 143196 73434
rect 142876 66434 143196 73198
rect 142876 66198 142918 66434
rect 143154 66198 143196 66434
rect 142876 59434 143196 66198
rect 142876 59198 142918 59434
rect 143154 59198 143196 59434
rect 142876 52434 143196 59198
rect 142876 52198 142918 52434
rect 143154 52198 143196 52434
rect 142876 45434 143196 52198
rect 142876 45198 142918 45434
rect 143154 45198 143196 45434
rect 142876 38434 143196 45198
rect 142876 38198 142918 38434
rect 143154 38198 143196 38434
rect 142876 31434 143196 38198
rect 142876 31198 142918 31434
rect 143154 31198 143196 31434
rect 142876 24434 143196 31198
rect 142876 24198 142918 24434
rect 143154 24198 143196 24434
rect 142876 17434 143196 24198
rect 142876 17198 142918 17434
rect 143154 17198 143196 17434
rect 142876 10434 143196 17198
rect 142876 10198 142918 10434
rect 143154 10198 143196 10434
rect 142876 3434 143196 10198
rect 142876 3198 142918 3434
rect 143154 3198 143196 3434
rect 142876 -1706 143196 3198
rect 142876 -1942 142918 -1706
rect 143154 -1942 143196 -1706
rect 142876 -2026 143196 -1942
rect 142876 -2262 142918 -2026
rect 143154 -2262 143196 -2026
rect 142876 -2294 143196 -2262
rect 148144 705238 148464 706230
rect 148144 705002 148186 705238
rect 148422 705002 148464 705238
rect 148144 704918 148464 705002
rect 148144 704682 148186 704918
rect 148422 704682 148464 704918
rect 148144 695494 148464 704682
rect 148144 695258 148186 695494
rect 148422 695258 148464 695494
rect 148144 688494 148464 695258
rect 148144 688258 148186 688494
rect 148422 688258 148464 688494
rect 148144 681494 148464 688258
rect 148144 681258 148186 681494
rect 148422 681258 148464 681494
rect 148144 674494 148464 681258
rect 148144 674258 148186 674494
rect 148422 674258 148464 674494
rect 148144 667494 148464 674258
rect 148144 667258 148186 667494
rect 148422 667258 148464 667494
rect 148144 660494 148464 667258
rect 148144 660258 148186 660494
rect 148422 660258 148464 660494
rect 148144 653494 148464 660258
rect 148144 653258 148186 653494
rect 148422 653258 148464 653494
rect 148144 646494 148464 653258
rect 148144 646258 148186 646494
rect 148422 646258 148464 646494
rect 148144 639494 148464 646258
rect 148144 639258 148186 639494
rect 148422 639258 148464 639494
rect 148144 632494 148464 639258
rect 148144 632258 148186 632494
rect 148422 632258 148464 632494
rect 148144 625494 148464 632258
rect 148144 625258 148186 625494
rect 148422 625258 148464 625494
rect 148144 618494 148464 625258
rect 148144 618258 148186 618494
rect 148422 618258 148464 618494
rect 148144 611494 148464 618258
rect 148144 611258 148186 611494
rect 148422 611258 148464 611494
rect 148144 604494 148464 611258
rect 148144 604258 148186 604494
rect 148422 604258 148464 604494
rect 148144 597494 148464 604258
rect 148144 597258 148186 597494
rect 148422 597258 148464 597494
rect 148144 590494 148464 597258
rect 148144 590258 148186 590494
rect 148422 590258 148464 590494
rect 148144 583494 148464 590258
rect 148144 583258 148186 583494
rect 148422 583258 148464 583494
rect 148144 576494 148464 583258
rect 148144 576258 148186 576494
rect 148422 576258 148464 576494
rect 148144 569494 148464 576258
rect 148144 569258 148186 569494
rect 148422 569258 148464 569494
rect 148144 562494 148464 569258
rect 148144 562258 148186 562494
rect 148422 562258 148464 562494
rect 148144 555494 148464 562258
rect 148144 555258 148186 555494
rect 148422 555258 148464 555494
rect 148144 548494 148464 555258
rect 148144 548258 148186 548494
rect 148422 548258 148464 548494
rect 148144 541494 148464 548258
rect 148144 541258 148186 541494
rect 148422 541258 148464 541494
rect 148144 534494 148464 541258
rect 148144 534258 148186 534494
rect 148422 534258 148464 534494
rect 148144 527494 148464 534258
rect 148144 527258 148186 527494
rect 148422 527258 148464 527494
rect 148144 520494 148464 527258
rect 148144 520258 148186 520494
rect 148422 520258 148464 520494
rect 148144 513494 148464 520258
rect 148144 513258 148186 513494
rect 148422 513258 148464 513494
rect 148144 506494 148464 513258
rect 148144 506258 148186 506494
rect 148422 506258 148464 506494
rect 148144 499494 148464 506258
rect 148144 499258 148186 499494
rect 148422 499258 148464 499494
rect 148144 492494 148464 499258
rect 148144 492258 148186 492494
rect 148422 492258 148464 492494
rect 148144 485494 148464 492258
rect 148144 485258 148186 485494
rect 148422 485258 148464 485494
rect 148144 478494 148464 485258
rect 148144 478258 148186 478494
rect 148422 478258 148464 478494
rect 148144 471494 148464 478258
rect 148144 471258 148186 471494
rect 148422 471258 148464 471494
rect 148144 464494 148464 471258
rect 148144 464258 148186 464494
rect 148422 464258 148464 464494
rect 148144 457494 148464 464258
rect 148144 457258 148186 457494
rect 148422 457258 148464 457494
rect 148144 450494 148464 457258
rect 148144 450258 148186 450494
rect 148422 450258 148464 450494
rect 148144 443494 148464 450258
rect 148144 443258 148186 443494
rect 148422 443258 148464 443494
rect 148144 436494 148464 443258
rect 148144 436258 148186 436494
rect 148422 436258 148464 436494
rect 148144 429494 148464 436258
rect 148144 429258 148186 429494
rect 148422 429258 148464 429494
rect 148144 422494 148464 429258
rect 148144 422258 148186 422494
rect 148422 422258 148464 422494
rect 148144 415494 148464 422258
rect 148144 415258 148186 415494
rect 148422 415258 148464 415494
rect 148144 408494 148464 415258
rect 148144 408258 148186 408494
rect 148422 408258 148464 408494
rect 148144 401494 148464 408258
rect 148144 401258 148186 401494
rect 148422 401258 148464 401494
rect 148144 394494 148464 401258
rect 148144 394258 148186 394494
rect 148422 394258 148464 394494
rect 148144 387494 148464 394258
rect 148144 387258 148186 387494
rect 148422 387258 148464 387494
rect 148144 380494 148464 387258
rect 148144 380258 148186 380494
rect 148422 380258 148464 380494
rect 148144 373494 148464 380258
rect 148144 373258 148186 373494
rect 148422 373258 148464 373494
rect 148144 366494 148464 373258
rect 148144 366258 148186 366494
rect 148422 366258 148464 366494
rect 148144 359494 148464 366258
rect 148144 359258 148186 359494
rect 148422 359258 148464 359494
rect 148144 352494 148464 359258
rect 148144 352258 148186 352494
rect 148422 352258 148464 352494
rect 148144 345494 148464 352258
rect 148144 345258 148186 345494
rect 148422 345258 148464 345494
rect 148144 338494 148464 345258
rect 148144 338258 148186 338494
rect 148422 338258 148464 338494
rect 148144 331494 148464 338258
rect 148144 331258 148186 331494
rect 148422 331258 148464 331494
rect 148144 324494 148464 331258
rect 148144 324258 148186 324494
rect 148422 324258 148464 324494
rect 148144 317494 148464 324258
rect 148144 317258 148186 317494
rect 148422 317258 148464 317494
rect 148144 310494 148464 317258
rect 148144 310258 148186 310494
rect 148422 310258 148464 310494
rect 148144 303494 148464 310258
rect 148144 303258 148186 303494
rect 148422 303258 148464 303494
rect 148144 296494 148464 303258
rect 148144 296258 148186 296494
rect 148422 296258 148464 296494
rect 148144 289494 148464 296258
rect 148144 289258 148186 289494
rect 148422 289258 148464 289494
rect 148144 282494 148464 289258
rect 148144 282258 148186 282494
rect 148422 282258 148464 282494
rect 148144 275494 148464 282258
rect 148144 275258 148186 275494
rect 148422 275258 148464 275494
rect 148144 268494 148464 275258
rect 148144 268258 148186 268494
rect 148422 268258 148464 268494
rect 148144 261494 148464 268258
rect 148144 261258 148186 261494
rect 148422 261258 148464 261494
rect 148144 254494 148464 261258
rect 148144 254258 148186 254494
rect 148422 254258 148464 254494
rect 148144 247494 148464 254258
rect 148144 247258 148186 247494
rect 148422 247258 148464 247494
rect 148144 240494 148464 247258
rect 148144 240258 148186 240494
rect 148422 240258 148464 240494
rect 148144 233494 148464 240258
rect 148144 233258 148186 233494
rect 148422 233258 148464 233494
rect 148144 226494 148464 233258
rect 148144 226258 148186 226494
rect 148422 226258 148464 226494
rect 148144 219494 148464 226258
rect 148144 219258 148186 219494
rect 148422 219258 148464 219494
rect 148144 212494 148464 219258
rect 148144 212258 148186 212494
rect 148422 212258 148464 212494
rect 148144 205494 148464 212258
rect 148144 205258 148186 205494
rect 148422 205258 148464 205494
rect 148144 198494 148464 205258
rect 148144 198258 148186 198494
rect 148422 198258 148464 198494
rect 148144 191494 148464 198258
rect 148144 191258 148186 191494
rect 148422 191258 148464 191494
rect 148144 184494 148464 191258
rect 148144 184258 148186 184494
rect 148422 184258 148464 184494
rect 148144 177494 148464 184258
rect 148144 177258 148186 177494
rect 148422 177258 148464 177494
rect 148144 170494 148464 177258
rect 148144 170258 148186 170494
rect 148422 170258 148464 170494
rect 148144 163494 148464 170258
rect 148144 163258 148186 163494
rect 148422 163258 148464 163494
rect 148144 156494 148464 163258
rect 148144 156258 148186 156494
rect 148422 156258 148464 156494
rect 148144 149494 148464 156258
rect 148144 149258 148186 149494
rect 148422 149258 148464 149494
rect 148144 142494 148464 149258
rect 148144 142258 148186 142494
rect 148422 142258 148464 142494
rect 148144 135494 148464 142258
rect 148144 135258 148186 135494
rect 148422 135258 148464 135494
rect 148144 128494 148464 135258
rect 148144 128258 148186 128494
rect 148422 128258 148464 128494
rect 148144 121494 148464 128258
rect 148144 121258 148186 121494
rect 148422 121258 148464 121494
rect 148144 114494 148464 121258
rect 148144 114258 148186 114494
rect 148422 114258 148464 114494
rect 148144 107494 148464 114258
rect 148144 107258 148186 107494
rect 148422 107258 148464 107494
rect 148144 100494 148464 107258
rect 148144 100258 148186 100494
rect 148422 100258 148464 100494
rect 148144 93494 148464 100258
rect 148144 93258 148186 93494
rect 148422 93258 148464 93494
rect 148144 86494 148464 93258
rect 148144 86258 148186 86494
rect 148422 86258 148464 86494
rect 148144 79494 148464 86258
rect 148144 79258 148186 79494
rect 148422 79258 148464 79494
rect 148144 72494 148464 79258
rect 148144 72258 148186 72494
rect 148422 72258 148464 72494
rect 148144 65494 148464 72258
rect 148144 65258 148186 65494
rect 148422 65258 148464 65494
rect 148144 58494 148464 65258
rect 148144 58258 148186 58494
rect 148422 58258 148464 58494
rect 148144 51494 148464 58258
rect 148144 51258 148186 51494
rect 148422 51258 148464 51494
rect 148144 44494 148464 51258
rect 148144 44258 148186 44494
rect 148422 44258 148464 44494
rect 148144 37494 148464 44258
rect 148144 37258 148186 37494
rect 148422 37258 148464 37494
rect 148144 30494 148464 37258
rect 148144 30258 148186 30494
rect 148422 30258 148464 30494
rect 148144 23494 148464 30258
rect 148144 23258 148186 23494
rect 148422 23258 148464 23494
rect 148144 16494 148464 23258
rect 148144 16258 148186 16494
rect 148422 16258 148464 16494
rect 148144 9494 148464 16258
rect 148144 9258 148186 9494
rect 148422 9258 148464 9494
rect 148144 2494 148464 9258
rect 148144 2258 148186 2494
rect 148422 2258 148464 2494
rect 148144 -746 148464 2258
rect 148144 -982 148186 -746
rect 148422 -982 148464 -746
rect 148144 -1066 148464 -982
rect 148144 -1302 148186 -1066
rect 148422 -1302 148464 -1066
rect 148144 -2294 148464 -1302
rect 149876 706198 150196 706230
rect 149876 705962 149918 706198
rect 150154 705962 150196 706198
rect 149876 705878 150196 705962
rect 149876 705642 149918 705878
rect 150154 705642 150196 705878
rect 149876 696434 150196 705642
rect 149876 696198 149918 696434
rect 150154 696198 150196 696434
rect 149876 689434 150196 696198
rect 149876 689198 149918 689434
rect 150154 689198 150196 689434
rect 149876 682434 150196 689198
rect 149876 682198 149918 682434
rect 150154 682198 150196 682434
rect 149876 675434 150196 682198
rect 149876 675198 149918 675434
rect 150154 675198 150196 675434
rect 149876 668434 150196 675198
rect 149876 668198 149918 668434
rect 150154 668198 150196 668434
rect 149876 661434 150196 668198
rect 149876 661198 149918 661434
rect 150154 661198 150196 661434
rect 149876 654434 150196 661198
rect 149876 654198 149918 654434
rect 150154 654198 150196 654434
rect 149876 647434 150196 654198
rect 149876 647198 149918 647434
rect 150154 647198 150196 647434
rect 149876 640434 150196 647198
rect 149876 640198 149918 640434
rect 150154 640198 150196 640434
rect 149876 633434 150196 640198
rect 149876 633198 149918 633434
rect 150154 633198 150196 633434
rect 149876 626434 150196 633198
rect 149876 626198 149918 626434
rect 150154 626198 150196 626434
rect 149876 619434 150196 626198
rect 149876 619198 149918 619434
rect 150154 619198 150196 619434
rect 149876 612434 150196 619198
rect 149876 612198 149918 612434
rect 150154 612198 150196 612434
rect 149876 605434 150196 612198
rect 149876 605198 149918 605434
rect 150154 605198 150196 605434
rect 149876 598434 150196 605198
rect 149876 598198 149918 598434
rect 150154 598198 150196 598434
rect 149876 591434 150196 598198
rect 149876 591198 149918 591434
rect 150154 591198 150196 591434
rect 149876 584434 150196 591198
rect 149876 584198 149918 584434
rect 150154 584198 150196 584434
rect 149876 577434 150196 584198
rect 149876 577198 149918 577434
rect 150154 577198 150196 577434
rect 149876 570434 150196 577198
rect 149876 570198 149918 570434
rect 150154 570198 150196 570434
rect 149876 563434 150196 570198
rect 149876 563198 149918 563434
rect 150154 563198 150196 563434
rect 149876 556434 150196 563198
rect 149876 556198 149918 556434
rect 150154 556198 150196 556434
rect 149876 549434 150196 556198
rect 149876 549198 149918 549434
rect 150154 549198 150196 549434
rect 149876 542434 150196 549198
rect 149876 542198 149918 542434
rect 150154 542198 150196 542434
rect 149876 535434 150196 542198
rect 149876 535198 149918 535434
rect 150154 535198 150196 535434
rect 149876 528434 150196 535198
rect 149876 528198 149918 528434
rect 150154 528198 150196 528434
rect 149876 521434 150196 528198
rect 149876 521198 149918 521434
rect 150154 521198 150196 521434
rect 149876 514434 150196 521198
rect 149876 514198 149918 514434
rect 150154 514198 150196 514434
rect 149876 507434 150196 514198
rect 149876 507198 149918 507434
rect 150154 507198 150196 507434
rect 149876 500434 150196 507198
rect 149876 500198 149918 500434
rect 150154 500198 150196 500434
rect 149876 493434 150196 500198
rect 149876 493198 149918 493434
rect 150154 493198 150196 493434
rect 149876 486434 150196 493198
rect 149876 486198 149918 486434
rect 150154 486198 150196 486434
rect 149876 479434 150196 486198
rect 149876 479198 149918 479434
rect 150154 479198 150196 479434
rect 149876 472434 150196 479198
rect 149876 472198 149918 472434
rect 150154 472198 150196 472434
rect 149876 465434 150196 472198
rect 149876 465198 149918 465434
rect 150154 465198 150196 465434
rect 149876 458434 150196 465198
rect 149876 458198 149918 458434
rect 150154 458198 150196 458434
rect 149876 451434 150196 458198
rect 149876 451198 149918 451434
rect 150154 451198 150196 451434
rect 149876 444434 150196 451198
rect 149876 444198 149918 444434
rect 150154 444198 150196 444434
rect 149876 437434 150196 444198
rect 149876 437198 149918 437434
rect 150154 437198 150196 437434
rect 149876 430434 150196 437198
rect 149876 430198 149918 430434
rect 150154 430198 150196 430434
rect 149876 423434 150196 430198
rect 149876 423198 149918 423434
rect 150154 423198 150196 423434
rect 149876 416434 150196 423198
rect 149876 416198 149918 416434
rect 150154 416198 150196 416434
rect 149876 409434 150196 416198
rect 149876 409198 149918 409434
rect 150154 409198 150196 409434
rect 149876 402434 150196 409198
rect 149876 402198 149918 402434
rect 150154 402198 150196 402434
rect 149876 395434 150196 402198
rect 149876 395198 149918 395434
rect 150154 395198 150196 395434
rect 149876 388434 150196 395198
rect 149876 388198 149918 388434
rect 150154 388198 150196 388434
rect 149876 381434 150196 388198
rect 149876 381198 149918 381434
rect 150154 381198 150196 381434
rect 149876 374434 150196 381198
rect 149876 374198 149918 374434
rect 150154 374198 150196 374434
rect 149876 367434 150196 374198
rect 149876 367198 149918 367434
rect 150154 367198 150196 367434
rect 149876 360434 150196 367198
rect 149876 360198 149918 360434
rect 150154 360198 150196 360434
rect 149876 353434 150196 360198
rect 149876 353198 149918 353434
rect 150154 353198 150196 353434
rect 149876 346434 150196 353198
rect 149876 346198 149918 346434
rect 150154 346198 150196 346434
rect 149876 339434 150196 346198
rect 149876 339198 149918 339434
rect 150154 339198 150196 339434
rect 149876 332434 150196 339198
rect 149876 332198 149918 332434
rect 150154 332198 150196 332434
rect 149876 325434 150196 332198
rect 149876 325198 149918 325434
rect 150154 325198 150196 325434
rect 149876 318434 150196 325198
rect 149876 318198 149918 318434
rect 150154 318198 150196 318434
rect 149876 311434 150196 318198
rect 149876 311198 149918 311434
rect 150154 311198 150196 311434
rect 149876 304434 150196 311198
rect 149876 304198 149918 304434
rect 150154 304198 150196 304434
rect 149876 297434 150196 304198
rect 149876 297198 149918 297434
rect 150154 297198 150196 297434
rect 149876 290434 150196 297198
rect 149876 290198 149918 290434
rect 150154 290198 150196 290434
rect 149876 283434 150196 290198
rect 149876 283198 149918 283434
rect 150154 283198 150196 283434
rect 149876 276434 150196 283198
rect 149876 276198 149918 276434
rect 150154 276198 150196 276434
rect 149876 269434 150196 276198
rect 149876 269198 149918 269434
rect 150154 269198 150196 269434
rect 149876 262434 150196 269198
rect 149876 262198 149918 262434
rect 150154 262198 150196 262434
rect 149876 255434 150196 262198
rect 149876 255198 149918 255434
rect 150154 255198 150196 255434
rect 149876 248434 150196 255198
rect 149876 248198 149918 248434
rect 150154 248198 150196 248434
rect 149876 241434 150196 248198
rect 149876 241198 149918 241434
rect 150154 241198 150196 241434
rect 149876 234434 150196 241198
rect 149876 234198 149918 234434
rect 150154 234198 150196 234434
rect 149876 227434 150196 234198
rect 149876 227198 149918 227434
rect 150154 227198 150196 227434
rect 149876 220434 150196 227198
rect 149876 220198 149918 220434
rect 150154 220198 150196 220434
rect 149876 213434 150196 220198
rect 149876 213198 149918 213434
rect 150154 213198 150196 213434
rect 149876 206434 150196 213198
rect 149876 206198 149918 206434
rect 150154 206198 150196 206434
rect 149876 199434 150196 206198
rect 149876 199198 149918 199434
rect 150154 199198 150196 199434
rect 149876 192434 150196 199198
rect 149876 192198 149918 192434
rect 150154 192198 150196 192434
rect 149876 185434 150196 192198
rect 149876 185198 149918 185434
rect 150154 185198 150196 185434
rect 149876 178434 150196 185198
rect 149876 178198 149918 178434
rect 150154 178198 150196 178434
rect 149876 171434 150196 178198
rect 149876 171198 149918 171434
rect 150154 171198 150196 171434
rect 149876 164434 150196 171198
rect 149876 164198 149918 164434
rect 150154 164198 150196 164434
rect 149876 157434 150196 164198
rect 149876 157198 149918 157434
rect 150154 157198 150196 157434
rect 149876 150434 150196 157198
rect 149876 150198 149918 150434
rect 150154 150198 150196 150434
rect 149876 143434 150196 150198
rect 149876 143198 149918 143434
rect 150154 143198 150196 143434
rect 149876 136434 150196 143198
rect 149876 136198 149918 136434
rect 150154 136198 150196 136434
rect 149876 129434 150196 136198
rect 149876 129198 149918 129434
rect 150154 129198 150196 129434
rect 149876 122434 150196 129198
rect 149876 122198 149918 122434
rect 150154 122198 150196 122434
rect 149876 115434 150196 122198
rect 149876 115198 149918 115434
rect 150154 115198 150196 115434
rect 149876 108434 150196 115198
rect 149876 108198 149918 108434
rect 150154 108198 150196 108434
rect 149876 101434 150196 108198
rect 149876 101198 149918 101434
rect 150154 101198 150196 101434
rect 149876 94434 150196 101198
rect 149876 94198 149918 94434
rect 150154 94198 150196 94434
rect 149876 87434 150196 94198
rect 149876 87198 149918 87434
rect 150154 87198 150196 87434
rect 149876 80434 150196 87198
rect 149876 80198 149918 80434
rect 150154 80198 150196 80434
rect 149876 73434 150196 80198
rect 149876 73198 149918 73434
rect 150154 73198 150196 73434
rect 149876 66434 150196 73198
rect 149876 66198 149918 66434
rect 150154 66198 150196 66434
rect 149876 59434 150196 66198
rect 149876 59198 149918 59434
rect 150154 59198 150196 59434
rect 149876 52434 150196 59198
rect 149876 52198 149918 52434
rect 150154 52198 150196 52434
rect 149876 45434 150196 52198
rect 149876 45198 149918 45434
rect 150154 45198 150196 45434
rect 149876 38434 150196 45198
rect 149876 38198 149918 38434
rect 150154 38198 150196 38434
rect 149876 31434 150196 38198
rect 149876 31198 149918 31434
rect 150154 31198 150196 31434
rect 149876 24434 150196 31198
rect 149876 24198 149918 24434
rect 150154 24198 150196 24434
rect 149876 17434 150196 24198
rect 149876 17198 149918 17434
rect 150154 17198 150196 17434
rect 149876 10434 150196 17198
rect 149876 10198 149918 10434
rect 150154 10198 150196 10434
rect 149876 3434 150196 10198
rect 149876 3198 149918 3434
rect 150154 3198 150196 3434
rect 149876 -1706 150196 3198
rect 149876 -1942 149918 -1706
rect 150154 -1942 150196 -1706
rect 149876 -2026 150196 -1942
rect 149876 -2262 149918 -2026
rect 150154 -2262 150196 -2026
rect 149876 -2294 150196 -2262
rect 155144 705238 155464 706230
rect 155144 705002 155186 705238
rect 155422 705002 155464 705238
rect 155144 704918 155464 705002
rect 155144 704682 155186 704918
rect 155422 704682 155464 704918
rect 155144 695494 155464 704682
rect 155144 695258 155186 695494
rect 155422 695258 155464 695494
rect 155144 688494 155464 695258
rect 155144 688258 155186 688494
rect 155422 688258 155464 688494
rect 155144 681494 155464 688258
rect 155144 681258 155186 681494
rect 155422 681258 155464 681494
rect 155144 674494 155464 681258
rect 155144 674258 155186 674494
rect 155422 674258 155464 674494
rect 155144 667494 155464 674258
rect 155144 667258 155186 667494
rect 155422 667258 155464 667494
rect 155144 660494 155464 667258
rect 155144 660258 155186 660494
rect 155422 660258 155464 660494
rect 155144 653494 155464 660258
rect 155144 653258 155186 653494
rect 155422 653258 155464 653494
rect 155144 646494 155464 653258
rect 155144 646258 155186 646494
rect 155422 646258 155464 646494
rect 155144 639494 155464 646258
rect 155144 639258 155186 639494
rect 155422 639258 155464 639494
rect 155144 632494 155464 639258
rect 155144 632258 155186 632494
rect 155422 632258 155464 632494
rect 155144 625494 155464 632258
rect 155144 625258 155186 625494
rect 155422 625258 155464 625494
rect 155144 618494 155464 625258
rect 155144 618258 155186 618494
rect 155422 618258 155464 618494
rect 155144 611494 155464 618258
rect 155144 611258 155186 611494
rect 155422 611258 155464 611494
rect 155144 604494 155464 611258
rect 155144 604258 155186 604494
rect 155422 604258 155464 604494
rect 155144 597494 155464 604258
rect 155144 597258 155186 597494
rect 155422 597258 155464 597494
rect 155144 590494 155464 597258
rect 155144 590258 155186 590494
rect 155422 590258 155464 590494
rect 155144 583494 155464 590258
rect 155144 583258 155186 583494
rect 155422 583258 155464 583494
rect 155144 576494 155464 583258
rect 155144 576258 155186 576494
rect 155422 576258 155464 576494
rect 155144 569494 155464 576258
rect 155144 569258 155186 569494
rect 155422 569258 155464 569494
rect 155144 562494 155464 569258
rect 155144 562258 155186 562494
rect 155422 562258 155464 562494
rect 155144 555494 155464 562258
rect 155144 555258 155186 555494
rect 155422 555258 155464 555494
rect 155144 548494 155464 555258
rect 155144 548258 155186 548494
rect 155422 548258 155464 548494
rect 155144 541494 155464 548258
rect 155144 541258 155186 541494
rect 155422 541258 155464 541494
rect 155144 534494 155464 541258
rect 155144 534258 155186 534494
rect 155422 534258 155464 534494
rect 155144 527494 155464 534258
rect 155144 527258 155186 527494
rect 155422 527258 155464 527494
rect 155144 520494 155464 527258
rect 155144 520258 155186 520494
rect 155422 520258 155464 520494
rect 155144 513494 155464 520258
rect 155144 513258 155186 513494
rect 155422 513258 155464 513494
rect 155144 506494 155464 513258
rect 155144 506258 155186 506494
rect 155422 506258 155464 506494
rect 155144 499494 155464 506258
rect 155144 499258 155186 499494
rect 155422 499258 155464 499494
rect 155144 492494 155464 499258
rect 155144 492258 155186 492494
rect 155422 492258 155464 492494
rect 155144 485494 155464 492258
rect 155144 485258 155186 485494
rect 155422 485258 155464 485494
rect 155144 478494 155464 485258
rect 155144 478258 155186 478494
rect 155422 478258 155464 478494
rect 155144 471494 155464 478258
rect 155144 471258 155186 471494
rect 155422 471258 155464 471494
rect 155144 464494 155464 471258
rect 155144 464258 155186 464494
rect 155422 464258 155464 464494
rect 155144 457494 155464 464258
rect 155144 457258 155186 457494
rect 155422 457258 155464 457494
rect 155144 450494 155464 457258
rect 155144 450258 155186 450494
rect 155422 450258 155464 450494
rect 155144 443494 155464 450258
rect 155144 443258 155186 443494
rect 155422 443258 155464 443494
rect 155144 436494 155464 443258
rect 155144 436258 155186 436494
rect 155422 436258 155464 436494
rect 155144 429494 155464 436258
rect 155144 429258 155186 429494
rect 155422 429258 155464 429494
rect 155144 422494 155464 429258
rect 155144 422258 155186 422494
rect 155422 422258 155464 422494
rect 155144 415494 155464 422258
rect 155144 415258 155186 415494
rect 155422 415258 155464 415494
rect 155144 408494 155464 415258
rect 155144 408258 155186 408494
rect 155422 408258 155464 408494
rect 155144 401494 155464 408258
rect 155144 401258 155186 401494
rect 155422 401258 155464 401494
rect 155144 394494 155464 401258
rect 155144 394258 155186 394494
rect 155422 394258 155464 394494
rect 155144 387494 155464 394258
rect 155144 387258 155186 387494
rect 155422 387258 155464 387494
rect 155144 380494 155464 387258
rect 155144 380258 155186 380494
rect 155422 380258 155464 380494
rect 155144 373494 155464 380258
rect 155144 373258 155186 373494
rect 155422 373258 155464 373494
rect 155144 366494 155464 373258
rect 155144 366258 155186 366494
rect 155422 366258 155464 366494
rect 155144 359494 155464 366258
rect 155144 359258 155186 359494
rect 155422 359258 155464 359494
rect 155144 352494 155464 359258
rect 155144 352258 155186 352494
rect 155422 352258 155464 352494
rect 155144 345494 155464 352258
rect 155144 345258 155186 345494
rect 155422 345258 155464 345494
rect 155144 338494 155464 345258
rect 155144 338258 155186 338494
rect 155422 338258 155464 338494
rect 155144 331494 155464 338258
rect 155144 331258 155186 331494
rect 155422 331258 155464 331494
rect 155144 324494 155464 331258
rect 155144 324258 155186 324494
rect 155422 324258 155464 324494
rect 155144 317494 155464 324258
rect 155144 317258 155186 317494
rect 155422 317258 155464 317494
rect 155144 310494 155464 317258
rect 155144 310258 155186 310494
rect 155422 310258 155464 310494
rect 155144 303494 155464 310258
rect 155144 303258 155186 303494
rect 155422 303258 155464 303494
rect 155144 296494 155464 303258
rect 155144 296258 155186 296494
rect 155422 296258 155464 296494
rect 155144 289494 155464 296258
rect 155144 289258 155186 289494
rect 155422 289258 155464 289494
rect 155144 282494 155464 289258
rect 155144 282258 155186 282494
rect 155422 282258 155464 282494
rect 155144 275494 155464 282258
rect 155144 275258 155186 275494
rect 155422 275258 155464 275494
rect 155144 268494 155464 275258
rect 155144 268258 155186 268494
rect 155422 268258 155464 268494
rect 155144 261494 155464 268258
rect 155144 261258 155186 261494
rect 155422 261258 155464 261494
rect 155144 254494 155464 261258
rect 155144 254258 155186 254494
rect 155422 254258 155464 254494
rect 155144 247494 155464 254258
rect 155144 247258 155186 247494
rect 155422 247258 155464 247494
rect 155144 240494 155464 247258
rect 155144 240258 155186 240494
rect 155422 240258 155464 240494
rect 155144 233494 155464 240258
rect 155144 233258 155186 233494
rect 155422 233258 155464 233494
rect 155144 226494 155464 233258
rect 155144 226258 155186 226494
rect 155422 226258 155464 226494
rect 155144 219494 155464 226258
rect 155144 219258 155186 219494
rect 155422 219258 155464 219494
rect 155144 212494 155464 219258
rect 155144 212258 155186 212494
rect 155422 212258 155464 212494
rect 155144 205494 155464 212258
rect 155144 205258 155186 205494
rect 155422 205258 155464 205494
rect 155144 198494 155464 205258
rect 155144 198258 155186 198494
rect 155422 198258 155464 198494
rect 155144 191494 155464 198258
rect 155144 191258 155186 191494
rect 155422 191258 155464 191494
rect 155144 184494 155464 191258
rect 155144 184258 155186 184494
rect 155422 184258 155464 184494
rect 155144 177494 155464 184258
rect 155144 177258 155186 177494
rect 155422 177258 155464 177494
rect 155144 170494 155464 177258
rect 155144 170258 155186 170494
rect 155422 170258 155464 170494
rect 155144 163494 155464 170258
rect 155144 163258 155186 163494
rect 155422 163258 155464 163494
rect 155144 156494 155464 163258
rect 155144 156258 155186 156494
rect 155422 156258 155464 156494
rect 155144 149494 155464 156258
rect 155144 149258 155186 149494
rect 155422 149258 155464 149494
rect 155144 142494 155464 149258
rect 155144 142258 155186 142494
rect 155422 142258 155464 142494
rect 155144 135494 155464 142258
rect 155144 135258 155186 135494
rect 155422 135258 155464 135494
rect 155144 128494 155464 135258
rect 155144 128258 155186 128494
rect 155422 128258 155464 128494
rect 155144 121494 155464 128258
rect 155144 121258 155186 121494
rect 155422 121258 155464 121494
rect 155144 114494 155464 121258
rect 155144 114258 155186 114494
rect 155422 114258 155464 114494
rect 155144 107494 155464 114258
rect 155144 107258 155186 107494
rect 155422 107258 155464 107494
rect 155144 100494 155464 107258
rect 155144 100258 155186 100494
rect 155422 100258 155464 100494
rect 155144 93494 155464 100258
rect 155144 93258 155186 93494
rect 155422 93258 155464 93494
rect 155144 86494 155464 93258
rect 155144 86258 155186 86494
rect 155422 86258 155464 86494
rect 155144 79494 155464 86258
rect 155144 79258 155186 79494
rect 155422 79258 155464 79494
rect 155144 72494 155464 79258
rect 155144 72258 155186 72494
rect 155422 72258 155464 72494
rect 155144 65494 155464 72258
rect 155144 65258 155186 65494
rect 155422 65258 155464 65494
rect 155144 58494 155464 65258
rect 155144 58258 155186 58494
rect 155422 58258 155464 58494
rect 155144 51494 155464 58258
rect 155144 51258 155186 51494
rect 155422 51258 155464 51494
rect 155144 44494 155464 51258
rect 155144 44258 155186 44494
rect 155422 44258 155464 44494
rect 155144 37494 155464 44258
rect 155144 37258 155186 37494
rect 155422 37258 155464 37494
rect 155144 30494 155464 37258
rect 155144 30258 155186 30494
rect 155422 30258 155464 30494
rect 155144 23494 155464 30258
rect 155144 23258 155186 23494
rect 155422 23258 155464 23494
rect 155144 16494 155464 23258
rect 155144 16258 155186 16494
rect 155422 16258 155464 16494
rect 155144 9494 155464 16258
rect 155144 9258 155186 9494
rect 155422 9258 155464 9494
rect 155144 2494 155464 9258
rect 155144 2258 155186 2494
rect 155422 2258 155464 2494
rect 155144 -746 155464 2258
rect 155144 -982 155186 -746
rect 155422 -982 155464 -746
rect 155144 -1066 155464 -982
rect 155144 -1302 155186 -1066
rect 155422 -1302 155464 -1066
rect 155144 -2294 155464 -1302
rect 156876 706198 157196 706230
rect 156876 705962 156918 706198
rect 157154 705962 157196 706198
rect 156876 705878 157196 705962
rect 156876 705642 156918 705878
rect 157154 705642 157196 705878
rect 156876 696434 157196 705642
rect 156876 696198 156918 696434
rect 157154 696198 157196 696434
rect 156876 689434 157196 696198
rect 156876 689198 156918 689434
rect 157154 689198 157196 689434
rect 156876 682434 157196 689198
rect 156876 682198 156918 682434
rect 157154 682198 157196 682434
rect 156876 675434 157196 682198
rect 156876 675198 156918 675434
rect 157154 675198 157196 675434
rect 156876 668434 157196 675198
rect 156876 668198 156918 668434
rect 157154 668198 157196 668434
rect 156876 661434 157196 668198
rect 156876 661198 156918 661434
rect 157154 661198 157196 661434
rect 156876 654434 157196 661198
rect 156876 654198 156918 654434
rect 157154 654198 157196 654434
rect 156876 647434 157196 654198
rect 156876 647198 156918 647434
rect 157154 647198 157196 647434
rect 156876 640434 157196 647198
rect 156876 640198 156918 640434
rect 157154 640198 157196 640434
rect 156876 633434 157196 640198
rect 156876 633198 156918 633434
rect 157154 633198 157196 633434
rect 156876 626434 157196 633198
rect 156876 626198 156918 626434
rect 157154 626198 157196 626434
rect 156876 619434 157196 626198
rect 156876 619198 156918 619434
rect 157154 619198 157196 619434
rect 156876 612434 157196 619198
rect 156876 612198 156918 612434
rect 157154 612198 157196 612434
rect 156876 605434 157196 612198
rect 156876 605198 156918 605434
rect 157154 605198 157196 605434
rect 156876 598434 157196 605198
rect 156876 598198 156918 598434
rect 157154 598198 157196 598434
rect 156876 591434 157196 598198
rect 156876 591198 156918 591434
rect 157154 591198 157196 591434
rect 156876 584434 157196 591198
rect 156876 584198 156918 584434
rect 157154 584198 157196 584434
rect 156876 577434 157196 584198
rect 156876 577198 156918 577434
rect 157154 577198 157196 577434
rect 156876 570434 157196 577198
rect 156876 570198 156918 570434
rect 157154 570198 157196 570434
rect 156876 563434 157196 570198
rect 156876 563198 156918 563434
rect 157154 563198 157196 563434
rect 156876 556434 157196 563198
rect 156876 556198 156918 556434
rect 157154 556198 157196 556434
rect 156876 549434 157196 556198
rect 156876 549198 156918 549434
rect 157154 549198 157196 549434
rect 156876 542434 157196 549198
rect 156876 542198 156918 542434
rect 157154 542198 157196 542434
rect 156876 535434 157196 542198
rect 156876 535198 156918 535434
rect 157154 535198 157196 535434
rect 156876 528434 157196 535198
rect 156876 528198 156918 528434
rect 157154 528198 157196 528434
rect 156876 521434 157196 528198
rect 156876 521198 156918 521434
rect 157154 521198 157196 521434
rect 156876 514434 157196 521198
rect 156876 514198 156918 514434
rect 157154 514198 157196 514434
rect 156876 507434 157196 514198
rect 156876 507198 156918 507434
rect 157154 507198 157196 507434
rect 156876 500434 157196 507198
rect 156876 500198 156918 500434
rect 157154 500198 157196 500434
rect 156876 493434 157196 500198
rect 156876 493198 156918 493434
rect 157154 493198 157196 493434
rect 156876 486434 157196 493198
rect 156876 486198 156918 486434
rect 157154 486198 157196 486434
rect 156876 479434 157196 486198
rect 156876 479198 156918 479434
rect 157154 479198 157196 479434
rect 156876 472434 157196 479198
rect 156876 472198 156918 472434
rect 157154 472198 157196 472434
rect 156876 465434 157196 472198
rect 156876 465198 156918 465434
rect 157154 465198 157196 465434
rect 156876 458434 157196 465198
rect 156876 458198 156918 458434
rect 157154 458198 157196 458434
rect 156876 451434 157196 458198
rect 156876 451198 156918 451434
rect 157154 451198 157196 451434
rect 156876 444434 157196 451198
rect 156876 444198 156918 444434
rect 157154 444198 157196 444434
rect 156876 437434 157196 444198
rect 156876 437198 156918 437434
rect 157154 437198 157196 437434
rect 156876 430434 157196 437198
rect 156876 430198 156918 430434
rect 157154 430198 157196 430434
rect 156876 423434 157196 430198
rect 156876 423198 156918 423434
rect 157154 423198 157196 423434
rect 156876 416434 157196 423198
rect 156876 416198 156918 416434
rect 157154 416198 157196 416434
rect 156876 409434 157196 416198
rect 156876 409198 156918 409434
rect 157154 409198 157196 409434
rect 156876 402434 157196 409198
rect 156876 402198 156918 402434
rect 157154 402198 157196 402434
rect 156876 395434 157196 402198
rect 156876 395198 156918 395434
rect 157154 395198 157196 395434
rect 156876 388434 157196 395198
rect 156876 388198 156918 388434
rect 157154 388198 157196 388434
rect 156876 381434 157196 388198
rect 156876 381198 156918 381434
rect 157154 381198 157196 381434
rect 156876 374434 157196 381198
rect 156876 374198 156918 374434
rect 157154 374198 157196 374434
rect 156876 367434 157196 374198
rect 156876 367198 156918 367434
rect 157154 367198 157196 367434
rect 156876 360434 157196 367198
rect 156876 360198 156918 360434
rect 157154 360198 157196 360434
rect 156876 353434 157196 360198
rect 156876 353198 156918 353434
rect 157154 353198 157196 353434
rect 156876 346434 157196 353198
rect 156876 346198 156918 346434
rect 157154 346198 157196 346434
rect 156876 339434 157196 346198
rect 156876 339198 156918 339434
rect 157154 339198 157196 339434
rect 156876 332434 157196 339198
rect 156876 332198 156918 332434
rect 157154 332198 157196 332434
rect 156876 325434 157196 332198
rect 156876 325198 156918 325434
rect 157154 325198 157196 325434
rect 156876 318434 157196 325198
rect 156876 318198 156918 318434
rect 157154 318198 157196 318434
rect 156876 311434 157196 318198
rect 156876 311198 156918 311434
rect 157154 311198 157196 311434
rect 156876 304434 157196 311198
rect 156876 304198 156918 304434
rect 157154 304198 157196 304434
rect 156876 297434 157196 304198
rect 156876 297198 156918 297434
rect 157154 297198 157196 297434
rect 156876 290434 157196 297198
rect 156876 290198 156918 290434
rect 157154 290198 157196 290434
rect 156876 283434 157196 290198
rect 156876 283198 156918 283434
rect 157154 283198 157196 283434
rect 156876 276434 157196 283198
rect 156876 276198 156918 276434
rect 157154 276198 157196 276434
rect 156876 269434 157196 276198
rect 156876 269198 156918 269434
rect 157154 269198 157196 269434
rect 156876 262434 157196 269198
rect 156876 262198 156918 262434
rect 157154 262198 157196 262434
rect 156876 255434 157196 262198
rect 156876 255198 156918 255434
rect 157154 255198 157196 255434
rect 156876 248434 157196 255198
rect 156876 248198 156918 248434
rect 157154 248198 157196 248434
rect 156876 241434 157196 248198
rect 156876 241198 156918 241434
rect 157154 241198 157196 241434
rect 156876 234434 157196 241198
rect 156876 234198 156918 234434
rect 157154 234198 157196 234434
rect 156876 227434 157196 234198
rect 156876 227198 156918 227434
rect 157154 227198 157196 227434
rect 156876 220434 157196 227198
rect 156876 220198 156918 220434
rect 157154 220198 157196 220434
rect 156876 213434 157196 220198
rect 156876 213198 156918 213434
rect 157154 213198 157196 213434
rect 156876 206434 157196 213198
rect 156876 206198 156918 206434
rect 157154 206198 157196 206434
rect 156876 199434 157196 206198
rect 156876 199198 156918 199434
rect 157154 199198 157196 199434
rect 156876 192434 157196 199198
rect 156876 192198 156918 192434
rect 157154 192198 157196 192434
rect 156876 185434 157196 192198
rect 156876 185198 156918 185434
rect 157154 185198 157196 185434
rect 156876 178434 157196 185198
rect 156876 178198 156918 178434
rect 157154 178198 157196 178434
rect 156876 171434 157196 178198
rect 156876 171198 156918 171434
rect 157154 171198 157196 171434
rect 156876 164434 157196 171198
rect 156876 164198 156918 164434
rect 157154 164198 157196 164434
rect 156876 157434 157196 164198
rect 156876 157198 156918 157434
rect 157154 157198 157196 157434
rect 156876 150434 157196 157198
rect 156876 150198 156918 150434
rect 157154 150198 157196 150434
rect 156876 143434 157196 150198
rect 156876 143198 156918 143434
rect 157154 143198 157196 143434
rect 156876 136434 157196 143198
rect 156876 136198 156918 136434
rect 157154 136198 157196 136434
rect 156876 129434 157196 136198
rect 156876 129198 156918 129434
rect 157154 129198 157196 129434
rect 156876 122434 157196 129198
rect 156876 122198 156918 122434
rect 157154 122198 157196 122434
rect 156876 115434 157196 122198
rect 156876 115198 156918 115434
rect 157154 115198 157196 115434
rect 156876 108434 157196 115198
rect 156876 108198 156918 108434
rect 157154 108198 157196 108434
rect 156876 101434 157196 108198
rect 156876 101198 156918 101434
rect 157154 101198 157196 101434
rect 156876 94434 157196 101198
rect 156876 94198 156918 94434
rect 157154 94198 157196 94434
rect 156876 87434 157196 94198
rect 156876 87198 156918 87434
rect 157154 87198 157196 87434
rect 156876 80434 157196 87198
rect 156876 80198 156918 80434
rect 157154 80198 157196 80434
rect 156876 73434 157196 80198
rect 156876 73198 156918 73434
rect 157154 73198 157196 73434
rect 156876 66434 157196 73198
rect 156876 66198 156918 66434
rect 157154 66198 157196 66434
rect 156876 59434 157196 66198
rect 156876 59198 156918 59434
rect 157154 59198 157196 59434
rect 156876 52434 157196 59198
rect 156876 52198 156918 52434
rect 157154 52198 157196 52434
rect 156876 45434 157196 52198
rect 156876 45198 156918 45434
rect 157154 45198 157196 45434
rect 156876 38434 157196 45198
rect 156876 38198 156918 38434
rect 157154 38198 157196 38434
rect 156876 31434 157196 38198
rect 156876 31198 156918 31434
rect 157154 31198 157196 31434
rect 156876 24434 157196 31198
rect 156876 24198 156918 24434
rect 157154 24198 157196 24434
rect 156876 17434 157196 24198
rect 156876 17198 156918 17434
rect 157154 17198 157196 17434
rect 156876 10434 157196 17198
rect 156876 10198 156918 10434
rect 157154 10198 157196 10434
rect 156876 3434 157196 10198
rect 156876 3198 156918 3434
rect 157154 3198 157196 3434
rect 156876 -1706 157196 3198
rect 156876 -1942 156918 -1706
rect 157154 -1942 157196 -1706
rect 156876 -2026 157196 -1942
rect 156876 -2262 156918 -2026
rect 157154 -2262 157196 -2026
rect 156876 -2294 157196 -2262
rect 162144 705238 162464 706230
rect 162144 705002 162186 705238
rect 162422 705002 162464 705238
rect 162144 704918 162464 705002
rect 162144 704682 162186 704918
rect 162422 704682 162464 704918
rect 162144 695494 162464 704682
rect 162144 695258 162186 695494
rect 162422 695258 162464 695494
rect 162144 688494 162464 695258
rect 162144 688258 162186 688494
rect 162422 688258 162464 688494
rect 162144 681494 162464 688258
rect 162144 681258 162186 681494
rect 162422 681258 162464 681494
rect 162144 674494 162464 681258
rect 162144 674258 162186 674494
rect 162422 674258 162464 674494
rect 162144 667494 162464 674258
rect 162144 667258 162186 667494
rect 162422 667258 162464 667494
rect 162144 660494 162464 667258
rect 162144 660258 162186 660494
rect 162422 660258 162464 660494
rect 162144 653494 162464 660258
rect 162144 653258 162186 653494
rect 162422 653258 162464 653494
rect 162144 646494 162464 653258
rect 162144 646258 162186 646494
rect 162422 646258 162464 646494
rect 162144 639494 162464 646258
rect 162144 639258 162186 639494
rect 162422 639258 162464 639494
rect 162144 632494 162464 639258
rect 162144 632258 162186 632494
rect 162422 632258 162464 632494
rect 162144 625494 162464 632258
rect 162144 625258 162186 625494
rect 162422 625258 162464 625494
rect 162144 618494 162464 625258
rect 162144 618258 162186 618494
rect 162422 618258 162464 618494
rect 162144 611494 162464 618258
rect 162144 611258 162186 611494
rect 162422 611258 162464 611494
rect 162144 604494 162464 611258
rect 162144 604258 162186 604494
rect 162422 604258 162464 604494
rect 162144 597494 162464 604258
rect 162144 597258 162186 597494
rect 162422 597258 162464 597494
rect 162144 590494 162464 597258
rect 162144 590258 162186 590494
rect 162422 590258 162464 590494
rect 162144 583494 162464 590258
rect 162144 583258 162186 583494
rect 162422 583258 162464 583494
rect 162144 576494 162464 583258
rect 162144 576258 162186 576494
rect 162422 576258 162464 576494
rect 162144 569494 162464 576258
rect 162144 569258 162186 569494
rect 162422 569258 162464 569494
rect 162144 562494 162464 569258
rect 162144 562258 162186 562494
rect 162422 562258 162464 562494
rect 162144 555494 162464 562258
rect 162144 555258 162186 555494
rect 162422 555258 162464 555494
rect 162144 548494 162464 555258
rect 162144 548258 162186 548494
rect 162422 548258 162464 548494
rect 162144 541494 162464 548258
rect 162144 541258 162186 541494
rect 162422 541258 162464 541494
rect 162144 534494 162464 541258
rect 162144 534258 162186 534494
rect 162422 534258 162464 534494
rect 162144 527494 162464 534258
rect 162144 527258 162186 527494
rect 162422 527258 162464 527494
rect 162144 520494 162464 527258
rect 162144 520258 162186 520494
rect 162422 520258 162464 520494
rect 162144 513494 162464 520258
rect 162144 513258 162186 513494
rect 162422 513258 162464 513494
rect 162144 506494 162464 513258
rect 162144 506258 162186 506494
rect 162422 506258 162464 506494
rect 162144 499494 162464 506258
rect 162144 499258 162186 499494
rect 162422 499258 162464 499494
rect 162144 492494 162464 499258
rect 162144 492258 162186 492494
rect 162422 492258 162464 492494
rect 162144 485494 162464 492258
rect 162144 485258 162186 485494
rect 162422 485258 162464 485494
rect 162144 478494 162464 485258
rect 162144 478258 162186 478494
rect 162422 478258 162464 478494
rect 162144 471494 162464 478258
rect 162144 471258 162186 471494
rect 162422 471258 162464 471494
rect 162144 464494 162464 471258
rect 162144 464258 162186 464494
rect 162422 464258 162464 464494
rect 162144 457494 162464 464258
rect 162144 457258 162186 457494
rect 162422 457258 162464 457494
rect 162144 450494 162464 457258
rect 162144 450258 162186 450494
rect 162422 450258 162464 450494
rect 162144 443494 162464 450258
rect 162144 443258 162186 443494
rect 162422 443258 162464 443494
rect 162144 436494 162464 443258
rect 162144 436258 162186 436494
rect 162422 436258 162464 436494
rect 162144 429494 162464 436258
rect 162144 429258 162186 429494
rect 162422 429258 162464 429494
rect 162144 422494 162464 429258
rect 162144 422258 162186 422494
rect 162422 422258 162464 422494
rect 162144 415494 162464 422258
rect 162144 415258 162186 415494
rect 162422 415258 162464 415494
rect 162144 408494 162464 415258
rect 162144 408258 162186 408494
rect 162422 408258 162464 408494
rect 162144 401494 162464 408258
rect 162144 401258 162186 401494
rect 162422 401258 162464 401494
rect 162144 394494 162464 401258
rect 162144 394258 162186 394494
rect 162422 394258 162464 394494
rect 162144 387494 162464 394258
rect 162144 387258 162186 387494
rect 162422 387258 162464 387494
rect 162144 380494 162464 387258
rect 162144 380258 162186 380494
rect 162422 380258 162464 380494
rect 162144 373494 162464 380258
rect 162144 373258 162186 373494
rect 162422 373258 162464 373494
rect 162144 366494 162464 373258
rect 162144 366258 162186 366494
rect 162422 366258 162464 366494
rect 162144 359494 162464 366258
rect 162144 359258 162186 359494
rect 162422 359258 162464 359494
rect 162144 352494 162464 359258
rect 162144 352258 162186 352494
rect 162422 352258 162464 352494
rect 162144 345494 162464 352258
rect 162144 345258 162186 345494
rect 162422 345258 162464 345494
rect 162144 338494 162464 345258
rect 162144 338258 162186 338494
rect 162422 338258 162464 338494
rect 162144 331494 162464 338258
rect 162144 331258 162186 331494
rect 162422 331258 162464 331494
rect 162144 324494 162464 331258
rect 162144 324258 162186 324494
rect 162422 324258 162464 324494
rect 162144 317494 162464 324258
rect 162144 317258 162186 317494
rect 162422 317258 162464 317494
rect 162144 310494 162464 317258
rect 162144 310258 162186 310494
rect 162422 310258 162464 310494
rect 162144 303494 162464 310258
rect 162144 303258 162186 303494
rect 162422 303258 162464 303494
rect 162144 296494 162464 303258
rect 162144 296258 162186 296494
rect 162422 296258 162464 296494
rect 162144 289494 162464 296258
rect 162144 289258 162186 289494
rect 162422 289258 162464 289494
rect 162144 282494 162464 289258
rect 162144 282258 162186 282494
rect 162422 282258 162464 282494
rect 162144 275494 162464 282258
rect 162144 275258 162186 275494
rect 162422 275258 162464 275494
rect 162144 268494 162464 275258
rect 162144 268258 162186 268494
rect 162422 268258 162464 268494
rect 162144 261494 162464 268258
rect 162144 261258 162186 261494
rect 162422 261258 162464 261494
rect 162144 254494 162464 261258
rect 162144 254258 162186 254494
rect 162422 254258 162464 254494
rect 162144 247494 162464 254258
rect 162144 247258 162186 247494
rect 162422 247258 162464 247494
rect 162144 240494 162464 247258
rect 162144 240258 162186 240494
rect 162422 240258 162464 240494
rect 162144 233494 162464 240258
rect 162144 233258 162186 233494
rect 162422 233258 162464 233494
rect 162144 226494 162464 233258
rect 162144 226258 162186 226494
rect 162422 226258 162464 226494
rect 162144 219494 162464 226258
rect 162144 219258 162186 219494
rect 162422 219258 162464 219494
rect 162144 212494 162464 219258
rect 162144 212258 162186 212494
rect 162422 212258 162464 212494
rect 162144 205494 162464 212258
rect 162144 205258 162186 205494
rect 162422 205258 162464 205494
rect 162144 198494 162464 205258
rect 162144 198258 162186 198494
rect 162422 198258 162464 198494
rect 162144 191494 162464 198258
rect 162144 191258 162186 191494
rect 162422 191258 162464 191494
rect 162144 184494 162464 191258
rect 162144 184258 162186 184494
rect 162422 184258 162464 184494
rect 162144 177494 162464 184258
rect 162144 177258 162186 177494
rect 162422 177258 162464 177494
rect 162144 170494 162464 177258
rect 162144 170258 162186 170494
rect 162422 170258 162464 170494
rect 162144 163494 162464 170258
rect 162144 163258 162186 163494
rect 162422 163258 162464 163494
rect 162144 156494 162464 163258
rect 162144 156258 162186 156494
rect 162422 156258 162464 156494
rect 162144 149494 162464 156258
rect 162144 149258 162186 149494
rect 162422 149258 162464 149494
rect 162144 142494 162464 149258
rect 162144 142258 162186 142494
rect 162422 142258 162464 142494
rect 162144 135494 162464 142258
rect 162144 135258 162186 135494
rect 162422 135258 162464 135494
rect 162144 128494 162464 135258
rect 162144 128258 162186 128494
rect 162422 128258 162464 128494
rect 162144 121494 162464 128258
rect 162144 121258 162186 121494
rect 162422 121258 162464 121494
rect 162144 114494 162464 121258
rect 162144 114258 162186 114494
rect 162422 114258 162464 114494
rect 162144 107494 162464 114258
rect 162144 107258 162186 107494
rect 162422 107258 162464 107494
rect 162144 100494 162464 107258
rect 162144 100258 162186 100494
rect 162422 100258 162464 100494
rect 162144 93494 162464 100258
rect 162144 93258 162186 93494
rect 162422 93258 162464 93494
rect 162144 86494 162464 93258
rect 162144 86258 162186 86494
rect 162422 86258 162464 86494
rect 162144 79494 162464 86258
rect 162144 79258 162186 79494
rect 162422 79258 162464 79494
rect 162144 72494 162464 79258
rect 162144 72258 162186 72494
rect 162422 72258 162464 72494
rect 162144 65494 162464 72258
rect 162144 65258 162186 65494
rect 162422 65258 162464 65494
rect 162144 58494 162464 65258
rect 162144 58258 162186 58494
rect 162422 58258 162464 58494
rect 162144 51494 162464 58258
rect 162144 51258 162186 51494
rect 162422 51258 162464 51494
rect 162144 44494 162464 51258
rect 162144 44258 162186 44494
rect 162422 44258 162464 44494
rect 162144 37494 162464 44258
rect 162144 37258 162186 37494
rect 162422 37258 162464 37494
rect 162144 30494 162464 37258
rect 162144 30258 162186 30494
rect 162422 30258 162464 30494
rect 162144 23494 162464 30258
rect 162144 23258 162186 23494
rect 162422 23258 162464 23494
rect 162144 16494 162464 23258
rect 162144 16258 162186 16494
rect 162422 16258 162464 16494
rect 162144 9494 162464 16258
rect 162144 9258 162186 9494
rect 162422 9258 162464 9494
rect 162144 2494 162464 9258
rect 162144 2258 162186 2494
rect 162422 2258 162464 2494
rect 162144 -746 162464 2258
rect 162144 -982 162186 -746
rect 162422 -982 162464 -746
rect 162144 -1066 162464 -982
rect 162144 -1302 162186 -1066
rect 162422 -1302 162464 -1066
rect 162144 -2294 162464 -1302
rect 163876 706198 164196 706230
rect 163876 705962 163918 706198
rect 164154 705962 164196 706198
rect 163876 705878 164196 705962
rect 163876 705642 163918 705878
rect 164154 705642 164196 705878
rect 163876 696434 164196 705642
rect 163876 696198 163918 696434
rect 164154 696198 164196 696434
rect 163876 689434 164196 696198
rect 163876 689198 163918 689434
rect 164154 689198 164196 689434
rect 163876 682434 164196 689198
rect 163876 682198 163918 682434
rect 164154 682198 164196 682434
rect 163876 675434 164196 682198
rect 163876 675198 163918 675434
rect 164154 675198 164196 675434
rect 163876 668434 164196 675198
rect 163876 668198 163918 668434
rect 164154 668198 164196 668434
rect 163876 661434 164196 668198
rect 163876 661198 163918 661434
rect 164154 661198 164196 661434
rect 163876 654434 164196 661198
rect 163876 654198 163918 654434
rect 164154 654198 164196 654434
rect 163876 647434 164196 654198
rect 163876 647198 163918 647434
rect 164154 647198 164196 647434
rect 163876 640434 164196 647198
rect 163876 640198 163918 640434
rect 164154 640198 164196 640434
rect 163876 633434 164196 640198
rect 163876 633198 163918 633434
rect 164154 633198 164196 633434
rect 163876 626434 164196 633198
rect 163876 626198 163918 626434
rect 164154 626198 164196 626434
rect 163876 619434 164196 626198
rect 163876 619198 163918 619434
rect 164154 619198 164196 619434
rect 163876 612434 164196 619198
rect 163876 612198 163918 612434
rect 164154 612198 164196 612434
rect 163876 605434 164196 612198
rect 163876 605198 163918 605434
rect 164154 605198 164196 605434
rect 163876 598434 164196 605198
rect 163876 598198 163918 598434
rect 164154 598198 164196 598434
rect 163876 591434 164196 598198
rect 163876 591198 163918 591434
rect 164154 591198 164196 591434
rect 163876 584434 164196 591198
rect 163876 584198 163918 584434
rect 164154 584198 164196 584434
rect 163876 577434 164196 584198
rect 163876 577198 163918 577434
rect 164154 577198 164196 577434
rect 163876 570434 164196 577198
rect 163876 570198 163918 570434
rect 164154 570198 164196 570434
rect 163876 563434 164196 570198
rect 163876 563198 163918 563434
rect 164154 563198 164196 563434
rect 163876 556434 164196 563198
rect 163876 556198 163918 556434
rect 164154 556198 164196 556434
rect 163876 549434 164196 556198
rect 163876 549198 163918 549434
rect 164154 549198 164196 549434
rect 163876 542434 164196 549198
rect 163876 542198 163918 542434
rect 164154 542198 164196 542434
rect 163876 535434 164196 542198
rect 163876 535198 163918 535434
rect 164154 535198 164196 535434
rect 163876 528434 164196 535198
rect 163876 528198 163918 528434
rect 164154 528198 164196 528434
rect 163876 521434 164196 528198
rect 163876 521198 163918 521434
rect 164154 521198 164196 521434
rect 163876 514434 164196 521198
rect 163876 514198 163918 514434
rect 164154 514198 164196 514434
rect 163876 507434 164196 514198
rect 163876 507198 163918 507434
rect 164154 507198 164196 507434
rect 163876 500434 164196 507198
rect 163876 500198 163918 500434
rect 164154 500198 164196 500434
rect 163876 493434 164196 500198
rect 163876 493198 163918 493434
rect 164154 493198 164196 493434
rect 163876 486434 164196 493198
rect 163876 486198 163918 486434
rect 164154 486198 164196 486434
rect 163876 479434 164196 486198
rect 163876 479198 163918 479434
rect 164154 479198 164196 479434
rect 163876 472434 164196 479198
rect 163876 472198 163918 472434
rect 164154 472198 164196 472434
rect 163876 465434 164196 472198
rect 163876 465198 163918 465434
rect 164154 465198 164196 465434
rect 163876 458434 164196 465198
rect 163876 458198 163918 458434
rect 164154 458198 164196 458434
rect 163876 451434 164196 458198
rect 163876 451198 163918 451434
rect 164154 451198 164196 451434
rect 163876 444434 164196 451198
rect 163876 444198 163918 444434
rect 164154 444198 164196 444434
rect 163876 437434 164196 444198
rect 163876 437198 163918 437434
rect 164154 437198 164196 437434
rect 163876 430434 164196 437198
rect 163876 430198 163918 430434
rect 164154 430198 164196 430434
rect 163876 423434 164196 430198
rect 163876 423198 163918 423434
rect 164154 423198 164196 423434
rect 163876 416434 164196 423198
rect 163876 416198 163918 416434
rect 164154 416198 164196 416434
rect 163876 409434 164196 416198
rect 163876 409198 163918 409434
rect 164154 409198 164196 409434
rect 163876 402434 164196 409198
rect 163876 402198 163918 402434
rect 164154 402198 164196 402434
rect 163876 395434 164196 402198
rect 163876 395198 163918 395434
rect 164154 395198 164196 395434
rect 163876 388434 164196 395198
rect 163876 388198 163918 388434
rect 164154 388198 164196 388434
rect 163876 381434 164196 388198
rect 163876 381198 163918 381434
rect 164154 381198 164196 381434
rect 163876 374434 164196 381198
rect 163876 374198 163918 374434
rect 164154 374198 164196 374434
rect 163876 367434 164196 374198
rect 163876 367198 163918 367434
rect 164154 367198 164196 367434
rect 163876 360434 164196 367198
rect 163876 360198 163918 360434
rect 164154 360198 164196 360434
rect 163876 353434 164196 360198
rect 163876 353198 163918 353434
rect 164154 353198 164196 353434
rect 163876 346434 164196 353198
rect 163876 346198 163918 346434
rect 164154 346198 164196 346434
rect 163876 339434 164196 346198
rect 163876 339198 163918 339434
rect 164154 339198 164196 339434
rect 163876 332434 164196 339198
rect 163876 332198 163918 332434
rect 164154 332198 164196 332434
rect 163876 325434 164196 332198
rect 163876 325198 163918 325434
rect 164154 325198 164196 325434
rect 163876 318434 164196 325198
rect 163876 318198 163918 318434
rect 164154 318198 164196 318434
rect 163876 311434 164196 318198
rect 163876 311198 163918 311434
rect 164154 311198 164196 311434
rect 163876 304434 164196 311198
rect 163876 304198 163918 304434
rect 164154 304198 164196 304434
rect 163876 297434 164196 304198
rect 163876 297198 163918 297434
rect 164154 297198 164196 297434
rect 163876 290434 164196 297198
rect 163876 290198 163918 290434
rect 164154 290198 164196 290434
rect 163876 283434 164196 290198
rect 163876 283198 163918 283434
rect 164154 283198 164196 283434
rect 163876 276434 164196 283198
rect 163876 276198 163918 276434
rect 164154 276198 164196 276434
rect 163876 269434 164196 276198
rect 163876 269198 163918 269434
rect 164154 269198 164196 269434
rect 163876 262434 164196 269198
rect 163876 262198 163918 262434
rect 164154 262198 164196 262434
rect 163876 255434 164196 262198
rect 163876 255198 163918 255434
rect 164154 255198 164196 255434
rect 163876 248434 164196 255198
rect 163876 248198 163918 248434
rect 164154 248198 164196 248434
rect 163876 241434 164196 248198
rect 163876 241198 163918 241434
rect 164154 241198 164196 241434
rect 163876 234434 164196 241198
rect 163876 234198 163918 234434
rect 164154 234198 164196 234434
rect 163876 227434 164196 234198
rect 163876 227198 163918 227434
rect 164154 227198 164196 227434
rect 163876 220434 164196 227198
rect 163876 220198 163918 220434
rect 164154 220198 164196 220434
rect 163876 213434 164196 220198
rect 163876 213198 163918 213434
rect 164154 213198 164196 213434
rect 163876 206434 164196 213198
rect 163876 206198 163918 206434
rect 164154 206198 164196 206434
rect 163876 199434 164196 206198
rect 163876 199198 163918 199434
rect 164154 199198 164196 199434
rect 163876 192434 164196 199198
rect 163876 192198 163918 192434
rect 164154 192198 164196 192434
rect 163876 185434 164196 192198
rect 163876 185198 163918 185434
rect 164154 185198 164196 185434
rect 163876 178434 164196 185198
rect 163876 178198 163918 178434
rect 164154 178198 164196 178434
rect 163876 171434 164196 178198
rect 163876 171198 163918 171434
rect 164154 171198 164196 171434
rect 163876 164434 164196 171198
rect 163876 164198 163918 164434
rect 164154 164198 164196 164434
rect 163876 157434 164196 164198
rect 163876 157198 163918 157434
rect 164154 157198 164196 157434
rect 163876 150434 164196 157198
rect 163876 150198 163918 150434
rect 164154 150198 164196 150434
rect 163876 143434 164196 150198
rect 163876 143198 163918 143434
rect 164154 143198 164196 143434
rect 163876 136434 164196 143198
rect 163876 136198 163918 136434
rect 164154 136198 164196 136434
rect 163876 129434 164196 136198
rect 163876 129198 163918 129434
rect 164154 129198 164196 129434
rect 163876 122434 164196 129198
rect 163876 122198 163918 122434
rect 164154 122198 164196 122434
rect 163876 115434 164196 122198
rect 163876 115198 163918 115434
rect 164154 115198 164196 115434
rect 163876 108434 164196 115198
rect 163876 108198 163918 108434
rect 164154 108198 164196 108434
rect 163876 101434 164196 108198
rect 163876 101198 163918 101434
rect 164154 101198 164196 101434
rect 163876 94434 164196 101198
rect 163876 94198 163918 94434
rect 164154 94198 164196 94434
rect 163876 87434 164196 94198
rect 163876 87198 163918 87434
rect 164154 87198 164196 87434
rect 163876 80434 164196 87198
rect 163876 80198 163918 80434
rect 164154 80198 164196 80434
rect 163876 73434 164196 80198
rect 163876 73198 163918 73434
rect 164154 73198 164196 73434
rect 163876 66434 164196 73198
rect 163876 66198 163918 66434
rect 164154 66198 164196 66434
rect 163876 59434 164196 66198
rect 163876 59198 163918 59434
rect 164154 59198 164196 59434
rect 163876 52434 164196 59198
rect 163876 52198 163918 52434
rect 164154 52198 164196 52434
rect 163876 45434 164196 52198
rect 163876 45198 163918 45434
rect 164154 45198 164196 45434
rect 163876 38434 164196 45198
rect 163876 38198 163918 38434
rect 164154 38198 164196 38434
rect 163876 31434 164196 38198
rect 163876 31198 163918 31434
rect 164154 31198 164196 31434
rect 163876 24434 164196 31198
rect 163876 24198 163918 24434
rect 164154 24198 164196 24434
rect 163876 17434 164196 24198
rect 163876 17198 163918 17434
rect 164154 17198 164196 17434
rect 163876 10434 164196 17198
rect 163876 10198 163918 10434
rect 164154 10198 164196 10434
rect 163876 3434 164196 10198
rect 163876 3198 163918 3434
rect 164154 3198 164196 3434
rect 163876 -1706 164196 3198
rect 163876 -1942 163918 -1706
rect 164154 -1942 164196 -1706
rect 163876 -2026 164196 -1942
rect 163876 -2262 163918 -2026
rect 164154 -2262 164196 -2026
rect 163876 -2294 164196 -2262
rect 169144 705238 169464 706230
rect 169144 705002 169186 705238
rect 169422 705002 169464 705238
rect 169144 704918 169464 705002
rect 169144 704682 169186 704918
rect 169422 704682 169464 704918
rect 169144 695494 169464 704682
rect 169144 695258 169186 695494
rect 169422 695258 169464 695494
rect 169144 688494 169464 695258
rect 169144 688258 169186 688494
rect 169422 688258 169464 688494
rect 169144 681494 169464 688258
rect 169144 681258 169186 681494
rect 169422 681258 169464 681494
rect 169144 674494 169464 681258
rect 169144 674258 169186 674494
rect 169422 674258 169464 674494
rect 169144 667494 169464 674258
rect 169144 667258 169186 667494
rect 169422 667258 169464 667494
rect 169144 660494 169464 667258
rect 169144 660258 169186 660494
rect 169422 660258 169464 660494
rect 169144 653494 169464 660258
rect 169144 653258 169186 653494
rect 169422 653258 169464 653494
rect 169144 646494 169464 653258
rect 169144 646258 169186 646494
rect 169422 646258 169464 646494
rect 169144 639494 169464 646258
rect 169144 639258 169186 639494
rect 169422 639258 169464 639494
rect 169144 632494 169464 639258
rect 169144 632258 169186 632494
rect 169422 632258 169464 632494
rect 169144 625494 169464 632258
rect 169144 625258 169186 625494
rect 169422 625258 169464 625494
rect 169144 618494 169464 625258
rect 169144 618258 169186 618494
rect 169422 618258 169464 618494
rect 169144 611494 169464 618258
rect 169144 611258 169186 611494
rect 169422 611258 169464 611494
rect 169144 604494 169464 611258
rect 169144 604258 169186 604494
rect 169422 604258 169464 604494
rect 169144 597494 169464 604258
rect 169144 597258 169186 597494
rect 169422 597258 169464 597494
rect 169144 590494 169464 597258
rect 169144 590258 169186 590494
rect 169422 590258 169464 590494
rect 169144 583494 169464 590258
rect 169144 583258 169186 583494
rect 169422 583258 169464 583494
rect 169144 576494 169464 583258
rect 169144 576258 169186 576494
rect 169422 576258 169464 576494
rect 169144 569494 169464 576258
rect 169144 569258 169186 569494
rect 169422 569258 169464 569494
rect 169144 562494 169464 569258
rect 169144 562258 169186 562494
rect 169422 562258 169464 562494
rect 169144 555494 169464 562258
rect 169144 555258 169186 555494
rect 169422 555258 169464 555494
rect 169144 548494 169464 555258
rect 169144 548258 169186 548494
rect 169422 548258 169464 548494
rect 169144 541494 169464 548258
rect 169144 541258 169186 541494
rect 169422 541258 169464 541494
rect 169144 534494 169464 541258
rect 169144 534258 169186 534494
rect 169422 534258 169464 534494
rect 169144 527494 169464 534258
rect 169144 527258 169186 527494
rect 169422 527258 169464 527494
rect 169144 520494 169464 527258
rect 169144 520258 169186 520494
rect 169422 520258 169464 520494
rect 169144 513494 169464 520258
rect 169144 513258 169186 513494
rect 169422 513258 169464 513494
rect 169144 506494 169464 513258
rect 169144 506258 169186 506494
rect 169422 506258 169464 506494
rect 169144 499494 169464 506258
rect 169144 499258 169186 499494
rect 169422 499258 169464 499494
rect 169144 492494 169464 499258
rect 169144 492258 169186 492494
rect 169422 492258 169464 492494
rect 169144 485494 169464 492258
rect 169144 485258 169186 485494
rect 169422 485258 169464 485494
rect 169144 478494 169464 485258
rect 169144 478258 169186 478494
rect 169422 478258 169464 478494
rect 169144 471494 169464 478258
rect 169144 471258 169186 471494
rect 169422 471258 169464 471494
rect 169144 464494 169464 471258
rect 169144 464258 169186 464494
rect 169422 464258 169464 464494
rect 169144 457494 169464 464258
rect 169144 457258 169186 457494
rect 169422 457258 169464 457494
rect 169144 450494 169464 457258
rect 169144 450258 169186 450494
rect 169422 450258 169464 450494
rect 169144 443494 169464 450258
rect 169144 443258 169186 443494
rect 169422 443258 169464 443494
rect 169144 436494 169464 443258
rect 169144 436258 169186 436494
rect 169422 436258 169464 436494
rect 169144 429494 169464 436258
rect 169144 429258 169186 429494
rect 169422 429258 169464 429494
rect 169144 422494 169464 429258
rect 169144 422258 169186 422494
rect 169422 422258 169464 422494
rect 169144 415494 169464 422258
rect 169144 415258 169186 415494
rect 169422 415258 169464 415494
rect 169144 408494 169464 415258
rect 169144 408258 169186 408494
rect 169422 408258 169464 408494
rect 169144 401494 169464 408258
rect 169144 401258 169186 401494
rect 169422 401258 169464 401494
rect 169144 394494 169464 401258
rect 169144 394258 169186 394494
rect 169422 394258 169464 394494
rect 169144 387494 169464 394258
rect 169144 387258 169186 387494
rect 169422 387258 169464 387494
rect 169144 380494 169464 387258
rect 169144 380258 169186 380494
rect 169422 380258 169464 380494
rect 169144 373494 169464 380258
rect 169144 373258 169186 373494
rect 169422 373258 169464 373494
rect 169144 366494 169464 373258
rect 169144 366258 169186 366494
rect 169422 366258 169464 366494
rect 169144 359494 169464 366258
rect 169144 359258 169186 359494
rect 169422 359258 169464 359494
rect 169144 352494 169464 359258
rect 169144 352258 169186 352494
rect 169422 352258 169464 352494
rect 169144 345494 169464 352258
rect 169144 345258 169186 345494
rect 169422 345258 169464 345494
rect 169144 338494 169464 345258
rect 169144 338258 169186 338494
rect 169422 338258 169464 338494
rect 169144 331494 169464 338258
rect 169144 331258 169186 331494
rect 169422 331258 169464 331494
rect 169144 324494 169464 331258
rect 169144 324258 169186 324494
rect 169422 324258 169464 324494
rect 169144 317494 169464 324258
rect 169144 317258 169186 317494
rect 169422 317258 169464 317494
rect 169144 310494 169464 317258
rect 169144 310258 169186 310494
rect 169422 310258 169464 310494
rect 169144 303494 169464 310258
rect 169144 303258 169186 303494
rect 169422 303258 169464 303494
rect 169144 296494 169464 303258
rect 169144 296258 169186 296494
rect 169422 296258 169464 296494
rect 169144 289494 169464 296258
rect 169144 289258 169186 289494
rect 169422 289258 169464 289494
rect 169144 282494 169464 289258
rect 169144 282258 169186 282494
rect 169422 282258 169464 282494
rect 169144 275494 169464 282258
rect 169144 275258 169186 275494
rect 169422 275258 169464 275494
rect 169144 268494 169464 275258
rect 169144 268258 169186 268494
rect 169422 268258 169464 268494
rect 169144 261494 169464 268258
rect 169144 261258 169186 261494
rect 169422 261258 169464 261494
rect 169144 254494 169464 261258
rect 169144 254258 169186 254494
rect 169422 254258 169464 254494
rect 169144 247494 169464 254258
rect 169144 247258 169186 247494
rect 169422 247258 169464 247494
rect 169144 240494 169464 247258
rect 169144 240258 169186 240494
rect 169422 240258 169464 240494
rect 169144 233494 169464 240258
rect 169144 233258 169186 233494
rect 169422 233258 169464 233494
rect 169144 226494 169464 233258
rect 169144 226258 169186 226494
rect 169422 226258 169464 226494
rect 169144 219494 169464 226258
rect 169144 219258 169186 219494
rect 169422 219258 169464 219494
rect 169144 212494 169464 219258
rect 169144 212258 169186 212494
rect 169422 212258 169464 212494
rect 169144 205494 169464 212258
rect 169144 205258 169186 205494
rect 169422 205258 169464 205494
rect 169144 198494 169464 205258
rect 169144 198258 169186 198494
rect 169422 198258 169464 198494
rect 169144 191494 169464 198258
rect 169144 191258 169186 191494
rect 169422 191258 169464 191494
rect 169144 184494 169464 191258
rect 169144 184258 169186 184494
rect 169422 184258 169464 184494
rect 169144 177494 169464 184258
rect 169144 177258 169186 177494
rect 169422 177258 169464 177494
rect 169144 170494 169464 177258
rect 169144 170258 169186 170494
rect 169422 170258 169464 170494
rect 169144 163494 169464 170258
rect 169144 163258 169186 163494
rect 169422 163258 169464 163494
rect 169144 156494 169464 163258
rect 169144 156258 169186 156494
rect 169422 156258 169464 156494
rect 169144 149494 169464 156258
rect 169144 149258 169186 149494
rect 169422 149258 169464 149494
rect 169144 142494 169464 149258
rect 169144 142258 169186 142494
rect 169422 142258 169464 142494
rect 169144 135494 169464 142258
rect 169144 135258 169186 135494
rect 169422 135258 169464 135494
rect 169144 128494 169464 135258
rect 169144 128258 169186 128494
rect 169422 128258 169464 128494
rect 169144 121494 169464 128258
rect 169144 121258 169186 121494
rect 169422 121258 169464 121494
rect 169144 114494 169464 121258
rect 169144 114258 169186 114494
rect 169422 114258 169464 114494
rect 169144 107494 169464 114258
rect 169144 107258 169186 107494
rect 169422 107258 169464 107494
rect 169144 100494 169464 107258
rect 169144 100258 169186 100494
rect 169422 100258 169464 100494
rect 169144 93494 169464 100258
rect 169144 93258 169186 93494
rect 169422 93258 169464 93494
rect 169144 86494 169464 93258
rect 169144 86258 169186 86494
rect 169422 86258 169464 86494
rect 169144 79494 169464 86258
rect 169144 79258 169186 79494
rect 169422 79258 169464 79494
rect 169144 72494 169464 79258
rect 169144 72258 169186 72494
rect 169422 72258 169464 72494
rect 169144 65494 169464 72258
rect 169144 65258 169186 65494
rect 169422 65258 169464 65494
rect 169144 58494 169464 65258
rect 169144 58258 169186 58494
rect 169422 58258 169464 58494
rect 169144 51494 169464 58258
rect 169144 51258 169186 51494
rect 169422 51258 169464 51494
rect 169144 44494 169464 51258
rect 169144 44258 169186 44494
rect 169422 44258 169464 44494
rect 169144 37494 169464 44258
rect 169144 37258 169186 37494
rect 169422 37258 169464 37494
rect 169144 30494 169464 37258
rect 169144 30258 169186 30494
rect 169422 30258 169464 30494
rect 169144 23494 169464 30258
rect 169144 23258 169186 23494
rect 169422 23258 169464 23494
rect 169144 16494 169464 23258
rect 169144 16258 169186 16494
rect 169422 16258 169464 16494
rect 169144 9494 169464 16258
rect 169144 9258 169186 9494
rect 169422 9258 169464 9494
rect 169144 2494 169464 9258
rect 169144 2258 169186 2494
rect 169422 2258 169464 2494
rect 169144 -746 169464 2258
rect 169144 -982 169186 -746
rect 169422 -982 169464 -746
rect 169144 -1066 169464 -982
rect 169144 -1302 169186 -1066
rect 169422 -1302 169464 -1066
rect 169144 -2294 169464 -1302
rect 170876 706198 171196 706230
rect 170876 705962 170918 706198
rect 171154 705962 171196 706198
rect 170876 705878 171196 705962
rect 170876 705642 170918 705878
rect 171154 705642 171196 705878
rect 170876 696434 171196 705642
rect 170876 696198 170918 696434
rect 171154 696198 171196 696434
rect 170876 689434 171196 696198
rect 170876 689198 170918 689434
rect 171154 689198 171196 689434
rect 170876 682434 171196 689198
rect 170876 682198 170918 682434
rect 171154 682198 171196 682434
rect 170876 675434 171196 682198
rect 170876 675198 170918 675434
rect 171154 675198 171196 675434
rect 170876 668434 171196 675198
rect 170876 668198 170918 668434
rect 171154 668198 171196 668434
rect 170876 661434 171196 668198
rect 170876 661198 170918 661434
rect 171154 661198 171196 661434
rect 170876 654434 171196 661198
rect 170876 654198 170918 654434
rect 171154 654198 171196 654434
rect 170876 647434 171196 654198
rect 170876 647198 170918 647434
rect 171154 647198 171196 647434
rect 170876 640434 171196 647198
rect 170876 640198 170918 640434
rect 171154 640198 171196 640434
rect 170876 633434 171196 640198
rect 170876 633198 170918 633434
rect 171154 633198 171196 633434
rect 170876 626434 171196 633198
rect 170876 626198 170918 626434
rect 171154 626198 171196 626434
rect 170876 619434 171196 626198
rect 170876 619198 170918 619434
rect 171154 619198 171196 619434
rect 170876 612434 171196 619198
rect 170876 612198 170918 612434
rect 171154 612198 171196 612434
rect 170876 605434 171196 612198
rect 170876 605198 170918 605434
rect 171154 605198 171196 605434
rect 170876 598434 171196 605198
rect 170876 598198 170918 598434
rect 171154 598198 171196 598434
rect 170876 591434 171196 598198
rect 170876 591198 170918 591434
rect 171154 591198 171196 591434
rect 170876 584434 171196 591198
rect 170876 584198 170918 584434
rect 171154 584198 171196 584434
rect 170876 577434 171196 584198
rect 170876 577198 170918 577434
rect 171154 577198 171196 577434
rect 170876 570434 171196 577198
rect 170876 570198 170918 570434
rect 171154 570198 171196 570434
rect 170876 563434 171196 570198
rect 170876 563198 170918 563434
rect 171154 563198 171196 563434
rect 170876 556434 171196 563198
rect 170876 556198 170918 556434
rect 171154 556198 171196 556434
rect 170876 549434 171196 556198
rect 170876 549198 170918 549434
rect 171154 549198 171196 549434
rect 170876 542434 171196 549198
rect 170876 542198 170918 542434
rect 171154 542198 171196 542434
rect 170876 535434 171196 542198
rect 170876 535198 170918 535434
rect 171154 535198 171196 535434
rect 170876 528434 171196 535198
rect 170876 528198 170918 528434
rect 171154 528198 171196 528434
rect 170876 521434 171196 528198
rect 170876 521198 170918 521434
rect 171154 521198 171196 521434
rect 170876 514434 171196 521198
rect 170876 514198 170918 514434
rect 171154 514198 171196 514434
rect 170876 507434 171196 514198
rect 170876 507198 170918 507434
rect 171154 507198 171196 507434
rect 170876 500434 171196 507198
rect 170876 500198 170918 500434
rect 171154 500198 171196 500434
rect 170876 493434 171196 500198
rect 170876 493198 170918 493434
rect 171154 493198 171196 493434
rect 170876 486434 171196 493198
rect 170876 486198 170918 486434
rect 171154 486198 171196 486434
rect 170876 479434 171196 486198
rect 170876 479198 170918 479434
rect 171154 479198 171196 479434
rect 170876 472434 171196 479198
rect 170876 472198 170918 472434
rect 171154 472198 171196 472434
rect 170876 465434 171196 472198
rect 170876 465198 170918 465434
rect 171154 465198 171196 465434
rect 170876 458434 171196 465198
rect 170876 458198 170918 458434
rect 171154 458198 171196 458434
rect 170876 451434 171196 458198
rect 170876 451198 170918 451434
rect 171154 451198 171196 451434
rect 170876 444434 171196 451198
rect 170876 444198 170918 444434
rect 171154 444198 171196 444434
rect 170876 437434 171196 444198
rect 170876 437198 170918 437434
rect 171154 437198 171196 437434
rect 170876 430434 171196 437198
rect 170876 430198 170918 430434
rect 171154 430198 171196 430434
rect 170876 423434 171196 430198
rect 170876 423198 170918 423434
rect 171154 423198 171196 423434
rect 170876 416434 171196 423198
rect 170876 416198 170918 416434
rect 171154 416198 171196 416434
rect 170876 409434 171196 416198
rect 170876 409198 170918 409434
rect 171154 409198 171196 409434
rect 170876 402434 171196 409198
rect 170876 402198 170918 402434
rect 171154 402198 171196 402434
rect 170876 395434 171196 402198
rect 170876 395198 170918 395434
rect 171154 395198 171196 395434
rect 170876 388434 171196 395198
rect 170876 388198 170918 388434
rect 171154 388198 171196 388434
rect 170876 381434 171196 388198
rect 170876 381198 170918 381434
rect 171154 381198 171196 381434
rect 170876 374434 171196 381198
rect 170876 374198 170918 374434
rect 171154 374198 171196 374434
rect 170876 367434 171196 374198
rect 170876 367198 170918 367434
rect 171154 367198 171196 367434
rect 170876 360434 171196 367198
rect 170876 360198 170918 360434
rect 171154 360198 171196 360434
rect 170876 353434 171196 360198
rect 170876 353198 170918 353434
rect 171154 353198 171196 353434
rect 170876 346434 171196 353198
rect 170876 346198 170918 346434
rect 171154 346198 171196 346434
rect 170876 339434 171196 346198
rect 170876 339198 170918 339434
rect 171154 339198 171196 339434
rect 170876 332434 171196 339198
rect 170876 332198 170918 332434
rect 171154 332198 171196 332434
rect 170876 325434 171196 332198
rect 170876 325198 170918 325434
rect 171154 325198 171196 325434
rect 170876 318434 171196 325198
rect 170876 318198 170918 318434
rect 171154 318198 171196 318434
rect 170876 311434 171196 318198
rect 170876 311198 170918 311434
rect 171154 311198 171196 311434
rect 170876 304434 171196 311198
rect 170876 304198 170918 304434
rect 171154 304198 171196 304434
rect 170876 297434 171196 304198
rect 170876 297198 170918 297434
rect 171154 297198 171196 297434
rect 170876 290434 171196 297198
rect 170876 290198 170918 290434
rect 171154 290198 171196 290434
rect 170876 283434 171196 290198
rect 170876 283198 170918 283434
rect 171154 283198 171196 283434
rect 170876 276434 171196 283198
rect 170876 276198 170918 276434
rect 171154 276198 171196 276434
rect 170876 269434 171196 276198
rect 170876 269198 170918 269434
rect 171154 269198 171196 269434
rect 170876 262434 171196 269198
rect 170876 262198 170918 262434
rect 171154 262198 171196 262434
rect 170876 255434 171196 262198
rect 170876 255198 170918 255434
rect 171154 255198 171196 255434
rect 170876 248434 171196 255198
rect 170876 248198 170918 248434
rect 171154 248198 171196 248434
rect 170876 241434 171196 248198
rect 170876 241198 170918 241434
rect 171154 241198 171196 241434
rect 170876 234434 171196 241198
rect 170876 234198 170918 234434
rect 171154 234198 171196 234434
rect 170876 227434 171196 234198
rect 170876 227198 170918 227434
rect 171154 227198 171196 227434
rect 170876 220434 171196 227198
rect 170876 220198 170918 220434
rect 171154 220198 171196 220434
rect 170876 213434 171196 220198
rect 170876 213198 170918 213434
rect 171154 213198 171196 213434
rect 170876 206434 171196 213198
rect 170876 206198 170918 206434
rect 171154 206198 171196 206434
rect 170876 199434 171196 206198
rect 170876 199198 170918 199434
rect 171154 199198 171196 199434
rect 170876 192434 171196 199198
rect 170876 192198 170918 192434
rect 171154 192198 171196 192434
rect 170876 185434 171196 192198
rect 170876 185198 170918 185434
rect 171154 185198 171196 185434
rect 170876 178434 171196 185198
rect 170876 178198 170918 178434
rect 171154 178198 171196 178434
rect 170876 171434 171196 178198
rect 170876 171198 170918 171434
rect 171154 171198 171196 171434
rect 170876 164434 171196 171198
rect 170876 164198 170918 164434
rect 171154 164198 171196 164434
rect 170876 157434 171196 164198
rect 170876 157198 170918 157434
rect 171154 157198 171196 157434
rect 170876 150434 171196 157198
rect 170876 150198 170918 150434
rect 171154 150198 171196 150434
rect 170876 143434 171196 150198
rect 170876 143198 170918 143434
rect 171154 143198 171196 143434
rect 170876 136434 171196 143198
rect 170876 136198 170918 136434
rect 171154 136198 171196 136434
rect 170876 129434 171196 136198
rect 170876 129198 170918 129434
rect 171154 129198 171196 129434
rect 170876 122434 171196 129198
rect 170876 122198 170918 122434
rect 171154 122198 171196 122434
rect 170876 115434 171196 122198
rect 170876 115198 170918 115434
rect 171154 115198 171196 115434
rect 170876 108434 171196 115198
rect 170876 108198 170918 108434
rect 171154 108198 171196 108434
rect 170876 101434 171196 108198
rect 170876 101198 170918 101434
rect 171154 101198 171196 101434
rect 170876 94434 171196 101198
rect 170876 94198 170918 94434
rect 171154 94198 171196 94434
rect 170876 87434 171196 94198
rect 170876 87198 170918 87434
rect 171154 87198 171196 87434
rect 170876 80434 171196 87198
rect 170876 80198 170918 80434
rect 171154 80198 171196 80434
rect 170876 73434 171196 80198
rect 170876 73198 170918 73434
rect 171154 73198 171196 73434
rect 170876 66434 171196 73198
rect 170876 66198 170918 66434
rect 171154 66198 171196 66434
rect 170876 59434 171196 66198
rect 170876 59198 170918 59434
rect 171154 59198 171196 59434
rect 170876 52434 171196 59198
rect 170876 52198 170918 52434
rect 171154 52198 171196 52434
rect 170876 45434 171196 52198
rect 170876 45198 170918 45434
rect 171154 45198 171196 45434
rect 170876 38434 171196 45198
rect 170876 38198 170918 38434
rect 171154 38198 171196 38434
rect 170876 31434 171196 38198
rect 170876 31198 170918 31434
rect 171154 31198 171196 31434
rect 170876 24434 171196 31198
rect 170876 24198 170918 24434
rect 171154 24198 171196 24434
rect 170876 17434 171196 24198
rect 170876 17198 170918 17434
rect 171154 17198 171196 17434
rect 170876 10434 171196 17198
rect 170876 10198 170918 10434
rect 171154 10198 171196 10434
rect 170876 3434 171196 10198
rect 170876 3198 170918 3434
rect 171154 3198 171196 3434
rect 170876 -1706 171196 3198
rect 170876 -1942 170918 -1706
rect 171154 -1942 171196 -1706
rect 170876 -2026 171196 -1942
rect 170876 -2262 170918 -2026
rect 171154 -2262 171196 -2026
rect 170876 -2294 171196 -2262
rect 176144 705238 176464 706230
rect 176144 705002 176186 705238
rect 176422 705002 176464 705238
rect 176144 704918 176464 705002
rect 176144 704682 176186 704918
rect 176422 704682 176464 704918
rect 176144 695494 176464 704682
rect 176144 695258 176186 695494
rect 176422 695258 176464 695494
rect 176144 688494 176464 695258
rect 176144 688258 176186 688494
rect 176422 688258 176464 688494
rect 176144 681494 176464 688258
rect 176144 681258 176186 681494
rect 176422 681258 176464 681494
rect 176144 674494 176464 681258
rect 176144 674258 176186 674494
rect 176422 674258 176464 674494
rect 176144 667494 176464 674258
rect 176144 667258 176186 667494
rect 176422 667258 176464 667494
rect 176144 660494 176464 667258
rect 176144 660258 176186 660494
rect 176422 660258 176464 660494
rect 176144 653494 176464 660258
rect 176144 653258 176186 653494
rect 176422 653258 176464 653494
rect 176144 646494 176464 653258
rect 176144 646258 176186 646494
rect 176422 646258 176464 646494
rect 176144 639494 176464 646258
rect 176144 639258 176186 639494
rect 176422 639258 176464 639494
rect 176144 632494 176464 639258
rect 176144 632258 176186 632494
rect 176422 632258 176464 632494
rect 176144 625494 176464 632258
rect 176144 625258 176186 625494
rect 176422 625258 176464 625494
rect 176144 618494 176464 625258
rect 176144 618258 176186 618494
rect 176422 618258 176464 618494
rect 176144 611494 176464 618258
rect 176144 611258 176186 611494
rect 176422 611258 176464 611494
rect 176144 604494 176464 611258
rect 176144 604258 176186 604494
rect 176422 604258 176464 604494
rect 176144 597494 176464 604258
rect 176144 597258 176186 597494
rect 176422 597258 176464 597494
rect 176144 590494 176464 597258
rect 176144 590258 176186 590494
rect 176422 590258 176464 590494
rect 176144 583494 176464 590258
rect 176144 583258 176186 583494
rect 176422 583258 176464 583494
rect 176144 576494 176464 583258
rect 176144 576258 176186 576494
rect 176422 576258 176464 576494
rect 176144 569494 176464 576258
rect 176144 569258 176186 569494
rect 176422 569258 176464 569494
rect 176144 562494 176464 569258
rect 176144 562258 176186 562494
rect 176422 562258 176464 562494
rect 176144 555494 176464 562258
rect 176144 555258 176186 555494
rect 176422 555258 176464 555494
rect 176144 548494 176464 555258
rect 176144 548258 176186 548494
rect 176422 548258 176464 548494
rect 176144 541494 176464 548258
rect 176144 541258 176186 541494
rect 176422 541258 176464 541494
rect 176144 534494 176464 541258
rect 176144 534258 176186 534494
rect 176422 534258 176464 534494
rect 176144 527494 176464 534258
rect 176144 527258 176186 527494
rect 176422 527258 176464 527494
rect 176144 520494 176464 527258
rect 176144 520258 176186 520494
rect 176422 520258 176464 520494
rect 176144 513494 176464 520258
rect 176144 513258 176186 513494
rect 176422 513258 176464 513494
rect 176144 506494 176464 513258
rect 176144 506258 176186 506494
rect 176422 506258 176464 506494
rect 176144 499494 176464 506258
rect 176144 499258 176186 499494
rect 176422 499258 176464 499494
rect 176144 492494 176464 499258
rect 176144 492258 176186 492494
rect 176422 492258 176464 492494
rect 176144 485494 176464 492258
rect 176144 485258 176186 485494
rect 176422 485258 176464 485494
rect 176144 478494 176464 485258
rect 176144 478258 176186 478494
rect 176422 478258 176464 478494
rect 176144 471494 176464 478258
rect 176144 471258 176186 471494
rect 176422 471258 176464 471494
rect 176144 464494 176464 471258
rect 176144 464258 176186 464494
rect 176422 464258 176464 464494
rect 176144 457494 176464 464258
rect 176144 457258 176186 457494
rect 176422 457258 176464 457494
rect 176144 450494 176464 457258
rect 176144 450258 176186 450494
rect 176422 450258 176464 450494
rect 176144 443494 176464 450258
rect 176144 443258 176186 443494
rect 176422 443258 176464 443494
rect 176144 436494 176464 443258
rect 176144 436258 176186 436494
rect 176422 436258 176464 436494
rect 176144 429494 176464 436258
rect 176144 429258 176186 429494
rect 176422 429258 176464 429494
rect 176144 422494 176464 429258
rect 176144 422258 176186 422494
rect 176422 422258 176464 422494
rect 176144 415494 176464 422258
rect 176144 415258 176186 415494
rect 176422 415258 176464 415494
rect 176144 408494 176464 415258
rect 176144 408258 176186 408494
rect 176422 408258 176464 408494
rect 176144 401494 176464 408258
rect 176144 401258 176186 401494
rect 176422 401258 176464 401494
rect 176144 394494 176464 401258
rect 176144 394258 176186 394494
rect 176422 394258 176464 394494
rect 176144 387494 176464 394258
rect 176144 387258 176186 387494
rect 176422 387258 176464 387494
rect 176144 380494 176464 387258
rect 176144 380258 176186 380494
rect 176422 380258 176464 380494
rect 176144 373494 176464 380258
rect 176144 373258 176186 373494
rect 176422 373258 176464 373494
rect 176144 366494 176464 373258
rect 176144 366258 176186 366494
rect 176422 366258 176464 366494
rect 176144 359494 176464 366258
rect 176144 359258 176186 359494
rect 176422 359258 176464 359494
rect 176144 352494 176464 359258
rect 176144 352258 176186 352494
rect 176422 352258 176464 352494
rect 176144 345494 176464 352258
rect 176144 345258 176186 345494
rect 176422 345258 176464 345494
rect 176144 338494 176464 345258
rect 176144 338258 176186 338494
rect 176422 338258 176464 338494
rect 176144 331494 176464 338258
rect 176144 331258 176186 331494
rect 176422 331258 176464 331494
rect 176144 324494 176464 331258
rect 176144 324258 176186 324494
rect 176422 324258 176464 324494
rect 176144 317494 176464 324258
rect 176144 317258 176186 317494
rect 176422 317258 176464 317494
rect 176144 310494 176464 317258
rect 176144 310258 176186 310494
rect 176422 310258 176464 310494
rect 176144 303494 176464 310258
rect 176144 303258 176186 303494
rect 176422 303258 176464 303494
rect 176144 296494 176464 303258
rect 176144 296258 176186 296494
rect 176422 296258 176464 296494
rect 176144 289494 176464 296258
rect 176144 289258 176186 289494
rect 176422 289258 176464 289494
rect 176144 282494 176464 289258
rect 176144 282258 176186 282494
rect 176422 282258 176464 282494
rect 176144 275494 176464 282258
rect 176144 275258 176186 275494
rect 176422 275258 176464 275494
rect 176144 268494 176464 275258
rect 176144 268258 176186 268494
rect 176422 268258 176464 268494
rect 176144 261494 176464 268258
rect 176144 261258 176186 261494
rect 176422 261258 176464 261494
rect 176144 254494 176464 261258
rect 176144 254258 176186 254494
rect 176422 254258 176464 254494
rect 176144 247494 176464 254258
rect 176144 247258 176186 247494
rect 176422 247258 176464 247494
rect 176144 240494 176464 247258
rect 176144 240258 176186 240494
rect 176422 240258 176464 240494
rect 176144 233494 176464 240258
rect 176144 233258 176186 233494
rect 176422 233258 176464 233494
rect 176144 226494 176464 233258
rect 176144 226258 176186 226494
rect 176422 226258 176464 226494
rect 176144 219494 176464 226258
rect 176144 219258 176186 219494
rect 176422 219258 176464 219494
rect 176144 212494 176464 219258
rect 176144 212258 176186 212494
rect 176422 212258 176464 212494
rect 176144 205494 176464 212258
rect 176144 205258 176186 205494
rect 176422 205258 176464 205494
rect 176144 198494 176464 205258
rect 176144 198258 176186 198494
rect 176422 198258 176464 198494
rect 176144 191494 176464 198258
rect 176144 191258 176186 191494
rect 176422 191258 176464 191494
rect 176144 184494 176464 191258
rect 176144 184258 176186 184494
rect 176422 184258 176464 184494
rect 176144 177494 176464 184258
rect 176144 177258 176186 177494
rect 176422 177258 176464 177494
rect 176144 170494 176464 177258
rect 176144 170258 176186 170494
rect 176422 170258 176464 170494
rect 176144 163494 176464 170258
rect 176144 163258 176186 163494
rect 176422 163258 176464 163494
rect 176144 156494 176464 163258
rect 176144 156258 176186 156494
rect 176422 156258 176464 156494
rect 176144 149494 176464 156258
rect 176144 149258 176186 149494
rect 176422 149258 176464 149494
rect 176144 142494 176464 149258
rect 176144 142258 176186 142494
rect 176422 142258 176464 142494
rect 176144 135494 176464 142258
rect 176144 135258 176186 135494
rect 176422 135258 176464 135494
rect 176144 128494 176464 135258
rect 176144 128258 176186 128494
rect 176422 128258 176464 128494
rect 176144 121494 176464 128258
rect 176144 121258 176186 121494
rect 176422 121258 176464 121494
rect 176144 114494 176464 121258
rect 176144 114258 176186 114494
rect 176422 114258 176464 114494
rect 176144 107494 176464 114258
rect 176144 107258 176186 107494
rect 176422 107258 176464 107494
rect 176144 100494 176464 107258
rect 176144 100258 176186 100494
rect 176422 100258 176464 100494
rect 176144 93494 176464 100258
rect 176144 93258 176186 93494
rect 176422 93258 176464 93494
rect 176144 86494 176464 93258
rect 176144 86258 176186 86494
rect 176422 86258 176464 86494
rect 176144 79494 176464 86258
rect 176144 79258 176186 79494
rect 176422 79258 176464 79494
rect 176144 72494 176464 79258
rect 176144 72258 176186 72494
rect 176422 72258 176464 72494
rect 176144 65494 176464 72258
rect 176144 65258 176186 65494
rect 176422 65258 176464 65494
rect 176144 58494 176464 65258
rect 176144 58258 176186 58494
rect 176422 58258 176464 58494
rect 176144 51494 176464 58258
rect 176144 51258 176186 51494
rect 176422 51258 176464 51494
rect 176144 44494 176464 51258
rect 176144 44258 176186 44494
rect 176422 44258 176464 44494
rect 176144 37494 176464 44258
rect 176144 37258 176186 37494
rect 176422 37258 176464 37494
rect 176144 30494 176464 37258
rect 176144 30258 176186 30494
rect 176422 30258 176464 30494
rect 176144 23494 176464 30258
rect 176144 23258 176186 23494
rect 176422 23258 176464 23494
rect 176144 16494 176464 23258
rect 176144 16258 176186 16494
rect 176422 16258 176464 16494
rect 176144 9494 176464 16258
rect 176144 9258 176186 9494
rect 176422 9258 176464 9494
rect 176144 2494 176464 9258
rect 176144 2258 176186 2494
rect 176422 2258 176464 2494
rect 176144 -746 176464 2258
rect 176144 -982 176186 -746
rect 176422 -982 176464 -746
rect 176144 -1066 176464 -982
rect 176144 -1302 176186 -1066
rect 176422 -1302 176464 -1066
rect 176144 -2294 176464 -1302
rect 177876 706198 178196 706230
rect 177876 705962 177918 706198
rect 178154 705962 178196 706198
rect 177876 705878 178196 705962
rect 177876 705642 177918 705878
rect 178154 705642 178196 705878
rect 177876 696434 178196 705642
rect 177876 696198 177918 696434
rect 178154 696198 178196 696434
rect 177876 689434 178196 696198
rect 177876 689198 177918 689434
rect 178154 689198 178196 689434
rect 177876 682434 178196 689198
rect 177876 682198 177918 682434
rect 178154 682198 178196 682434
rect 177876 675434 178196 682198
rect 177876 675198 177918 675434
rect 178154 675198 178196 675434
rect 177876 668434 178196 675198
rect 177876 668198 177918 668434
rect 178154 668198 178196 668434
rect 177876 661434 178196 668198
rect 177876 661198 177918 661434
rect 178154 661198 178196 661434
rect 177876 654434 178196 661198
rect 177876 654198 177918 654434
rect 178154 654198 178196 654434
rect 177876 647434 178196 654198
rect 177876 647198 177918 647434
rect 178154 647198 178196 647434
rect 177876 640434 178196 647198
rect 177876 640198 177918 640434
rect 178154 640198 178196 640434
rect 177876 633434 178196 640198
rect 177876 633198 177918 633434
rect 178154 633198 178196 633434
rect 177876 626434 178196 633198
rect 177876 626198 177918 626434
rect 178154 626198 178196 626434
rect 177876 619434 178196 626198
rect 177876 619198 177918 619434
rect 178154 619198 178196 619434
rect 177876 612434 178196 619198
rect 177876 612198 177918 612434
rect 178154 612198 178196 612434
rect 177876 605434 178196 612198
rect 177876 605198 177918 605434
rect 178154 605198 178196 605434
rect 177876 598434 178196 605198
rect 177876 598198 177918 598434
rect 178154 598198 178196 598434
rect 177876 591434 178196 598198
rect 177876 591198 177918 591434
rect 178154 591198 178196 591434
rect 177876 584434 178196 591198
rect 177876 584198 177918 584434
rect 178154 584198 178196 584434
rect 177876 577434 178196 584198
rect 177876 577198 177918 577434
rect 178154 577198 178196 577434
rect 177876 570434 178196 577198
rect 177876 570198 177918 570434
rect 178154 570198 178196 570434
rect 177876 563434 178196 570198
rect 177876 563198 177918 563434
rect 178154 563198 178196 563434
rect 177876 556434 178196 563198
rect 177876 556198 177918 556434
rect 178154 556198 178196 556434
rect 177876 549434 178196 556198
rect 177876 549198 177918 549434
rect 178154 549198 178196 549434
rect 177876 542434 178196 549198
rect 177876 542198 177918 542434
rect 178154 542198 178196 542434
rect 177876 535434 178196 542198
rect 177876 535198 177918 535434
rect 178154 535198 178196 535434
rect 177876 528434 178196 535198
rect 177876 528198 177918 528434
rect 178154 528198 178196 528434
rect 177876 521434 178196 528198
rect 177876 521198 177918 521434
rect 178154 521198 178196 521434
rect 177876 514434 178196 521198
rect 177876 514198 177918 514434
rect 178154 514198 178196 514434
rect 177876 507434 178196 514198
rect 177876 507198 177918 507434
rect 178154 507198 178196 507434
rect 177876 500434 178196 507198
rect 177876 500198 177918 500434
rect 178154 500198 178196 500434
rect 177876 493434 178196 500198
rect 177876 493198 177918 493434
rect 178154 493198 178196 493434
rect 177876 486434 178196 493198
rect 177876 486198 177918 486434
rect 178154 486198 178196 486434
rect 177876 479434 178196 486198
rect 177876 479198 177918 479434
rect 178154 479198 178196 479434
rect 177876 472434 178196 479198
rect 177876 472198 177918 472434
rect 178154 472198 178196 472434
rect 177876 465434 178196 472198
rect 177876 465198 177918 465434
rect 178154 465198 178196 465434
rect 177876 458434 178196 465198
rect 177876 458198 177918 458434
rect 178154 458198 178196 458434
rect 177876 451434 178196 458198
rect 177876 451198 177918 451434
rect 178154 451198 178196 451434
rect 177876 444434 178196 451198
rect 177876 444198 177918 444434
rect 178154 444198 178196 444434
rect 177876 437434 178196 444198
rect 177876 437198 177918 437434
rect 178154 437198 178196 437434
rect 177876 430434 178196 437198
rect 177876 430198 177918 430434
rect 178154 430198 178196 430434
rect 177876 423434 178196 430198
rect 177876 423198 177918 423434
rect 178154 423198 178196 423434
rect 177876 416434 178196 423198
rect 177876 416198 177918 416434
rect 178154 416198 178196 416434
rect 177876 409434 178196 416198
rect 177876 409198 177918 409434
rect 178154 409198 178196 409434
rect 177876 402434 178196 409198
rect 177876 402198 177918 402434
rect 178154 402198 178196 402434
rect 177876 395434 178196 402198
rect 177876 395198 177918 395434
rect 178154 395198 178196 395434
rect 177876 388434 178196 395198
rect 177876 388198 177918 388434
rect 178154 388198 178196 388434
rect 177876 381434 178196 388198
rect 177876 381198 177918 381434
rect 178154 381198 178196 381434
rect 177876 374434 178196 381198
rect 177876 374198 177918 374434
rect 178154 374198 178196 374434
rect 177876 367434 178196 374198
rect 177876 367198 177918 367434
rect 178154 367198 178196 367434
rect 177876 360434 178196 367198
rect 177876 360198 177918 360434
rect 178154 360198 178196 360434
rect 177876 353434 178196 360198
rect 177876 353198 177918 353434
rect 178154 353198 178196 353434
rect 177876 346434 178196 353198
rect 177876 346198 177918 346434
rect 178154 346198 178196 346434
rect 177876 339434 178196 346198
rect 177876 339198 177918 339434
rect 178154 339198 178196 339434
rect 177876 332434 178196 339198
rect 177876 332198 177918 332434
rect 178154 332198 178196 332434
rect 177876 325434 178196 332198
rect 177876 325198 177918 325434
rect 178154 325198 178196 325434
rect 177876 318434 178196 325198
rect 177876 318198 177918 318434
rect 178154 318198 178196 318434
rect 177876 311434 178196 318198
rect 177876 311198 177918 311434
rect 178154 311198 178196 311434
rect 177876 304434 178196 311198
rect 177876 304198 177918 304434
rect 178154 304198 178196 304434
rect 177876 297434 178196 304198
rect 177876 297198 177918 297434
rect 178154 297198 178196 297434
rect 177876 290434 178196 297198
rect 177876 290198 177918 290434
rect 178154 290198 178196 290434
rect 177876 283434 178196 290198
rect 177876 283198 177918 283434
rect 178154 283198 178196 283434
rect 177876 276434 178196 283198
rect 177876 276198 177918 276434
rect 178154 276198 178196 276434
rect 177876 269434 178196 276198
rect 177876 269198 177918 269434
rect 178154 269198 178196 269434
rect 177876 262434 178196 269198
rect 177876 262198 177918 262434
rect 178154 262198 178196 262434
rect 177876 255434 178196 262198
rect 177876 255198 177918 255434
rect 178154 255198 178196 255434
rect 177876 248434 178196 255198
rect 177876 248198 177918 248434
rect 178154 248198 178196 248434
rect 177876 241434 178196 248198
rect 177876 241198 177918 241434
rect 178154 241198 178196 241434
rect 177876 234434 178196 241198
rect 177876 234198 177918 234434
rect 178154 234198 178196 234434
rect 177876 227434 178196 234198
rect 177876 227198 177918 227434
rect 178154 227198 178196 227434
rect 177876 220434 178196 227198
rect 177876 220198 177918 220434
rect 178154 220198 178196 220434
rect 177876 213434 178196 220198
rect 177876 213198 177918 213434
rect 178154 213198 178196 213434
rect 177876 206434 178196 213198
rect 177876 206198 177918 206434
rect 178154 206198 178196 206434
rect 177876 199434 178196 206198
rect 177876 199198 177918 199434
rect 178154 199198 178196 199434
rect 177876 192434 178196 199198
rect 177876 192198 177918 192434
rect 178154 192198 178196 192434
rect 177876 185434 178196 192198
rect 177876 185198 177918 185434
rect 178154 185198 178196 185434
rect 177876 178434 178196 185198
rect 177876 178198 177918 178434
rect 178154 178198 178196 178434
rect 177876 171434 178196 178198
rect 177876 171198 177918 171434
rect 178154 171198 178196 171434
rect 177876 164434 178196 171198
rect 177876 164198 177918 164434
rect 178154 164198 178196 164434
rect 177876 157434 178196 164198
rect 177876 157198 177918 157434
rect 178154 157198 178196 157434
rect 177876 150434 178196 157198
rect 177876 150198 177918 150434
rect 178154 150198 178196 150434
rect 177876 143434 178196 150198
rect 177876 143198 177918 143434
rect 178154 143198 178196 143434
rect 177876 136434 178196 143198
rect 177876 136198 177918 136434
rect 178154 136198 178196 136434
rect 177876 129434 178196 136198
rect 177876 129198 177918 129434
rect 178154 129198 178196 129434
rect 177876 122434 178196 129198
rect 177876 122198 177918 122434
rect 178154 122198 178196 122434
rect 177876 115434 178196 122198
rect 177876 115198 177918 115434
rect 178154 115198 178196 115434
rect 177876 108434 178196 115198
rect 177876 108198 177918 108434
rect 178154 108198 178196 108434
rect 177876 101434 178196 108198
rect 177876 101198 177918 101434
rect 178154 101198 178196 101434
rect 177876 94434 178196 101198
rect 177876 94198 177918 94434
rect 178154 94198 178196 94434
rect 177876 87434 178196 94198
rect 177876 87198 177918 87434
rect 178154 87198 178196 87434
rect 177876 80434 178196 87198
rect 177876 80198 177918 80434
rect 178154 80198 178196 80434
rect 177876 73434 178196 80198
rect 177876 73198 177918 73434
rect 178154 73198 178196 73434
rect 177876 66434 178196 73198
rect 177876 66198 177918 66434
rect 178154 66198 178196 66434
rect 177876 59434 178196 66198
rect 177876 59198 177918 59434
rect 178154 59198 178196 59434
rect 177876 52434 178196 59198
rect 177876 52198 177918 52434
rect 178154 52198 178196 52434
rect 177876 45434 178196 52198
rect 177876 45198 177918 45434
rect 178154 45198 178196 45434
rect 177876 38434 178196 45198
rect 177876 38198 177918 38434
rect 178154 38198 178196 38434
rect 177876 31434 178196 38198
rect 177876 31198 177918 31434
rect 178154 31198 178196 31434
rect 177876 24434 178196 31198
rect 177876 24198 177918 24434
rect 178154 24198 178196 24434
rect 177876 17434 178196 24198
rect 177876 17198 177918 17434
rect 178154 17198 178196 17434
rect 177876 10434 178196 17198
rect 177876 10198 177918 10434
rect 178154 10198 178196 10434
rect 177876 3434 178196 10198
rect 177876 3198 177918 3434
rect 178154 3198 178196 3434
rect 177876 -1706 178196 3198
rect 177876 -1942 177918 -1706
rect 178154 -1942 178196 -1706
rect 177876 -2026 178196 -1942
rect 177876 -2262 177918 -2026
rect 178154 -2262 178196 -2026
rect 177876 -2294 178196 -2262
rect 183144 705238 183464 706230
rect 183144 705002 183186 705238
rect 183422 705002 183464 705238
rect 183144 704918 183464 705002
rect 183144 704682 183186 704918
rect 183422 704682 183464 704918
rect 183144 695494 183464 704682
rect 183144 695258 183186 695494
rect 183422 695258 183464 695494
rect 183144 688494 183464 695258
rect 183144 688258 183186 688494
rect 183422 688258 183464 688494
rect 183144 681494 183464 688258
rect 183144 681258 183186 681494
rect 183422 681258 183464 681494
rect 183144 674494 183464 681258
rect 183144 674258 183186 674494
rect 183422 674258 183464 674494
rect 183144 667494 183464 674258
rect 183144 667258 183186 667494
rect 183422 667258 183464 667494
rect 183144 660494 183464 667258
rect 183144 660258 183186 660494
rect 183422 660258 183464 660494
rect 183144 653494 183464 660258
rect 183144 653258 183186 653494
rect 183422 653258 183464 653494
rect 183144 646494 183464 653258
rect 183144 646258 183186 646494
rect 183422 646258 183464 646494
rect 183144 639494 183464 646258
rect 183144 639258 183186 639494
rect 183422 639258 183464 639494
rect 183144 632494 183464 639258
rect 183144 632258 183186 632494
rect 183422 632258 183464 632494
rect 183144 625494 183464 632258
rect 183144 625258 183186 625494
rect 183422 625258 183464 625494
rect 183144 618494 183464 625258
rect 183144 618258 183186 618494
rect 183422 618258 183464 618494
rect 183144 611494 183464 618258
rect 183144 611258 183186 611494
rect 183422 611258 183464 611494
rect 183144 604494 183464 611258
rect 183144 604258 183186 604494
rect 183422 604258 183464 604494
rect 183144 597494 183464 604258
rect 183144 597258 183186 597494
rect 183422 597258 183464 597494
rect 183144 590494 183464 597258
rect 183144 590258 183186 590494
rect 183422 590258 183464 590494
rect 183144 583494 183464 590258
rect 183144 583258 183186 583494
rect 183422 583258 183464 583494
rect 183144 576494 183464 583258
rect 183144 576258 183186 576494
rect 183422 576258 183464 576494
rect 183144 569494 183464 576258
rect 183144 569258 183186 569494
rect 183422 569258 183464 569494
rect 183144 562494 183464 569258
rect 183144 562258 183186 562494
rect 183422 562258 183464 562494
rect 183144 555494 183464 562258
rect 183144 555258 183186 555494
rect 183422 555258 183464 555494
rect 183144 548494 183464 555258
rect 183144 548258 183186 548494
rect 183422 548258 183464 548494
rect 183144 541494 183464 548258
rect 183144 541258 183186 541494
rect 183422 541258 183464 541494
rect 183144 534494 183464 541258
rect 183144 534258 183186 534494
rect 183422 534258 183464 534494
rect 183144 527494 183464 534258
rect 183144 527258 183186 527494
rect 183422 527258 183464 527494
rect 183144 520494 183464 527258
rect 183144 520258 183186 520494
rect 183422 520258 183464 520494
rect 183144 513494 183464 520258
rect 183144 513258 183186 513494
rect 183422 513258 183464 513494
rect 183144 506494 183464 513258
rect 183144 506258 183186 506494
rect 183422 506258 183464 506494
rect 183144 499494 183464 506258
rect 183144 499258 183186 499494
rect 183422 499258 183464 499494
rect 183144 492494 183464 499258
rect 183144 492258 183186 492494
rect 183422 492258 183464 492494
rect 183144 485494 183464 492258
rect 183144 485258 183186 485494
rect 183422 485258 183464 485494
rect 183144 478494 183464 485258
rect 183144 478258 183186 478494
rect 183422 478258 183464 478494
rect 183144 471494 183464 478258
rect 183144 471258 183186 471494
rect 183422 471258 183464 471494
rect 183144 464494 183464 471258
rect 183144 464258 183186 464494
rect 183422 464258 183464 464494
rect 183144 457494 183464 464258
rect 183144 457258 183186 457494
rect 183422 457258 183464 457494
rect 183144 450494 183464 457258
rect 183144 450258 183186 450494
rect 183422 450258 183464 450494
rect 183144 443494 183464 450258
rect 183144 443258 183186 443494
rect 183422 443258 183464 443494
rect 183144 436494 183464 443258
rect 183144 436258 183186 436494
rect 183422 436258 183464 436494
rect 183144 429494 183464 436258
rect 183144 429258 183186 429494
rect 183422 429258 183464 429494
rect 183144 422494 183464 429258
rect 183144 422258 183186 422494
rect 183422 422258 183464 422494
rect 183144 415494 183464 422258
rect 183144 415258 183186 415494
rect 183422 415258 183464 415494
rect 183144 408494 183464 415258
rect 183144 408258 183186 408494
rect 183422 408258 183464 408494
rect 183144 401494 183464 408258
rect 183144 401258 183186 401494
rect 183422 401258 183464 401494
rect 183144 394494 183464 401258
rect 183144 394258 183186 394494
rect 183422 394258 183464 394494
rect 183144 387494 183464 394258
rect 183144 387258 183186 387494
rect 183422 387258 183464 387494
rect 183144 380494 183464 387258
rect 183144 380258 183186 380494
rect 183422 380258 183464 380494
rect 183144 373494 183464 380258
rect 183144 373258 183186 373494
rect 183422 373258 183464 373494
rect 183144 366494 183464 373258
rect 183144 366258 183186 366494
rect 183422 366258 183464 366494
rect 183144 359494 183464 366258
rect 183144 359258 183186 359494
rect 183422 359258 183464 359494
rect 183144 352494 183464 359258
rect 183144 352258 183186 352494
rect 183422 352258 183464 352494
rect 183144 345494 183464 352258
rect 183144 345258 183186 345494
rect 183422 345258 183464 345494
rect 183144 338494 183464 345258
rect 183144 338258 183186 338494
rect 183422 338258 183464 338494
rect 183144 331494 183464 338258
rect 183144 331258 183186 331494
rect 183422 331258 183464 331494
rect 183144 324494 183464 331258
rect 183144 324258 183186 324494
rect 183422 324258 183464 324494
rect 183144 317494 183464 324258
rect 183144 317258 183186 317494
rect 183422 317258 183464 317494
rect 183144 310494 183464 317258
rect 183144 310258 183186 310494
rect 183422 310258 183464 310494
rect 183144 303494 183464 310258
rect 183144 303258 183186 303494
rect 183422 303258 183464 303494
rect 183144 296494 183464 303258
rect 183144 296258 183186 296494
rect 183422 296258 183464 296494
rect 183144 289494 183464 296258
rect 183144 289258 183186 289494
rect 183422 289258 183464 289494
rect 183144 282494 183464 289258
rect 183144 282258 183186 282494
rect 183422 282258 183464 282494
rect 183144 275494 183464 282258
rect 183144 275258 183186 275494
rect 183422 275258 183464 275494
rect 183144 268494 183464 275258
rect 183144 268258 183186 268494
rect 183422 268258 183464 268494
rect 183144 261494 183464 268258
rect 183144 261258 183186 261494
rect 183422 261258 183464 261494
rect 183144 254494 183464 261258
rect 183144 254258 183186 254494
rect 183422 254258 183464 254494
rect 183144 247494 183464 254258
rect 183144 247258 183186 247494
rect 183422 247258 183464 247494
rect 183144 240494 183464 247258
rect 183144 240258 183186 240494
rect 183422 240258 183464 240494
rect 183144 233494 183464 240258
rect 183144 233258 183186 233494
rect 183422 233258 183464 233494
rect 183144 226494 183464 233258
rect 183144 226258 183186 226494
rect 183422 226258 183464 226494
rect 183144 219494 183464 226258
rect 183144 219258 183186 219494
rect 183422 219258 183464 219494
rect 183144 212494 183464 219258
rect 183144 212258 183186 212494
rect 183422 212258 183464 212494
rect 183144 205494 183464 212258
rect 183144 205258 183186 205494
rect 183422 205258 183464 205494
rect 183144 198494 183464 205258
rect 183144 198258 183186 198494
rect 183422 198258 183464 198494
rect 183144 191494 183464 198258
rect 183144 191258 183186 191494
rect 183422 191258 183464 191494
rect 183144 184494 183464 191258
rect 183144 184258 183186 184494
rect 183422 184258 183464 184494
rect 183144 177494 183464 184258
rect 183144 177258 183186 177494
rect 183422 177258 183464 177494
rect 183144 170494 183464 177258
rect 183144 170258 183186 170494
rect 183422 170258 183464 170494
rect 183144 163494 183464 170258
rect 183144 163258 183186 163494
rect 183422 163258 183464 163494
rect 183144 156494 183464 163258
rect 183144 156258 183186 156494
rect 183422 156258 183464 156494
rect 183144 149494 183464 156258
rect 183144 149258 183186 149494
rect 183422 149258 183464 149494
rect 183144 142494 183464 149258
rect 183144 142258 183186 142494
rect 183422 142258 183464 142494
rect 183144 135494 183464 142258
rect 183144 135258 183186 135494
rect 183422 135258 183464 135494
rect 183144 128494 183464 135258
rect 183144 128258 183186 128494
rect 183422 128258 183464 128494
rect 183144 121494 183464 128258
rect 183144 121258 183186 121494
rect 183422 121258 183464 121494
rect 183144 114494 183464 121258
rect 183144 114258 183186 114494
rect 183422 114258 183464 114494
rect 183144 107494 183464 114258
rect 183144 107258 183186 107494
rect 183422 107258 183464 107494
rect 183144 100494 183464 107258
rect 183144 100258 183186 100494
rect 183422 100258 183464 100494
rect 183144 93494 183464 100258
rect 183144 93258 183186 93494
rect 183422 93258 183464 93494
rect 183144 86494 183464 93258
rect 183144 86258 183186 86494
rect 183422 86258 183464 86494
rect 183144 79494 183464 86258
rect 183144 79258 183186 79494
rect 183422 79258 183464 79494
rect 183144 72494 183464 79258
rect 183144 72258 183186 72494
rect 183422 72258 183464 72494
rect 183144 65494 183464 72258
rect 183144 65258 183186 65494
rect 183422 65258 183464 65494
rect 183144 58494 183464 65258
rect 183144 58258 183186 58494
rect 183422 58258 183464 58494
rect 183144 51494 183464 58258
rect 183144 51258 183186 51494
rect 183422 51258 183464 51494
rect 183144 44494 183464 51258
rect 183144 44258 183186 44494
rect 183422 44258 183464 44494
rect 183144 37494 183464 44258
rect 183144 37258 183186 37494
rect 183422 37258 183464 37494
rect 183144 30494 183464 37258
rect 183144 30258 183186 30494
rect 183422 30258 183464 30494
rect 183144 23494 183464 30258
rect 183144 23258 183186 23494
rect 183422 23258 183464 23494
rect 183144 16494 183464 23258
rect 183144 16258 183186 16494
rect 183422 16258 183464 16494
rect 183144 9494 183464 16258
rect 183144 9258 183186 9494
rect 183422 9258 183464 9494
rect 183144 2494 183464 9258
rect 183144 2258 183186 2494
rect 183422 2258 183464 2494
rect 183144 -746 183464 2258
rect 183144 -982 183186 -746
rect 183422 -982 183464 -746
rect 183144 -1066 183464 -982
rect 183144 -1302 183186 -1066
rect 183422 -1302 183464 -1066
rect 183144 -2294 183464 -1302
rect 184876 706198 185196 706230
rect 184876 705962 184918 706198
rect 185154 705962 185196 706198
rect 184876 705878 185196 705962
rect 184876 705642 184918 705878
rect 185154 705642 185196 705878
rect 184876 696434 185196 705642
rect 184876 696198 184918 696434
rect 185154 696198 185196 696434
rect 184876 689434 185196 696198
rect 184876 689198 184918 689434
rect 185154 689198 185196 689434
rect 184876 682434 185196 689198
rect 184876 682198 184918 682434
rect 185154 682198 185196 682434
rect 184876 675434 185196 682198
rect 184876 675198 184918 675434
rect 185154 675198 185196 675434
rect 184876 668434 185196 675198
rect 184876 668198 184918 668434
rect 185154 668198 185196 668434
rect 184876 661434 185196 668198
rect 184876 661198 184918 661434
rect 185154 661198 185196 661434
rect 184876 654434 185196 661198
rect 184876 654198 184918 654434
rect 185154 654198 185196 654434
rect 184876 647434 185196 654198
rect 184876 647198 184918 647434
rect 185154 647198 185196 647434
rect 184876 640434 185196 647198
rect 184876 640198 184918 640434
rect 185154 640198 185196 640434
rect 184876 633434 185196 640198
rect 184876 633198 184918 633434
rect 185154 633198 185196 633434
rect 184876 626434 185196 633198
rect 184876 626198 184918 626434
rect 185154 626198 185196 626434
rect 184876 619434 185196 626198
rect 184876 619198 184918 619434
rect 185154 619198 185196 619434
rect 184876 612434 185196 619198
rect 184876 612198 184918 612434
rect 185154 612198 185196 612434
rect 184876 605434 185196 612198
rect 184876 605198 184918 605434
rect 185154 605198 185196 605434
rect 184876 598434 185196 605198
rect 184876 598198 184918 598434
rect 185154 598198 185196 598434
rect 184876 591434 185196 598198
rect 184876 591198 184918 591434
rect 185154 591198 185196 591434
rect 184876 584434 185196 591198
rect 184876 584198 184918 584434
rect 185154 584198 185196 584434
rect 184876 577434 185196 584198
rect 184876 577198 184918 577434
rect 185154 577198 185196 577434
rect 184876 570434 185196 577198
rect 184876 570198 184918 570434
rect 185154 570198 185196 570434
rect 184876 563434 185196 570198
rect 184876 563198 184918 563434
rect 185154 563198 185196 563434
rect 184876 556434 185196 563198
rect 184876 556198 184918 556434
rect 185154 556198 185196 556434
rect 184876 549434 185196 556198
rect 184876 549198 184918 549434
rect 185154 549198 185196 549434
rect 184876 542434 185196 549198
rect 184876 542198 184918 542434
rect 185154 542198 185196 542434
rect 184876 535434 185196 542198
rect 184876 535198 184918 535434
rect 185154 535198 185196 535434
rect 184876 528434 185196 535198
rect 184876 528198 184918 528434
rect 185154 528198 185196 528434
rect 184876 521434 185196 528198
rect 184876 521198 184918 521434
rect 185154 521198 185196 521434
rect 184876 514434 185196 521198
rect 184876 514198 184918 514434
rect 185154 514198 185196 514434
rect 184876 507434 185196 514198
rect 184876 507198 184918 507434
rect 185154 507198 185196 507434
rect 184876 500434 185196 507198
rect 184876 500198 184918 500434
rect 185154 500198 185196 500434
rect 184876 493434 185196 500198
rect 184876 493198 184918 493434
rect 185154 493198 185196 493434
rect 184876 486434 185196 493198
rect 184876 486198 184918 486434
rect 185154 486198 185196 486434
rect 184876 479434 185196 486198
rect 184876 479198 184918 479434
rect 185154 479198 185196 479434
rect 184876 472434 185196 479198
rect 184876 472198 184918 472434
rect 185154 472198 185196 472434
rect 184876 465434 185196 472198
rect 184876 465198 184918 465434
rect 185154 465198 185196 465434
rect 184876 458434 185196 465198
rect 184876 458198 184918 458434
rect 185154 458198 185196 458434
rect 184876 451434 185196 458198
rect 184876 451198 184918 451434
rect 185154 451198 185196 451434
rect 184876 444434 185196 451198
rect 184876 444198 184918 444434
rect 185154 444198 185196 444434
rect 184876 437434 185196 444198
rect 184876 437198 184918 437434
rect 185154 437198 185196 437434
rect 184876 430434 185196 437198
rect 184876 430198 184918 430434
rect 185154 430198 185196 430434
rect 184876 423434 185196 430198
rect 184876 423198 184918 423434
rect 185154 423198 185196 423434
rect 184876 416434 185196 423198
rect 184876 416198 184918 416434
rect 185154 416198 185196 416434
rect 184876 409434 185196 416198
rect 184876 409198 184918 409434
rect 185154 409198 185196 409434
rect 184876 402434 185196 409198
rect 184876 402198 184918 402434
rect 185154 402198 185196 402434
rect 184876 395434 185196 402198
rect 184876 395198 184918 395434
rect 185154 395198 185196 395434
rect 184876 388434 185196 395198
rect 184876 388198 184918 388434
rect 185154 388198 185196 388434
rect 184876 381434 185196 388198
rect 184876 381198 184918 381434
rect 185154 381198 185196 381434
rect 184876 374434 185196 381198
rect 184876 374198 184918 374434
rect 185154 374198 185196 374434
rect 184876 367434 185196 374198
rect 184876 367198 184918 367434
rect 185154 367198 185196 367434
rect 184876 360434 185196 367198
rect 184876 360198 184918 360434
rect 185154 360198 185196 360434
rect 184876 353434 185196 360198
rect 184876 353198 184918 353434
rect 185154 353198 185196 353434
rect 184876 346434 185196 353198
rect 184876 346198 184918 346434
rect 185154 346198 185196 346434
rect 184876 339434 185196 346198
rect 184876 339198 184918 339434
rect 185154 339198 185196 339434
rect 184876 332434 185196 339198
rect 184876 332198 184918 332434
rect 185154 332198 185196 332434
rect 184876 325434 185196 332198
rect 184876 325198 184918 325434
rect 185154 325198 185196 325434
rect 184876 318434 185196 325198
rect 184876 318198 184918 318434
rect 185154 318198 185196 318434
rect 184876 311434 185196 318198
rect 184876 311198 184918 311434
rect 185154 311198 185196 311434
rect 184876 304434 185196 311198
rect 184876 304198 184918 304434
rect 185154 304198 185196 304434
rect 184876 297434 185196 304198
rect 184876 297198 184918 297434
rect 185154 297198 185196 297434
rect 184876 290434 185196 297198
rect 184876 290198 184918 290434
rect 185154 290198 185196 290434
rect 184876 283434 185196 290198
rect 184876 283198 184918 283434
rect 185154 283198 185196 283434
rect 184876 276434 185196 283198
rect 184876 276198 184918 276434
rect 185154 276198 185196 276434
rect 184876 269434 185196 276198
rect 184876 269198 184918 269434
rect 185154 269198 185196 269434
rect 184876 262434 185196 269198
rect 184876 262198 184918 262434
rect 185154 262198 185196 262434
rect 184876 255434 185196 262198
rect 184876 255198 184918 255434
rect 185154 255198 185196 255434
rect 184876 248434 185196 255198
rect 184876 248198 184918 248434
rect 185154 248198 185196 248434
rect 184876 241434 185196 248198
rect 184876 241198 184918 241434
rect 185154 241198 185196 241434
rect 184876 234434 185196 241198
rect 184876 234198 184918 234434
rect 185154 234198 185196 234434
rect 184876 227434 185196 234198
rect 184876 227198 184918 227434
rect 185154 227198 185196 227434
rect 184876 220434 185196 227198
rect 184876 220198 184918 220434
rect 185154 220198 185196 220434
rect 184876 213434 185196 220198
rect 184876 213198 184918 213434
rect 185154 213198 185196 213434
rect 184876 206434 185196 213198
rect 184876 206198 184918 206434
rect 185154 206198 185196 206434
rect 184876 199434 185196 206198
rect 184876 199198 184918 199434
rect 185154 199198 185196 199434
rect 184876 192434 185196 199198
rect 184876 192198 184918 192434
rect 185154 192198 185196 192434
rect 184876 185434 185196 192198
rect 184876 185198 184918 185434
rect 185154 185198 185196 185434
rect 184876 178434 185196 185198
rect 184876 178198 184918 178434
rect 185154 178198 185196 178434
rect 184876 171434 185196 178198
rect 184876 171198 184918 171434
rect 185154 171198 185196 171434
rect 184876 164434 185196 171198
rect 184876 164198 184918 164434
rect 185154 164198 185196 164434
rect 184876 157434 185196 164198
rect 184876 157198 184918 157434
rect 185154 157198 185196 157434
rect 184876 150434 185196 157198
rect 184876 150198 184918 150434
rect 185154 150198 185196 150434
rect 184876 143434 185196 150198
rect 184876 143198 184918 143434
rect 185154 143198 185196 143434
rect 184876 136434 185196 143198
rect 184876 136198 184918 136434
rect 185154 136198 185196 136434
rect 184876 129434 185196 136198
rect 184876 129198 184918 129434
rect 185154 129198 185196 129434
rect 184876 122434 185196 129198
rect 184876 122198 184918 122434
rect 185154 122198 185196 122434
rect 184876 115434 185196 122198
rect 184876 115198 184918 115434
rect 185154 115198 185196 115434
rect 184876 108434 185196 115198
rect 184876 108198 184918 108434
rect 185154 108198 185196 108434
rect 184876 101434 185196 108198
rect 184876 101198 184918 101434
rect 185154 101198 185196 101434
rect 184876 94434 185196 101198
rect 184876 94198 184918 94434
rect 185154 94198 185196 94434
rect 184876 87434 185196 94198
rect 184876 87198 184918 87434
rect 185154 87198 185196 87434
rect 184876 80434 185196 87198
rect 184876 80198 184918 80434
rect 185154 80198 185196 80434
rect 184876 73434 185196 80198
rect 184876 73198 184918 73434
rect 185154 73198 185196 73434
rect 184876 66434 185196 73198
rect 184876 66198 184918 66434
rect 185154 66198 185196 66434
rect 184876 59434 185196 66198
rect 184876 59198 184918 59434
rect 185154 59198 185196 59434
rect 184876 52434 185196 59198
rect 184876 52198 184918 52434
rect 185154 52198 185196 52434
rect 184876 45434 185196 52198
rect 184876 45198 184918 45434
rect 185154 45198 185196 45434
rect 184876 38434 185196 45198
rect 184876 38198 184918 38434
rect 185154 38198 185196 38434
rect 184876 31434 185196 38198
rect 184876 31198 184918 31434
rect 185154 31198 185196 31434
rect 184876 24434 185196 31198
rect 184876 24198 184918 24434
rect 185154 24198 185196 24434
rect 184876 17434 185196 24198
rect 184876 17198 184918 17434
rect 185154 17198 185196 17434
rect 184876 10434 185196 17198
rect 184876 10198 184918 10434
rect 185154 10198 185196 10434
rect 184876 3434 185196 10198
rect 184876 3198 184918 3434
rect 185154 3198 185196 3434
rect 184876 -1706 185196 3198
rect 184876 -1942 184918 -1706
rect 185154 -1942 185196 -1706
rect 184876 -2026 185196 -1942
rect 184876 -2262 184918 -2026
rect 185154 -2262 185196 -2026
rect 184876 -2294 185196 -2262
rect 190144 705238 190464 706230
rect 190144 705002 190186 705238
rect 190422 705002 190464 705238
rect 190144 704918 190464 705002
rect 190144 704682 190186 704918
rect 190422 704682 190464 704918
rect 190144 695494 190464 704682
rect 190144 695258 190186 695494
rect 190422 695258 190464 695494
rect 190144 688494 190464 695258
rect 190144 688258 190186 688494
rect 190422 688258 190464 688494
rect 190144 681494 190464 688258
rect 190144 681258 190186 681494
rect 190422 681258 190464 681494
rect 190144 674494 190464 681258
rect 190144 674258 190186 674494
rect 190422 674258 190464 674494
rect 190144 667494 190464 674258
rect 190144 667258 190186 667494
rect 190422 667258 190464 667494
rect 190144 660494 190464 667258
rect 190144 660258 190186 660494
rect 190422 660258 190464 660494
rect 190144 653494 190464 660258
rect 190144 653258 190186 653494
rect 190422 653258 190464 653494
rect 190144 646494 190464 653258
rect 190144 646258 190186 646494
rect 190422 646258 190464 646494
rect 190144 639494 190464 646258
rect 190144 639258 190186 639494
rect 190422 639258 190464 639494
rect 190144 632494 190464 639258
rect 190144 632258 190186 632494
rect 190422 632258 190464 632494
rect 190144 625494 190464 632258
rect 190144 625258 190186 625494
rect 190422 625258 190464 625494
rect 190144 618494 190464 625258
rect 190144 618258 190186 618494
rect 190422 618258 190464 618494
rect 190144 611494 190464 618258
rect 190144 611258 190186 611494
rect 190422 611258 190464 611494
rect 190144 604494 190464 611258
rect 190144 604258 190186 604494
rect 190422 604258 190464 604494
rect 190144 597494 190464 604258
rect 190144 597258 190186 597494
rect 190422 597258 190464 597494
rect 190144 590494 190464 597258
rect 190144 590258 190186 590494
rect 190422 590258 190464 590494
rect 190144 583494 190464 590258
rect 190144 583258 190186 583494
rect 190422 583258 190464 583494
rect 190144 576494 190464 583258
rect 190144 576258 190186 576494
rect 190422 576258 190464 576494
rect 190144 569494 190464 576258
rect 190144 569258 190186 569494
rect 190422 569258 190464 569494
rect 190144 562494 190464 569258
rect 190144 562258 190186 562494
rect 190422 562258 190464 562494
rect 190144 555494 190464 562258
rect 190144 555258 190186 555494
rect 190422 555258 190464 555494
rect 190144 548494 190464 555258
rect 190144 548258 190186 548494
rect 190422 548258 190464 548494
rect 190144 541494 190464 548258
rect 190144 541258 190186 541494
rect 190422 541258 190464 541494
rect 190144 534494 190464 541258
rect 190144 534258 190186 534494
rect 190422 534258 190464 534494
rect 190144 527494 190464 534258
rect 190144 527258 190186 527494
rect 190422 527258 190464 527494
rect 190144 520494 190464 527258
rect 190144 520258 190186 520494
rect 190422 520258 190464 520494
rect 190144 513494 190464 520258
rect 190144 513258 190186 513494
rect 190422 513258 190464 513494
rect 190144 506494 190464 513258
rect 190144 506258 190186 506494
rect 190422 506258 190464 506494
rect 190144 499494 190464 506258
rect 190144 499258 190186 499494
rect 190422 499258 190464 499494
rect 190144 492494 190464 499258
rect 190144 492258 190186 492494
rect 190422 492258 190464 492494
rect 190144 485494 190464 492258
rect 190144 485258 190186 485494
rect 190422 485258 190464 485494
rect 190144 478494 190464 485258
rect 190144 478258 190186 478494
rect 190422 478258 190464 478494
rect 190144 471494 190464 478258
rect 190144 471258 190186 471494
rect 190422 471258 190464 471494
rect 190144 464494 190464 471258
rect 190144 464258 190186 464494
rect 190422 464258 190464 464494
rect 190144 457494 190464 464258
rect 190144 457258 190186 457494
rect 190422 457258 190464 457494
rect 190144 450494 190464 457258
rect 190144 450258 190186 450494
rect 190422 450258 190464 450494
rect 190144 443494 190464 450258
rect 190144 443258 190186 443494
rect 190422 443258 190464 443494
rect 190144 436494 190464 443258
rect 190144 436258 190186 436494
rect 190422 436258 190464 436494
rect 190144 429494 190464 436258
rect 190144 429258 190186 429494
rect 190422 429258 190464 429494
rect 190144 422494 190464 429258
rect 190144 422258 190186 422494
rect 190422 422258 190464 422494
rect 190144 415494 190464 422258
rect 190144 415258 190186 415494
rect 190422 415258 190464 415494
rect 190144 408494 190464 415258
rect 190144 408258 190186 408494
rect 190422 408258 190464 408494
rect 190144 401494 190464 408258
rect 190144 401258 190186 401494
rect 190422 401258 190464 401494
rect 190144 394494 190464 401258
rect 190144 394258 190186 394494
rect 190422 394258 190464 394494
rect 190144 387494 190464 394258
rect 190144 387258 190186 387494
rect 190422 387258 190464 387494
rect 190144 380494 190464 387258
rect 190144 380258 190186 380494
rect 190422 380258 190464 380494
rect 190144 373494 190464 380258
rect 190144 373258 190186 373494
rect 190422 373258 190464 373494
rect 190144 366494 190464 373258
rect 190144 366258 190186 366494
rect 190422 366258 190464 366494
rect 190144 359494 190464 366258
rect 190144 359258 190186 359494
rect 190422 359258 190464 359494
rect 190144 352494 190464 359258
rect 190144 352258 190186 352494
rect 190422 352258 190464 352494
rect 190144 345494 190464 352258
rect 190144 345258 190186 345494
rect 190422 345258 190464 345494
rect 190144 338494 190464 345258
rect 190144 338258 190186 338494
rect 190422 338258 190464 338494
rect 190144 331494 190464 338258
rect 190144 331258 190186 331494
rect 190422 331258 190464 331494
rect 190144 324494 190464 331258
rect 190144 324258 190186 324494
rect 190422 324258 190464 324494
rect 190144 317494 190464 324258
rect 190144 317258 190186 317494
rect 190422 317258 190464 317494
rect 190144 310494 190464 317258
rect 190144 310258 190186 310494
rect 190422 310258 190464 310494
rect 190144 303494 190464 310258
rect 190144 303258 190186 303494
rect 190422 303258 190464 303494
rect 190144 296494 190464 303258
rect 190144 296258 190186 296494
rect 190422 296258 190464 296494
rect 190144 289494 190464 296258
rect 190144 289258 190186 289494
rect 190422 289258 190464 289494
rect 190144 282494 190464 289258
rect 190144 282258 190186 282494
rect 190422 282258 190464 282494
rect 190144 275494 190464 282258
rect 190144 275258 190186 275494
rect 190422 275258 190464 275494
rect 190144 268494 190464 275258
rect 190144 268258 190186 268494
rect 190422 268258 190464 268494
rect 190144 261494 190464 268258
rect 190144 261258 190186 261494
rect 190422 261258 190464 261494
rect 190144 254494 190464 261258
rect 190144 254258 190186 254494
rect 190422 254258 190464 254494
rect 190144 247494 190464 254258
rect 190144 247258 190186 247494
rect 190422 247258 190464 247494
rect 190144 240494 190464 247258
rect 190144 240258 190186 240494
rect 190422 240258 190464 240494
rect 190144 233494 190464 240258
rect 190144 233258 190186 233494
rect 190422 233258 190464 233494
rect 190144 226494 190464 233258
rect 190144 226258 190186 226494
rect 190422 226258 190464 226494
rect 190144 219494 190464 226258
rect 190144 219258 190186 219494
rect 190422 219258 190464 219494
rect 190144 212494 190464 219258
rect 190144 212258 190186 212494
rect 190422 212258 190464 212494
rect 190144 205494 190464 212258
rect 190144 205258 190186 205494
rect 190422 205258 190464 205494
rect 190144 198494 190464 205258
rect 190144 198258 190186 198494
rect 190422 198258 190464 198494
rect 190144 191494 190464 198258
rect 190144 191258 190186 191494
rect 190422 191258 190464 191494
rect 190144 184494 190464 191258
rect 190144 184258 190186 184494
rect 190422 184258 190464 184494
rect 190144 177494 190464 184258
rect 190144 177258 190186 177494
rect 190422 177258 190464 177494
rect 190144 170494 190464 177258
rect 190144 170258 190186 170494
rect 190422 170258 190464 170494
rect 190144 163494 190464 170258
rect 190144 163258 190186 163494
rect 190422 163258 190464 163494
rect 190144 156494 190464 163258
rect 190144 156258 190186 156494
rect 190422 156258 190464 156494
rect 190144 149494 190464 156258
rect 190144 149258 190186 149494
rect 190422 149258 190464 149494
rect 190144 142494 190464 149258
rect 190144 142258 190186 142494
rect 190422 142258 190464 142494
rect 190144 135494 190464 142258
rect 190144 135258 190186 135494
rect 190422 135258 190464 135494
rect 190144 128494 190464 135258
rect 190144 128258 190186 128494
rect 190422 128258 190464 128494
rect 190144 121494 190464 128258
rect 190144 121258 190186 121494
rect 190422 121258 190464 121494
rect 190144 114494 190464 121258
rect 190144 114258 190186 114494
rect 190422 114258 190464 114494
rect 190144 107494 190464 114258
rect 190144 107258 190186 107494
rect 190422 107258 190464 107494
rect 190144 100494 190464 107258
rect 190144 100258 190186 100494
rect 190422 100258 190464 100494
rect 190144 93494 190464 100258
rect 190144 93258 190186 93494
rect 190422 93258 190464 93494
rect 190144 86494 190464 93258
rect 190144 86258 190186 86494
rect 190422 86258 190464 86494
rect 190144 79494 190464 86258
rect 190144 79258 190186 79494
rect 190422 79258 190464 79494
rect 190144 72494 190464 79258
rect 190144 72258 190186 72494
rect 190422 72258 190464 72494
rect 190144 65494 190464 72258
rect 190144 65258 190186 65494
rect 190422 65258 190464 65494
rect 190144 58494 190464 65258
rect 190144 58258 190186 58494
rect 190422 58258 190464 58494
rect 190144 51494 190464 58258
rect 190144 51258 190186 51494
rect 190422 51258 190464 51494
rect 190144 44494 190464 51258
rect 190144 44258 190186 44494
rect 190422 44258 190464 44494
rect 190144 37494 190464 44258
rect 190144 37258 190186 37494
rect 190422 37258 190464 37494
rect 190144 30494 190464 37258
rect 190144 30258 190186 30494
rect 190422 30258 190464 30494
rect 190144 23494 190464 30258
rect 190144 23258 190186 23494
rect 190422 23258 190464 23494
rect 190144 16494 190464 23258
rect 190144 16258 190186 16494
rect 190422 16258 190464 16494
rect 190144 9494 190464 16258
rect 190144 9258 190186 9494
rect 190422 9258 190464 9494
rect 190144 2494 190464 9258
rect 190144 2258 190186 2494
rect 190422 2258 190464 2494
rect 190144 -746 190464 2258
rect 190144 -982 190186 -746
rect 190422 -982 190464 -746
rect 190144 -1066 190464 -982
rect 190144 -1302 190186 -1066
rect 190422 -1302 190464 -1066
rect 190144 -2294 190464 -1302
rect 191876 706198 192196 706230
rect 191876 705962 191918 706198
rect 192154 705962 192196 706198
rect 191876 705878 192196 705962
rect 191876 705642 191918 705878
rect 192154 705642 192196 705878
rect 191876 696434 192196 705642
rect 191876 696198 191918 696434
rect 192154 696198 192196 696434
rect 191876 689434 192196 696198
rect 191876 689198 191918 689434
rect 192154 689198 192196 689434
rect 191876 682434 192196 689198
rect 191876 682198 191918 682434
rect 192154 682198 192196 682434
rect 191876 675434 192196 682198
rect 191876 675198 191918 675434
rect 192154 675198 192196 675434
rect 191876 668434 192196 675198
rect 191876 668198 191918 668434
rect 192154 668198 192196 668434
rect 191876 661434 192196 668198
rect 191876 661198 191918 661434
rect 192154 661198 192196 661434
rect 191876 654434 192196 661198
rect 191876 654198 191918 654434
rect 192154 654198 192196 654434
rect 191876 647434 192196 654198
rect 191876 647198 191918 647434
rect 192154 647198 192196 647434
rect 191876 640434 192196 647198
rect 191876 640198 191918 640434
rect 192154 640198 192196 640434
rect 191876 633434 192196 640198
rect 191876 633198 191918 633434
rect 192154 633198 192196 633434
rect 191876 626434 192196 633198
rect 191876 626198 191918 626434
rect 192154 626198 192196 626434
rect 191876 619434 192196 626198
rect 191876 619198 191918 619434
rect 192154 619198 192196 619434
rect 191876 612434 192196 619198
rect 191876 612198 191918 612434
rect 192154 612198 192196 612434
rect 191876 605434 192196 612198
rect 191876 605198 191918 605434
rect 192154 605198 192196 605434
rect 191876 598434 192196 605198
rect 191876 598198 191918 598434
rect 192154 598198 192196 598434
rect 191876 591434 192196 598198
rect 191876 591198 191918 591434
rect 192154 591198 192196 591434
rect 191876 584434 192196 591198
rect 191876 584198 191918 584434
rect 192154 584198 192196 584434
rect 191876 577434 192196 584198
rect 191876 577198 191918 577434
rect 192154 577198 192196 577434
rect 191876 570434 192196 577198
rect 191876 570198 191918 570434
rect 192154 570198 192196 570434
rect 191876 563434 192196 570198
rect 191876 563198 191918 563434
rect 192154 563198 192196 563434
rect 191876 556434 192196 563198
rect 191876 556198 191918 556434
rect 192154 556198 192196 556434
rect 191876 549434 192196 556198
rect 191876 549198 191918 549434
rect 192154 549198 192196 549434
rect 191876 542434 192196 549198
rect 191876 542198 191918 542434
rect 192154 542198 192196 542434
rect 191876 535434 192196 542198
rect 191876 535198 191918 535434
rect 192154 535198 192196 535434
rect 191876 528434 192196 535198
rect 191876 528198 191918 528434
rect 192154 528198 192196 528434
rect 191876 521434 192196 528198
rect 191876 521198 191918 521434
rect 192154 521198 192196 521434
rect 191876 514434 192196 521198
rect 191876 514198 191918 514434
rect 192154 514198 192196 514434
rect 191876 507434 192196 514198
rect 191876 507198 191918 507434
rect 192154 507198 192196 507434
rect 191876 500434 192196 507198
rect 191876 500198 191918 500434
rect 192154 500198 192196 500434
rect 191876 493434 192196 500198
rect 191876 493198 191918 493434
rect 192154 493198 192196 493434
rect 191876 486434 192196 493198
rect 191876 486198 191918 486434
rect 192154 486198 192196 486434
rect 191876 479434 192196 486198
rect 191876 479198 191918 479434
rect 192154 479198 192196 479434
rect 191876 472434 192196 479198
rect 191876 472198 191918 472434
rect 192154 472198 192196 472434
rect 191876 465434 192196 472198
rect 191876 465198 191918 465434
rect 192154 465198 192196 465434
rect 191876 458434 192196 465198
rect 191876 458198 191918 458434
rect 192154 458198 192196 458434
rect 191876 451434 192196 458198
rect 191876 451198 191918 451434
rect 192154 451198 192196 451434
rect 191876 444434 192196 451198
rect 191876 444198 191918 444434
rect 192154 444198 192196 444434
rect 191876 437434 192196 444198
rect 191876 437198 191918 437434
rect 192154 437198 192196 437434
rect 191876 430434 192196 437198
rect 191876 430198 191918 430434
rect 192154 430198 192196 430434
rect 191876 423434 192196 430198
rect 191876 423198 191918 423434
rect 192154 423198 192196 423434
rect 191876 416434 192196 423198
rect 191876 416198 191918 416434
rect 192154 416198 192196 416434
rect 191876 409434 192196 416198
rect 191876 409198 191918 409434
rect 192154 409198 192196 409434
rect 191876 402434 192196 409198
rect 191876 402198 191918 402434
rect 192154 402198 192196 402434
rect 191876 395434 192196 402198
rect 191876 395198 191918 395434
rect 192154 395198 192196 395434
rect 191876 388434 192196 395198
rect 191876 388198 191918 388434
rect 192154 388198 192196 388434
rect 191876 381434 192196 388198
rect 191876 381198 191918 381434
rect 192154 381198 192196 381434
rect 191876 374434 192196 381198
rect 191876 374198 191918 374434
rect 192154 374198 192196 374434
rect 191876 367434 192196 374198
rect 191876 367198 191918 367434
rect 192154 367198 192196 367434
rect 191876 360434 192196 367198
rect 191876 360198 191918 360434
rect 192154 360198 192196 360434
rect 191876 353434 192196 360198
rect 191876 353198 191918 353434
rect 192154 353198 192196 353434
rect 191876 346434 192196 353198
rect 191876 346198 191918 346434
rect 192154 346198 192196 346434
rect 191876 339434 192196 346198
rect 191876 339198 191918 339434
rect 192154 339198 192196 339434
rect 191876 332434 192196 339198
rect 191876 332198 191918 332434
rect 192154 332198 192196 332434
rect 191876 325434 192196 332198
rect 191876 325198 191918 325434
rect 192154 325198 192196 325434
rect 191876 318434 192196 325198
rect 191876 318198 191918 318434
rect 192154 318198 192196 318434
rect 191876 311434 192196 318198
rect 191876 311198 191918 311434
rect 192154 311198 192196 311434
rect 191876 304434 192196 311198
rect 191876 304198 191918 304434
rect 192154 304198 192196 304434
rect 191876 297434 192196 304198
rect 191876 297198 191918 297434
rect 192154 297198 192196 297434
rect 191876 290434 192196 297198
rect 191876 290198 191918 290434
rect 192154 290198 192196 290434
rect 191876 283434 192196 290198
rect 191876 283198 191918 283434
rect 192154 283198 192196 283434
rect 191876 276434 192196 283198
rect 191876 276198 191918 276434
rect 192154 276198 192196 276434
rect 191876 269434 192196 276198
rect 191876 269198 191918 269434
rect 192154 269198 192196 269434
rect 191876 262434 192196 269198
rect 191876 262198 191918 262434
rect 192154 262198 192196 262434
rect 191876 255434 192196 262198
rect 191876 255198 191918 255434
rect 192154 255198 192196 255434
rect 191876 248434 192196 255198
rect 191876 248198 191918 248434
rect 192154 248198 192196 248434
rect 191876 241434 192196 248198
rect 191876 241198 191918 241434
rect 192154 241198 192196 241434
rect 191876 234434 192196 241198
rect 191876 234198 191918 234434
rect 192154 234198 192196 234434
rect 191876 227434 192196 234198
rect 191876 227198 191918 227434
rect 192154 227198 192196 227434
rect 191876 220434 192196 227198
rect 191876 220198 191918 220434
rect 192154 220198 192196 220434
rect 191876 213434 192196 220198
rect 191876 213198 191918 213434
rect 192154 213198 192196 213434
rect 191876 206434 192196 213198
rect 191876 206198 191918 206434
rect 192154 206198 192196 206434
rect 191876 199434 192196 206198
rect 191876 199198 191918 199434
rect 192154 199198 192196 199434
rect 191876 192434 192196 199198
rect 191876 192198 191918 192434
rect 192154 192198 192196 192434
rect 191876 185434 192196 192198
rect 191876 185198 191918 185434
rect 192154 185198 192196 185434
rect 191876 178434 192196 185198
rect 191876 178198 191918 178434
rect 192154 178198 192196 178434
rect 191876 171434 192196 178198
rect 191876 171198 191918 171434
rect 192154 171198 192196 171434
rect 191876 164434 192196 171198
rect 191876 164198 191918 164434
rect 192154 164198 192196 164434
rect 191876 157434 192196 164198
rect 191876 157198 191918 157434
rect 192154 157198 192196 157434
rect 191876 150434 192196 157198
rect 191876 150198 191918 150434
rect 192154 150198 192196 150434
rect 191876 143434 192196 150198
rect 191876 143198 191918 143434
rect 192154 143198 192196 143434
rect 191876 136434 192196 143198
rect 191876 136198 191918 136434
rect 192154 136198 192196 136434
rect 191876 129434 192196 136198
rect 191876 129198 191918 129434
rect 192154 129198 192196 129434
rect 191876 122434 192196 129198
rect 191876 122198 191918 122434
rect 192154 122198 192196 122434
rect 191876 115434 192196 122198
rect 191876 115198 191918 115434
rect 192154 115198 192196 115434
rect 191876 108434 192196 115198
rect 191876 108198 191918 108434
rect 192154 108198 192196 108434
rect 191876 101434 192196 108198
rect 191876 101198 191918 101434
rect 192154 101198 192196 101434
rect 191876 94434 192196 101198
rect 191876 94198 191918 94434
rect 192154 94198 192196 94434
rect 191876 87434 192196 94198
rect 191876 87198 191918 87434
rect 192154 87198 192196 87434
rect 191876 80434 192196 87198
rect 191876 80198 191918 80434
rect 192154 80198 192196 80434
rect 191876 73434 192196 80198
rect 191876 73198 191918 73434
rect 192154 73198 192196 73434
rect 191876 66434 192196 73198
rect 191876 66198 191918 66434
rect 192154 66198 192196 66434
rect 191876 59434 192196 66198
rect 191876 59198 191918 59434
rect 192154 59198 192196 59434
rect 191876 52434 192196 59198
rect 191876 52198 191918 52434
rect 192154 52198 192196 52434
rect 191876 45434 192196 52198
rect 191876 45198 191918 45434
rect 192154 45198 192196 45434
rect 191876 38434 192196 45198
rect 191876 38198 191918 38434
rect 192154 38198 192196 38434
rect 191876 31434 192196 38198
rect 191876 31198 191918 31434
rect 192154 31198 192196 31434
rect 191876 24434 192196 31198
rect 191876 24198 191918 24434
rect 192154 24198 192196 24434
rect 191876 17434 192196 24198
rect 191876 17198 191918 17434
rect 192154 17198 192196 17434
rect 191876 10434 192196 17198
rect 191876 10198 191918 10434
rect 192154 10198 192196 10434
rect 191876 3434 192196 10198
rect 191876 3198 191918 3434
rect 192154 3198 192196 3434
rect 191876 -1706 192196 3198
rect 191876 -1942 191918 -1706
rect 192154 -1942 192196 -1706
rect 191876 -2026 192196 -1942
rect 191876 -2262 191918 -2026
rect 192154 -2262 192196 -2026
rect 191876 -2294 192196 -2262
rect 197144 705238 197464 706230
rect 197144 705002 197186 705238
rect 197422 705002 197464 705238
rect 197144 704918 197464 705002
rect 197144 704682 197186 704918
rect 197422 704682 197464 704918
rect 197144 695494 197464 704682
rect 197144 695258 197186 695494
rect 197422 695258 197464 695494
rect 197144 688494 197464 695258
rect 197144 688258 197186 688494
rect 197422 688258 197464 688494
rect 197144 681494 197464 688258
rect 197144 681258 197186 681494
rect 197422 681258 197464 681494
rect 197144 674494 197464 681258
rect 197144 674258 197186 674494
rect 197422 674258 197464 674494
rect 197144 667494 197464 674258
rect 197144 667258 197186 667494
rect 197422 667258 197464 667494
rect 197144 660494 197464 667258
rect 197144 660258 197186 660494
rect 197422 660258 197464 660494
rect 197144 653494 197464 660258
rect 197144 653258 197186 653494
rect 197422 653258 197464 653494
rect 197144 646494 197464 653258
rect 197144 646258 197186 646494
rect 197422 646258 197464 646494
rect 197144 639494 197464 646258
rect 197144 639258 197186 639494
rect 197422 639258 197464 639494
rect 197144 632494 197464 639258
rect 197144 632258 197186 632494
rect 197422 632258 197464 632494
rect 197144 625494 197464 632258
rect 197144 625258 197186 625494
rect 197422 625258 197464 625494
rect 197144 618494 197464 625258
rect 197144 618258 197186 618494
rect 197422 618258 197464 618494
rect 197144 611494 197464 618258
rect 197144 611258 197186 611494
rect 197422 611258 197464 611494
rect 197144 604494 197464 611258
rect 197144 604258 197186 604494
rect 197422 604258 197464 604494
rect 197144 597494 197464 604258
rect 197144 597258 197186 597494
rect 197422 597258 197464 597494
rect 197144 590494 197464 597258
rect 197144 590258 197186 590494
rect 197422 590258 197464 590494
rect 197144 583494 197464 590258
rect 197144 583258 197186 583494
rect 197422 583258 197464 583494
rect 197144 576494 197464 583258
rect 197144 576258 197186 576494
rect 197422 576258 197464 576494
rect 197144 569494 197464 576258
rect 197144 569258 197186 569494
rect 197422 569258 197464 569494
rect 197144 562494 197464 569258
rect 197144 562258 197186 562494
rect 197422 562258 197464 562494
rect 197144 555494 197464 562258
rect 197144 555258 197186 555494
rect 197422 555258 197464 555494
rect 197144 548494 197464 555258
rect 197144 548258 197186 548494
rect 197422 548258 197464 548494
rect 197144 541494 197464 548258
rect 197144 541258 197186 541494
rect 197422 541258 197464 541494
rect 197144 534494 197464 541258
rect 197144 534258 197186 534494
rect 197422 534258 197464 534494
rect 197144 527494 197464 534258
rect 197144 527258 197186 527494
rect 197422 527258 197464 527494
rect 197144 520494 197464 527258
rect 197144 520258 197186 520494
rect 197422 520258 197464 520494
rect 197144 513494 197464 520258
rect 197144 513258 197186 513494
rect 197422 513258 197464 513494
rect 197144 506494 197464 513258
rect 197144 506258 197186 506494
rect 197422 506258 197464 506494
rect 197144 499494 197464 506258
rect 197144 499258 197186 499494
rect 197422 499258 197464 499494
rect 197144 492494 197464 499258
rect 197144 492258 197186 492494
rect 197422 492258 197464 492494
rect 197144 485494 197464 492258
rect 197144 485258 197186 485494
rect 197422 485258 197464 485494
rect 197144 478494 197464 485258
rect 197144 478258 197186 478494
rect 197422 478258 197464 478494
rect 197144 471494 197464 478258
rect 197144 471258 197186 471494
rect 197422 471258 197464 471494
rect 197144 464494 197464 471258
rect 197144 464258 197186 464494
rect 197422 464258 197464 464494
rect 197144 457494 197464 464258
rect 197144 457258 197186 457494
rect 197422 457258 197464 457494
rect 197144 450494 197464 457258
rect 197144 450258 197186 450494
rect 197422 450258 197464 450494
rect 197144 443494 197464 450258
rect 197144 443258 197186 443494
rect 197422 443258 197464 443494
rect 197144 436494 197464 443258
rect 197144 436258 197186 436494
rect 197422 436258 197464 436494
rect 197144 429494 197464 436258
rect 197144 429258 197186 429494
rect 197422 429258 197464 429494
rect 197144 422494 197464 429258
rect 197144 422258 197186 422494
rect 197422 422258 197464 422494
rect 197144 415494 197464 422258
rect 197144 415258 197186 415494
rect 197422 415258 197464 415494
rect 197144 408494 197464 415258
rect 197144 408258 197186 408494
rect 197422 408258 197464 408494
rect 197144 401494 197464 408258
rect 197144 401258 197186 401494
rect 197422 401258 197464 401494
rect 197144 394494 197464 401258
rect 197144 394258 197186 394494
rect 197422 394258 197464 394494
rect 197144 387494 197464 394258
rect 197144 387258 197186 387494
rect 197422 387258 197464 387494
rect 197144 380494 197464 387258
rect 197144 380258 197186 380494
rect 197422 380258 197464 380494
rect 197144 373494 197464 380258
rect 197144 373258 197186 373494
rect 197422 373258 197464 373494
rect 197144 366494 197464 373258
rect 197144 366258 197186 366494
rect 197422 366258 197464 366494
rect 197144 359494 197464 366258
rect 197144 359258 197186 359494
rect 197422 359258 197464 359494
rect 197144 352494 197464 359258
rect 197144 352258 197186 352494
rect 197422 352258 197464 352494
rect 197144 345494 197464 352258
rect 197144 345258 197186 345494
rect 197422 345258 197464 345494
rect 197144 338494 197464 345258
rect 197144 338258 197186 338494
rect 197422 338258 197464 338494
rect 197144 331494 197464 338258
rect 197144 331258 197186 331494
rect 197422 331258 197464 331494
rect 197144 324494 197464 331258
rect 197144 324258 197186 324494
rect 197422 324258 197464 324494
rect 197144 317494 197464 324258
rect 197144 317258 197186 317494
rect 197422 317258 197464 317494
rect 197144 310494 197464 317258
rect 197144 310258 197186 310494
rect 197422 310258 197464 310494
rect 197144 303494 197464 310258
rect 197144 303258 197186 303494
rect 197422 303258 197464 303494
rect 197144 296494 197464 303258
rect 197144 296258 197186 296494
rect 197422 296258 197464 296494
rect 197144 289494 197464 296258
rect 197144 289258 197186 289494
rect 197422 289258 197464 289494
rect 197144 282494 197464 289258
rect 197144 282258 197186 282494
rect 197422 282258 197464 282494
rect 197144 275494 197464 282258
rect 197144 275258 197186 275494
rect 197422 275258 197464 275494
rect 197144 268494 197464 275258
rect 197144 268258 197186 268494
rect 197422 268258 197464 268494
rect 197144 261494 197464 268258
rect 197144 261258 197186 261494
rect 197422 261258 197464 261494
rect 197144 254494 197464 261258
rect 197144 254258 197186 254494
rect 197422 254258 197464 254494
rect 197144 247494 197464 254258
rect 197144 247258 197186 247494
rect 197422 247258 197464 247494
rect 197144 240494 197464 247258
rect 197144 240258 197186 240494
rect 197422 240258 197464 240494
rect 197144 233494 197464 240258
rect 197144 233258 197186 233494
rect 197422 233258 197464 233494
rect 197144 226494 197464 233258
rect 197144 226258 197186 226494
rect 197422 226258 197464 226494
rect 197144 219494 197464 226258
rect 197144 219258 197186 219494
rect 197422 219258 197464 219494
rect 197144 212494 197464 219258
rect 197144 212258 197186 212494
rect 197422 212258 197464 212494
rect 197144 205494 197464 212258
rect 197144 205258 197186 205494
rect 197422 205258 197464 205494
rect 197144 198494 197464 205258
rect 197144 198258 197186 198494
rect 197422 198258 197464 198494
rect 197144 191494 197464 198258
rect 197144 191258 197186 191494
rect 197422 191258 197464 191494
rect 197144 184494 197464 191258
rect 197144 184258 197186 184494
rect 197422 184258 197464 184494
rect 197144 177494 197464 184258
rect 197144 177258 197186 177494
rect 197422 177258 197464 177494
rect 197144 170494 197464 177258
rect 197144 170258 197186 170494
rect 197422 170258 197464 170494
rect 197144 163494 197464 170258
rect 197144 163258 197186 163494
rect 197422 163258 197464 163494
rect 197144 156494 197464 163258
rect 197144 156258 197186 156494
rect 197422 156258 197464 156494
rect 197144 149494 197464 156258
rect 197144 149258 197186 149494
rect 197422 149258 197464 149494
rect 197144 142494 197464 149258
rect 197144 142258 197186 142494
rect 197422 142258 197464 142494
rect 197144 135494 197464 142258
rect 197144 135258 197186 135494
rect 197422 135258 197464 135494
rect 197144 128494 197464 135258
rect 197144 128258 197186 128494
rect 197422 128258 197464 128494
rect 197144 121494 197464 128258
rect 197144 121258 197186 121494
rect 197422 121258 197464 121494
rect 197144 114494 197464 121258
rect 197144 114258 197186 114494
rect 197422 114258 197464 114494
rect 197144 107494 197464 114258
rect 197144 107258 197186 107494
rect 197422 107258 197464 107494
rect 197144 100494 197464 107258
rect 197144 100258 197186 100494
rect 197422 100258 197464 100494
rect 197144 93494 197464 100258
rect 197144 93258 197186 93494
rect 197422 93258 197464 93494
rect 197144 86494 197464 93258
rect 197144 86258 197186 86494
rect 197422 86258 197464 86494
rect 197144 79494 197464 86258
rect 197144 79258 197186 79494
rect 197422 79258 197464 79494
rect 197144 72494 197464 79258
rect 197144 72258 197186 72494
rect 197422 72258 197464 72494
rect 197144 65494 197464 72258
rect 197144 65258 197186 65494
rect 197422 65258 197464 65494
rect 197144 58494 197464 65258
rect 197144 58258 197186 58494
rect 197422 58258 197464 58494
rect 197144 51494 197464 58258
rect 197144 51258 197186 51494
rect 197422 51258 197464 51494
rect 197144 44494 197464 51258
rect 197144 44258 197186 44494
rect 197422 44258 197464 44494
rect 197144 37494 197464 44258
rect 197144 37258 197186 37494
rect 197422 37258 197464 37494
rect 197144 30494 197464 37258
rect 197144 30258 197186 30494
rect 197422 30258 197464 30494
rect 197144 23494 197464 30258
rect 197144 23258 197186 23494
rect 197422 23258 197464 23494
rect 197144 16494 197464 23258
rect 197144 16258 197186 16494
rect 197422 16258 197464 16494
rect 197144 9494 197464 16258
rect 197144 9258 197186 9494
rect 197422 9258 197464 9494
rect 197144 2494 197464 9258
rect 197144 2258 197186 2494
rect 197422 2258 197464 2494
rect 197144 -746 197464 2258
rect 197144 -982 197186 -746
rect 197422 -982 197464 -746
rect 197144 -1066 197464 -982
rect 197144 -1302 197186 -1066
rect 197422 -1302 197464 -1066
rect 197144 -2294 197464 -1302
rect 198876 706198 199196 706230
rect 198876 705962 198918 706198
rect 199154 705962 199196 706198
rect 198876 705878 199196 705962
rect 198876 705642 198918 705878
rect 199154 705642 199196 705878
rect 198876 696434 199196 705642
rect 198876 696198 198918 696434
rect 199154 696198 199196 696434
rect 198876 689434 199196 696198
rect 198876 689198 198918 689434
rect 199154 689198 199196 689434
rect 198876 682434 199196 689198
rect 198876 682198 198918 682434
rect 199154 682198 199196 682434
rect 198876 675434 199196 682198
rect 198876 675198 198918 675434
rect 199154 675198 199196 675434
rect 198876 668434 199196 675198
rect 198876 668198 198918 668434
rect 199154 668198 199196 668434
rect 198876 661434 199196 668198
rect 198876 661198 198918 661434
rect 199154 661198 199196 661434
rect 198876 654434 199196 661198
rect 198876 654198 198918 654434
rect 199154 654198 199196 654434
rect 198876 647434 199196 654198
rect 198876 647198 198918 647434
rect 199154 647198 199196 647434
rect 198876 640434 199196 647198
rect 198876 640198 198918 640434
rect 199154 640198 199196 640434
rect 198876 633434 199196 640198
rect 198876 633198 198918 633434
rect 199154 633198 199196 633434
rect 198876 626434 199196 633198
rect 198876 626198 198918 626434
rect 199154 626198 199196 626434
rect 198876 619434 199196 626198
rect 198876 619198 198918 619434
rect 199154 619198 199196 619434
rect 198876 612434 199196 619198
rect 198876 612198 198918 612434
rect 199154 612198 199196 612434
rect 198876 605434 199196 612198
rect 198876 605198 198918 605434
rect 199154 605198 199196 605434
rect 198876 598434 199196 605198
rect 198876 598198 198918 598434
rect 199154 598198 199196 598434
rect 198876 591434 199196 598198
rect 198876 591198 198918 591434
rect 199154 591198 199196 591434
rect 198876 584434 199196 591198
rect 198876 584198 198918 584434
rect 199154 584198 199196 584434
rect 198876 577434 199196 584198
rect 198876 577198 198918 577434
rect 199154 577198 199196 577434
rect 198876 570434 199196 577198
rect 198876 570198 198918 570434
rect 199154 570198 199196 570434
rect 198876 563434 199196 570198
rect 198876 563198 198918 563434
rect 199154 563198 199196 563434
rect 198876 556434 199196 563198
rect 198876 556198 198918 556434
rect 199154 556198 199196 556434
rect 198876 549434 199196 556198
rect 198876 549198 198918 549434
rect 199154 549198 199196 549434
rect 198876 542434 199196 549198
rect 198876 542198 198918 542434
rect 199154 542198 199196 542434
rect 198876 535434 199196 542198
rect 198876 535198 198918 535434
rect 199154 535198 199196 535434
rect 198876 528434 199196 535198
rect 198876 528198 198918 528434
rect 199154 528198 199196 528434
rect 198876 521434 199196 528198
rect 198876 521198 198918 521434
rect 199154 521198 199196 521434
rect 198876 514434 199196 521198
rect 198876 514198 198918 514434
rect 199154 514198 199196 514434
rect 198876 507434 199196 514198
rect 198876 507198 198918 507434
rect 199154 507198 199196 507434
rect 198876 500434 199196 507198
rect 198876 500198 198918 500434
rect 199154 500198 199196 500434
rect 198876 493434 199196 500198
rect 198876 493198 198918 493434
rect 199154 493198 199196 493434
rect 198876 486434 199196 493198
rect 198876 486198 198918 486434
rect 199154 486198 199196 486434
rect 198876 479434 199196 486198
rect 198876 479198 198918 479434
rect 199154 479198 199196 479434
rect 198876 472434 199196 479198
rect 198876 472198 198918 472434
rect 199154 472198 199196 472434
rect 198876 465434 199196 472198
rect 198876 465198 198918 465434
rect 199154 465198 199196 465434
rect 198876 458434 199196 465198
rect 198876 458198 198918 458434
rect 199154 458198 199196 458434
rect 198876 451434 199196 458198
rect 198876 451198 198918 451434
rect 199154 451198 199196 451434
rect 198876 444434 199196 451198
rect 198876 444198 198918 444434
rect 199154 444198 199196 444434
rect 198876 437434 199196 444198
rect 198876 437198 198918 437434
rect 199154 437198 199196 437434
rect 198876 430434 199196 437198
rect 198876 430198 198918 430434
rect 199154 430198 199196 430434
rect 198876 423434 199196 430198
rect 198876 423198 198918 423434
rect 199154 423198 199196 423434
rect 198876 416434 199196 423198
rect 198876 416198 198918 416434
rect 199154 416198 199196 416434
rect 198876 409434 199196 416198
rect 198876 409198 198918 409434
rect 199154 409198 199196 409434
rect 198876 402434 199196 409198
rect 198876 402198 198918 402434
rect 199154 402198 199196 402434
rect 198876 395434 199196 402198
rect 198876 395198 198918 395434
rect 199154 395198 199196 395434
rect 198876 388434 199196 395198
rect 198876 388198 198918 388434
rect 199154 388198 199196 388434
rect 198876 381434 199196 388198
rect 198876 381198 198918 381434
rect 199154 381198 199196 381434
rect 198876 374434 199196 381198
rect 198876 374198 198918 374434
rect 199154 374198 199196 374434
rect 198876 367434 199196 374198
rect 198876 367198 198918 367434
rect 199154 367198 199196 367434
rect 198876 360434 199196 367198
rect 198876 360198 198918 360434
rect 199154 360198 199196 360434
rect 198876 353434 199196 360198
rect 198876 353198 198918 353434
rect 199154 353198 199196 353434
rect 198876 346434 199196 353198
rect 198876 346198 198918 346434
rect 199154 346198 199196 346434
rect 198876 339434 199196 346198
rect 198876 339198 198918 339434
rect 199154 339198 199196 339434
rect 198876 332434 199196 339198
rect 198876 332198 198918 332434
rect 199154 332198 199196 332434
rect 198876 325434 199196 332198
rect 198876 325198 198918 325434
rect 199154 325198 199196 325434
rect 198876 318434 199196 325198
rect 198876 318198 198918 318434
rect 199154 318198 199196 318434
rect 198876 311434 199196 318198
rect 198876 311198 198918 311434
rect 199154 311198 199196 311434
rect 198876 304434 199196 311198
rect 198876 304198 198918 304434
rect 199154 304198 199196 304434
rect 198876 297434 199196 304198
rect 198876 297198 198918 297434
rect 199154 297198 199196 297434
rect 198876 290434 199196 297198
rect 198876 290198 198918 290434
rect 199154 290198 199196 290434
rect 198876 283434 199196 290198
rect 198876 283198 198918 283434
rect 199154 283198 199196 283434
rect 198876 276434 199196 283198
rect 198876 276198 198918 276434
rect 199154 276198 199196 276434
rect 198876 269434 199196 276198
rect 198876 269198 198918 269434
rect 199154 269198 199196 269434
rect 198876 262434 199196 269198
rect 198876 262198 198918 262434
rect 199154 262198 199196 262434
rect 198876 255434 199196 262198
rect 198876 255198 198918 255434
rect 199154 255198 199196 255434
rect 198876 248434 199196 255198
rect 198876 248198 198918 248434
rect 199154 248198 199196 248434
rect 198876 241434 199196 248198
rect 198876 241198 198918 241434
rect 199154 241198 199196 241434
rect 198876 234434 199196 241198
rect 198876 234198 198918 234434
rect 199154 234198 199196 234434
rect 198876 227434 199196 234198
rect 198876 227198 198918 227434
rect 199154 227198 199196 227434
rect 198876 220434 199196 227198
rect 198876 220198 198918 220434
rect 199154 220198 199196 220434
rect 198876 213434 199196 220198
rect 198876 213198 198918 213434
rect 199154 213198 199196 213434
rect 198876 206434 199196 213198
rect 198876 206198 198918 206434
rect 199154 206198 199196 206434
rect 198876 199434 199196 206198
rect 198876 199198 198918 199434
rect 199154 199198 199196 199434
rect 198876 192434 199196 199198
rect 198876 192198 198918 192434
rect 199154 192198 199196 192434
rect 198876 185434 199196 192198
rect 198876 185198 198918 185434
rect 199154 185198 199196 185434
rect 198876 178434 199196 185198
rect 198876 178198 198918 178434
rect 199154 178198 199196 178434
rect 198876 171434 199196 178198
rect 198876 171198 198918 171434
rect 199154 171198 199196 171434
rect 198876 164434 199196 171198
rect 198876 164198 198918 164434
rect 199154 164198 199196 164434
rect 198876 157434 199196 164198
rect 198876 157198 198918 157434
rect 199154 157198 199196 157434
rect 198876 150434 199196 157198
rect 198876 150198 198918 150434
rect 199154 150198 199196 150434
rect 198876 143434 199196 150198
rect 198876 143198 198918 143434
rect 199154 143198 199196 143434
rect 198876 136434 199196 143198
rect 198876 136198 198918 136434
rect 199154 136198 199196 136434
rect 198876 129434 199196 136198
rect 198876 129198 198918 129434
rect 199154 129198 199196 129434
rect 198876 122434 199196 129198
rect 198876 122198 198918 122434
rect 199154 122198 199196 122434
rect 198876 115434 199196 122198
rect 198876 115198 198918 115434
rect 199154 115198 199196 115434
rect 198876 108434 199196 115198
rect 198876 108198 198918 108434
rect 199154 108198 199196 108434
rect 198876 101434 199196 108198
rect 198876 101198 198918 101434
rect 199154 101198 199196 101434
rect 198876 94434 199196 101198
rect 198876 94198 198918 94434
rect 199154 94198 199196 94434
rect 198876 87434 199196 94198
rect 198876 87198 198918 87434
rect 199154 87198 199196 87434
rect 198876 80434 199196 87198
rect 198876 80198 198918 80434
rect 199154 80198 199196 80434
rect 198876 73434 199196 80198
rect 198876 73198 198918 73434
rect 199154 73198 199196 73434
rect 198876 66434 199196 73198
rect 198876 66198 198918 66434
rect 199154 66198 199196 66434
rect 198876 59434 199196 66198
rect 198876 59198 198918 59434
rect 199154 59198 199196 59434
rect 198876 52434 199196 59198
rect 198876 52198 198918 52434
rect 199154 52198 199196 52434
rect 198876 45434 199196 52198
rect 198876 45198 198918 45434
rect 199154 45198 199196 45434
rect 198876 38434 199196 45198
rect 198876 38198 198918 38434
rect 199154 38198 199196 38434
rect 198876 31434 199196 38198
rect 198876 31198 198918 31434
rect 199154 31198 199196 31434
rect 198876 24434 199196 31198
rect 198876 24198 198918 24434
rect 199154 24198 199196 24434
rect 198876 17434 199196 24198
rect 198876 17198 198918 17434
rect 199154 17198 199196 17434
rect 198876 10434 199196 17198
rect 198876 10198 198918 10434
rect 199154 10198 199196 10434
rect 198876 3434 199196 10198
rect 198876 3198 198918 3434
rect 199154 3198 199196 3434
rect 198876 -1706 199196 3198
rect 198876 -1942 198918 -1706
rect 199154 -1942 199196 -1706
rect 198876 -2026 199196 -1942
rect 198876 -2262 198918 -2026
rect 199154 -2262 199196 -2026
rect 198876 -2294 199196 -2262
rect 204144 705238 204464 706230
rect 204144 705002 204186 705238
rect 204422 705002 204464 705238
rect 204144 704918 204464 705002
rect 204144 704682 204186 704918
rect 204422 704682 204464 704918
rect 204144 695494 204464 704682
rect 204144 695258 204186 695494
rect 204422 695258 204464 695494
rect 204144 688494 204464 695258
rect 204144 688258 204186 688494
rect 204422 688258 204464 688494
rect 204144 681494 204464 688258
rect 204144 681258 204186 681494
rect 204422 681258 204464 681494
rect 204144 674494 204464 681258
rect 204144 674258 204186 674494
rect 204422 674258 204464 674494
rect 204144 667494 204464 674258
rect 204144 667258 204186 667494
rect 204422 667258 204464 667494
rect 204144 660494 204464 667258
rect 204144 660258 204186 660494
rect 204422 660258 204464 660494
rect 204144 653494 204464 660258
rect 204144 653258 204186 653494
rect 204422 653258 204464 653494
rect 204144 646494 204464 653258
rect 204144 646258 204186 646494
rect 204422 646258 204464 646494
rect 204144 639494 204464 646258
rect 204144 639258 204186 639494
rect 204422 639258 204464 639494
rect 204144 632494 204464 639258
rect 204144 632258 204186 632494
rect 204422 632258 204464 632494
rect 204144 625494 204464 632258
rect 204144 625258 204186 625494
rect 204422 625258 204464 625494
rect 204144 618494 204464 625258
rect 204144 618258 204186 618494
rect 204422 618258 204464 618494
rect 204144 611494 204464 618258
rect 204144 611258 204186 611494
rect 204422 611258 204464 611494
rect 204144 604494 204464 611258
rect 204144 604258 204186 604494
rect 204422 604258 204464 604494
rect 204144 597494 204464 604258
rect 204144 597258 204186 597494
rect 204422 597258 204464 597494
rect 204144 590494 204464 597258
rect 204144 590258 204186 590494
rect 204422 590258 204464 590494
rect 204144 583494 204464 590258
rect 204144 583258 204186 583494
rect 204422 583258 204464 583494
rect 204144 576494 204464 583258
rect 204144 576258 204186 576494
rect 204422 576258 204464 576494
rect 204144 569494 204464 576258
rect 204144 569258 204186 569494
rect 204422 569258 204464 569494
rect 204144 562494 204464 569258
rect 204144 562258 204186 562494
rect 204422 562258 204464 562494
rect 204144 555494 204464 562258
rect 204144 555258 204186 555494
rect 204422 555258 204464 555494
rect 204144 548494 204464 555258
rect 204144 548258 204186 548494
rect 204422 548258 204464 548494
rect 204144 541494 204464 548258
rect 204144 541258 204186 541494
rect 204422 541258 204464 541494
rect 204144 534494 204464 541258
rect 204144 534258 204186 534494
rect 204422 534258 204464 534494
rect 204144 527494 204464 534258
rect 204144 527258 204186 527494
rect 204422 527258 204464 527494
rect 204144 520494 204464 527258
rect 204144 520258 204186 520494
rect 204422 520258 204464 520494
rect 204144 513494 204464 520258
rect 204144 513258 204186 513494
rect 204422 513258 204464 513494
rect 204144 506494 204464 513258
rect 204144 506258 204186 506494
rect 204422 506258 204464 506494
rect 204144 499494 204464 506258
rect 204144 499258 204186 499494
rect 204422 499258 204464 499494
rect 204144 492494 204464 499258
rect 204144 492258 204186 492494
rect 204422 492258 204464 492494
rect 204144 485494 204464 492258
rect 204144 485258 204186 485494
rect 204422 485258 204464 485494
rect 204144 478494 204464 485258
rect 204144 478258 204186 478494
rect 204422 478258 204464 478494
rect 204144 471494 204464 478258
rect 204144 471258 204186 471494
rect 204422 471258 204464 471494
rect 204144 464494 204464 471258
rect 204144 464258 204186 464494
rect 204422 464258 204464 464494
rect 204144 457494 204464 464258
rect 204144 457258 204186 457494
rect 204422 457258 204464 457494
rect 204144 450494 204464 457258
rect 204144 450258 204186 450494
rect 204422 450258 204464 450494
rect 204144 443494 204464 450258
rect 204144 443258 204186 443494
rect 204422 443258 204464 443494
rect 204144 436494 204464 443258
rect 204144 436258 204186 436494
rect 204422 436258 204464 436494
rect 204144 429494 204464 436258
rect 204144 429258 204186 429494
rect 204422 429258 204464 429494
rect 204144 422494 204464 429258
rect 204144 422258 204186 422494
rect 204422 422258 204464 422494
rect 204144 415494 204464 422258
rect 204144 415258 204186 415494
rect 204422 415258 204464 415494
rect 204144 408494 204464 415258
rect 204144 408258 204186 408494
rect 204422 408258 204464 408494
rect 204144 401494 204464 408258
rect 204144 401258 204186 401494
rect 204422 401258 204464 401494
rect 204144 394494 204464 401258
rect 204144 394258 204186 394494
rect 204422 394258 204464 394494
rect 204144 387494 204464 394258
rect 204144 387258 204186 387494
rect 204422 387258 204464 387494
rect 204144 380494 204464 387258
rect 204144 380258 204186 380494
rect 204422 380258 204464 380494
rect 204144 373494 204464 380258
rect 204144 373258 204186 373494
rect 204422 373258 204464 373494
rect 204144 366494 204464 373258
rect 204144 366258 204186 366494
rect 204422 366258 204464 366494
rect 204144 359494 204464 366258
rect 204144 359258 204186 359494
rect 204422 359258 204464 359494
rect 204144 352494 204464 359258
rect 204144 352258 204186 352494
rect 204422 352258 204464 352494
rect 204144 345494 204464 352258
rect 204144 345258 204186 345494
rect 204422 345258 204464 345494
rect 204144 338494 204464 345258
rect 204144 338258 204186 338494
rect 204422 338258 204464 338494
rect 204144 331494 204464 338258
rect 204144 331258 204186 331494
rect 204422 331258 204464 331494
rect 204144 324494 204464 331258
rect 204144 324258 204186 324494
rect 204422 324258 204464 324494
rect 204144 317494 204464 324258
rect 204144 317258 204186 317494
rect 204422 317258 204464 317494
rect 204144 310494 204464 317258
rect 204144 310258 204186 310494
rect 204422 310258 204464 310494
rect 204144 303494 204464 310258
rect 204144 303258 204186 303494
rect 204422 303258 204464 303494
rect 204144 296494 204464 303258
rect 204144 296258 204186 296494
rect 204422 296258 204464 296494
rect 204144 289494 204464 296258
rect 204144 289258 204186 289494
rect 204422 289258 204464 289494
rect 204144 282494 204464 289258
rect 204144 282258 204186 282494
rect 204422 282258 204464 282494
rect 204144 275494 204464 282258
rect 204144 275258 204186 275494
rect 204422 275258 204464 275494
rect 204144 268494 204464 275258
rect 204144 268258 204186 268494
rect 204422 268258 204464 268494
rect 204144 261494 204464 268258
rect 204144 261258 204186 261494
rect 204422 261258 204464 261494
rect 204144 254494 204464 261258
rect 204144 254258 204186 254494
rect 204422 254258 204464 254494
rect 204144 247494 204464 254258
rect 204144 247258 204186 247494
rect 204422 247258 204464 247494
rect 204144 240494 204464 247258
rect 204144 240258 204186 240494
rect 204422 240258 204464 240494
rect 204144 233494 204464 240258
rect 204144 233258 204186 233494
rect 204422 233258 204464 233494
rect 204144 226494 204464 233258
rect 204144 226258 204186 226494
rect 204422 226258 204464 226494
rect 204144 219494 204464 226258
rect 204144 219258 204186 219494
rect 204422 219258 204464 219494
rect 204144 212494 204464 219258
rect 204144 212258 204186 212494
rect 204422 212258 204464 212494
rect 204144 205494 204464 212258
rect 204144 205258 204186 205494
rect 204422 205258 204464 205494
rect 204144 198494 204464 205258
rect 204144 198258 204186 198494
rect 204422 198258 204464 198494
rect 204144 191494 204464 198258
rect 204144 191258 204186 191494
rect 204422 191258 204464 191494
rect 204144 184494 204464 191258
rect 204144 184258 204186 184494
rect 204422 184258 204464 184494
rect 204144 177494 204464 184258
rect 204144 177258 204186 177494
rect 204422 177258 204464 177494
rect 204144 170494 204464 177258
rect 204144 170258 204186 170494
rect 204422 170258 204464 170494
rect 204144 163494 204464 170258
rect 204144 163258 204186 163494
rect 204422 163258 204464 163494
rect 204144 156494 204464 163258
rect 204144 156258 204186 156494
rect 204422 156258 204464 156494
rect 204144 149494 204464 156258
rect 204144 149258 204186 149494
rect 204422 149258 204464 149494
rect 204144 142494 204464 149258
rect 204144 142258 204186 142494
rect 204422 142258 204464 142494
rect 204144 135494 204464 142258
rect 204144 135258 204186 135494
rect 204422 135258 204464 135494
rect 204144 128494 204464 135258
rect 204144 128258 204186 128494
rect 204422 128258 204464 128494
rect 204144 121494 204464 128258
rect 204144 121258 204186 121494
rect 204422 121258 204464 121494
rect 204144 114494 204464 121258
rect 204144 114258 204186 114494
rect 204422 114258 204464 114494
rect 204144 107494 204464 114258
rect 204144 107258 204186 107494
rect 204422 107258 204464 107494
rect 204144 100494 204464 107258
rect 204144 100258 204186 100494
rect 204422 100258 204464 100494
rect 204144 93494 204464 100258
rect 204144 93258 204186 93494
rect 204422 93258 204464 93494
rect 204144 86494 204464 93258
rect 204144 86258 204186 86494
rect 204422 86258 204464 86494
rect 204144 79494 204464 86258
rect 204144 79258 204186 79494
rect 204422 79258 204464 79494
rect 204144 72494 204464 79258
rect 204144 72258 204186 72494
rect 204422 72258 204464 72494
rect 204144 65494 204464 72258
rect 204144 65258 204186 65494
rect 204422 65258 204464 65494
rect 204144 58494 204464 65258
rect 204144 58258 204186 58494
rect 204422 58258 204464 58494
rect 204144 51494 204464 58258
rect 204144 51258 204186 51494
rect 204422 51258 204464 51494
rect 204144 44494 204464 51258
rect 204144 44258 204186 44494
rect 204422 44258 204464 44494
rect 204144 37494 204464 44258
rect 204144 37258 204186 37494
rect 204422 37258 204464 37494
rect 204144 30494 204464 37258
rect 204144 30258 204186 30494
rect 204422 30258 204464 30494
rect 204144 23494 204464 30258
rect 204144 23258 204186 23494
rect 204422 23258 204464 23494
rect 204144 16494 204464 23258
rect 204144 16258 204186 16494
rect 204422 16258 204464 16494
rect 204144 9494 204464 16258
rect 204144 9258 204186 9494
rect 204422 9258 204464 9494
rect 204144 2494 204464 9258
rect 204144 2258 204186 2494
rect 204422 2258 204464 2494
rect 204144 -746 204464 2258
rect 204144 -982 204186 -746
rect 204422 -982 204464 -746
rect 204144 -1066 204464 -982
rect 204144 -1302 204186 -1066
rect 204422 -1302 204464 -1066
rect 204144 -2294 204464 -1302
rect 205876 706198 206196 706230
rect 205876 705962 205918 706198
rect 206154 705962 206196 706198
rect 205876 705878 206196 705962
rect 205876 705642 205918 705878
rect 206154 705642 206196 705878
rect 205876 696434 206196 705642
rect 205876 696198 205918 696434
rect 206154 696198 206196 696434
rect 205876 689434 206196 696198
rect 205876 689198 205918 689434
rect 206154 689198 206196 689434
rect 205876 682434 206196 689198
rect 205876 682198 205918 682434
rect 206154 682198 206196 682434
rect 205876 675434 206196 682198
rect 205876 675198 205918 675434
rect 206154 675198 206196 675434
rect 205876 668434 206196 675198
rect 205876 668198 205918 668434
rect 206154 668198 206196 668434
rect 205876 661434 206196 668198
rect 205876 661198 205918 661434
rect 206154 661198 206196 661434
rect 205876 654434 206196 661198
rect 205876 654198 205918 654434
rect 206154 654198 206196 654434
rect 205876 647434 206196 654198
rect 205876 647198 205918 647434
rect 206154 647198 206196 647434
rect 205876 640434 206196 647198
rect 205876 640198 205918 640434
rect 206154 640198 206196 640434
rect 205876 633434 206196 640198
rect 205876 633198 205918 633434
rect 206154 633198 206196 633434
rect 205876 626434 206196 633198
rect 205876 626198 205918 626434
rect 206154 626198 206196 626434
rect 205876 619434 206196 626198
rect 205876 619198 205918 619434
rect 206154 619198 206196 619434
rect 205876 612434 206196 619198
rect 205876 612198 205918 612434
rect 206154 612198 206196 612434
rect 205876 605434 206196 612198
rect 205876 605198 205918 605434
rect 206154 605198 206196 605434
rect 205876 598434 206196 605198
rect 205876 598198 205918 598434
rect 206154 598198 206196 598434
rect 205876 591434 206196 598198
rect 205876 591198 205918 591434
rect 206154 591198 206196 591434
rect 205876 584434 206196 591198
rect 205876 584198 205918 584434
rect 206154 584198 206196 584434
rect 205876 577434 206196 584198
rect 205876 577198 205918 577434
rect 206154 577198 206196 577434
rect 205876 570434 206196 577198
rect 205876 570198 205918 570434
rect 206154 570198 206196 570434
rect 205876 563434 206196 570198
rect 205876 563198 205918 563434
rect 206154 563198 206196 563434
rect 205876 556434 206196 563198
rect 205876 556198 205918 556434
rect 206154 556198 206196 556434
rect 205876 549434 206196 556198
rect 205876 549198 205918 549434
rect 206154 549198 206196 549434
rect 205876 542434 206196 549198
rect 205876 542198 205918 542434
rect 206154 542198 206196 542434
rect 205876 535434 206196 542198
rect 205876 535198 205918 535434
rect 206154 535198 206196 535434
rect 205876 528434 206196 535198
rect 205876 528198 205918 528434
rect 206154 528198 206196 528434
rect 205876 521434 206196 528198
rect 205876 521198 205918 521434
rect 206154 521198 206196 521434
rect 205876 514434 206196 521198
rect 205876 514198 205918 514434
rect 206154 514198 206196 514434
rect 205876 507434 206196 514198
rect 205876 507198 205918 507434
rect 206154 507198 206196 507434
rect 205876 500434 206196 507198
rect 205876 500198 205918 500434
rect 206154 500198 206196 500434
rect 205876 493434 206196 500198
rect 205876 493198 205918 493434
rect 206154 493198 206196 493434
rect 205876 486434 206196 493198
rect 205876 486198 205918 486434
rect 206154 486198 206196 486434
rect 205876 479434 206196 486198
rect 205876 479198 205918 479434
rect 206154 479198 206196 479434
rect 205876 472434 206196 479198
rect 205876 472198 205918 472434
rect 206154 472198 206196 472434
rect 205876 465434 206196 472198
rect 205876 465198 205918 465434
rect 206154 465198 206196 465434
rect 205876 458434 206196 465198
rect 205876 458198 205918 458434
rect 206154 458198 206196 458434
rect 205876 451434 206196 458198
rect 205876 451198 205918 451434
rect 206154 451198 206196 451434
rect 205876 444434 206196 451198
rect 205876 444198 205918 444434
rect 206154 444198 206196 444434
rect 205876 437434 206196 444198
rect 205876 437198 205918 437434
rect 206154 437198 206196 437434
rect 205876 430434 206196 437198
rect 205876 430198 205918 430434
rect 206154 430198 206196 430434
rect 205876 423434 206196 430198
rect 205876 423198 205918 423434
rect 206154 423198 206196 423434
rect 205876 416434 206196 423198
rect 205876 416198 205918 416434
rect 206154 416198 206196 416434
rect 205876 409434 206196 416198
rect 205876 409198 205918 409434
rect 206154 409198 206196 409434
rect 205876 402434 206196 409198
rect 205876 402198 205918 402434
rect 206154 402198 206196 402434
rect 205876 395434 206196 402198
rect 205876 395198 205918 395434
rect 206154 395198 206196 395434
rect 205876 388434 206196 395198
rect 205876 388198 205918 388434
rect 206154 388198 206196 388434
rect 205876 381434 206196 388198
rect 205876 381198 205918 381434
rect 206154 381198 206196 381434
rect 205876 374434 206196 381198
rect 205876 374198 205918 374434
rect 206154 374198 206196 374434
rect 205876 367434 206196 374198
rect 205876 367198 205918 367434
rect 206154 367198 206196 367434
rect 205876 360434 206196 367198
rect 205876 360198 205918 360434
rect 206154 360198 206196 360434
rect 205876 353434 206196 360198
rect 205876 353198 205918 353434
rect 206154 353198 206196 353434
rect 205876 346434 206196 353198
rect 205876 346198 205918 346434
rect 206154 346198 206196 346434
rect 205876 339434 206196 346198
rect 205876 339198 205918 339434
rect 206154 339198 206196 339434
rect 205876 332434 206196 339198
rect 205876 332198 205918 332434
rect 206154 332198 206196 332434
rect 205876 325434 206196 332198
rect 205876 325198 205918 325434
rect 206154 325198 206196 325434
rect 205876 318434 206196 325198
rect 205876 318198 205918 318434
rect 206154 318198 206196 318434
rect 205876 311434 206196 318198
rect 205876 311198 205918 311434
rect 206154 311198 206196 311434
rect 205876 304434 206196 311198
rect 205876 304198 205918 304434
rect 206154 304198 206196 304434
rect 205876 297434 206196 304198
rect 205876 297198 205918 297434
rect 206154 297198 206196 297434
rect 205876 290434 206196 297198
rect 205876 290198 205918 290434
rect 206154 290198 206196 290434
rect 205876 283434 206196 290198
rect 205876 283198 205918 283434
rect 206154 283198 206196 283434
rect 205876 276434 206196 283198
rect 205876 276198 205918 276434
rect 206154 276198 206196 276434
rect 205876 269434 206196 276198
rect 205876 269198 205918 269434
rect 206154 269198 206196 269434
rect 205876 262434 206196 269198
rect 205876 262198 205918 262434
rect 206154 262198 206196 262434
rect 205876 255434 206196 262198
rect 205876 255198 205918 255434
rect 206154 255198 206196 255434
rect 205876 248434 206196 255198
rect 205876 248198 205918 248434
rect 206154 248198 206196 248434
rect 205876 241434 206196 248198
rect 205876 241198 205918 241434
rect 206154 241198 206196 241434
rect 205876 234434 206196 241198
rect 205876 234198 205918 234434
rect 206154 234198 206196 234434
rect 205876 227434 206196 234198
rect 205876 227198 205918 227434
rect 206154 227198 206196 227434
rect 205876 220434 206196 227198
rect 205876 220198 205918 220434
rect 206154 220198 206196 220434
rect 205876 213434 206196 220198
rect 205876 213198 205918 213434
rect 206154 213198 206196 213434
rect 205876 206434 206196 213198
rect 205876 206198 205918 206434
rect 206154 206198 206196 206434
rect 205876 199434 206196 206198
rect 205876 199198 205918 199434
rect 206154 199198 206196 199434
rect 205876 192434 206196 199198
rect 205876 192198 205918 192434
rect 206154 192198 206196 192434
rect 205876 185434 206196 192198
rect 205876 185198 205918 185434
rect 206154 185198 206196 185434
rect 205876 178434 206196 185198
rect 205876 178198 205918 178434
rect 206154 178198 206196 178434
rect 205876 171434 206196 178198
rect 205876 171198 205918 171434
rect 206154 171198 206196 171434
rect 205876 164434 206196 171198
rect 205876 164198 205918 164434
rect 206154 164198 206196 164434
rect 205876 157434 206196 164198
rect 205876 157198 205918 157434
rect 206154 157198 206196 157434
rect 205876 150434 206196 157198
rect 205876 150198 205918 150434
rect 206154 150198 206196 150434
rect 205876 143434 206196 150198
rect 205876 143198 205918 143434
rect 206154 143198 206196 143434
rect 205876 136434 206196 143198
rect 205876 136198 205918 136434
rect 206154 136198 206196 136434
rect 205876 129434 206196 136198
rect 205876 129198 205918 129434
rect 206154 129198 206196 129434
rect 205876 122434 206196 129198
rect 205876 122198 205918 122434
rect 206154 122198 206196 122434
rect 205876 115434 206196 122198
rect 205876 115198 205918 115434
rect 206154 115198 206196 115434
rect 205876 108434 206196 115198
rect 205876 108198 205918 108434
rect 206154 108198 206196 108434
rect 205876 101434 206196 108198
rect 205876 101198 205918 101434
rect 206154 101198 206196 101434
rect 205876 94434 206196 101198
rect 205876 94198 205918 94434
rect 206154 94198 206196 94434
rect 205876 87434 206196 94198
rect 205876 87198 205918 87434
rect 206154 87198 206196 87434
rect 205876 80434 206196 87198
rect 205876 80198 205918 80434
rect 206154 80198 206196 80434
rect 205876 73434 206196 80198
rect 205876 73198 205918 73434
rect 206154 73198 206196 73434
rect 205876 66434 206196 73198
rect 205876 66198 205918 66434
rect 206154 66198 206196 66434
rect 205876 59434 206196 66198
rect 205876 59198 205918 59434
rect 206154 59198 206196 59434
rect 205876 52434 206196 59198
rect 205876 52198 205918 52434
rect 206154 52198 206196 52434
rect 205876 45434 206196 52198
rect 205876 45198 205918 45434
rect 206154 45198 206196 45434
rect 205876 38434 206196 45198
rect 205876 38198 205918 38434
rect 206154 38198 206196 38434
rect 205876 31434 206196 38198
rect 205876 31198 205918 31434
rect 206154 31198 206196 31434
rect 205876 24434 206196 31198
rect 205876 24198 205918 24434
rect 206154 24198 206196 24434
rect 205876 17434 206196 24198
rect 205876 17198 205918 17434
rect 206154 17198 206196 17434
rect 205876 10434 206196 17198
rect 205876 10198 205918 10434
rect 206154 10198 206196 10434
rect 205876 3434 206196 10198
rect 205876 3198 205918 3434
rect 206154 3198 206196 3434
rect 205876 -1706 206196 3198
rect 205876 -1942 205918 -1706
rect 206154 -1942 206196 -1706
rect 205876 -2026 206196 -1942
rect 205876 -2262 205918 -2026
rect 206154 -2262 206196 -2026
rect 205876 -2294 206196 -2262
rect 211144 705238 211464 706230
rect 211144 705002 211186 705238
rect 211422 705002 211464 705238
rect 211144 704918 211464 705002
rect 211144 704682 211186 704918
rect 211422 704682 211464 704918
rect 211144 695494 211464 704682
rect 211144 695258 211186 695494
rect 211422 695258 211464 695494
rect 211144 688494 211464 695258
rect 211144 688258 211186 688494
rect 211422 688258 211464 688494
rect 211144 681494 211464 688258
rect 211144 681258 211186 681494
rect 211422 681258 211464 681494
rect 211144 674494 211464 681258
rect 211144 674258 211186 674494
rect 211422 674258 211464 674494
rect 211144 667494 211464 674258
rect 211144 667258 211186 667494
rect 211422 667258 211464 667494
rect 211144 660494 211464 667258
rect 211144 660258 211186 660494
rect 211422 660258 211464 660494
rect 211144 653494 211464 660258
rect 211144 653258 211186 653494
rect 211422 653258 211464 653494
rect 211144 646494 211464 653258
rect 211144 646258 211186 646494
rect 211422 646258 211464 646494
rect 211144 639494 211464 646258
rect 211144 639258 211186 639494
rect 211422 639258 211464 639494
rect 211144 632494 211464 639258
rect 211144 632258 211186 632494
rect 211422 632258 211464 632494
rect 211144 625494 211464 632258
rect 211144 625258 211186 625494
rect 211422 625258 211464 625494
rect 211144 618494 211464 625258
rect 211144 618258 211186 618494
rect 211422 618258 211464 618494
rect 211144 611494 211464 618258
rect 211144 611258 211186 611494
rect 211422 611258 211464 611494
rect 211144 604494 211464 611258
rect 211144 604258 211186 604494
rect 211422 604258 211464 604494
rect 211144 597494 211464 604258
rect 211144 597258 211186 597494
rect 211422 597258 211464 597494
rect 211144 590494 211464 597258
rect 211144 590258 211186 590494
rect 211422 590258 211464 590494
rect 211144 583494 211464 590258
rect 211144 583258 211186 583494
rect 211422 583258 211464 583494
rect 211144 576494 211464 583258
rect 211144 576258 211186 576494
rect 211422 576258 211464 576494
rect 211144 569494 211464 576258
rect 211144 569258 211186 569494
rect 211422 569258 211464 569494
rect 211144 562494 211464 569258
rect 211144 562258 211186 562494
rect 211422 562258 211464 562494
rect 211144 555494 211464 562258
rect 211144 555258 211186 555494
rect 211422 555258 211464 555494
rect 211144 548494 211464 555258
rect 211144 548258 211186 548494
rect 211422 548258 211464 548494
rect 211144 541494 211464 548258
rect 211144 541258 211186 541494
rect 211422 541258 211464 541494
rect 211144 534494 211464 541258
rect 211144 534258 211186 534494
rect 211422 534258 211464 534494
rect 211144 527494 211464 534258
rect 211144 527258 211186 527494
rect 211422 527258 211464 527494
rect 211144 520494 211464 527258
rect 211144 520258 211186 520494
rect 211422 520258 211464 520494
rect 211144 513494 211464 520258
rect 211144 513258 211186 513494
rect 211422 513258 211464 513494
rect 211144 506494 211464 513258
rect 211144 506258 211186 506494
rect 211422 506258 211464 506494
rect 211144 499494 211464 506258
rect 211144 499258 211186 499494
rect 211422 499258 211464 499494
rect 211144 492494 211464 499258
rect 211144 492258 211186 492494
rect 211422 492258 211464 492494
rect 211144 485494 211464 492258
rect 211144 485258 211186 485494
rect 211422 485258 211464 485494
rect 211144 478494 211464 485258
rect 211144 478258 211186 478494
rect 211422 478258 211464 478494
rect 211144 471494 211464 478258
rect 211144 471258 211186 471494
rect 211422 471258 211464 471494
rect 211144 464494 211464 471258
rect 211144 464258 211186 464494
rect 211422 464258 211464 464494
rect 211144 457494 211464 464258
rect 211144 457258 211186 457494
rect 211422 457258 211464 457494
rect 211144 450494 211464 457258
rect 211144 450258 211186 450494
rect 211422 450258 211464 450494
rect 211144 443494 211464 450258
rect 211144 443258 211186 443494
rect 211422 443258 211464 443494
rect 211144 436494 211464 443258
rect 211144 436258 211186 436494
rect 211422 436258 211464 436494
rect 211144 429494 211464 436258
rect 211144 429258 211186 429494
rect 211422 429258 211464 429494
rect 211144 422494 211464 429258
rect 211144 422258 211186 422494
rect 211422 422258 211464 422494
rect 211144 415494 211464 422258
rect 211144 415258 211186 415494
rect 211422 415258 211464 415494
rect 211144 408494 211464 415258
rect 211144 408258 211186 408494
rect 211422 408258 211464 408494
rect 211144 401494 211464 408258
rect 211144 401258 211186 401494
rect 211422 401258 211464 401494
rect 211144 394494 211464 401258
rect 211144 394258 211186 394494
rect 211422 394258 211464 394494
rect 211144 387494 211464 394258
rect 211144 387258 211186 387494
rect 211422 387258 211464 387494
rect 211144 380494 211464 387258
rect 211144 380258 211186 380494
rect 211422 380258 211464 380494
rect 211144 373494 211464 380258
rect 211144 373258 211186 373494
rect 211422 373258 211464 373494
rect 211144 366494 211464 373258
rect 211144 366258 211186 366494
rect 211422 366258 211464 366494
rect 211144 359494 211464 366258
rect 211144 359258 211186 359494
rect 211422 359258 211464 359494
rect 211144 352494 211464 359258
rect 211144 352258 211186 352494
rect 211422 352258 211464 352494
rect 211144 345494 211464 352258
rect 211144 345258 211186 345494
rect 211422 345258 211464 345494
rect 211144 338494 211464 345258
rect 211144 338258 211186 338494
rect 211422 338258 211464 338494
rect 211144 331494 211464 338258
rect 211144 331258 211186 331494
rect 211422 331258 211464 331494
rect 211144 324494 211464 331258
rect 211144 324258 211186 324494
rect 211422 324258 211464 324494
rect 211144 317494 211464 324258
rect 211144 317258 211186 317494
rect 211422 317258 211464 317494
rect 211144 310494 211464 317258
rect 211144 310258 211186 310494
rect 211422 310258 211464 310494
rect 211144 303494 211464 310258
rect 211144 303258 211186 303494
rect 211422 303258 211464 303494
rect 211144 296494 211464 303258
rect 211144 296258 211186 296494
rect 211422 296258 211464 296494
rect 211144 289494 211464 296258
rect 211144 289258 211186 289494
rect 211422 289258 211464 289494
rect 211144 282494 211464 289258
rect 211144 282258 211186 282494
rect 211422 282258 211464 282494
rect 211144 275494 211464 282258
rect 211144 275258 211186 275494
rect 211422 275258 211464 275494
rect 211144 268494 211464 275258
rect 211144 268258 211186 268494
rect 211422 268258 211464 268494
rect 211144 261494 211464 268258
rect 211144 261258 211186 261494
rect 211422 261258 211464 261494
rect 211144 254494 211464 261258
rect 211144 254258 211186 254494
rect 211422 254258 211464 254494
rect 211144 247494 211464 254258
rect 211144 247258 211186 247494
rect 211422 247258 211464 247494
rect 211144 240494 211464 247258
rect 211144 240258 211186 240494
rect 211422 240258 211464 240494
rect 211144 233494 211464 240258
rect 211144 233258 211186 233494
rect 211422 233258 211464 233494
rect 211144 226494 211464 233258
rect 211144 226258 211186 226494
rect 211422 226258 211464 226494
rect 211144 219494 211464 226258
rect 211144 219258 211186 219494
rect 211422 219258 211464 219494
rect 211144 212494 211464 219258
rect 211144 212258 211186 212494
rect 211422 212258 211464 212494
rect 211144 205494 211464 212258
rect 211144 205258 211186 205494
rect 211422 205258 211464 205494
rect 211144 198494 211464 205258
rect 211144 198258 211186 198494
rect 211422 198258 211464 198494
rect 211144 191494 211464 198258
rect 211144 191258 211186 191494
rect 211422 191258 211464 191494
rect 211144 184494 211464 191258
rect 211144 184258 211186 184494
rect 211422 184258 211464 184494
rect 211144 177494 211464 184258
rect 211144 177258 211186 177494
rect 211422 177258 211464 177494
rect 211144 170494 211464 177258
rect 211144 170258 211186 170494
rect 211422 170258 211464 170494
rect 211144 163494 211464 170258
rect 211144 163258 211186 163494
rect 211422 163258 211464 163494
rect 211144 156494 211464 163258
rect 211144 156258 211186 156494
rect 211422 156258 211464 156494
rect 211144 149494 211464 156258
rect 211144 149258 211186 149494
rect 211422 149258 211464 149494
rect 211144 142494 211464 149258
rect 211144 142258 211186 142494
rect 211422 142258 211464 142494
rect 211144 135494 211464 142258
rect 211144 135258 211186 135494
rect 211422 135258 211464 135494
rect 211144 128494 211464 135258
rect 211144 128258 211186 128494
rect 211422 128258 211464 128494
rect 211144 121494 211464 128258
rect 211144 121258 211186 121494
rect 211422 121258 211464 121494
rect 211144 114494 211464 121258
rect 211144 114258 211186 114494
rect 211422 114258 211464 114494
rect 211144 107494 211464 114258
rect 211144 107258 211186 107494
rect 211422 107258 211464 107494
rect 211144 100494 211464 107258
rect 211144 100258 211186 100494
rect 211422 100258 211464 100494
rect 211144 93494 211464 100258
rect 211144 93258 211186 93494
rect 211422 93258 211464 93494
rect 211144 86494 211464 93258
rect 211144 86258 211186 86494
rect 211422 86258 211464 86494
rect 211144 79494 211464 86258
rect 211144 79258 211186 79494
rect 211422 79258 211464 79494
rect 211144 72494 211464 79258
rect 211144 72258 211186 72494
rect 211422 72258 211464 72494
rect 211144 65494 211464 72258
rect 211144 65258 211186 65494
rect 211422 65258 211464 65494
rect 211144 58494 211464 65258
rect 211144 58258 211186 58494
rect 211422 58258 211464 58494
rect 211144 51494 211464 58258
rect 211144 51258 211186 51494
rect 211422 51258 211464 51494
rect 211144 44494 211464 51258
rect 211144 44258 211186 44494
rect 211422 44258 211464 44494
rect 211144 37494 211464 44258
rect 211144 37258 211186 37494
rect 211422 37258 211464 37494
rect 211144 30494 211464 37258
rect 211144 30258 211186 30494
rect 211422 30258 211464 30494
rect 211144 23494 211464 30258
rect 211144 23258 211186 23494
rect 211422 23258 211464 23494
rect 211144 16494 211464 23258
rect 211144 16258 211186 16494
rect 211422 16258 211464 16494
rect 211144 9494 211464 16258
rect 211144 9258 211186 9494
rect 211422 9258 211464 9494
rect 211144 2494 211464 9258
rect 211144 2258 211186 2494
rect 211422 2258 211464 2494
rect 211144 -746 211464 2258
rect 211144 -982 211186 -746
rect 211422 -982 211464 -746
rect 211144 -1066 211464 -982
rect 211144 -1302 211186 -1066
rect 211422 -1302 211464 -1066
rect 211144 -2294 211464 -1302
rect 212876 706198 213196 706230
rect 212876 705962 212918 706198
rect 213154 705962 213196 706198
rect 212876 705878 213196 705962
rect 212876 705642 212918 705878
rect 213154 705642 213196 705878
rect 212876 696434 213196 705642
rect 212876 696198 212918 696434
rect 213154 696198 213196 696434
rect 212876 689434 213196 696198
rect 212876 689198 212918 689434
rect 213154 689198 213196 689434
rect 212876 682434 213196 689198
rect 212876 682198 212918 682434
rect 213154 682198 213196 682434
rect 212876 675434 213196 682198
rect 212876 675198 212918 675434
rect 213154 675198 213196 675434
rect 212876 668434 213196 675198
rect 212876 668198 212918 668434
rect 213154 668198 213196 668434
rect 212876 661434 213196 668198
rect 212876 661198 212918 661434
rect 213154 661198 213196 661434
rect 212876 654434 213196 661198
rect 212876 654198 212918 654434
rect 213154 654198 213196 654434
rect 212876 647434 213196 654198
rect 212876 647198 212918 647434
rect 213154 647198 213196 647434
rect 212876 640434 213196 647198
rect 212876 640198 212918 640434
rect 213154 640198 213196 640434
rect 212876 633434 213196 640198
rect 212876 633198 212918 633434
rect 213154 633198 213196 633434
rect 212876 626434 213196 633198
rect 212876 626198 212918 626434
rect 213154 626198 213196 626434
rect 212876 619434 213196 626198
rect 212876 619198 212918 619434
rect 213154 619198 213196 619434
rect 212876 612434 213196 619198
rect 212876 612198 212918 612434
rect 213154 612198 213196 612434
rect 212876 605434 213196 612198
rect 212876 605198 212918 605434
rect 213154 605198 213196 605434
rect 212876 598434 213196 605198
rect 212876 598198 212918 598434
rect 213154 598198 213196 598434
rect 212876 591434 213196 598198
rect 212876 591198 212918 591434
rect 213154 591198 213196 591434
rect 212876 584434 213196 591198
rect 212876 584198 212918 584434
rect 213154 584198 213196 584434
rect 212876 577434 213196 584198
rect 212876 577198 212918 577434
rect 213154 577198 213196 577434
rect 212876 570434 213196 577198
rect 212876 570198 212918 570434
rect 213154 570198 213196 570434
rect 212876 563434 213196 570198
rect 212876 563198 212918 563434
rect 213154 563198 213196 563434
rect 212876 556434 213196 563198
rect 212876 556198 212918 556434
rect 213154 556198 213196 556434
rect 212876 549434 213196 556198
rect 212876 549198 212918 549434
rect 213154 549198 213196 549434
rect 212876 542434 213196 549198
rect 212876 542198 212918 542434
rect 213154 542198 213196 542434
rect 212876 535434 213196 542198
rect 212876 535198 212918 535434
rect 213154 535198 213196 535434
rect 212876 528434 213196 535198
rect 212876 528198 212918 528434
rect 213154 528198 213196 528434
rect 212876 521434 213196 528198
rect 212876 521198 212918 521434
rect 213154 521198 213196 521434
rect 212876 514434 213196 521198
rect 212876 514198 212918 514434
rect 213154 514198 213196 514434
rect 212876 507434 213196 514198
rect 212876 507198 212918 507434
rect 213154 507198 213196 507434
rect 212876 500434 213196 507198
rect 212876 500198 212918 500434
rect 213154 500198 213196 500434
rect 212876 493434 213196 500198
rect 212876 493198 212918 493434
rect 213154 493198 213196 493434
rect 212876 486434 213196 493198
rect 212876 486198 212918 486434
rect 213154 486198 213196 486434
rect 212876 479434 213196 486198
rect 212876 479198 212918 479434
rect 213154 479198 213196 479434
rect 212876 472434 213196 479198
rect 212876 472198 212918 472434
rect 213154 472198 213196 472434
rect 212876 465434 213196 472198
rect 212876 465198 212918 465434
rect 213154 465198 213196 465434
rect 212876 458434 213196 465198
rect 212876 458198 212918 458434
rect 213154 458198 213196 458434
rect 212876 451434 213196 458198
rect 212876 451198 212918 451434
rect 213154 451198 213196 451434
rect 212876 444434 213196 451198
rect 212876 444198 212918 444434
rect 213154 444198 213196 444434
rect 212876 437434 213196 444198
rect 212876 437198 212918 437434
rect 213154 437198 213196 437434
rect 212876 430434 213196 437198
rect 212876 430198 212918 430434
rect 213154 430198 213196 430434
rect 212876 423434 213196 430198
rect 212876 423198 212918 423434
rect 213154 423198 213196 423434
rect 212876 416434 213196 423198
rect 212876 416198 212918 416434
rect 213154 416198 213196 416434
rect 212876 409434 213196 416198
rect 212876 409198 212918 409434
rect 213154 409198 213196 409434
rect 212876 402434 213196 409198
rect 212876 402198 212918 402434
rect 213154 402198 213196 402434
rect 212876 395434 213196 402198
rect 212876 395198 212918 395434
rect 213154 395198 213196 395434
rect 212876 388434 213196 395198
rect 212876 388198 212918 388434
rect 213154 388198 213196 388434
rect 212876 381434 213196 388198
rect 212876 381198 212918 381434
rect 213154 381198 213196 381434
rect 212876 374434 213196 381198
rect 212876 374198 212918 374434
rect 213154 374198 213196 374434
rect 212876 367434 213196 374198
rect 212876 367198 212918 367434
rect 213154 367198 213196 367434
rect 212876 360434 213196 367198
rect 212876 360198 212918 360434
rect 213154 360198 213196 360434
rect 212876 353434 213196 360198
rect 212876 353198 212918 353434
rect 213154 353198 213196 353434
rect 212876 346434 213196 353198
rect 212876 346198 212918 346434
rect 213154 346198 213196 346434
rect 212876 339434 213196 346198
rect 212876 339198 212918 339434
rect 213154 339198 213196 339434
rect 212876 332434 213196 339198
rect 212876 332198 212918 332434
rect 213154 332198 213196 332434
rect 212876 325434 213196 332198
rect 212876 325198 212918 325434
rect 213154 325198 213196 325434
rect 212876 318434 213196 325198
rect 212876 318198 212918 318434
rect 213154 318198 213196 318434
rect 212876 311434 213196 318198
rect 212876 311198 212918 311434
rect 213154 311198 213196 311434
rect 212876 304434 213196 311198
rect 212876 304198 212918 304434
rect 213154 304198 213196 304434
rect 212876 297434 213196 304198
rect 212876 297198 212918 297434
rect 213154 297198 213196 297434
rect 212876 290434 213196 297198
rect 212876 290198 212918 290434
rect 213154 290198 213196 290434
rect 212876 283434 213196 290198
rect 212876 283198 212918 283434
rect 213154 283198 213196 283434
rect 212876 276434 213196 283198
rect 212876 276198 212918 276434
rect 213154 276198 213196 276434
rect 212876 269434 213196 276198
rect 212876 269198 212918 269434
rect 213154 269198 213196 269434
rect 212876 262434 213196 269198
rect 212876 262198 212918 262434
rect 213154 262198 213196 262434
rect 212876 255434 213196 262198
rect 212876 255198 212918 255434
rect 213154 255198 213196 255434
rect 212876 248434 213196 255198
rect 212876 248198 212918 248434
rect 213154 248198 213196 248434
rect 212876 241434 213196 248198
rect 212876 241198 212918 241434
rect 213154 241198 213196 241434
rect 212876 234434 213196 241198
rect 212876 234198 212918 234434
rect 213154 234198 213196 234434
rect 212876 227434 213196 234198
rect 212876 227198 212918 227434
rect 213154 227198 213196 227434
rect 212876 220434 213196 227198
rect 212876 220198 212918 220434
rect 213154 220198 213196 220434
rect 212876 213434 213196 220198
rect 212876 213198 212918 213434
rect 213154 213198 213196 213434
rect 212876 206434 213196 213198
rect 212876 206198 212918 206434
rect 213154 206198 213196 206434
rect 212876 199434 213196 206198
rect 212876 199198 212918 199434
rect 213154 199198 213196 199434
rect 212876 192434 213196 199198
rect 212876 192198 212918 192434
rect 213154 192198 213196 192434
rect 212876 185434 213196 192198
rect 212876 185198 212918 185434
rect 213154 185198 213196 185434
rect 212876 178434 213196 185198
rect 212876 178198 212918 178434
rect 213154 178198 213196 178434
rect 212876 171434 213196 178198
rect 212876 171198 212918 171434
rect 213154 171198 213196 171434
rect 212876 164434 213196 171198
rect 212876 164198 212918 164434
rect 213154 164198 213196 164434
rect 212876 157434 213196 164198
rect 212876 157198 212918 157434
rect 213154 157198 213196 157434
rect 212876 150434 213196 157198
rect 212876 150198 212918 150434
rect 213154 150198 213196 150434
rect 212876 143434 213196 150198
rect 212876 143198 212918 143434
rect 213154 143198 213196 143434
rect 212876 136434 213196 143198
rect 212876 136198 212918 136434
rect 213154 136198 213196 136434
rect 212876 129434 213196 136198
rect 212876 129198 212918 129434
rect 213154 129198 213196 129434
rect 212876 122434 213196 129198
rect 212876 122198 212918 122434
rect 213154 122198 213196 122434
rect 212876 115434 213196 122198
rect 212876 115198 212918 115434
rect 213154 115198 213196 115434
rect 212876 108434 213196 115198
rect 212876 108198 212918 108434
rect 213154 108198 213196 108434
rect 212876 101434 213196 108198
rect 212876 101198 212918 101434
rect 213154 101198 213196 101434
rect 212876 94434 213196 101198
rect 212876 94198 212918 94434
rect 213154 94198 213196 94434
rect 212876 87434 213196 94198
rect 212876 87198 212918 87434
rect 213154 87198 213196 87434
rect 212876 80434 213196 87198
rect 212876 80198 212918 80434
rect 213154 80198 213196 80434
rect 212876 73434 213196 80198
rect 212876 73198 212918 73434
rect 213154 73198 213196 73434
rect 212876 66434 213196 73198
rect 212876 66198 212918 66434
rect 213154 66198 213196 66434
rect 212876 59434 213196 66198
rect 212876 59198 212918 59434
rect 213154 59198 213196 59434
rect 212876 52434 213196 59198
rect 212876 52198 212918 52434
rect 213154 52198 213196 52434
rect 212876 45434 213196 52198
rect 212876 45198 212918 45434
rect 213154 45198 213196 45434
rect 212876 38434 213196 45198
rect 212876 38198 212918 38434
rect 213154 38198 213196 38434
rect 212876 31434 213196 38198
rect 212876 31198 212918 31434
rect 213154 31198 213196 31434
rect 212876 24434 213196 31198
rect 212876 24198 212918 24434
rect 213154 24198 213196 24434
rect 212876 17434 213196 24198
rect 212876 17198 212918 17434
rect 213154 17198 213196 17434
rect 212876 10434 213196 17198
rect 212876 10198 212918 10434
rect 213154 10198 213196 10434
rect 212876 3434 213196 10198
rect 212876 3198 212918 3434
rect 213154 3198 213196 3434
rect 212876 -1706 213196 3198
rect 212876 -1942 212918 -1706
rect 213154 -1942 213196 -1706
rect 212876 -2026 213196 -1942
rect 212876 -2262 212918 -2026
rect 213154 -2262 213196 -2026
rect 212876 -2294 213196 -2262
rect 218144 705238 218464 706230
rect 218144 705002 218186 705238
rect 218422 705002 218464 705238
rect 218144 704918 218464 705002
rect 218144 704682 218186 704918
rect 218422 704682 218464 704918
rect 218144 695494 218464 704682
rect 218144 695258 218186 695494
rect 218422 695258 218464 695494
rect 218144 688494 218464 695258
rect 218144 688258 218186 688494
rect 218422 688258 218464 688494
rect 218144 681494 218464 688258
rect 218144 681258 218186 681494
rect 218422 681258 218464 681494
rect 218144 674494 218464 681258
rect 218144 674258 218186 674494
rect 218422 674258 218464 674494
rect 218144 667494 218464 674258
rect 218144 667258 218186 667494
rect 218422 667258 218464 667494
rect 218144 660494 218464 667258
rect 218144 660258 218186 660494
rect 218422 660258 218464 660494
rect 218144 653494 218464 660258
rect 218144 653258 218186 653494
rect 218422 653258 218464 653494
rect 218144 646494 218464 653258
rect 218144 646258 218186 646494
rect 218422 646258 218464 646494
rect 218144 639494 218464 646258
rect 218144 639258 218186 639494
rect 218422 639258 218464 639494
rect 218144 632494 218464 639258
rect 218144 632258 218186 632494
rect 218422 632258 218464 632494
rect 218144 625494 218464 632258
rect 218144 625258 218186 625494
rect 218422 625258 218464 625494
rect 218144 618494 218464 625258
rect 218144 618258 218186 618494
rect 218422 618258 218464 618494
rect 218144 611494 218464 618258
rect 218144 611258 218186 611494
rect 218422 611258 218464 611494
rect 218144 604494 218464 611258
rect 218144 604258 218186 604494
rect 218422 604258 218464 604494
rect 218144 597494 218464 604258
rect 218144 597258 218186 597494
rect 218422 597258 218464 597494
rect 218144 590494 218464 597258
rect 218144 590258 218186 590494
rect 218422 590258 218464 590494
rect 218144 583494 218464 590258
rect 218144 583258 218186 583494
rect 218422 583258 218464 583494
rect 218144 576494 218464 583258
rect 218144 576258 218186 576494
rect 218422 576258 218464 576494
rect 218144 569494 218464 576258
rect 218144 569258 218186 569494
rect 218422 569258 218464 569494
rect 218144 562494 218464 569258
rect 218144 562258 218186 562494
rect 218422 562258 218464 562494
rect 218144 555494 218464 562258
rect 218144 555258 218186 555494
rect 218422 555258 218464 555494
rect 218144 548494 218464 555258
rect 218144 548258 218186 548494
rect 218422 548258 218464 548494
rect 218144 541494 218464 548258
rect 218144 541258 218186 541494
rect 218422 541258 218464 541494
rect 218144 534494 218464 541258
rect 218144 534258 218186 534494
rect 218422 534258 218464 534494
rect 218144 527494 218464 534258
rect 218144 527258 218186 527494
rect 218422 527258 218464 527494
rect 218144 520494 218464 527258
rect 218144 520258 218186 520494
rect 218422 520258 218464 520494
rect 218144 513494 218464 520258
rect 218144 513258 218186 513494
rect 218422 513258 218464 513494
rect 218144 506494 218464 513258
rect 218144 506258 218186 506494
rect 218422 506258 218464 506494
rect 218144 499494 218464 506258
rect 218144 499258 218186 499494
rect 218422 499258 218464 499494
rect 218144 492494 218464 499258
rect 218144 492258 218186 492494
rect 218422 492258 218464 492494
rect 218144 485494 218464 492258
rect 218144 485258 218186 485494
rect 218422 485258 218464 485494
rect 218144 478494 218464 485258
rect 218144 478258 218186 478494
rect 218422 478258 218464 478494
rect 218144 471494 218464 478258
rect 218144 471258 218186 471494
rect 218422 471258 218464 471494
rect 218144 464494 218464 471258
rect 218144 464258 218186 464494
rect 218422 464258 218464 464494
rect 218144 457494 218464 464258
rect 218144 457258 218186 457494
rect 218422 457258 218464 457494
rect 218144 450494 218464 457258
rect 218144 450258 218186 450494
rect 218422 450258 218464 450494
rect 218144 443494 218464 450258
rect 218144 443258 218186 443494
rect 218422 443258 218464 443494
rect 218144 436494 218464 443258
rect 218144 436258 218186 436494
rect 218422 436258 218464 436494
rect 218144 429494 218464 436258
rect 218144 429258 218186 429494
rect 218422 429258 218464 429494
rect 218144 422494 218464 429258
rect 218144 422258 218186 422494
rect 218422 422258 218464 422494
rect 218144 415494 218464 422258
rect 218144 415258 218186 415494
rect 218422 415258 218464 415494
rect 218144 408494 218464 415258
rect 218144 408258 218186 408494
rect 218422 408258 218464 408494
rect 218144 401494 218464 408258
rect 218144 401258 218186 401494
rect 218422 401258 218464 401494
rect 218144 394494 218464 401258
rect 218144 394258 218186 394494
rect 218422 394258 218464 394494
rect 218144 387494 218464 394258
rect 218144 387258 218186 387494
rect 218422 387258 218464 387494
rect 218144 380494 218464 387258
rect 218144 380258 218186 380494
rect 218422 380258 218464 380494
rect 218144 373494 218464 380258
rect 218144 373258 218186 373494
rect 218422 373258 218464 373494
rect 218144 366494 218464 373258
rect 218144 366258 218186 366494
rect 218422 366258 218464 366494
rect 218144 359494 218464 366258
rect 218144 359258 218186 359494
rect 218422 359258 218464 359494
rect 218144 352494 218464 359258
rect 218144 352258 218186 352494
rect 218422 352258 218464 352494
rect 218144 345494 218464 352258
rect 218144 345258 218186 345494
rect 218422 345258 218464 345494
rect 218144 338494 218464 345258
rect 218144 338258 218186 338494
rect 218422 338258 218464 338494
rect 218144 331494 218464 338258
rect 218144 331258 218186 331494
rect 218422 331258 218464 331494
rect 218144 324494 218464 331258
rect 218144 324258 218186 324494
rect 218422 324258 218464 324494
rect 218144 317494 218464 324258
rect 218144 317258 218186 317494
rect 218422 317258 218464 317494
rect 218144 310494 218464 317258
rect 218144 310258 218186 310494
rect 218422 310258 218464 310494
rect 218144 303494 218464 310258
rect 218144 303258 218186 303494
rect 218422 303258 218464 303494
rect 218144 296494 218464 303258
rect 218144 296258 218186 296494
rect 218422 296258 218464 296494
rect 218144 289494 218464 296258
rect 218144 289258 218186 289494
rect 218422 289258 218464 289494
rect 218144 282494 218464 289258
rect 218144 282258 218186 282494
rect 218422 282258 218464 282494
rect 218144 275494 218464 282258
rect 218144 275258 218186 275494
rect 218422 275258 218464 275494
rect 218144 268494 218464 275258
rect 218144 268258 218186 268494
rect 218422 268258 218464 268494
rect 218144 261494 218464 268258
rect 218144 261258 218186 261494
rect 218422 261258 218464 261494
rect 218144 254494 218464 261258
rect 218144 254258 218186 254494
rect 218422 254258 218464 254494
rect 218144 247494 218464 254258
rect 218144 247258 218186 247494
rect 218422 247258 218464 247494
rect 218144 240494 218464 247258
rect 218144 240258 218186 240494
rect 218422 240258 218464 240494
rect 218144 233494 218464 240258
rect 218144 233258 218186 233494
rect 218422 233258 218464 233494
rect 218144 226494 218464 233258
rect 218144 226258 218186 226494
rect 218422 226258 218464 226494
rect 218144 219494 218464 226258
rect 218144 219258 218186 219494
rect 218422 219258 218464 219494
rect 218144 212494 218464 219258
rect 218144 212258 218186 212494
rect 218422 212258 218464 212494
rect 218144 205494 218464 212258
rect 218144 205258 218186 205494
rect 218422 205258 218464 205494
rect 218144 198494 218464 205258
rect 218144 198258 218186 198494
rect 218422 198258 218464 198494
rect 218144 191494 218464 198258
rect 218144 191258 218186 191494
rect 218422 191258 218464 191494
rect 218144 184494 218464 191258
rect 218144 184258 218186 184494
rect 218422 184258 218464 184494
rect 218144 177494 218464 184258
rect 218144 177258 218186 177494
rect 218422 177258 218464 177494
rect 218144 170494 218464 177258
rect 218144 170258 218186 170494
rect 218422 170258 218464 170494
rect 218144 163494 218464 170258
rect 218144 163258 218186 163494
rect 218422 163258 218464 163494
rect 218144 156494 218464 163258
rect 218144 156258 218186 156494
rect 218422 156258 218464 156494
rect 218144 149494 218464 156258
rect 218144 149258 218186 149494
rect 218422 149258 218464 149494
rect 218144 142494 218464 149258
rect 218144 142258 218186 142494
rect 218422 142258 218464 142494
rect 218144 135494 218464 142258
rect 218144 135258 218186 135494
rect 218422 135258 218464 135494
rect 218144 128494 218464 135258
rect 218144 128258 218186 128494
rect 218422 128258 218464 128494
rect 218144 121494 218464 128258
rect 218144 121258 218186 121494
rect 218422 121258 218464 121494
rect 218144 114494 218464 121258
rect 218144 114258 218186 114494
rect 218422 114258 218464 114494
rect 218144 107494 218464 114258
rect 218144 107258 218186 107494
rect 218422 107258 218464 107494
rect 218144 100494 218464 107258
rect 218144 100258 218186 100494
rect 218422 100258 218464 100494
rect 218144 93494 218464 100258
rect 218144 93258 218186 93494
rect 218422 93258 218464 93494
rect 218144 86494 218464 93258
rect 218144 86258 218186 86494
rect 218422 86258 218464 86494
rect 218144 79494 218464 86258
rect 218144 79258 218186 79494
rect 218422 79258 218464 79494
rect 218144 72494 218464 79258
rect 218144 72258 218186 72494
rect 218422 72258 218464 72494
rect 218144 65494 218464 72258
rect 218144 65258 218186 65494
rect 218422 65258 218464 65494
rect 218144 58494 218464 65258
rect 218144 58258 218186 58494
rect 218422 58258 218464 58494
rect 218144 51494 218464 58258
rect 218144 51258 218186 51494
rect 218422 51258 218464 51494
rect 218144 44494 218464 51258
rect 218144 44258 218186 44494
rect 218422 44258 218464 44494
rect 218144 37494 218464 44258
rect 218144 37258 218186 37494
rect 218422 37258 218464 37494
rect 218144 30494 218464 37258
rect 218144 30258 218186 30494
rect 218422 30258 218464 30494
rect 218144 23494 218464 30258
rect 218144 23258 218186 23494
rect 218422 23258 218464 23494
rect 218144 16494 218464 23258
rect 218144 16258 218186 16494
rect 218422 16258 218464 16494
rect 218144 9494 218464 16258
rect 218144 9258 218186 9494
rect 218422 9258 218464 9494
rect 218144 2494 218464 9258
rect 218144 2258 218186 2494
rect 218422 2258 218464 2494
rect 218144 -746 218464 2258
rect 218144 -982 218186 -746
rect 218422 -982 218464 -746
rect 218144 -1066 218464 -982
rect 218144 -1302 218186 -1066
rect 218422 -1302 218464 -1066
rect 218144 -2294 218464 -1302
rect 219876 706198 220196 706230
rect 219876 705962 219918 706198
rect 220154 705962 220196 706198
rect 219876 705878 220196 705962
rect 219876 705642 219918 705878
rect 220154 705642 220196 705878
rect 219876 696434 220196 705642
rect 219876 696198 219918 696434
rect 220154 696198 220196 696434
rect 219876 689434 220196 696198
rect 219876 689198 219918 689434
rect 220154 689198 220196 689434
rect 219876 682434 220196 689198
rect 219876 682198 219918 682434
rect 220154 682198 220196 682434
rect 219876 675434 220196 682198
rect 219876 675198 219918 675434
rect 220154 675198 220196 675434
rect 219876 668434 220196 675198
rect 219876 668198 219918 668434
rect 220154 668198 220196 668434
rect 219876 661434 220196 668198
rect 219876 661198 219918 661434
rect 220154 661198 220196 661434
rect 219876 654434 220196 661198
rect 219876 654198 219918 654434
rect 220154 654198 220196 654434
rect 219876 647434 220196 654198
rect 219876 647198 219918 647434
rect 220154 647198 220196 647434
rect 219876 640434 220196 647198
rect 219876 640198 219918 640434
rect 220154 640198 220196 640434
rect 219876 633434 220196 640198
rect 219876 633198 219918 633434
rect 220154 633198 220196 633434
rect 219876 626434 220196 633198
rect 219876 626198 219918 626434
rect 220154 626198 220196 626434
rect 219876 619434 220196 626198
rect 219876 619198 219918 619434
rect 220154 619198 220196 619434
rect 219876 612434 220196 619198
rect 219876 612198 219918 612434
rect 220154 612198 220196 612434
rect 219876 605434 220196 612198
rect 219876 605198 219918 605434
rect 220154 605198 220196 605434
rect 219876 598434 220196 605198
rect 219876 598198 219918 598434
rect 220154 598198 220196 598434
rect 219876 591434 220196 598198
rect 219876 591198 219918 591434
rect 220154 591198 220196 591434
rect 219876 584434 220196 591198
rect 219876 584198 219918 584434
rect 220154 584198 220196 584434
rect 219876 577434 220196 584198
rect 219876 577198 219918 577434
rect 220154 577198 220196 577434
rect 219876 570434 220196 577198
rect 219876 570198 219918 570434
rect 220154 570198 220196 570434
rect 219876 563434 220196 570198
rect 219876 563198 219918 563434
rect 220154 563198 220196 563434
rect 219876 556434 220196 563198
rect 219876 556198 219918 556434
rect 220154 556198 220196 556434
rect 219876 549434 220196 556198
rect 219876 549198 219918 549434
rect 220154 549198 220196 549434
rect 219876 542434 220196 549198
rect 219876 542198 219918 542434
rect 220154 542198 220196 542434
rect 219876 535434 220196 542198
rect 219876 535198 219918 535434
rect 220154 535198 220196 535434
rect 219876 528434 220196 535198
rect 219876 528198 219918 528434
rect 220154 528198 220196 528434
rect 219876 521434 220196 528198
rect 219876 521198 219918 521434
rect 220154 521198 220196 521434
rect 219876 514434 220196 521198
rect 219876 514198 219918 514434
rect 220154 514198 220196 514434
rect 219876 507434 220196 514198
rect 219876 507198 219918 507434
rect 220154 507198 220196 507434
rect 219876 500434 220196 507198
rect 219876 500198 219918 500434
rect 220154 500198 220196 500434
rect 219876 493434 220196 500198
rect 219876 493198 219918 493434
rect 220154 493198 220196 493434
rect 219876 486434 220196 493198
rect 219876 486198 219918 486434
rect 220154 486198 220196 486434
rect 219876 479434 220196 486198
rect 219876 479198 219918 479434
rect 220154 479198 220196 479434
rect 219876 472434 220196 479198
rect 219876 472198 219918 472434
rect 220154 472198 220196 472434
rect 219876 465434 220196 472198
rect 219876 465198 219918 465434
rect 220154 465198 220196 465434
rect 219876 458434 220196 465198
rect 219876 458198 219918 458434
rect 220154 458198 220196 458434
rect 219876 451434 220196 458198
rect 219876 451198 219918 451434
rect 220154 451198 220196 451434
rect 219876 444434 220196 451198
rect 219876 444198 219918 444434
rect 220154 444198 220196 444434
rect 219876 437434 220196 444198
rect 219876 437198 219918 437434
rect 220154 437198 220196 437434
rect 219876 430434 220196 437198
rect 219876 430198 219918 430434
rect 220154 430198 220196 430434
rect 219876 423434 220196 430198
rect 219876 423198 219918 423434
rect 220154 423198 220196 423434
rect 219876 416434 220196 423198
rect 219876 416198 219918 416434
rect 220154 416198 220196 416434
rect 219876 409434 220196 416198
rect 219876 409198 219918 409434
rect 220154 409198 220196 409434
rect 219876 402434 220196 409198
rect 219876 402198 219918 402434
rect 220154 402198 220196 402434
rect 219876 395434 220196 402198
rect 219876 395198 219918 395434
rect 220154 395198 220196 395434
rect 219876 388434 220196 395198
rect 219876 388198 219918 388434
rect 220154 388198 220196 388434
rect 219876 381434 220196 388198
rect 219876 381198 219918 381434
rect 220154 381198 220196 381434
rect 219876 374434 220196 381198
rect 219876 374198 219918 374434
rect 220154 374198 220196 374434
rect 219876 367434 220196 374198
rect 219876 367198 219918 367434
rect 220154 367198 220196 367434
rect 219876 360434 220196 367198
rect 219876 360198 219918 360434
rect 220154 360198 220196 360434
rect 219876 353434 220196 360198
rect 219876 353198 219918 353434
rect 220154 353198 220196 353434
rect 219876 346434 220196 353198
rect 219876 346198 219918 346434
rect 220154 346198 220196 346434
rect 219876 339434 220196 346198
rect 219876 339198 219918 339434
rect 220154 339198 220196 339434
rect 219876 332434 220196 339198
rect 219876 332198 219918 332434
rect 220154 332198 220196 332434
rect 219876 325434 220196 332198
rect 219876 325198 219918 325434
rect 220154 325198 220196 325434
rect 219876 318434 220196 325198
rect 219876 318198 219918 318434
rect 220154 318198 220196 318434
rect 219876 311434 220196 318198
rect 219876 311198 219918 311434
rect 220154 311198 220196 311434
rect 219876 304434 220196 311198
rect 219876 304198 219918 304434
rect 220154 304198 220196 304434
rect 219876 297434 220196 304198
rect 219876 297198 219918 297434
rect 220154 297198 220196 297434
rect 219876 290434 220196 297198
rect 219876 290198 219918 290434
rect 220154 290198 220196 290434
rect 219876 283434 220196 290198
rect 219876 283198 219918 283434
rect 220154 283198 220196 283434
rect 219876 276434 220196 283198
rect 219876 276198 219918 276434
rect 220154 276198 220196 276434
rect 219876 269434 220196 276198
rect 219876 269198 219918 269434
rect 220154 269198 220196 269434
rect 219876 262434 220196 269198
rect 219876 262198 219918 262434
rect 220154 262198 220196 262434
rect 219876 255434 220196 262198
rect 219876 255198 219918 255434
rect 220154 255198 220196 255434
rect 219876 248434 220196 255198
rect 219876 248198 219918 248434
rect 220154 248198 220196 248434
rect 219876 241434 220196 248198
rect 219876 241198 219918 241434
rect 220154 241198 220196 241434
rect 219876 234434 220196 241198
rect 219876 234198 219918 234434
rect 220154 234198 220196 234434
rect 219876 227434 220196 234198
rect 219876 227198 219918 227434
rect 220154 227198 220196 227434
rect 219876 220434 220196 227198
rect 219876 220198 219918 220434
rect 220154 220198 220196 220434
rect 219876 213434 220196 220198
rect 219876 213198 219918 213434
rect 220154 213198 220196 213434
rect 219876 206434 220196 213198
rect 219876 206198 219918 206434
rect 220154 206198 220196 206434
rect 219876 199434 220196 206198
rect 219876 199198 219918 199434
rect 220154 199198 220196 199434
rect 219876 192434 220196 199198
rect 219876 192198 219918 192434
rect 220154 192198 220196 192434
rect 219876 185434 220196 192198
rect 219876 185198 219918 185434
rect 220154 185198 220196 185434
rect 219876 178434 220196 185198
rect 219876 178198 219918 178434
rect 220154 178198 220196 178434
rect 219876 171434 220196 178198
rect 219876 171198 219918 171434
rect 220154 171198 220196 171434
rect 219876 164434 220196 171198
rect 219876 164198 219918 164434
rect 220154 164198 220196 164434
rect 219876 157434 220196 164198
rect 219876 157198 219918 157434
rect 220154 157198 220196 157434
rect 219876 150434 220196 157198
rect 219876 150198 219918 150434
rect 220154 150198 220196 150434
rect 219876 143434 220196 150198
rect 219876 143198 219918 143434
rect 220154 143198 220196 143434
rect 219876 136434 220196 143198
rect 219876 136198 219918 136434
rect 220154 136198 220196 136434
rect 219876 129434 220196 136198
rect 219876 129198 219918 129434
rect 220154 129198 220196 129434
rect 219876 122434 220196 129198
rect 219876 122198 219918 122434
rect 220154 122198 220196 122434
rect 219876 115434 220196 122198
rect 219876 115198 219918 115434
rect 220154 115198 220196 115434
rect 219876 108434 220196 115198
rect 219876 108198 219918 108434
rect 220154 108198 220196 108434
rect 219876 101434 220196 108198
rect 219876 101198 219918 101434
rect 220154 101198 220196 101434
rect 219876 94434 220196 101198
rect 219876 94198 219918 94434
rect 220154 94198 220196 94434
rect 219876 87434 220196 94198
rect 219876 87198 219918 87434
rect 220154 87198 220196 87434
rect 219876 80434 220196 87198
rect 219876 80198 219918 80434
rect 220154 80198 220196 80434
rect 219876 73434 220196 80198
rect 219876 73198 219918 73434
rect 220154 73198 220196 73434
rect 219876 66434 220196 73198
rect 219876 66198 219918 66434
rect 220154 66198 220196 66434
rect 219876 59434 220196 66198
rect 219876 59198 219918 59434
rect 220154 59198 220196 59434
rect 219876 52434 220196 59198
rect 219876 52198 219918 52434
rect 220154 52198 220196 52434
rect 219876 45434 220196 52198
rect 219876 45198 219918 45434
rect 220154 45198 220196 45434
rect 219876 38434 220196 45198
rect 219876 38198 219918 38434
rect 220154 38198 220196 38434
rect 219876 31434 220196 38198
rect 219876 31198 219918 31434
rect 220154 31198 220196 31434
rect 219876 24434 220196 31198
rect 219876 24198 219918 24434
rect 220154 24198 220196 24434
rect 219876 17434 220196 24198
rect 219876 17198 219918 17434
rect 220154 17198 220196 17434
rect 219876 10434 220196 17198
rect 219876 10198 219918 10434
rect 220154 10198 220196 10434
rect 219876 3434 220196 10198
rect 219876 3198 219918 3434
rect 220154 3198 220196 3434
rect 219876 -1706 220196 3198
rect 219876 -1942 219918 -1706
rect 220154 -1942 220196 -1706
rect 219876 -2026 220196 -1942
rect 219876 -2262 219918 -2026
rect 220154 -2262 220196 -2026
rect 219876 -2294 220196 -2262
rect 225144 705238 225464 706230
rect 225144 705002 225186 705238
rect 225422 705002 225464 705238
rect 225144 704918 225464 705002
rect 225144 704682 225186 704918
rect 225422 704682 225464 704918
rect 225144 695494 225464 704682
rect 225144 695258 225186 695494
rect 225422 695258 225464 695494
rect 225144 688494 225464 695258
rect 225144 688258 225186 688494
rect 225422 688258 225464 688494
rect 225144 681494 225464 688258
rect 225144 681258 225186 681494
rect 225422 681258 225464 681494
rect 225144 674494 225464 681258
rect 225144 674258 225186 674494
rect 225422 674258 225464 674494
rect 225144 667494 225464 674258
rect 225144 667258 225186 667494
rect 225422 667258 225464 667494
rect 225144 660494 225464 667258
rect 225144 660258 225186 660494
rect 225422 660258 225464 660494
rect 225144 653494 225464 660258
rect 225144 653258 225186 653494
rect 225422 653258 225464 653494
rect 225144 646494 225464 653258
rect 225144 646258 225186 646494
rect 225422 646258 225464 646494
rect 225144 639494 225464 646258
rect 225144 639258 225186 639494
rect 225422 639258 225464 639494
rect 225144 632494 225464 639258
rect 225144 632258 225186 632494
rect 225422 632258 225464 632494
rect 225144 625494 225464 632258
rect 225144 625258 225186 625494
rect 225422 625258 225464 625494
rect 225144 618494 225464 625258
rect 225144 618258 225186 618494
rect 225422 618258 225464 618494
rect 225144 611494 225464 618258
rect 225144 611258 225186 611494
rect 225422 611258 225464 611494
rect 225144 604494 225464 611258
rect 225144 604258 225186 604494
rect 225422 604258 225464 604494
rect 225144 597494 225464 604258
rect 225144 597258 225186 597494
rect 225422 597258 225464 597494
rect 225144 590494 225464 597258
rect 225144 590258 225186 590494
rect 225422 590258 225464 590494
rect 225144 583494 225464 590258
rect 225144 583258 225186 583494
rect 225422 583258 225464 583494
rect 225144 576494 225464 583258
rect 225144 576258 225186 576494
rect 225422 576258 225464 576494
rect 225144 569494 225464 576258
rect 225144 569258 225186 569494
rect 225422 569258 225464 569494
rect 225144 562494 225464 569258
rect 225144 562258 225186 562494
rect 225422 562258 225464 562494
rect 225144 555494 225464 562258
rect 225144 555258 225186 555494
rect 225422 555258 225464 555494
rect 225144 548494 225464 555258
rect 225144 548258 225186 548494
rect 225422 548258 225464 548494
rect 225144 541494 225464 548258
rect 225144 541258 225186 541494
rect 225422 541258 225464 541494
rect 225144 534494 225464 541258
rect 225144 534258 225186 534494
rect 225422 534258 225464 534494
rect 225144 527494 225464 534258
rect 225144 527258 225186 527494
rect 225422 527258 225464 527494
rect 225144 520494 225464 527258
rect 225144 520258 225186 520494
rect 225422 520258 225464 520494
rect 225144 513494 225464 520258
rect 225144 513258 225186 513494
rect 225422 513258 225464 513494
rect 225144 506494 225464 513258
rect 225144 506258 225186 506494
rect 225422 506258 225464 506494
rect 225144 499494 225464 506258
rect 225144 499258 225186 499494
rect 225422 499258 225464 499494
rect 225144 492494 225464 499258
rect 225144 492258 225186 492494
rect 225422 492258 225464 492494
rect 225144 485494 225464 492258
rect 225144 485258 225186 485494
rect 225422 485258 225464 485494
rect 225144 478494 225464 485258
rect 225144 478258 225186 478494
rect 225422 478258 225464 478494
rect 225144 471494 225464 478258
rect 225144 471258 225186 471494
rect 225422 471258 225464 471494
rect 225144 464494 225464 471258
rect 225144 464258 225186 464494
rect 225422 464258 225464 464494
rect 225144 457494 225464 464258
rect 225144 457258 225186 457494
rect 225422 457258 225464 457494
rect 225144 450494 225464 457258
rect 225144 450258 225186 450494
rect 225422 450258 225464 450494
rect 225144 443494 225464 450258
rect 225144 443258 225186 443494
rect 225422 443258 225464 443494
rect 225144 436494 225464 443258
rect 225144 436258 225186 436494
rect 225422 436258 225464 436494
rect 225144 429494 225464 436258
rect 225144 429258 225186 429494
rect 225422 429258 225464 429494
rect 225144 422494 225464 429258
rect 225144 422258 225186 422494
rect 225422 422258 225464 422494
rect 225144 415494 225464 422258
rect 225144 415258 225186 415494
rect 225422 415258 225464 415494
rect 225144 408494 225464 415258
rect 225144 408258 225186 408494
rect 225422 408258 225464 408494
rect 225144 401494 225464 408258
rect 225144 401258 225186 401494
rect 225422 401258 225464 401494
rect 225144 394494 225464 401258
rect 225144 394258 225186 394494
rect 225422 394258 225464 394494
rect 225144 387494 225464 394258
rect 225144 387258 225186 387494
rect 225422 387258 225464 387494
rect 225144 380494 225464 387258
rect 225144 380258 225186 380494
rect 225422 380258 225464 380494
rect 225144 373494 225464 380258
rect 225144 373258 225186 373494
rect 225422 373258 225464 373494
rect 225144 366494 225464 373258
rect 225144 366258 225186 366494
rect 225422 366258 225464 366494
rect 225144 359494 225464 366258
rect 225144 359258 225186 359494
rect 225422 359258 225464 359494
rect 225144 352494 225464 359258
rect 225144 352258 225186 352494
rect 225422 352258 225464 352494
rect 225144 345494 225464 352258
rect 225144 345258 225186 345494
rect 225422 345258 225464 345494
rect 225144 338494 225464 345258
rect 225144 338258 225186 338494
rect 225422 338258 225464 338494
rect 225144 331494 225464 338258
rect 225144 331258 225186 331494
rect 225422 331258 225464 331494
rect 225144 324494 225464 331258
rect 225144 324258 225186 324494
rect 225422 324258 225464 324494
rect 225144 317494 225464 324258
rect 225144 317258 225186 317494
rect 225422 317258 225464 317494
rect 225144 310494 225464 317258
rect 225144 310258 225186 310494
rect 225422 310258 225464 310494
rect 225144 303494 225464 310258
rect 225144 303258 225186 303494
rect 225422 303258 225464 303494
rect 225144 296494 225464 303258
rect 225144 296258 225186 296494
rect 225422 296258 225464 296494
rect 225144 289494 225464 296258
rect 225144 289258 225186 289494
rect 225422 289258 225464 289494
rect 225144 282494 225464 289258
rect 225144 282258 225186 282494
rect 225422 282258 225464 282494
rect 225144 275494 225464 282258
rect 225144 275258 225186 275494
rect 225422 275258 225464 275494
rect 225144 268494 225464 275258
rect 225144 268258 225186 268494
rect 225422 268258 225464 268494
rect 225144 261494 225464 268258
rect 225144 261258 225186 261494
rect 225422 261258 225464 261494
rect 225144 254494 225464 261258
rect 225144 254258 225186 254494
rect 225422 254258 225464 254494
rect 225144 247494 225464 254258
rect 225144 247258 225186 247494
rect 225422 247258 225464 247494
rect 225144 240494 225464 247258
rect 225144 240258 225186 240494
rect 225422 240258 225464 240494
rect 225144 233494 225464 240258
rect 225144 233258 225186 233494
rect 225422 233258 225464 233494
rect 225144 226494 225464 233258
rect 225144 226258 225186 226494
rect 225422 226258 225464 226494
rect 225144 219494 225464 226258
rect 225144 219258 225186 219494
rect 225422 219258 225464 219494
rect 225144 212494 225464 219258
rect 225144 212258 225186 212494
rect 225422 212258 225464 212494
rect 225144 205494 225464 212258
rect 225144 205258 225186 205494
rect 225422 205258 225464 205494
rect 225144 198494 225464 205258
rect 225144 198258 225186 198494
rect 225422 198258 225464 198494
rect 225144 191494 225464 198258
rect 225144 191258 225186 191494
rect 225422 191258 225464 191494
rect 225144 184494 225464 191258
rect 225144 184258 225186 184494
rect 225422 184258 225464 184494
rect 225144 177494 225464 184258
rect 225144 177258 225186 177494
rect 225422 177258 225464 177494
rect 225144 170494 225464 177258
rect 225144 170258 225186 170494
rect 225422 170258 225464 170494
rect 225144 163494 225464 170258
rect 225144 163258 225186 163494
rect 225422 163258 225464 163494
rect 225144 156494 225464 163258
rect 225144 156258 225186 156494
rect 225422 156258 225464 156494
rect 225144 149494 225464 156258
rect 225144 149258 225186 149494
rect 225422 149258 225464 149494
rect 225144 142494 225464 149258
rect 225144 142258 225186 142494
rect 225422 142258 225464 142494
rect 225144 135494 225464 142258
rect 225144 135258 225186 135494
rect 225422 135258 225464 135494
rect 225144 128494 225464 135258
rect 225144 128258 225186 128494
rect 225422 128258 225464 128494
rect 225144 121494 225464 128258
rect 225144 121258 225186 121494
rect 225422 121258 225464 121494
rect 225144 114494 225464 121258
rect 225144 114258 225186 114494
rect 225422 114258 225464 114494
rect 225144 107494 225464 114258
rect 225144 107258 225186 107494
rect 225422 107258 225464 107494
rect 225144 100494 225464 107258
rect 225144 100258 225186 100494
rect 225422 100258 225464 100494
rect 225144 93494 225464 100258
rect 225144 93258 225186 93494
rect 225422 93258 225464 93494
rect 225144 86494 225464 93258
rect 225144 86258 225186 86494
rect 225422 86258 225464 86494
rect 225144 79494 225464 86258
rect 225144 79258 225186 79494
rect 225422 79258 225464 79494
rect 225144 72494 225464 79258
rect 225144 72258 225186 72494
rect 225422 72258 225464 72494
rect 225144 65494 225464 72258
rect 225144 65258 225186 65494
rect 225422 65258 225464 65494
rect 225144 58494 225464 65258
rect 225144 58258 225186 58494
rect 225422 58258 225464 58494
rect 225144 51494 225464 58258
rect 225144 51258 225186 51494
rect 225422 51258 225464 51494
rect 225144 44494 225464 51258
rect 225144 44258 225186 44494
rect 225422 44258 225464 44494
rect 225144 37494 225464 44258
rect 225144 37258 225186 37494
rect 225422 37258 225464 37494
rect 225144 30494 225464 37258
rect 225144 30258 225186 30494
rect 225422 30258 225464 30494
rect 225144 23494 225464 30258
rect 225144 23258 225186 23494
rect 225422 23258 225464 23494
rect 225144 16494 225464 23258
rect 225144 16258 225186 16494
rect 225422 16258 225464 16494
rect 225144 9494 225464 16258
rect 225144 9258 225186 9494
rect 225422 9258 225464 9494
rect 225144 2494 225464 9258
rect 225144 2258 225186 2494
rect 225422 2258 225464 2494
rect 225144 -746 225464 2258
rect 225144 -982 225186 -746
rect 225422 -982 225464 -746
rect 225144 -1066 225464 -982
rect 225144 -1302 225186 -1066
rect 225422 -1302 225464 -1066
rect 225144 -2294 225464 -1302
rect 226876 706198 227196 706230
rect 226876 705962 226918 706198
rect 227154 705962 227196 706198
rect 226876 705878 227196 705962
rect 226876 705642 226918 705878
rect 227154 705642 227196 705878
rect 226876 696434 227196 705642
rect 226876 696198 226918 696434
rect 227154 696198 227196 696434
rect 226876 689434 227196 696198
rect 226876 689198 226918 689434
rect 227154 689198 227196 689434
rect 226876 682434 227196 689198
rect 226876 682198 226918 682434
rect 227154 682198 227196 682434
rect 226876 675434 227196 682198
rect 226876 675198 226918 675434
rect 227154 675198 227196 675434
rect 226876 668434 227196 675198
rect 226876 668198 226918 668434
rect 227154 668198 227196 668434
rect 226876 661434 227196 668198
rect 226876 661198 226918 661434
rect 227154 661198 227196 661434
rect 226876 654434 227196 661198
rect 226876 654198 226918 654434
rect 227154 654198 227196 654434
rect 226876 647434 227196 654198
rect 226876 647198 226918 647434
rect 227154 647198 227196 647434
rect 226876 640434 227196 647198
rect 226876 640198 226918 640434
rect 227154 640198 227196 640434
rect 226876 633434 227196 640198
rect 226876 633198 226918 633434
rect 227154 633198 227196 633434
rect 226876 626434 227196 633198
rect 226876 626198 226918 626434
rect 227154 626198 227196 626434
rect 226876 619434 227196 626198
rect 226876 619198 226918 619434
rect 227154 619198 227196 619434
rect 226876 612434 227196 619198
rect 226876 612198 226918 612434
rect 227154 612198 227196 612434
rect 226876 605434 227196 612198
rect 226876 605198 226918 605434
rect 227154 605198 227196 605434
rect 226876 598434 227196 605198
rect 226876 598198 226918 598434
rect 227154 598198 227196 598434
rect 226876 591434 227196 598198
rect 226876 591198 226918 591434
rect 227154 591198 227196 591434
rect 226876 584434 227196 591198
rect 226876 584198 226918 584434
rect 227154 584198 227196 584434
rect 226876 577434 227196 584198
rect 226876 577198 226918 577434
rect 227154 577198 227196 577434
rect 226876 570434 227196 577198
rect 226876 570198 226918 570434
rect 227154 570198 227196 570434
rect 226876 563434 227196 570198
rect 226876 563198 226918 563434
rect 227154 563198 227196 563434
rect 226876 556434 227196 563198
rect 226876 556198 226918 556434
rect 227154 556198 227196 556434
rect 226876 549434 227196 556198
rect 226876 549198 226918 549434
rect 227154 549198 227196 549434
rect 226876 542434 227196 549198
rect 226876 542198 226918 542434
rect 227154 542198 227196 542434
rect 226876 535434 227196 542198
rect 226876 535198 226918 535434
rect 227154 535198 227196 535434
rect 226876 528434 227196 535198
rect 226876 528198 226918 528434
rect 227154 528198 227196 528434
rect 226876 521434 227196 528198
rect 226876 521198 226918 521434
rect 227154 521198 227196 521434
rect 226876 514434 227196 521198
rect 226876 514198 226918 514434
rect 227154 514198 227196 514434
rect 226876 507434 227196 514198
rect 226876 507198 226918 507434
rect 227154 507198 227196 507434
rect 226876 500434 227196 507198
rect 226876 500198 226918 500434
rect 227154 500198 227196 500434
rect 226876 493434 227196 500198
rect 226876 493198 226918 493434
rect 227154 493198 227196 493434
rect 226876 486434 227196 493198
rect 226876 486198 226918 486434
rect 227154 486198 227196 486434
rect 226876 479434 227196 486198
rect 226876 479198 226918 479434
rect 227154 479198 227196 479434
rect 226876 472434 227196 479198
rect 226876 472198 226918 472434
rect 227154 472198 227196 472434
rect 226876 465434 227196 472198
rect 226876 465198 226918 465434
rect 227154 465198 227196 465434
rect 226876 458434 227196 465198
rect 226876 458198 226918 458434
rect 227154 458198 227196 458434
rect 226876 451434 227196 458198
rect 226876 451198 226918 451434
rect 227154 451198 227196 451434
rect 226876 444434 227196 451198
rect 226876 444198 226918 444434
rect 227154 444198 227196 444434
rect 226876 437434 227196 444198
rect 226876 437198 226918 437434
rect 227154 437198 227196 437434
rect 226876 430434 227196 437198
rect 226876 430198 226918 430434
rect 227154 430198 227196 430434
rect 226876 423434 227196 430198
rect 226876 423198 226918 423434
rect 227154 423198 227196 423434
rect 226876 416434 227196 423198
rect 226876 416198 226918 416434
rect 227154 416198 227196 416434
rect 226876 409434 227196 416198
rect 226876 409198 226918 409434
rect 227154 409198 227196 409434
rect 226876 402434 227196 409198
rect 226876 402198 226918 402434
rect 227154 402198 227196 402434
rect 226876 395434 227196 402198
rect 226876 395198 226918 395434
rect 227154 395198 227196 395434
rect 226876 388434 227196 395198
rect 226876 388198 226918 388434
rect 227154 388198 227196 388434
rect 226876 381434 227196 388198
rect 226876 381198 226918 381434
rect 227154 381198 227196 381434
rect 226876 374434 227196 381198
rect 226876 374198 226918 374434
rect 227154 374198 227196 374434
rect 226876 367434 227196 374198
rect 226876 367198 226918 367434
rect 227154 367198 227196 367434
rect 226876 360434 227196 367198
rect 226876 360198 226918 360434
rect 227154 360198 227196 360434
rect 226876 353434 227196 360198
rect 226876 353198 226918 353434
rect 227154 353198 227196 353434
rect 226876 346434 227196 353198
rect 226876 346198 226918 346434
rect 227154 346198 227196 346434
rect 226876 339434 227196 346198
rect 226876 339198 226918 339434
rect 227154 339198 227196 339434
rect 226876 332434 227196 339198
rect 226876 332198 226918 332434
rect 227154 332198 227196 332434
rect 226876 325434 227196 332198
rect 226876 325198 226918 325434
rect 227154 325198 227196 325434
rect 226876 318434 227196 325198
rect 226876 318198 226918 318434
rect 227154 318198 227196 318434
rect 226876 311434 227196 318198
rect 226876 311198 226918 311434
rect 227154 311198 227196 311434
rect 226876 304434 227196 311198
rect 226876 304198 226918 304434
rect 227154 304198 227196 304434
rect 226876 297434 227196 304198
rect 226876 297198 226918 297434
rect 227154 297198 227196 297434
rect 226876 290434 227196 297198
rect 226876 290198 226918 290434
rect 227154 290198 227196 290434
rect 226876 283434 227196 290198
rect 226876 283198 226918 283434
rect 227154 283198 227196 283434
rect 226876 276434 227196 283198
rect 226876 276198 226918 276434
rect 227154 276198 227196 276434
rect 226876 269434 227196 276198
rect 226876 269198 226918 269434
rect 227154 269198 227196 269434
rect 226876 262434 227196 269198
rect 226876 262198 226918 262434
rect 227154 262198 227196 262434
rect 226876 255434 227196 262198
rect 226876 255198 226918 255434
rect 227154 255198 227196 255434
rect 226876 248434 227196 255198
rect 226876 248198 226918 248434
rect 227154 248198 227196 248434
rect 226876 241434 227196 248198
rect 226876 241198 226918 241434
rect 227154 241198 227196 241434
rect 226876 234434 227196 241198
rect 226876 234198 226918 234434
rect 227154 234198 227196 234434
rect 226876 227434 227196 234198
rect 226876 227198 226918 227434
rect 227154 227198 227196 227434
rect 226876 220434 227196 227198
rect 226876 220198 226918 220434
rect 227154 220198 227196 220434
rect 226876 213434 227196 220198
rect 226876 213198 226918 213434
rect 227154 213198 227196 213434
rect 226876 206434 227196 213198
rect 226876 206198 226918 206434
rect 227154 206198 227196 206434
rect 226876 199434 227196 206198
rect 226876 199198 226918 199434
rect 227154 199198 227196 199434
rect 226876 192434 227196 199198
rect 226876 192198 226918 192434
rect 227154 192198 227196 192434
rect 226876 185434 227196 192198
rect 226876 185198 226918 185434
rect 227154 185198 227196 185434
rect 226876 178434 227196 185198
rect 226876 178198 226918 178434
rect 227154 178198 227196 178434
rect 226876 171434 227196 178198
rect 226876 171198 226918 171434
rect 227154 171198 227196 171434
rect 226876 164434 227196 171198
rect 226876 164198 226918 164434
rect 227154 164198 227196 164434
rect 226876 157434 227196 164198
rect 226876 157198 226918 157434
rect 227154 157198 227196 157434
rect 226876 150434 227196 157198
rect 226876 150198 226918 150434
rect 227154 150198 227196 150434
rect 226876 143434 227196 150198
rect 226876 143198 226918 143434
rect 227154 143198 227196 143434
rect 226876 136434 227196 143198
rect 226876 136198 226918 136434
rect 227154 136198 227196 136434
rect 226876 129434 227196 136198
rect 226876 129198 226918 129434
rect 227154 129198 227196 129434
rect 226876 122434 227196 129198
rect 226876 122198 226918 122434
rect 227154 122198 227196 122434
rect 226876 115434 227196 122198
rect 226876 115198 226918 115434
rect 227154 115198 227196 115434
rect 226876 108434 227196 115198
rect 226876 108198 226918 108434
rect 227154 108198 227196 108434
rect 226876 101434 227196 108198
rect 226876 101198 226918 101434
rect 227154 101198 227196 101434
rect 226876 94434 227196 101198
rect 226876 94198 226918 94434
rect 227154 94198 227196 94434
rect 226876 87434 227196 94198
rect 226876 87198 226918 87434
rect 227154 87198 227196 87434
rect 226876 80434 227196 87198
rect 226876 80198 226918 80434
rect 227154 80198 227196 80434
rect 226876 73434 227196 80198
rect 226876 73198 226918 73434
rect 227154 73198 227196 73434
rect 226876 66434 227196 73198
rect 226876 66198 226918 66434
rect 227154 66198 227196 66434
rect 226876 59434 227196 66198
rect 226876 59198 226918 59434
rect 227154 59198 227196 59434
rect 226876 52434 227196 59198
rect 226876 52198 226918 52434
rect 227154 52198 227196 52434
rect 226876 45434 227196 52198
rect 226876 45198 226918 45434
rect 227154 45198 227196 45434
rect 226876 38434 227196 45198
rect 226876 38198 226918 38434
rect 227154 38198 227196 38434
rect 226876 31434 227196 38198
rect 226876 31198 226918 31434
rect 227154 31198 227196 31434
rect 226876 24434 227196 31198
rect 226876 24198 226918 24434
rect 227154 24198 227196 24434
rect 226876 17434 227196 24198
rect 226876 17198 226918 17434
rect 227154 17198 227196 17434
rect 226876 10434 227196 17198
rect 226876 10198 226918 10434
rect 227154 10198 227196 10434
rect 226876 3434 227196 10198
rect 226876 3198 226918 3434
rect 227154 3198 227196 3434
rect 226876 -1706 227196 3198
rect 226876 -1942 226918 -1706
rect 227154 -1942 227196 -1706
rect 226876 -2026 227196 -1942
rect 226876 -2262 226918 -2026
rect 227154 -2262 227196 -2026
rect 226876 -2294 227196 -2262
rect 232144 705238 232464 706230
rect 232144 705002 232186 705238
rect 232422 705002 232464 705238
rect 232144 704918 232464 705002
rect 232144 704682 232186 704918
rect 232422 704682 232464 704918
rect 232144 695494 232464 704682
rect 232144 695258 232186 695494
rect 232422 695258 232464 695494
rect 232144 688494 232464 695258
rect 232144 688258 232186 688494
rect 232422 688258 232464 688494
rect 232144 681494 232464 688258
rect 232144 681258 232186 681494
rect 232422 681258 232464 681494
rect 232144 674494 232464 681258
rect 232144 674258 232186 674494
rect 232422 674258 232464 674494
rect 232144 667494 232464 674258
rect 232144 667258 232186 667494
rect 232422 667258 232464 667494
rect 232144 660494 232464 667258
rect 232144 660258 232186 660494
rect 232422 660258 232464 660494
rect 232144 653494 232464 660258
rect 232144 653258 232186 653494
rect 232422 653258 232464 653494
rect 232144 646494 232464 653258
rect 232144 646258 232186 646494
rect 232422 646258 232464 646494
rect 232144 639494 232464 646258
rect 232144 639258 232186 639494
rect 232422 639258 232464 639494
rect 232144 632494 232464 639258
rect 232144 632258 232186 632494
rect 232422 632258 232464 632494
rect 232144 625494 232464 632258
rect 232144 625258 232186 625494
rect 232422 625258 232464 625494
rect 232144 618494 232464 625258
rect 232144 618258 232186 618494
rect 232422 618258 232464 618494
rect 232144 611494 232464 618258
rect 232144 611258 232186 611494
rect 232422 611258 232464 611494
rect 232144 604494 232464 611258
rect 232144 604258 232186 604494
rect 232422 604258 232464 604494
rect 232144 597494 232464 604258
rect 232144 597258 232186 597494
rect 232422 597258 232464 597494
rect 232144 590494 232464 597258
rect 232144 590258 232186 590494
rect 232422 590258 232464 590494
rect 232144 583494 232464 590258
rect 232144 583258 232186 583494
rect 232422 583258 232464 583494
rect 232144 576494 232464 583258
rect 232144 576258 232186 576494
rect 232422 576258 232464 576494
rect 232144 569494 232464 576258
rect 232144 569258 232186 569494
rect 232422 569258 232464 569494
rect 232144 562494 232464 569258
rect 232144 562258 232186 562494
rect 232422 562258 232464 562494
rect 232144 555494 232464 562258
rect 232144 555258 232186 555494
rect 232422 555258 232464 555494
rect 232144 548494 232464 555258
rect 232144 548258 232186 548494
rect 232422 548258 232464 548494
rect 232144 541494 232464 548258
rect 232144 541258 232186 541494
rect 232422 541258 232464 541494
rect 232144 534494 232464 541258
rect 232144 534258 232186 534494
rect 232422 534258 232464 534494
rect 232144 527494 232464 534258
rect 232144 527258 232186 527494
rect 232422 527258 232464 527494
rect 232144 520494 232464 527258
rect 232144 520258 232186 520494
rect 232422 520258 232464 520494
rect 232144 513494 232464 520258
rect 232144 513258 232186 513494
rect 232422 513258 232464 513494
rect 232144 506494 232464 513258
rect 232144 506258 232186 506494
rect 232422 506258 232464 506494
rect 232144 499494 232464 506258
rect 232144 499258 232186 499494
rect 232422 499258 232464 499494
rect 232144 492494 232464 499258
rect 232144 492258 232186 492494
rect 232422 492258 232464 492494
rect 232144 485494 232464 492258
rect 232144 485258 232186 485494
rect 232422 485258 232464 485494
rect 232144 478494 232464 485258
rect 232144 478258 232186 478494
rect 232422 478258 232464 478494
rect 232144 471494 232464 478258
rect 232144 471258 232186 471494
rect 232422 471258 232464 471494
rect 232144 464494 232464 471258
rect 232144 464258 232186 464494
rect 232422 464258 232464 464494
rect 232144 457494 232464 464258
rect 232144 457258 232186 457494
rect 232422 457258 232464 457494
rect 232144 450494 232464 457258
rect 232144 450258 232186 450494
rect 232422 450258 232464 450494
rect 232144 443494 232464 450258
rect 232144 443258 232186 443494
rect 232422 443258 232464 443494
rect 232144 436494 232464 443258
rect 232144 436258 232186 436494
rect 232422 436258 232464 436494
rect 232144 429494 232464 436258
rect 232144 429258 232186 429494
rect 232422 429258 232464 429494
rect 232144 422494 232464 429258
rect 232144 422258 232186 422494
rect 232422 422258 232464 422494
rect 232144 415494 232464 422258
rect 232144 415258 232186 415494
rect 232422 415258 232464 415494
rect 232144 408494 232464 415258
rect 232144 408258 232186 408494
rect 232422 408258 232464 408494
rect 232144 401494 232464 408258
rect 232144 401258 232186 401494
rect 232422 401258 232464 401494
rect 232144 394494 232464 401258
rect 232144 394258 232186 394494
rect 232422 394258 232464 394494
rect 232144 387494 232464 394258
rect 232144 387258 232186 387494
rect 232422 387258 232464 387494
rect 232144 380494 232464 387258
rect 232144 380258 232186 380494
rect 232422 380258 232464 380494
rect 232144 373494 232464 380258
rect 232144 373258 232186 373494
rect 232422 373258 232464 373494
rect 232144 366494 232464 373258
rect 232144 366258 232186 366494
rect 232422 366258 232464 366494
rect 232144 359494 232464 366258
rect 232144 359258 232186 359494
rect 232422 359258 232464 359494
rect 232144 352494 232464 359258
rect 232144 352258 232186 352494
rect 232422 352258 232464 352494
rect 232144 345494 232464 352258
rect 232144 345258 232186 345494
rect 232422 345258 232464 345494
rect 232144 338494 232464 345258
rect 232144 338258 232186 338494
rect 232422 338258 232464 338494
rect 232144 331494 232464 338258
rect 232144 331258 232186 331494
rect 232422 331258 232464 331494
rect 232144 324494 232464 331258
rect 232144 324258 232186 324494
rect 232422 324258 232464 324494
rect 232144 317494 232464 324258
rect 232144 317258 232186 317494
rect 232422 317258 232464 317494
rect 232144 310494 232464 317258
rect 232144 310258 232186 310494
rect 232422 310258 232464 310494
rect 232144 303494 232464 310258
rect 232144 303258 232186 303494
rect 232422 303258 232464 303494
rect 232144 296494 232464 303258
rect 232144 296258 232186 296494
rect 232422 296258 232464 296494
rect 232144 289494 232464 296258
rect 232144 289258 232186 289494
rect 232422 289258 232464 289494
rect 232144 282494 232464 289258
rect 232144 282258 232186 282494
rect 232422 282258 232464 282494
rect 232144 275494 232464 282258
rect 232144 275258 232186 275494
rect 232422 275258 232464 275494
rect 232144 268494 232464 275258
rect 232144 268258 232186 268494
rect 232422 268258 232464 268494
rect 232144 261494 232464 268258
rect 232144 261258 232186 261494
rect 232422 261258 232464 261494
rect 232144 254494 232464 261258
rect 232144 254258 232186 254494
rect 232422 254258 232464 254494
rect 232144 247494 232464 254258
rect 232144 247258 232186 247494
rect 232422 247258 232464 247494
rect 232144 240494 232464 247258
rect 232144 240258 232186 240494
rect 232422 240258 232464 240494
rect 232144 233494 232464 240258
rect 232144 233258 232186 233494
rect 232422 233258 232464 233494
rect 232144 226494 232464 233258
rect 232144 226258 232186 226494
rect 232422 226258 232464 226494
rect 232144 219494 232464 226258
rect 232144 219258 232186 219494
rect 232422 219258 232464 219494
rect 232144 212494 232464 219258
rect 232144 212258 232186 212494
rect 232422 212258 232464 212494
rect 232144 205494 232464 212258
rect 232144 205258 232186 205494
rect 232422 205258 232464 205494
rect 232144 198494 232464 205258
rect 232144 198258 232186 198494
rect 232422 198258 232464 198494
rect 232144 191494 232464 198258
rect 232144 191258 232186 191494
rect 232422 191258 232464 191494
rect 232144 184494 232464 191258
rect 232144 184258 232186 184494
rect 232422 184258 232464 184494
rect 232144 177494 232464 184258
rect 232144 177258 232186 177494
rect 232422 177258 232464 177494
rect 232144 170494 232464 177258
rect 232144 170258 232186 170494
rect 232422 170258 232464 170494
rect 232144 163494 232464 170258
rect 232144 163258 232186 163494
rect 232422 163258 232464 163494
rect 232144 156494 232464 163258
rect 232144 156258 232186 156494
rect 232422 156258 232464 156494
rect 232144 149494 232464 156258
rect 232144 149258 232186 149494
rect 232422 149258 232464 149494
rect 232144 142494 232464 149258
rect 232144 142258 232186 142494
rect 232422 142258 232464 142494
rect 232144 135494 232464 142258
rect 232144 135258 232186 135494
rect 232422 135258 232464 135494
rect 232144 128494 232464 135258
rect 232144 128258 232186 128494
rect 232422 128258 232464 128494
rect 232144 121494 232464 128258
rect 232144 121258 232186 121494
rect 232422 121258 232464 121494
rect 232144 114494 232464 121258
rect 232144 114258 232186 114494
rect 232422 114258 232464 114494
rect 232144 107494 232464 114258
rect 232144 107258 232186 107494
rect 232422 107258 232464 107494
rect 232144 100494 232464 107258
rect 232144 100258 232186 100494
rect 232422 100258 232464 100494
rect 232144 93494 232464 100258
rect 232144 93258 232186 93494
rect 232422 93258 232464 93494
rect 232144 86494 232464 93258
rect 232144 86258 232186 86494
rect 232422 86258 232464 86494
rect 232144 79494 232464 86258
rect 232144 79258 232186 79494
rect 232422 79258 232464 79494
rect 232144 72494 232464 79258
rect 232144 72258 232186 72494
rect 232422 72258 232464 72494
rect 232144 65494 232464 72258
rect 232144 65258 232186 65494
rect 232422 65258 232464 65494
rect 232144 58494 232464 65258
rect 232144 58258 232186 58494
rect 232422 58258 232464 58494
rect 232144 51494 232464 58258
rect 232144 51258 232186 51494
rect 232422 51258 232464 51494
rect 232144 44494 232464 51258
rect 232144 44258 232186 44494
rect 232422 44258 232464 44494
rect 232144 37494 232464 44258
rect 232144 37258 232186 37494
rect 232422 37258 232464 37494
rect 232144 30494 232464 37258
rect 232144 30258 232186 30494
rect 232422 30258 232464 30494
rect 232144 23494 232464 30258
rect 232144 23258 232186 23494
rect 232422 23258 232464 23494
rect 232144 16494 232464 23258
rect 232144 16258 232186 16494
rect 232422 16258 232464 16494
rect 232144 9494 232464 16258
rect 232144 9258 232186 9494
rect 232422 9258 232464 9494
rect 232144 2494 232464 9258
rect 232144 2258 232186 2494
rect 232422 2258 232464 2494
rect 232144 -746 232464 2258
rect 232144 -982 232186 -746
rect 232422 -982 232464 -746
rect 232144 -1066 232464 -982
rect 232144 -1302 232186 -1066
rect 232422 -1302 232464 -1066
rect 232144 -2294 232464 -1302
rect 233876 706198 234196 706230
rect 233876 705962 233918 706198
rect 234154 705962 234196 706198
rect 233876 705878 234196 705962
rect 233876 705642 233918 705878
rect 234154 705642 234196 705878
rect 233876 696434 234196 705642
rect 233876 696198 233918 696434
rect 234154 696198 234196 696434
rect 233876 689434 234196 696198
rect 233876 689198 233918 689434
rect 234154 689198 234196 689434
rect 233876 682434 234196 689198
rect 233876 682198 233918 682434
rect 234154 682198 234196 682434
rect 233876 675434 234196 682198
rect 233876 675198 233918 675434
rect 234154 675198 234196 675434
rect 233876 668434 234196 675198
rect 233876 668198 233918 668434
rect 234154 668198 234196 668434
rect 233876 661434 234196 668198
rect 233876 661198 233918 661434
rect 234154 661198 234196 661434
rect 233876 654434 234196 661198
rect 233876 654198 233918 654434
rect 234154 654198 234196 654434
rect 233876 647434 234196 654198
rect 233876 647198 233918 647434
rect 234154 647198 234196 647434
rect 233876 640434 234196 647198
rect 233876 640198 233918 640434
rect 234154 640198 234196 640434
rect 233876 633434 234196 640198
rect 233876 633198 233918 633434
rect 234154 633198 234196 633434
rect 233876 626434 234196 633198
rect 233876 626198 233918 626434
rect 234154 626198 234196 626434
rect 233876 619434 234196 626198
rect 233876 619198 233918 619434
rect 234154 619198 234196 619434
rect 233876 612434 234196 619198
rect 233876 612198 233918 612434
rect 234154 612198 234196 612434
rect 233876 605434 234196 612198
rect 233876 605198 233918 605434
rect 234154 605198 234196 605434
rect 233876 598434 234196 605198
rect 233876 598198 233918 598434
rect 234154 598198 234196 598434
rect 233876 591434 234196 598198
rect 233876 591198 233918 591434
rect 234154 591198 234196 591434
rect 233876 584434 234196 591198
rect 233876 584198 233918 584434
rect 234154 584198 234196 584434
rect 233876 577434 234196 584198
rect 233876 577198 233918 577434
rect 234154 577198 234196 577434
rect 233876 570434 234196 577198
rect 233876 570198 233918 570434
rect 234154 570198 234196 570434
rect 233876 563434 234196 570198
rect 233876 563198 233918 563434
rect 234154 563198 234196 563434
rect 233876 556434 234196 563198
rect 233876 556198 233918 556434
rect 234154 556198 234196 556434
rect 233876 549434 234196 556198
rect 233876 549198 233918 549434
rect 234154 549198 234196 549434
rect 233876 542434 234196 549198
rect 233876 542198 233918 542434
rect 234154 542198 234196 542434
rect 233876 535434 234196 542198
rect 233876 535198 233918 535434
rect 234154 535198 234196 535434
rect 233876 528434 234196 535198
rect 233876 528198 233918 528434
rect 234154 528198 234196 528434
rect 233876 521434 234196 528198
rect 233876 521198 233918 521434
rect 234154 521198 234196 521434
rect 233876 514434 234196 521198
rect 233876 514198 233918 514434
rect 234154 514198 234196 514434
rect 233876 507434 234196 514198
rect 233876 507198 233918 507434
rect 234154 507198 234196 507434
rect 233876 500434 234196 507198
rect 233876 500198 233918 500434
rect 234154 500198 234196 500434
rect 233876 493434 234196 500198
rect 233876 493198 233918 493434
rect 234154 493198 234196 493434
rect 233876 486434 234196 493198
rect 233876 486198 233918 486434
rect 234154 486198 234196 486434
rect 233876 479434 234196 486198
rect 233876 479198 233918 479434
rect 234154 479198 234196 479434
rect 233876 472434 234196 479198
rect 233876 472198 233918 472434
rect 234154 472198 234196 472434
rect 233876 465434 234196 472198
rect 233876 465198 233918 465434
rect 234154 465198 234196 465434
rect 233876 458434 234196 465198
rect 233876 458198 233918 458434
rect 234154 458198 234196 458434
rect 233876 451434 234196 458198
rect 233876 451198 233918 451434
rect 234154 451198 234196 451434
rect 233876 444434 234196 451198
rect 233876 444198 233918 444434
rect 234154 444198 234196 444434
rect 233876 437434 234196 444198
rect 233876 437198 233918 437434
rect 234154 437198 234196 437434
rect 233876 430434 234196 437198
rect 233876 430198 233918 430434
rect 234154 430198 234196 430434
rect 233876 423434 234196 430198
rect 233876 423198 233918 423434
rect 234154 423198 234196 423434
rect 233876 416434 234196 423198
rect 233876 416198 233918 416434
rect 234154 416198 234196 416434
rect 233876 409434 234196 416198
rect 233876 409198 233918 409434
rect 234154 409198 234196 409434
rect 233876 402434 234196 409198
rect 233876 402198 233918 402434
rect 234154 402198 234196 402434
rect 233876 395434 234196 402198
rect 233876 395198 233918 395434
rect 234154 395198 234196 395434
rect 233876 388434 234196 395198
rect 233876 388198 233918 388434
rect 234154 388198 234196 388434
rect 233876 381434 234196 388198
rect 233876 381198 233918 381434
rect 234154 381198 234196 381434
rect 233876 374434 234196 381198
rect 233876 374198 233918 374434
rect 234154 374198 234196 374434
rect 233876 367434 234196 374198
rect 233876 367198 233918 367434
rect 234154 367198 234196 367434
rect 233876 360434 234196 367198
rect 233876 360198 233918 360434
rect 234154 360198 234196 360434
rect 233876 353434 234196 360198
rect 233876 353198 233918 353434
rect 234154 353198 234196 353434
rect 233876 346434 234196 353198
rect 233876 346198 233918 346434
rect 234154 346198 234196 346434
rect 233876 339434 234196 346198
rect 233876 339198 233918 339434
rect 234154 339198 234196 339434
rect 233876 332434 234196 339198
rect 233876 332198 233918 332434
rect 234154 332198 234196 332434
rect 233876 325434 234196 332198
rect 233876 325198 233918 325434
rect 234154 325198 234196 325434
rect 233876 318434 234196 325198
rect 233876 318198 233918 318434
rect 234154 318198 234196 318434
rect 233876 311434 234196 318198
rect 233876 311198 233918 311434
rect 234154 311198 234196 311434
rect 233876 304434 234196 311198
rect 233876 304198 233918 304434
rect 234154 304198 234196 304434
rect 233876 297434 234196 304198
rect 233876 297198 233918 297434
rect 234154 297198 234196 297434
rect 233876 290434 234196 297198
rect 233876 290198 233918 290434
rect 234154 290198 234196 290434
rect 233876 283434 234196 290198
rect 233876 283198 233918 283434
rect 234154 283198 234196 283434
rect 233876 276434 234196 283198
rect 233876 276198 233918 276434
rect 234154 276198 234196 276434
rect 233876 269434 234196 276198
rect 233876 269198 233918 269434
rect 234154 269198 234196 269434
rect 233876 262434 234196 269198
rect 233876 262198 233918 262434
rect 234154 262198 234196 262434
rect 233876 255434 234196 262198
rect 233876 255198 233918 255434
rect 234154 255198 234196 255434
rect 233876 248434 234196 255198
rect 233876 248198 233918 248434
rect 234154 248198 234196 248434
rect 233876 241434 234196 248198
rect 233876 241198 233918 241434
rect 234154 241198 234196 241434
rect 233876 234434 234196 241198
rect 233876 234198 233918 234434
rect 234154 234198 234196 234434
rect 233876 227434 234196 234198
rect 233876 227198 233918 227434
rect 234154 227198 234196 227434
rect 233876 220434 234196 227198
rect 233876 220198 233918 220434
rect 234154 220198 234196 220434
rect 233876 213434 234196 220198
rect 233876 213198 233918 213434
rect 234154 213198 234196 213434
rect 233876 206434 234196 213198
rect 233876 206198 233918 206434
rect 234154 206198 234196 206434
rect 233876 199434 234196 206198
rect 233876 199198 233918 199434
rect 234154 199198 234196 199434
rect 233876 192434 234196 199198
rect 233876 192198 233918 192434
rect 234154 192198 234196 192434
rect 233876 185434 234196 192198
rect 233876 185198 233918 185434
rect 234154 185198 234196 185434
rect 233876 178434 234196 185198
rect 233876 178198 233918 178434
rect 234154 178198 234196 178434
rect 233876 171434 234196 178198
rect 233876 171198 233918 171434
rect 234154 171198 234196 171434
rect 233876 164434 234196 171198
rect 233876 164198 233918 164434
rect 234154 164198 234196 164434
rect 233876 157434 234196 164198
rect 233876 157198 233918 157434
rect 234154 157198 234196 157434
rect 233876 150434 234196 157198
rect 233876 150198 233918 150434
rect 234154 150198 234196 150434
rect 233876 143434 234196 150198
rect 233876 143198 233918 143434
rect 234154 143198 234196 143434
rect 233876 136434 234196 143198
rect 233876 136198 233918 136434
rect 234154 136198 234196 136434
rect 233876 129434 234196 136198
rect 233876 129198 233918 129434
rect 234154 129198 234196 129434
rect 233876 122434 234196 129198
rect 233876 122198 233918 122434
rect 234154 122198 234196 122434
rect 233876 115434 234196 122198
rect 233876 115198 233918 115434
rect 234154 115198 234196 115434
rect 233876 108434 234196 115198
rect 233876 108198 233918 108434
rect 234154 108198 234196 108434
rect 233876 101434 234196 108198
rect 233876 101198 233918 101434
rect 234154 101198 234196 101434
rect 233876 94434 234196 101198
rect 233876 94198 233918 94434
rect 234154 94198 234196 94434
rect 233876 87434 234196 94198
rect 233876 87198 233918 87434
rect 234154 87198 234196 87434
rect 233876 80434 234196 87198
rect 233876 80198 233918 80434
rect 234154 80198 234196 80434
rect 233876 73434 234196 80198
rect 233876 73198 233918 73434
rect 234154 73198 234196 73434
rect 233876 66434 234196 73198
rect 233876 66198 233918 66434
rect 234154 66198 234196 66434
rect 233876 59434 234196 66198
rect 233876 59198 233918 59434
rect 234154 59198 234196 59434
rect 233876 52434 234196 59198
rect 233876 52198 233918 52434
rect 234154 52198 234196 52434
rect 233876 45434 234196 52198
rect 233876 45198 233918 45434
rect 234154 45198 234196 45434
rect 233876 38434 234196 45198
rect 233876 38198 233918 38434
rect 234154 38198 234196 38434
rect 233876 31434 234196 38198
rect 233876 31198 233918 31434
rect 234154 31198 234196 31434
rect 233876 24434 234196 31198
rect 233876 24198 233918 24434
rect 234154 24198 234196 24434
rect 233876 17434 234196 24198
rect 233876 17198 233918 17434
rect 234154 17198 234196 17434
rect 233876 10434 234196 17198
rect 233876 10198 233918 10434
rect 234154 10198 234196 10434
rect 233876 3434 234196 10198
rect 233876 3198 233918 3434
rect 234154 3198 234196 3434
rect 233876 -1706 234196 3198
rect 233876 -1942 233918 -1706
rect 234154 -1942 234196 -1706
rect 233876 -2026 234196 -1942
rect 233876 -2262 233918 -2026
rect 234154 -2262 234196 -2026
rect 233876 -2294 234196 -2262
rect 239144 705238 239464 706230
rect 239144 705002 239186 705238
rect 239422 705002 239464 705238
rect 239144 704918 239464 705002
rect 239144 704682 239186 704918
rect 239422 704682 239464 704918
rect 239144 695494 239464 704682
rect 239144 695258 239186 695494
rect 239422 695258 239464 695494
rect 239144 688494 239464 695258
rect 239144 688258 239186 688494
rect 239422 688258 239464 688494
rect 239144 681494 239464 688258
rect 239144 681258 239186 681494
rect 239422 681258 239464 681494
rect 239144 674494 239464 681258
rect 239144 674258 239186 674494
rect 239422 674258 239464 674494
rect 239144 667494 239464 674258
rect 239144 667258 239186 667494
rect 239422 667258 239464 667494
rect 239144 660494 239464 667258
rect 239144 660258 239186 660494
rect 239422 660258 239464 660494
rect 239144 653494 239464 660258
rect 239144 653258 239186 653494
rect 239422 653258 239464 653494
rect 239144 646494 239464 653258
rect 239144 646258 239186 646494
rect 239422 646258 239464 646494
rect 239144 639494 239464 646258
rect 239144 639258 239186 639494
rect 239422 639258 239464 639494
rect 239144 632494 239464 639258
rect 239144 632258 239186 632494
rect 239422 632258 239464 632494
rect 239144 625494 239464 632258
rect 239144 625258 239186 625494
rect 239422 625258 239464 625494
rect 239144 618494 239464 625258
rect 239144 618258 239186 618494
rect 239422 618258 239464 618494
rect 239144 611494 239464 618258
rect 239144 611258 239186 611494
rect 239422 611258 239464 611494
rect 239144 604494 239464 611258
rect 239144 604258 239186 604494
rect 239422 604258 239464 604494
rect 239144 597494 239464 604258
rect 239144 597258 239186 597494
rect 239422 597258 239464 597494
rect 239144 590494 239464 597258
rect 239144 590258 239186 590494
rect 239422 590258 239464 590494
rect 239144 583494 239464 590258
rect 239144 583258 239186 583494
rect 239422 583258 239464 583494
rect 239144 576494 239464 583258
rect 239144 576258 239186 576494
rect 239422 576258 239464 576494
rect 239144 569494 239464 576258
rect 239144 569258 239186 569494
rect 239422 569258 239464 569494
rect 239144 562494 239464 569258
rect 239144 562258 239186 562494
rect 239422 562258 239464 562494
rect 239144 555494 239464 562258
rect 239144 555258 239186 555494
rect 239422 555258 239464 555494
rect 239144 548494 239464 555258
rect 239144 548258 239186 548494
rect 239422 548258 239464 548494
rect 239144 541494 239464 548258
rect 239144 541258 239186 541494
rect 239422 541258 239464 541494
rect 239144 534494 239464 541258
rect 239144 534258 239186 534494
rect 239422 534258 239464 534494
rect 239144 527494 239464 534258
rect 239144 527258 239186 527494
rect 239422 527258 239464 527494
rect 239144 520494 239464 527258
rect 239144 520258 239186 520494
rect 239422 520258 239464 520494
rect 239144 513494 239464 520258
rect 239144 513258 239186 513494
rect 239422 513258 239464 513494
rect 239144 506494 239464 513258
rect 239144 506258 239186 506494
rect 239422 506258 239464 506494
rect 239144 499494 239464 506258
rect 239144 499258 239186 499494
rect 239422 499258 239464 499494
rect 239144 492494 239464 499258
rect 239144 492258 239186 492494
rect 239422 492258 239464 492494
rect 239144 485494 239464 492258
rect 239144 485258 239186 485494
rect 239422 485258 239464 485494
rect 239144 478494 239464 485258
rect 239144 478258 239186 478494
rect 239422 478258 239464 478494
rect 239144 471494 239464 478258
rect 239144 471258 239186 471494
rect 239422 471258 239464 471494
rect 239144 464494 239464 471258
rect 239144 464258 239186 464494
rect 239422 464258 239464 464494
rect 239144 457494 239464 464258
rect 239144 457258 239186 457494
rect 239422 457258 239464 457494
rect 239144 450494 239464 457258
rect 239144 450258 239186 450494
rect 239422 450258 239464 450494
rect 239144 443494 239464 450258
rect 239144 443258 239186 443494
rect 239422 443258 239464 443494
rect 239144 436494 239464 443258
rect 239144 436258 239186 436494
rect 239422 436258 239464 436494
rect 239144 429494 239464 436258
rect 239144 429258 239186 429494
rect 239422 429258 239464 429494
rect 239144 422494 239464 429258
rect 239144 422258 239186 422494
rect 239422 422258 239464 422494
rect 239144 415494 239464 422258
rect 239144 415258 239186 415494
rect 239422 415258 239464 415494
rect 239144 408494 239464 415258
rect 239144 408258 239186 408494
rect 239422 408258 239464 408494
rect 239144 401494 239464 408258
rect 239144 401258 239186 401494
rect 239422 401258 239464 401494
rect 239144 394494 239464 401258
rect 239144 394258 239186 394494
rect 239422 394258 239464 394494
rect 239144 387494 239464 394258
rect 239144 387258 239186 387494
rect 239422 387258 239464 387494
rect 239144 380494 239464 387258
rect 239144 380258 239186 380494
rect 239422 380258 239464 380494
rect 239144 373494 239464 380258
rect 239144 373258 239186 373494
rect 239422 373258 239464 373494
rect 239144 366494 239464 373258
rect 239144 366258 239186 366494
rect 239422 366258 239464 366494
rect 239144 359494 239464 366258
rect 239144 359258 239186 359494
rect 239422 359258 239464 359494
rect 239144 352494 239464 359258
rect 239144 352258 239186 352494
rect 239422 352258 239464 352494
rect 239144 345494 239464 352258
rect 239144 345258 239186 345494
rect 239422 345258 239464 345494
rect 239144 338494 239464 345258
rect 239144 338258 239186 338494
rect 239422 338258 239464 338494
rect 239144 331494 239464 338258
rect 239144 331258 239186 331494
rect 239422 331258 239464 331494
rect 239144 324494 239464 331258
rect 239144 324258 239186 324494
rect 239422 324258 239464 324494
rect 239144 317494 239464 324258
rect 239144 317258 239186 317494
rect 239422 317258 239464 317494
rect 239144 310494 239464 317258
rect 239144 310258 239186 310494
rect 239422 310258 239464 310494
rect 239144 303494 239464 310258
rect 239144 303258 239186 303494
rect 239422 303258 239464 303494
rect 239144 296494 239464 303258
rect 239144 296258 239186 296494
rect 239422 296258 239464 296494
rect 239144 289494 239464 296258
rect 239144 289258 239186 289494
rect 239422 289258 239464 289494
rect 239144 282494 239464 289258
rect 239144 282258 239186 282494
rect 239422 282258 239464 282494
rect 239144 275494 239464 282258
rect 239144 275258 239186 275494
rect 239422 275258 239464 275494
rect 239144 268494 239464 275258
rect 239144 268258 239186 268494
rect 239422 268258 239464 268494
rect 239144 261494 239464 268258
rect 239144 261258 239186 261494
rect 239422 261258 239464 261494
rect 239144 254494 239464 261258
rect 239144 254258 239186 254494
rect 239422 254258 239464 254494
rect 239144 247494 239464 254258
rect 239144 247258 239186 247494
rect 239422 247258 239464 247494
rect 239144 240494 239464 247258
rect 239144 240258 239186 240494
rect 239422 240258 239464 240494
rect 239144 233494 239464 240258
rect 239144 233258 239186 233494
rect 239422 233258 239464 233494
rect 239144 226494 239464 233258
rect 239144 226258 239186 226494
rect 239422 226258 239464 226494
rect 239144 219494 239464 226258
rect 239144 219258 239186 219494
rect 239422 219258 239464 219494
rect 239144 212494 239464 219258
rect 239144 212258 239186 212494
rect 239422 212258 239464 212494
rect 239144 205494 239464 212258
rect 239144 205258 239186 205494
rect 239422 205258 239464 205494
rect 239144 198494 239464 205258
rect 239144 198258 239186 198494
rect 239422 198258 239464 198494
rect 239144 191494 239464 198258
rect 239144 191258 239186 191494
rect 239422 191258 239464 191494
rect 239144 184494 239464 191258
rect 239144 184258 239186 184494
rect 239422 184258 239464 184494
rect 239144 177494 239464 184258
rect 239144 177258 239186 177494
rect 239422 177258 239464 177494
rect 239144 170494 239464 177258
rect 239144 170258 239186 170494
rect 239422 170258 239464 170494
rect 239144 163494 239464 170258
rect 239144 163258 239186 163494
rect 239422 163258 239464 163494
rect 239144 156494 239464 163258
rect 239144 156258 239186 156494
rect 239422 156258 239464 156494
rect 239144 149494 239464 156258
rect 239144 149258 239186 149494
rect 239422 149258 239464 149494
rect 239144 142494 239464 149258
rect 239144 142258 239186 142494
rect 239422 142258 239464 142494
rect 239144 135494 239464 142258
rect 239144 135258 239186 135494
rect 239422 135258 239464 135494
rect 239144 128494 239464 135258
rect 239144 128258 239186 128494
rect 239422 128258 239464 128494
rect 239144 121494 239464 128258
rect 239144 121258 239186 121494
rect 239422 121258 239464 121494
rect 239144 114494 239464 121258
rect 239144 114258 239186 114494
rect 239422 114258 239464 114494
rect 239144 107494 239464 114258
rect 239144 107258 239186 107494
rect 239422 107258 239464 107494
rect 239144 100494 239464 107258
rect 239144 100258 239186 100494
rect 239422 100258 239464 100494
rect 239144 93494 239464 100258
rect 239144 93258 239186 93494
rect 239422 93258 239464 93494
rect 239144 86494 239464 93258
rect 239144 86258 239186 86494
rect 239422 86258 239464 86494
rect 239144 79494 239464 86258
rect 239144 79258 239186 79494
rect 239422 79258 239464 79494
rect 239144 72494 239464 79258
rect 239144 72258 239186 72494
rect 239422 72258 239464 72494
rect 239144 65494 239464 72258
rect 239144 65258 239186 65494
rect 239422 65258 239464 65494
rect 239144 58494 239464 65258
rect 239144 58258 239186 58494
rect 239422 58258 239464 58494
rect 239144 51494 239464 58258
rect 239144 51258 239186 51494
rect 239422 51258 239464 51494
rect 239144 44494 239464 51258
rect 239144 44258 239186 44494
rect 239422 44258 239464 44494
rect 239144 37494 239464 44258
rect 239144 37258 239186 37494
rect 239422 37258 239464 37494
rect 239144 30494 239464 37258
rect 239144 30258 239186 30494
rect 239422 30258 239464 30494
rect 239144 23494 239464 30258
rect 239144 23258 239186 23494
rect 239422 23258 239464 23494
rect 239144 16494 239464 23258
rect 239144 16258 239186 16494
rect 239422 16258 239464 16494
rect 239144 9494 239464 16258
rect 239144 9258 239186 9494
rect 239422 9258 239464 9494
rect 239144 2494 239464 9258
rect 239144 2258 239186 2494
rect 239422 2258 239464 2494
rect 239144 -746 239464 2258
rect 239144 -982 239186 -746
rect 239422 -982 239464 -746
rect 239144 -1066 239464 -982
rect 239144 -1302 239186 -1066
rect 239422 -1302 239464 -1066
rect 239144 -2294 239464 -1302
rect 240876 706198 241196 706230
rect 240876 705962 240918 706198
rect 241154 705962 241196 706198
rect 240876 705878 241196 705962
rect 240876 705642 240918 705878
rect 241154 705642 241196 705878
rect 240876 696434 241196 705642
rect 240876 696198 240918 696434
rect 241154 696198 241196 696434
rect 240876 689434 241196 696198
rect 240876 689198 240918 689434
rect 241154 689198 241196 689434
rect 240876 682434 241196 689198
rect 240876 682198 240918 682434
rect 241154 682198 241196 682434
rect 240876 675434 241196 682198
rect 240876 675198 240918 675434
rect 241154 675198 241196 675434
rect 240876 668434 241196 675198
rect 240876 668198 240918 668434
rect 241154 668198 241196 668434
rect 240876 661434 241196 668198
rect 240876 661198 240918 661434
rect 241154 661198 241196 661434
rect 240876 654434 241196 661198
rect 240876 654198 240918 654434
rect 241154 654198 241196 654434
rect 240876 647434 241196 654198
rect 240876 647198 240918 647434
rect 241154 647198 241196 647434
rect 240876 640434 241196 647198
rect 240876 640198 240918 640434
rect 241154 640198 241196 640434
rect 240876 633434 241196 640198
rect 240876 633198 240918 633434
rect 241154 633198 241196 633434
rect 240876 626434 241196 633198
rect 240876 626198 240918 626434
rect 241154 626198 241196 626434
rect 240876 619434 241196 626198
rect 240876 619198 240918 619434
rect 241154 619198 241196 619434
rect 240876 612434 241196 619198
rect 240876 612198 240918 612434
rect 241154 612198 241196 612434
rect 240876 605434 241196 612198
rect 240876 605198 240918 605434
rect 241154 605198 241196 605434
rect 240876 598434 241196 605198
rect 240876 598198 240918 598434
rect 241154 598198 241196 598434
rect 240876 591434 241196 598198
rect 240876 591198 240918 591434
rect 241154 591198 241196 591434
rect 240876 584434 241196 591198
rect 240876 584198 240918 584434
rect 241154 584198 241196 584434
rect 240876 577434 241196 584198
rect 240876 577198 240918 577434
rect 241154 577198 241196 577434
rect 240876 570434 241196 577198
rect 240876 570198 240918 570434
rect 241154 570198 241196 570434
rect 240876 563434 241196 570198
rect 240876 563198 240918 563434
rect 241154 563198 241196 563434
rect 240876 556434 241196 563198
rect 240876 556198 240918 556434
rect 241154 556198 241196 556434
rect 240876 549434 241196 556198
rect 240876 549198 240918 549434
rect 241154 549198 241196 549434
rect 240876 542434 241196 549198
rect 240876 542198 240918 542434
rect 241154 542198 241196 542434
rect 240876 535434 241196 542198
rect 240876 535198 240918 535434
rect 241154 535198 241196 535434
rect 240876 528434 241196 535198
rect 240876 528198 240918 528434
rect 241154 528198 241196 528434
rect 240876 521434 241196 528198
rect 240876 521198 240918 521434
rect 241154 521198 241196 521434
rect 240876 514434 241196 521198
rect 240876 514198 240918 514434
rect 241154 514198 241196 514434
rect 240876 507434 241196 514198
rect 240876 507198 240918 507434
rect 241154 507198 241196 507434
rect 240876 500434 241196 507198
rect 240876 500198 240918 500434
rect 241154 500198 241196 500434
rect 240876 493434 241196 500198
rect 240876 493198 240918 493434
rect 241154 493198 241196 493434
rect 240876 486434 241196 493198
rect 240876 486198 240918 486434
rect 241154 486198 241196 486434
rect 240876 479434 241196 486198
rect 240876 479198 240918 479434
rect 241154 479198 241196 479434
rect 240876 472434 241196 479198
rect 240876 472198 240918 472434
rect 241154 472198 241196 472434
rect 240876 465434 241196 472198
rect 240876 465198 240918 465434
rect 241154 465198 241196 465434
rect 240876 458434 241196 465198
rect 240876 458198 240918 458434
rect 241154 458198 241196 458434
rect 240876 451434 241196 458198
rect 240876 451198 240918 451434
rect 241154 451198 241196 451434
rect 240876 444434 241196 451198
rect 240876 444198 240918 444434
rect 241154 444198 241196 444434
rect 240876 437434 241196 444198
rect 240876 437198 240918 437434
rect 241154 437198 241196 437434
rect 240876 430434 241196 437198
rect 240876 430198 240918 430434
rect 241154 430198 241196 430434
rect 240876 423434 241196 430198
rect 240876 423198 240918 423434
rect 241154 423198 241196 423434
rect 240876 416434 241196 423198
rect 240876 416198 240918 416434
rect 241154 416198 241196 416434
rect 240876 409434 241196 416198
rect 240876 409198 240918 409434
rect 241154 409198 241196 409434
rect 240876 402434 241196 409198
rect 240876 402198 240918 402434
rect 241154 402198 241196 402434
rect 240876 395434 241196 402198
rect 240876 395198 240918 395434
rect 241154 395198 241196 395434
rect 240876 388434 241196 395198
rect 240876 388198 240918 388434
rect 241154 388198 241196 388434
rect 240876 381434 241196 388198
rect 240876 381198 240918 381434
rect 241154 381198 241196 381434
rect 240876 374434 241196 381198
rect 240876 374198 240918 374434
rect 241154 374198 241196 374434
rect 240876 367434 241196 374198
rect 240876 367198 240918 367434
rect 241154 367198 241196 367434
rect 240876 360434 241196 367198
rect 240876 360198 240918 360434
rect 241154 360198 241196 360434
rect 240876 353434 241196 360198
rect 240876 353198 240918 353434
rect 241154 353198 241196 353434
rect 240876 346434 241196 353198
rect 240876 346198 240918 346434
rect 241154 346198 241196 346434
rect 240876 339434 241196 346198
rect 240876 339198 240918 339434
rect 241154 339198 241196 339434
rect 240876 332434 241196 339198
rect 240876 332198 240918 332434
rect 241154 332198 241196 332434
rect 240876 325434 241196 332198
rect 240876 325198 240918 325434
rect 241154 325198 241196 325434
rect 240876 318434 241196 325198
rect 240876 318198 240918 318434
rect 241154 318198 241196 318434
rect 240876 311434 241196 318198
rect 240876 311198 240918 311434
rect 241154 311198 241196 311434
rect 240876 304434 241196 311198
rect 240876 304198 240918 304434
rect 241154 304198 241196 304434
rect 240876 297434 241196 304198
rect 240876 297198 240918 297434
rect 241154 297198 241196 297434
rect 240876 290434 241196 297198
rect 240876 290198 240918 290434
rect 241154 290198 241196 290434
rect 240876 283434 241196 290198
rect 240876 283198 240918 283434
rect 241154 283198 241196 283434
rect 240876 276434 241196 283198
rect 240876 276198 240918 276434
rect 241154 276198 241196 276434
rect 240876 269434 241196 276198
rect 240876 269198 240918 269434
rect 241154 269198 241196 269434
rect 240876 262434 241196 269198
rect 240876 262198 240918 262434
rect 241154 262198 241196 262434
rect 240876 255434 241196 262198
rect 240876 255198 240918 255434
rect 241154 255198 241196 255434
rect 240876 248434 241196 255198
rect 240876 248198 240918 248434
rect 241154 248198 241196 248434
rect 240876 241434 241196 248198
rect 240876 241198 240918 241434
rect 241154 241198 241196 241434
rect 240876 234434 241196 241198
rect 240876 234198 240918 234434
rect 241154 234198 241196 234434
rect 240876 227434 241196 234198
rect 240876 227198 240918 227434
rect 241154 227198 241196 227434
rect 240876 220434 241196 227198
rect 240876 220198 240918 220434
rect 241154 220198 241196 220434
rect 240876 213434 241196 220198
rect 240876 213198 240918 213434
rect 241154 213198 241196 213434
rect 240876 206434 241196 213198
rect 240876 206198 240918 206434
rect 241154 206198 241196 206434
rect 240876 199434 241196 206198
rect 240876 199198 240918 199434
rect 241154 199198 241196 199434
rect 240876 192434 241196 199198
rect 240876 192198 240918 192434
rect 241154 192198 241196 192434
rect 240876 185434 241196 192198
rect 240876 185198 240918 185434
rect 241154 185198 241196 185434
rect 240876 178434 241196 185198
rect 240876 178198 240918 178434
rect 241154 178198 241196 178434
rect 240876 171434 241196 178198
rect 240876 171198 240918 171434
rect 241154 171198 241196 171434
rect 240876 164434 241196 171198
rect 240876 164198 240918 164434
rect 241154 164198 241196 164434
rect 240876 157434 241196 164198
rect 240876 157198 240918 157434
rect 241154 157198 241196 157434
rect 240876 150434 241196 157198
rect 240876 150198 240918 150434
rect 241154 150198 241196 150434
rect 240876 143434 241196 150198
rect 240876 143198 240918 143434
rect 241154 143198 241196 143434
rect 240876 136434 241196 143198
rect 240876 136198 240918 136434
rect 241154 136198 241196 136434
rect 240876 129434 241196 136198
rect 240876 129198 240918 129434
rect 241154 129198 241196 129434
rect 240876 122434 241196 129198
rect 240876 122198 240918 122434
rect 241154 122198 241196 122434
rect 240876 115434 241196 122198
rect 240876 115198 240918 115434
rect 241154 115198 241196 115434
rect 240876 108434 241196 115198
rect 240876 108198 240918 108434
rect 241154 108198 241196 108434
rect 240876 101434 241196 108198
rect 240876 101198 240918 101434
rect 241154 101198 241196 101434
rect 240876 94434 241196 101198
rect 240876 94198 240918 94434
rect 241154 94198 241196 94434
rect 240876 87434 241196 94198
rect 240876 87198 240918 87434
rect 241154 87198 241196 87434
rect 240876 80434 241196 87198
rect 240876 80198 240918 80434
rect 241154 80198 241196 80434
rect 240876 73434 241196 80198
rect 240876 73198 240918 73434
rect 241154 73198 241196 73434
rect 240876 66434 241196 73198
rect 240876 66198 240918 66434
rect 241154 66198 241196 66434
rect 240876 59434 241196 66198
rect 240876 59198 240918 59434
rect 241154 59198 241196 59434
rect 240876 52434 241196 59198
rect 240876 52198 240918 52434
rect 241154 52198 241196 52434
rect 240876 45434 241196 52198
rect 240876 45198 240918 45434
rect 241154 45198 241196 45434
rect 240876 38434 241196 45198
rect 240876 38198 240918 38434
rect 241154 38198 241196 38434
rect 240876 31434 241196 38198
rect 240876 31198 240918 31434
rect 241154 31198 241196 31434
rect 240876 24434 241196 31198
rect 240876 24198 240918 24434
rect 241154 24198 241196 24434
rect 240876 17434 241196 24198
rect 240876 17198 240918 17434
rect 241154 17198 241196 17434
rect 240876 10434 241196 17198
rect 240876 10198 240918 10434
rect 241154 10198 241196 10434
rect 240876 3434 241196 10198
rect 240876 3198 240918 3434
rect 241154 3198 241196 3434
rect 240876 -1706 241196 3198
rect 240876 -1942 240918 -1706
rect 241154 -1942 241196 -1706
rect 240876 -2026 241196 -1942
rect 240876 -2262 240918 -2026
rect 241154 -2262 241196 -2026
rect 240876 -2294 241196 -2262
rect 246144 705238 246464 706230
rect 246144 705002 246186 705238
rect 246422 705002 246464 705238
rect 246144 704918 246464 705002
rect 246144 704682 246186 704918
rect 246422 704682 246464 704918
rect 246144 695494 246464 704682
rect 246144 695258 246186 695494
rect 246422 695258 246464 695494
rect 246144 688494 246464 695258
rect 246144 688258 246186 688494
rect 246422 688258 246464 688494
rect 246144 681494 246464 688258
rect 246144 681258 246186 681494
rect 246422 681258 246464 681494
rect 246144 674494 246464 681258
rect 246144 674258 246186 674494
rect 246422 674258 246464 674494
rect 246144 667494 246464 674258
rect 246144 667258 246186 667494
rect 246422 667258 246464 667494
rect 246144 660494 246464 667258
rect 246144 660258 246186 660494
rect 246422 660258 246464 660494
rect 246144 653494 246464 660258
rect 246144 653258 246186 653494
rect 246422 653258 246464 653494
rect 246144 646494 246464 653258
rect 246144 646258 246186 646494
rect 246422 646258 246464 646494
rect 246144 639494 246464 646258
rect 246144 639258 246186 639494
rect 246422 639258 246464 639494
rect 246144 632494 246464 639258
rect 246144 632258 246186 632494
rect 246422 632258 246464 632494
rect 246144 625494 246464 632258
rect 246144 625258 246186 625494
rect 246422 625258 246464 625494
rect 246144 618494 246464 625258
rect 246144 618258 246186 618494
rect 246422 618258 246464 618494
rect 246144 611494 246464 618258
rect 246144 611258 246186 611494
rect 246422 611258 246464 611494
rect 246144 604494 246464 611258
rect 246144 604258 246186 604494
rect 246422 604258 246464 604494
rect 246144 597494 246464 604258
rect 246144 597258 246186 597494
rect 246422 597258 246464 597494
rect 246144 590494 246464 597258
rect 246144 590258 246186 590494
rect 246422 590258 246464 590494
rect 246144 583494 246464 590258
rect 246144 583258 246186 583494
rect 246422 583258 246464 583494
rect 246144 576494 246464 583258
rect 246144 576258 246186 576494
rect 246422 576258 246464 576494
rect 246144 569494 246464 576258
rect 246144 569258 246186 569494
rect 246422 569258 246464 569494
rect 246144 562494 246464 569258
rect 246144 562258 246186 562494
rect 246422 562258 246464 562494
rect 246144 555494 246464 562258
rect 246144 555258 246186 555494
rect 246422 555258 246464 555494
rect 246144 548494 246464 555258
rect 246144 548258 246186 548494
rect 246422 548258 246464 548494
rect 246144 541494 246464 548258
rect 246144 541258 246186 541494
rect 246422 541258 246464 541494
rect 246144 534494 246464 541258
rect 246144 534258 246186 534494
rect 246422 534258 246464 534494
rect 246144 527494 246464 534258
rect 246144 527258 246186 527494
rect 246422 527258 246464 527494
rect 246144 520494 246464 527258
rect 246144 520258 246186 520494
rect 246422 520258 246464 520494
rect 246144 513494 246464 520258
rect 246144 513258 246186 513494
rect 246422 513258 246464 513494
rect 246144 506494 246464 513258
rect 246144 506258 246186 506494
rect 246422 506258 246464 506494
rect 246144 499494 246464 506258
rect 246144 499258 246186 499494
rect 246422 499258 246464 499494
rect 246144 492494 246464 499258
rect 246144 492258 246186 492494
rect 246422 492258 246464 492494
rect 246144 485494 246464 492258
rect 246144 485258 246186 485494
rect 246422 485258 246464 485494
rect 246144 478494 246464 485258
rect 246144 478258 246186 478494
rect 246422 478258 246464 478494
rect 246144 471494 246464 478258
rect 246144 471258 246186 471494
rect 246422 471258 246464 471494
rect 246144 464494 246464 471258
rect 246144 464258 246186 464494
rect 246422 464258 246464 464494
rect 246144 457494 246464 464258
rect 246144 457258 246186 457494
rect 246422 457258 246464 457494
rect 246144 450494 246464 457258
rect 246144 450258 246186 450494
rect 246422 450258 246464 450494
rect 246144 443494 246464 450258
rect 246144 443258 246186 443494
rect 246422 443258 246464 443494
rect 246144 436494 246464 443258
rect 246144 436258 246186 436494
rect 246422 436258 246464 436494
rect 246144 429494 246464 436258
rect 246144 429258 246186 429494
rect 246422 429258 246464 429494
rect 246144 422494 246464 429258
rect 246144 422258 246186 422494
rect 246422 422258 246464 422494
rect 246144 415494 246464 422258
rect 246144 415258 246186 415494
rect 246422 415258 246464 415494
rect 246144 408494 246464 415258
rect 246144 408258 246186 408494
rect 246422 408258 246464 408494
rect 246144 401494 246464 408258
rect 246144 401258 246186 401494
rect 246422 401258 246464 401494
rect 246144 394494 246464 401258
rect 246144 394258 246186 394494
rect 246422 394258 246464 394494
rect 246144 387494 246464 394258
rect 246144 387258 246186 387494
rect 246422 387258 246464 387494
rect 246144 380494 246464 387258
rect 246144 380258 246186 380494
rect 246422 380258 246464 380494
rect 246144 373494 246464 380258
rect 246144 373258 246186 373494
rect 246422 373258 246464 373494
rect 246144 366494 246464 373258
rect 246144 366258 246186 366494
rect 246422 366258 246464 366494
rect 246144 359494 246464 366258
rect 246144 359258 246186 359494
rect 246422 359258 246464 359494
rect 246144 352494 246464 359258
rect 246144 352258 246186 352494
rect 246422 352258 246464 352494
rect 246144 345494 246464 352258
rect 246144 345258 246186 345494
rect 246422 345258 246464 345494
rect 246144 338494 246464 345258
rect 246144 338258 246186 338494
rect 246422 338258 246464 338494
rect 246144 331494 246464 338258
rect 246144 331258 246186 331494
rect 246422 331258 246464 331494
rect 246144 324494 246464 331258
rect 246144 324258 246186 324494
rect 246422 324258 246464 324494
rect 246144 317494 246464 324258
rect 246144 317258 246186 317494
rect 246422 317258 246464 317494
rect 246144 310494 246464 317258
rect 246144 310258 246186 310494
rect 246422 310258 246464 310494
rect 246144 303494 246464 310258
rect 246144 303258 246186 303494
rect 246422 303258 246464 303494
rect 246144 296494 246464 303258
rect 246144 296258 246186 296494
rect 246422 296258 246464 296494
rect 246144 289494 246464 296258
rect 246144 289258 246186 289494
rect 246422 289258 246464 289494
rect 246144 282494 246464 289258
rect 246144 282258 246186 282494
rect 246422 282258 246464 282494
rect 246144 275494 246464 282258
rect 246144 275258 246186 275494
rect 246422 275258 246464 275494
rect 246144 268494 246464 275258
rect 246144 268258 246186 268494
rect 246422 268258 246464 268494
rect 246144 261494 246464 268258
rect 246144 261258 246186 261494
rect 246422 261258 246464 261494
rect 246144 254494 246464 261258
rect 246144 254258 246186 254494
rect 246422 254258 246464 254494
rect 246144 247494 246464 254258
rect 246144 247258 246186 247494
rect 246422 247258 246464 247494
rect 246144 240494 246464 247258
rect 246144 240258 246186 240494
rect 246422 240258 246464 240494
rect 246144 233494 246464 240258
rect 246144 233258 246186 233494
rect 246422 233258 246464 233494
rect 246144 226494 246464 233258
rect 246144 226258 246186 226494
rect 246422 226258 246464 226494
rect 246144 219494 246464 226258
rect 246144 219258 246186 219494
rect 246422 219258 246464 219494
rect 246144 212494 246464 219258
rect 246144 212258 246186 212494
rect 246422 212258 246464 212494
rect 246144 205494 246464 212258
rect 246144 205258 246186 205494
rect 246422 205258 246464 205494
rect 246144 198494 246464 205258
rect 246144 198258 246186 198494
rect 246422 198258 246464 198494
rect 246144 191494 246464 198258
rect 246144 191258 246186 191494
rect 246422 191258 246464 191494
rect 246144 184494 246464 191258
rect 246144 184258 246186 184494
rect 246422 184258 246464 184494
rect 246144 177494 246464 184258
rect 246144 177258 246186 177494
rect 246422 177258 246464 177494
rect 246144 170494 246464 177258
rect 246144 170258 246186 170494
rect 246422 170258 246464 170494
rect 246144 163494 246464 170258
rect 246144 163258 246186 163494
rect 246422 163258 246464 163494
rect 246144 156494 246464 163258
rect 246144 156258 246186 156494
rect 246422 156258 246464 156494
rect 246144 149494 246464 156258
rect 246144 149258 246186 149494
rect 246422 149258 246464 149494
rect 246144 142494 246464 149258
rect 246144 142258 246186 142494
rect 246422 142258 246464 142494
rect 246144 135494 246464 142258
rect 246144 135258 246186 135494
rect 246422 135258 246464 135494
rect 246144 128494 246464 135258
rect 246144 128258 246186 128494
rect 246422 128258 246464 128494
rect 246144 121494 246464 128258
rect 246144 121258 246186 121494
rect 246422 121258 246464 121494
rect 246144 114494 246464 121258
rect 246144 114258 246186 114494
rect 246422 114258 246464 114494
rect 246144 107494 246464 114258
rect 246144 107258 246186 107494
rect 246422 107258 246464 107494
rect 246144 100494 246464 107258
rect 246144 100258 246186 100494
rect 246422 100258 246464 100494
rect 246144 93494 246464 100258
rect 246144 93258 246186 93494
rect 246422 93258 246464 93494
rect 246144 86494 246464 93258
rect 246144 86258 246186 86494
rect 246422 86258 246464 86494
rect 246144 79494 246464 86258
rect 246144 79258 246186 79494
rect 246422 79258 246464 79494
rect 246144 72494 246464 79258
rect 246144 72258 246186 72494
rect 246422 72258 246464 72494
rect 246144 65494 246464 72258
rect 246144 65258 246186 65494
rect 246422 65258 246464 65494
rect 246144 58494 246464 65258
rect 246144 58258 246186 58494
rect 246422 58258 246464 58494
rect 246144 51494 246464 58258
rect 246144 51258 246186 51494
rect 246422 51258 246464 51494
rect 246144 44494 246464 51258
rect 246144 44258 246186 44494
rect 246422 44258 246464 44494
rect 246144 37494 246464 44258
rect 246144 37258 246186 37494
rect 246422 37258 246464 37494
rect 246144 30494 246464 37258
rect 246144 30258 246186 30494
rect 246422 30258 246464 30494
rect 246144 23494 246464 30258
rect 246144 23258 246186 23494
rect 246422 23258 246464 23494
rect 246144 16494 246464 23258
rect 246144 16258 246186 16494
rect 246422 16258 246464 16494
rect 246144 9494 246464 16258
rect 246144 9258 246186 9494
rect 246422 9258 246464 9494
rect 246144 2494 246464 9258
rect 246144 2258 246186 2494
rect 246422 2258 246464 2494
rect 246144 -746 246464 2258
rect 246144 -982 246186 -746
rect 246422 -982 246464 -746
rect 246144 -1066 246464 -982
rect 246144 -1302 246186 -1066
rect 246422 -1302 246464 -1066
rect 246144 -2294 246464 -1302
rect 247876 706198 248196 706230
rect 247876 705962 247918 706198
rect 248154 705962 248196 706198
rect 247876 705878 248196 705962
rect 247876 705642 247918 705878
rect 248154 705642 248196 705878
rect 247876 696434 248196 705642
rect 247876 696198 247918 696434
rect 248154 696198 248196 696434
rect 247876 689434 248196 696198
rect 247876 689198 247918 689434
rect 248154 689198 248196 689434
rect 247876 682434 248196 689198
rect 247876 682198 247918 682434
rect 248154 682198 248196 682434
rect 247876 675434 248196 682198
rect 247876 675198 247918 675434
rect 248154 675198 248196 675434
rect 247876 668434 248196 675198
rect 247876 668198 247918 668434
rect 248154 668198 248196 668434
rect 247876 661434 248196 668198
rect 247876 661198 247918 661434
rect 248154 661198 248196 661434
rect 247876 654434 248196 661198
rect 247876 654198 247918 654434
rect 248154 654198 248196 654434
rect 247876 647434 248196 654198
rect 247876 647198 247918 647434
rect 248154 647198 248196 647434
rect 247876 640434 248196 647198
rect 247876 640198 247918 640434
rect 248154 640198 248196 640434
rect 247876 633434 248196 640198
rect 247876 633198 247918 633434
rect 248154 633198 248196 633434
rect 247876 626434 248196 633198
rect 247876 626198 247918 626434
rect 248154 626198 248196 626434
rect 247876 619434 248196 626198
rect 247876 619198 247918 619434
rect 248154 619198 248196 619434
rect 247876 612434 248196 619198
rect 247876 612198 247918 612434
rect 248154 612198 248196 612434
rect 247876 605434 248196 612198
rect 247876 605198 247918 605434
rect 248154 605198 248196 605434
rect 247876 598434 248196 605198
rect 247876 598198 247918 598434
rect 248154 598198 248196 598434
rect 247876 591434 248196 598198
rect 247876 591198 247918 591434
rect 248154 591198 248196 591434
rect 247876 584434 248196 591198
rect 247876 584198 247918 584434
rect 248154 584198 248196 584434
rect 247876 577434 248196 584198
rect 247876 577198 247918 577434
rect 248154 577198 248196 577434
rect 247876 570434 248196 577198
rect 247876 570198 247918 570434
rect 248154 570198 248196 570434
rect 247876 563434 248196 570198
rect 247876 563198 247918 563434
rect 248154 563198 248196 563434
rect 247876 556434 248196 563198
rect 247876 556198 247918 556434
rect 248154 556198 248196 556434
rect 247876 549434 248196 556198
rect 247876 549198 247918 549434
rect 248154 549198 248196 549434
rect 247876 542434 248196 549198
rect 247876 542198 247918 542434
rect 248154 542198 248196 542434
rect 247876 535434 248196 542198
rect 247876 535198 247918 535434
rect 248154 535198 248196 535434
rect 247876 528434 248196 535198
rect 247876 528198 247918 528434
rect 248154 528198 248196 528434
rect 247876 521434 248196 528198
rect 247876 521198 247918 521434
rect 248154 521198 248196 521434
rect 247876 514434 248196 521198
rect 247876 514198 247918 514434
rect 248154 514198 248196 514434
rect 247876 507434 248196 514198
rect 247876 507198 247918 507434
rect 248154 507198 248196 507434
rect 247876 500434 248196 507198
rect 247876 500198 247918 500434
rect 248154 500198 248196 500434
rect 247876 493434 248196 500198
rect 247876 493198 247918 493434
rect 248154 493198 248196 493434
rect 247876 486434 248196 493198
rect 247876 486198 247918 486434
rect 248154 486198 248196 486434
rect 247876 479434 248196 486198
rect 247876 479198 247918 479434
rect 248154 479198 248196 479434
rect 247876 472434 248196 479198
rect 247876 472198 247918 472434
rect 248154 472198 248196 472434
rect 247876 465434 248196 472198
rect 247876 465198 247918 465434
rect 248154 465198 248196 465434
rect 247876 458434 248196 465198
rect 247876 458198 247918 458434
rect 248154 458198 248196 458434
rect 247876 451434 248196 458198
rect 247876 451198 247918 451434
rect 248154 451198 248196 451434
rect 247876 444434 248196 451198
rect 247876 444198 247918 444434
rect 248154 444198 248196 444434
rect 247876 437434 248196 444198
rect 247876 437198 247918 437434
rect 248154 437198 248196 437434
rect 247876 430434 248196 437198
rect 247876 430198 247918 430434
rect 248154 430198 248196 430434
rect 247876 423434 248196 430198
rect 247876 423198 247918 423434
rect 248154 423198 248196 423434
rect 247876 416434 248196 423198
rect 247876 416198 247918 416434
rect 248154 416198 248196 416434
rect 247876 409434 248196 416198
rect 247876 409198 247918 409434
rect 248154 409198 248196 409434
rect 247876 402434 248196 409198
rect 247876 402198 247918 402434
rect 248154 402198 248196 402434
rect 247876 395434 248196 402198
rect 247876 395198 247918 395434
rect 248154 395198 248196 395434
rect 247876 388434 248196 395198
rect 247876 388198 247918 388434
rect 248154 388198 248196 388434
rect 247876 381434 248196 388198
rect 247876 381198 247918 381434
rect 248154 381198 248196 381434
rect 247876 374434 248196 381198
rect 247876 374198 247918 374434
rect 248154 374198 248196 374434
rect 247876 367434 248196 374198
rect 247876 367198 247918 367434
rect 248154 367198 248196 367434
rect 247876 360434 248196 367198
rect 247876 360198 247918 360434
rect 248154 360198 248196 360434
rect 247876 353434 248196 360198
rect 247876 353198 247918 353434
rect 248154 353198 248196 353434
rect 247876 346434 248196 353198
rect 247876 346198 247918 346434
rect 248154 346198 248196 346434
rect 247876 339434 248196 346198
rect 247876 339198 247918 339434
rect 248154 339198 248196 339434
rect 247876 332434 248196 339198
rect 247876 332198 247918 332434
rect 248154 332198 248196 332434
rect 247876 325434 248196 332198
rect 247876 325198 247918 325434
rect 248154 325198 248196 325434
rect 247876 318434 248196 325198
rect 247876 318198 247918 318434
rect 248154 318198 248196 318434
rect 247876 311434 248196 318198
rect 247876 311198 247918 311434
rect 248154 311198 248196 311434
rect 247876 304434 248196 311198
rect 247876 304198 247918 304434
rect 248154 304198 248196 304434
rect 247876 297434 248196 304198
rect 247876 297198 247918 297434
rect 248154 297198 248196 297434
rect 247876 290434 248196 297198
rect 247876 290198 247918 290434
rect 248154 290198 248196 290434
rect 247876 283434 248196 290198
rect 247876 283198 247918 283434
rect 248154 283198 248196 283434
rect 247876 276434 248196 283198
rect 247876 276198 247918 276434
rect 248154 276198 248196 276434
rect 247876 269434 248196 276198
rect 247876 269198 247918 269434
rect 248154 269198 248196 269434
rect 247876 262434 248196 269198
rect 247876 262198 247918 262434
rect 248154 262198 248196 262434
rect 247876 255434 248196 262198
rect 247876 255198 247918 255434
rect 248154 255198 248196 255434
rect 247876 248434 248196 255198
rect 247876 248198 247918 248434
rect 248154 248198 248196 248434
rect 247876 241434 248196 248198
rect 247876 241198 247918 241434
rect 248154 241198 248196 241434
rect 247876 234434 248196 241198
rect 247876 234198 247918 234434
rect 248154 234198 248196 234434
rect 247876 227434 248196 234198
rect 247876 227198 247918 227434
rect 248154 227198 248196 227434
rect 247876 220434 248196 227198
rect 247876 220198 247918 220434
rect 248154 220198 248196 220434
rect 247876 213434 248196 220198
rect 247876 213198 247918 213434
rect 248154 213198 248196 213434
rect 247876 206434 248196 213198
rect 247876 206198 247918 206434
rect 248154 206198 248196 206434
rect 247876 199434 248196 206198
rect 247876 199198 247918 199434
rect 248154 199198 248196 199434
rect 247876 192434 248196 199198
rect 247876 192198 247918 192434
rect 248154 192198 248196 192434
rect 247876 185434 248196 192198
rect 247876 185198 247918 185434
rect 248154 185198 248196 185434
rect 247876 178434 248196 185198
rect 247876 178198 247918 178434
rect 248154 178198 248196 178434
rect 247876 171434 248196 178198
rect 247876 171198 247918 171434
rect 248154 171198 248196 171434
rect 247876 164434 248196 171198
rect 247876 164198 247918 164434
rect 248154 164198 248196 164434
rect 247876 157434 248196 164198
rect 247876 157198 247918 157434
rect 248154 157198 248196 157434
rect 247876 150434 248196 157198
rect 247876 150198 247918 150434
rect 248154 150198 248196 150434
rect 247876 143434 248196 150198
rect 247876 143198 247918 143434
rect 248154 143198 248196 143434
rect 247876 136434 248196 143198
rect 247876 136198 247918 136434
rect 248154 136198 248196 136434
rect 247876 129434 248196 136198
rect 247876 129198 247918 129434
rect 248154 129198 248196 129434
rect 247876 122434 248196 129198
rect 247876 122198 247918 122434
rect 248154 122198 248196 122434
rect 247876 115434 248196 122198
rect 247876 115198 247918 115434
rect 248154 115198 248196 115434
rect 247876 108434 248196 115198
rect 247876 108198 247918 108434
rect 248154 108198 248196 108434
rect 247876 101434 248196 108198
rect 247876 101198 247918 101434
rect 248154 101198 248196 101434
rect 247876 94434 248196 101198
rect 247876 94198 247918 94434
rect 248154 94198 248196 94434
rect 247876 87434 248196 94198
rect 247876 87198 247918 87434
rect 248154 87198 248196 87434
rect 247876 80434 248196 87198
rect 247876 80198 247918 80434
rect 248154 80198 248196 80434
rect 247876 73434 248196 80198
rect 247876 73198 247918 73434
rect 248154 73198 248196 73434
rect 247876 66434 248196 73198
rect 247876 66198 247918 66434
rect 248154 66198 248196 66434
rect 247876 59434 248196 66198
rect 247876 59198 247918 59434
rect 248154 59198 248196 59434
rect 247876 52434 248196 59198
rect 247876 52198 247918 52434
rect 248154 52198 248196 52434
rect 247876 45434 248196 52198
rect 247876 45198 247918 45434
rect 248154 45198 248196 45434
rect 247876 38434 248196 45198
rect 247876 38198 247918 38434
rect 248154 38198 248196 38434
rect 247876 31434 248196 38198
rect 247876 31198 247918 31434
rect 248154 31198 248196 31434
rect 247876 24434 248196 31198
rect 247876 24198 247918 24434
rect 248154 24198 248196 24434
rect 247876 17434 248196 24198
rect 247876 17198 247918 17434
rect 248154 17198 248196 17434
rect 247876 10434 248196 17198
rect 247876 10198 247918 10434
rect 248154 10198 248196 10434
rect 247876 3434 248196 10198
rect 247876 3198 247918 3434
rect 248154 3198 248196 3434
rect 247876 -1706 248196 3198
rect 247876 -1942 247918 -1706
rect 248154 -1942 248196 -1706
rect 247876 -2026 248196 -1942
rect 247876 -2262 247918 -2026
rect 248154 -2262 248196 -2026
rect 247876 -2294 248196 -2262
rect 253144 705238 253464 706230
rect 253144 705002 253186 705238
rect 253422 705002 253464 705238
rect 253144 704918 253464 705002
rect 253144 704682 253186 704918
rect 253422 704682 253464 704918
rect 253144 695494 253464 704682
rect 253144 695258 253186 695494
rect 253422 695258 253464 695494
rect 253144 688494 253464 695258
rect 253144 688258 253186 688494
rect 253422 688258 253464 688494
rect 253144 681494 253464 688258
rect 253144 681258 253186 681494
rect 253422 681258 253464 681494
rect 253144 674494 253464 681258
rect 253144 674258 253186 674494
rect 253422 674258 253464 674494
rect 253144 667494 253464 674258
rect 253144 667258 253186 667494
rect 253422 667258 253464 667494
rect 253144 660494 253464 667258
rect 253144 660258 253186 660494
rect 253422 660258 253464 660494
rect 253144 653494 253464 660258
rect 253144 653258 253186 653494
rect 253422 653258 253464 653494
rect 253144 646494 253464 653258
rect 253144 646258 253186 646494
rect 253422 646258 253464 646494
rect 253144 639494 253464 646258
rect 253144 639258 253186 639494
rect 253422 639258 253464 639494
rect 253144 632494 253464 639258
rect 253144 632258 253186 632494
rect 253422 632258 253464 632494
rect 253144 625494 253464 632258
rect 253144 625258 253186 625494
rect 253422 625258 253464 625494
rect 253144 618494 253464 625258
rect 253144 618258 253186 618494
rect 253422 618258 253464 618494
rect 253144 611494 253464 618258
rect 253144 611258 253186 611494
rect 253422 611258 253464 611494
rect 253144 604494 253464 611258
rect 253144 604258 253186 604494
rect 253422 604258 253464 604494
rect 253144 597494 253464 604258
rect 253144 597258 253186 597494
rect 253422 597258 253464 597494
rect 253144 590494 253464 597258
rect 253144 590258 253186 590494
rect 253422 590258 253464 590494
rect 253144 583494 253464 590258
rect 253144 583258 253186 583494
rect 253422 583258 253464 583494
rect 253144 576494 253464 583258
rect 253144 576258 253186 576494
rect 253422 576258 253464 576494
rect 253144 569494 253464 576258
rect 253144 569258 253186 569494
rect 253422 569258 253464 569494
rect 253144 562494 253464 569258
rect 253144 562258 253186 562494
rect 253422 562258 253464 562494
rect 253144 555494 253464 562258
rect 253144 555258 253186 555494
rect 253422 555258 253464 555494
rect 253144 548494 253464 555258
rect 253144 548258 253186 548494
rect 253422 548258 253464 548494
rect 253144 541494 253464 548258
rect 253144 541258 253186 541494
rect 253422 541258 253464 541494
rect 253144 534494 253464 541258
rect 253144 534258 253186 534494
rect 253422 534258 253464 534494
rect 253144 527494 253464 534258
rect 253144 527258 253186 527494
rect 253422 527258 253464 527494
rect 253144 520494 253464 527258
rect 253144 520258 253186 520494
rect 253422 520258 253464 520494
rect 253144 513494 253464 520258
rect 253144 513258 253186 513494
rect 253422 513258 253464 513494
rect 253144 506494 253464 513258
rect 253144 506258 253186 506494
rect 253422 506258 253464 506494
rect 253144 499494 253464 506258
rect 253144 499258 253186 499494
rect 253422 499258 253464 499494
rect 253144 492494 253464 499258
rect 253144 492258 253186 492494
rect 253422 492258 253464 492494
rect 253144 485494 253464 492258
rect 253144 485258 253186 485494
rect 253422 485258 253464 485494
rect 253144 478494 253464 485258
rect 253144 478258 253186 478494
rect 253422 478258 253464 478494
rect 253144 471494 253464 478258
rect 253144 471258 253186 471494
rect 253422 471258 253464 471494
rect 253144 464494 253464 471258
rect 253144 464258 253186 464494
rect 253422 464258 253464 464494
rect 253144 457494 253464 464258
rect 253144 457258 253186 457494
rect 253422 457258 253464 457494
rect 253144 450494 253464 457258
rect 253144 450258 253186 450494
rect 253422 450258 253464 450494
rect 253144 443494 253464 450258
rect 253144 443258 253186 443494
rect 253422 443258 253464 443494
rect 253144 436494 253464 443258
rect 253144 436258 253186 436494
rect 253422 436258 253464 436494
rect 253144 429494 253464 436258
rect 253144 429258 253186 429494
rect 253422 429258 253464 429494
rect 253144 422494 253464 429258
rect 253144 422258 253186 422494
rect 253422 422258 253464 422494
rect 253144 415494 253464 422258
rect 253144 415258 253186 415494
rect 253422 415258 253464 415494
rect 253144 408494 253464 415258
rect 253144 408258 253186 408494
rect 253422 408258 253464 408494
rect 253144 401494 253464 408258
rect 253144 401258 253186 401494
rect 253422 401258 253464 401494
rect 253144 394494 253464 401258
rect 253144 394258 253186 394494
rect 253422 394258 253464 394494
rect 253144 387494 253464 394258
rect 253144 387258 253186 387494
rect 253422 387258 253464 387494
rect 253144 380494 253464 387258
rect 253144 380258 253186 380494
rect 253422 380258 253464 380494
rect 253144 373494 253464 380258
rect 253144 373258 253186 373494
rect 253422 373258 253464 373494
rect 253144 366494 253464 373258
rect 253144 366258 253186 366494
rect 253422 366258 253464 366494
rect 253144 359494 253464 366258
rect 253144 359258 253186 359494
rect 253422 359258 253464 359494
rect 253144 352494 253464 359258
rect 253144 352258 253186 352494
rect 253422 352258 253464 352494
rect 253144 345494 253464 352258
rect 253144 345258 253186 345494
rect 253422 345258 253464 345494
rect 253144 338494 253464 345258
rect 253144 338258 253186 338494
rect 253422 338258 253464 338494
rect 253144 331494 253464 338258
rect 253144 331258 253186 331494
rect 253422 331258 253464 331494
rect 253144 324494 253464 331258
rect 253144 324258 253186 324494
rect 253422 324258 253464 324494
rect 253144 317494 253464 324258
rect 253144 317258 253186 317494
rect 253422 317258 253464 317494
rect 253144 310494 253464 317258
rect 253144 310258 253186 310494
rect 253422 310258 253464 310494
rect 253144 303494 253464 310258
rect 253144 303258 253186 303494
rect 253422 303258 253464 303494
rect 253144 296494 253464 303258
rect 253144 296258 253186 296494
rect 253422 296258 253464 296494
rect 253144 289494 253464 296258
rect 253144 289258 253186 289494
rect 253422 289258 253464 289494
rect 253144 282494 253464 289258
rect 253144 282258 253186 282494
rect 253422 282258 253464 282494
rect 253144 275494 253464 282258
rect 253144 275258 253186 275494
rect 253422 275258 253464 275494
rect 253144 268494 253464 275258
rect 253144 268258 253186 268494
rect 253422 268258 253464 268494
rect 253144 261494 253464 268258
rect 253144 261258 253186 261494
rect 253422 261258 253464 261494
rect 253144 254494 253464 261258
rect 253144 254258 253186 254494
rect 253422 254258 253464 254494
rect 253144 247494 253464 254258
rect 253144 247258 253186 247494
rect 253422 247258 253464 247494
rect 253144 240494 253464 247258
rect 253144 240258 253186 240494
rect 253422 240258 253464 240494
rect 253144 233494 253464 240258
rect 253144 233258 253186 233494
rect 253422 233258 253464 233494
rect 253144 226494 253464 233258
rect 253144 226258 253186 226494
rect 253422 226258 253464 226494
rect 253144 219494 253464 226258
rect 253144 219258 253186 219494
rect 253422 219258 253464 219494
rect 253144 212494 253464 219258
rect 253144 212258 253186 212494
rect 253422 212258 253464 212494
rect 253144 205494 253464 212258
rect 253144 205258 253186 205494
rect 253422 205258 253464 205494
rect 253144 198494 253464 205258
rect 253144 198258 253186 198494
rect 253422 198258 253464 198494
rect 253144 191494 253464 198258
rect 253144 191258 253186 191494
rect 253422 191258 253464 191494
rect 253144 184494 253464 191258
rect 253144 184258 253186 184494
rect 253422 184258 253464 184494
rect 253144 177494 253464 184258
rect 253144 177258 253186 177494
rect 253422 177258 253464 177494
rect 253144 170494 253464 177258
rect 253144 170258 253186 170494
rect 253422 170258 253464 170494
rect 253144 163494 253464 170258
rect 253144 163258 253186 163494
rect 253422 163258 253464 163494
rect 253144 156494 253464 163258
rect 253144 156258 253186 156494
rect 253422 156258 253464 156494
rect 253144 149494 253464 156258
rect 253144 149258 253186 149494
rect 253422 149258 253464 149494
rect 253144 142494 253464 149258
rect 253144 142258 253186 142494
rect 253422 142258 253464 142494
rect 253144 135494 253464 142258
rect 253144 135258 253186 135494
rect 253422 135258 253464 135494
rect 253144 128494 253464 135258
rect 253144 128258 253186 128494
rect 253422 128258 253464 128494
rect 253144 121494 253464 128258
rect 253144 121258 253186 121494
rect 253422 121258 253464 121494
rect 253144 114494 253464 121258
rect 253144 114258 253186 114494
rect 253422 114258 253464 114494
rect 253144 107494 253464 114258
rect 253144 107258 253186 107494
rect 253422 107258 253464 107494
rect 253144 100494 253464 107258
rect 253144 100258 253186 100494
rect 253422 100258 253464 100494
rect 253144 93494 253464 100258
rect 253144 93258 253186 93494
rect 253422 93258 253464 93494
rect 253144 86494 253464 93258
rect 253144 86258 253186 86494
rect 253422 86258 253464 86494
rect 253144 79494 253464 86258
rect 253144 79258 253186 79494
rect 253422 79258 253464 79494
rect 253144 72494 253464 79258
rect 253144 72258 253186 72494
rect 253422 72258 253464 72494
rect 253144 65494 253464 72258
rect 253144 65258 253186 65494
rect 253422 65258 253464 65494
rect 253144 58494 253464 65258
rect 253144 58258 253186 58494
rect 253422 58258 253464 58494
rect 253144 51494 253464 58258
rect 253144 51258 253186 51494
rect 253422 51258 253464 51494
rect 253144 44494 253464 51258
rect 253144 44258 253186 44494
rect 253422 44258 253464 44494
rect 253144 37494 253464 44258
rect 253144 37258 253186 37494
rect 253422 37258 253464 37494
rect 253144 30494 253464 37258
rect 253144 30258 253186 30494
rect 253422 30258 253464 30494
rect 253144 23494 253464 30258
rect 253144 23258 253186 23494
rect 253422 23258 253464 23494
rect 253144 16494 253464 23258
rect 253144 16258 253186 16494
rect 253422 16258 253464 16494
rect 253144 9494 253464 16258
rect 253144 9258 253186 9494
rect 253422 9258 253464 9494
rect 253144 2494 253464 9258
rect 253144 2258 253186 2494
rect 253422 2258 253464 2494
rect 253144 -746 253464 2258
rect 253144 -982 253186 -746
rect 253422 -982 253464 -746
rect 253144 -1066 253464 -982
rect 253144 -1302 253186 -1066
rect 253422 -1302 253464 -1066
rect 253144 -2294 253464 -1302
rect 254876 706198 255196 706230
rect 254876 705962 254918 706198
rect 255154 705962 255196 706198
rect 254876 705878 255196 705962
rect 254876 705642 254918 705878
rect 255154 705642 255196 705878
rect 254876 696434 255196 705642
rect 254876 696198 254918 696434
rect 255154 696198 255196 696434
rect 254876 689434 255196 696198
rect 254876 689198 254918 689434
rect 255154 689198 255196 689434
rect 254876 682434 255196 689198
rect 254876 682198 254918 682434
rect 255154 682198 255196 682434
rect 254876 675434 255196 682198
rect 254876 675198 254918 675434
rect 255154 675198 255196 675434
rect 254876 668434 255196 675198
rect 254876 668198 254918 668434
rect 255154 668198 255196 668434
rect 254876 661434 255196 668198
rect 254876 661198 254918 661434
rect 255154 661198 255196 661434
rect 254876 654434 255196 661198
rect 254876 654198 254918 654434
rect 255154 654198 255196 654434
rect 254876 647434 255196 654198
rect 254876 647198 254918 647434
rect 255154 647198 255196 647434
rect 254876 640434 255196 647198
rect 254876 640198 254918 640434
rect 255154 640198 255196 640434
rect 254876 633434 255196 640198
rect 254876 633198 254918 633434
rect 255154 633198 255196 633434
rect 254876 626434 255196 633198
rect 254876 626198 254918 626434
rect 255154 626198 255196 626434
rect 254876 619434 255196 626198
rect 254876 619198 254918 619434
rect 255154 619198 255196 619434
rect 254876 612434 255196 619198
rect 254876 612198 254918 612434
rect 255154 612198 255196 612434
rect 254876 605434 255196 612198
rect 254876 605198 254918 605434
rect 255154 605198 255196 605434
rect 254876 598434 255196 605198
rect 254876 598198 254918 598434
rect 255154 598198 255196 598434
rect 254876 591434 255196 598198
rect 254876 591198 254918 591434
rect 255154 591198 255196 591434
rect 254876 584434 255196 591198
rect 254876 584198 254918 584434
rect 255154 584198 255196 584434
rect 254876 577434 255196 584198
rect 254876 577198 254918 577434
rect 255154 577198 255196 577434
rect 254876 570434 255196 577198
rect 254876 570198 254918 570434
rect 255154 570198 255196 570434
rect 254876 563434 255196 570198
rect 254876 563198 254918 563434
rect 255154 563198 255196 563434
rect 254876 556434 255196 563198
rect 254876 556198 254918 556434
rect 255154 556198 255196 556434
rect 254876 549434 255196 556198
rect 254876 549198 254918 549434
rect 255154 549198 255196 549434
rect 254876 542434 255196 549198
rect 254876 542198 254918 542434
rect 255154 542198 255196 542434
rect 254876 535434 255196 542198
rect 254876 535198 254918 535434
rect 255154 535198 255196 535434
rect 254876 528434 255196 535198
rect 254876 528198 254918 528434
rect 255154 528198 255196 528434
rect 254876 521434 255196 528198
rect 254876 521198 254918 521434
rect 255154 521198 255196 521434
rect 254876 514434 255196 521198
rect 254876 514198 254918 514434
rect 255154 514198 255196 514434
rect 254876 507434 255196 514198
rect 254876 507198 254918 507434
rect 255154 507198 255196 507434
rect 254876 500434 255196 507198
rect 254876 500198 254918 500434
rect 255154 500198 255196 500434
rect 254876 493434 255196 500198
rect 254876 493198 254918 493434
rect 255154 493198 255196 493434
rect 254876 486434 255196 493198
rect 254876 486198 254918 486434
rect 255154 486198 255196 486434
rect 254876 479434 255196 486198
rect 254876 479198 254918 479434
rect 255154 479198 255196 479434
rect 254876 472434 255196 479198
rect 254876 472198 254918 472434
rect 255154 472198 255196 472434
rect 254876 465434 255196 472198
rect 254876 465198 254918 465434
rect 255154 465198 255196 465434
rect 254876 458434 255196 465198
rect 254876 458198 254918 458434
rect 255154 458198 255196 458434
rect 254876 451434 255196 458198
rect 254876 451198 254918 451434
rect 255154 451198 255196 451434
rect 254876 444434 255196 451198
rect 254876 444198 254918 444434
rect 255154 444198 255196 444434
rect 254876 437434 255196 444198
rect 254876 437198 254918 437434
rect 255154 437198 255196 437434
rect 254876 430434 255196 437198
rect 254876 430198 254918 430434
rect 255154 430198 255196 430434
rect 254876 423434 255196 430198
rect 254876 423198 254918 423434
rect 255154 423198 255196 423434
rect 254876 416434 255196 423198
rect 254876 416198 254918 416434
rect 255154 416198 255196 416434
rect 254876 409434 255196 416198
rect 254876 409198 254918 409434
rect 255154 409198 255196 409434
rect 254876 402434 255196 409198
rect 254876 402198 254918 402434
rect 255154 402198 255196 402434
rect 254876 395434 255196 402198
rect 254876 395198 254918 395434
rect 255154 395198 255196 395434
rect 254876 388434 255196 395198
rect 254876 388198 254918 388434
rect 255154 388198 255196 388434
rect 254876 381434 255196 388198
rect 254876 381198 254918 381434
rect 255154 381198 255196 381434
rect 254876 374434 255196 381198
rect 254876 374198 254918 374434
rect 255154 374198 255196 374434
rect 254876 367434 255196 374198
rect 254876 367198 254918 367434
rect 255154 367198 255196 367434
rect 254876 360434 255196 367198
rect 254876 360198 254918 360434
rect 255154 360198 255196 360434
rect 254876 353434 255196 360198
rect 254876 353198 254918 353434
rect 255154 353198 255196 353434
rect 254876 346434 255196 353198
rect 254876 346198 254918 346434
rect 255154 346198 255196 346434
rect 254876 339434 255196 346198
rect 254876 339198 254918 339434
rect 255154 339198 255196 339434
rect 254876 332434 255196 339198
rect 254876 332198 254918 332434
rect 255154 332198 255196 332434
rect 254876 325434 255196 332198
rect 254876 325198 254918 325434
rect 255154 325198 255196 325434
rect 254876 318434 255196 325198
rect 254876 318198 254918 318434
rect 255154 318198 255196 318434
rect 254876 311434 255196 318198
rect 254876 311198 254918 311434
rect 255154 311198 255196 311434
rect 254876 304434 255196 311198
rect 254876 304198 254918 304434
rect 255154 304198 255196 304434
rect 254876 297434 255196 304198
rect 254876 297198 254918 297434
rect 255154 297198 255196 297434
rect 254876 290434 255196 297198
rect 254876 290198 254918 290434
rect 255154 290198 255196 290434
rect 254876 283434 255196 290198
rect 254876 283198 254918 283434
rect 255154 283198 255196 283434
rect 254876 276434 255196 283198
rect 254876 276198 254918 276434
rect 255154 276198 255196 276434
rect 254876 269434 255196 276198
rect 254876 269198 254918 269434
rect 255154 269198 255196 269434
rect 254876 262434 255196 269198
rect 254876 262198 254918 262434
rect 255154 262198 255196 262434
rect 254876 255434 255196 262198
rect 254876 255198 254918 255434
rect 255154 255198 255196 255434
rect 254876 248434 255196 255198
rect 254876 248198 254918 248434
rect 255154 248198 255196 248434
rect 254876 241434 255196 248198
rect 254876 241198 254918 241434
rect 255154 241198 255196 241434
rect 254876 234434 255196 241198
rect 254876 234198 254918 234434
rect 255154 234198 255196 234434
rect 254876 227434 255196 234198
rect 254876 227198 254918 227434
rect 255154 227198 255196 227434
rect 254876 220434 255196 227198
rect 254876 220198 254918 220434
rect 255154 220198 255196 220434
rect 254876 213434 255196 220198
rect 254876 213198 254918 213434
rect 255154 213198 255196 213434
rect 254876 206434 255196 213198
rect 254876 206198 254918 206434
rect 255154 206198 255196 206434
rect 254876 199434 255196 206198
rect 254876 199198 254918 199434
rect 255154 199198 255196 199434
rect 254876 192434 255196 199198
rect 254876 192198 254918 192434
rect 255154 192198 255196 192434
rect 254876 185434 255196 192198
rect 254876 185198 254918 185434
rect 255154 185198 255196 185434
rect 254876 178434 255196 185198
rect 254876 178198 254918 178434
rect 255154 178198 255196 178434
rect 254876 171434 255196 178198
rect 254876 171198 254918 171434
rect 255154 171198 255196 171434
rect 254876 164434 255196 171198
rect 254876 164198 254918 164434
rect 255154 164198 255196 164434
rect 254876 157434 255196 164198
rect 254876 157198 254918 157434
rect 255154 157198 255196 157434
rect 254876 150434 255196 157198
rect 254876 150198 254918 150434
rect 255154 150198 255196 150434
rect 254876 143434 255196 150198
rect 254876 143198 254918 143434
rect 255154 143198 255196 143434
rect 254876 136434 255196 143198
rect 254876 136198 254918 136434
rect 255154 136198 255196 136434
rect 254876 129434 255196 136198
rect 254876 129198 254918 129434
rect 255154 129198 255196 129434
rect 254876 122434 255196 129198
rect 254876 122198 254918 122434
rect 255154 122198 255196 122434
rect 254876 115434 255196 122198
rect 254876 115198 254918 115434
rect 255154 115198 255196 115434
rect 254876 108434 255196 115198
rect 254876 108198 254918 108434
rect 255154 108198 255196 108434
rect 254876 101434 255196 108198
rect 254876 101198 254918 101434
rect 255154 101198 255196 101434
rect 254876 94434 255196 101198
rect 254876 94198 254918 94434
rect 255154 94198 255196 94434
rect 254876 87434 255196 94198
rect 254876 87198 254918 87434
rect 255154 87198 255196 87434
rect 254876 80434 255196 87198
rect 254876 80198 254918 80434
rect 255154 80198 255196 80434
rect 254876 73434 255196 80198
rect 254876 73198 254918 73434
rect 255154 73198 255196 73434
rect 254876 66434 255196 73198
rect 254876 66198 254918 66434
rect 255154 66198 255196 66434
rect 254876 59434 255196 66198
rect 254876 59198 254918 59434
rect 255154 59198 255196 59434
rect 254876 52434 255196 59198
rect 254876 52198 254918 52434
rect 255154 52198 255196 52434
rect 254876 45434 255196 52198
rect 254876 45198 254918 45434
rect 255154 45198 255196 45434
rect 254876 38434 255196 45198
rect 254876 38198 254918 38434
rect 255154 38198 255196 38434
rect 254876 31434 255196 38198
rect 254876 31198 254918 31434
rect 255154 31198 255196 31434
rect 254876 24434 255196 31198
rect 254876 24198 254918 24434
rect 255154 24198 255196 24434
rect 254876 17434 255196 24198
rect 254876 17198 254918 17434
rect 255154 17198 255196 17434
rect 254876 10434 255196 17198
rect 254876 10198 254918 10434
rect 255154 10198 255196 10434
rect 254876 3434 255196 10198
rect 254876 3198 254918 3434
rect 255154 3198 255196 3434
rect 254876 -1706 255196 3198
rect 254876 -1942 254918 -1706
rect 255154 -1942 255196 -1706
rect 254876 -2026 255196 -1942
rect 254876 -2262 254918 -2026
rect 255154 -2262 255196 -2026
rect 254876 -2294 255196 -2262
rect 260144 705238 260464 706230
rect 260144 705002 260186 705238
rect 260422 705002 260464 705238
rect 260144 704918 260464 705002
rect 260144 704682 260186 704918
rect 260422 704682 260464 704918
rect 260144 695494 260464 704682
rect 260144 695258 260186 695494
rect 260422 695258 260464 695494
rect 260144 688494 260464 695258
rect 260144 688258 260186 688494
rect 260422 688258 260464 688494
rect 260144 681494 260464 688258
rect 260144 681258 260186 681494
rect 260422 681258 260464 681494
rect 260144 674494 260464 681258
rect 260144 674258 260186 674494
rect 260422 674258 260464 674494
rect 260144 667494 260464 674258
rect 260144 667258 260186 667494
rect 260422 667258 260464 667494
rect 260144 660494 260464 667258
rect 260144 660258 260186 660494
rect 260422 660258 260464 660494
rect 260144 653494 260464 660258
rect 260144 653258 260186 653494
rect 260422 653258 260464 653494
rect 260144 646494 260464 653258
rect 260144 646258 260186 646494
rect 260422 646258 260464 646494
rect 260144 639494 260464 646258
rect 260144 639258 260186 639494
rect 260422 639258 260464 639494
rect 260144 632494 260464 639258
rect 260144 632258 260186 632494
rect 260422 632258 260464 632494
rect 260144 625494 260464 632258
rect 260144 625258 260186 625494
rect 260422 625258 260464 625494
rect 260144 618494 260464 625258
rect 260144 618258 260186 618494
rect 260422 618258 260464 618494
rect 260144 611494 260464 618258
rect 260144 611258 260186 611494
rect 260422 611258 260464 611494
rect 260144 604494 260464 611258
rect 260144 604258 260186 604494
rect 260422 604258 260464 604494
rect 260144 597494 260464 604258
rect 260144 597258 260186 597494
rect 260422 597258 260464 597494
rect 260144 590494 260464 597258
rect 260144 590258 260186 590494
rect 260422 590258 260464 590494
rect 260144 583494 260464 590258
rect 260144 583258 260186 583494
rect 260422 583258 260464 583494
rect 260144 576494 260464 583258
rect 260144 576258 260186 576494
rect 260422 576258 260464 576494
rect 260144 569494 260464 576258
rect 260144 569258 260186 569494
rect 260422 569258 260464 569494
rect 260144 562494 260464 569258
rect 260144 562258 260186 562494
rect 260422 562258 260464 562494
rect 260144 555494 260464 562258
rect 260144 555258 260186 555494
rect 260422 555258 260464 555494
rect 260144 548494 260464 555258
rect 260144 548258 260186 548494
rect 260422 548258 260464 548494
rect 260144 541494 260464 548258
rect 260144 541258 260186 541494
rect 260422 541258 260464 541494
rect 260144 534494 260464 541258
rect 260144 534258 260186 534494
rect 260422 534258 260464 534494
rect 260144 527494 260464 534258
rect 260144 527258 260186 527494
rect 260422 527258 260464 527494
rect 260144 520494 260464 527258
rect 260144 520258 260186 520494
rect 260422 520258 260464 520494
rect 260144 513494 260464 520258
rect 260144 513258 260186 513494
rect 260422 513258 260464 513494
rect 260144 506494 260464 513258
rect 260144 506258 260186 506494
rect 260422 506258 260464 506494
rect 260144 499494 260464 506258
rect 260144 499258 260186 499494
rect 260422 499258 260464 499494
rect 260144 492494 260464 499258
rect 260144 492258 260186 492494
rect 260422 492258 260464 492494
rect 260144 485494 260464 492258
rect 260144 485258 260186 485494
rect 260422 485258 260464 485494
rect 260144 478494 260464 485258
rect 260144 478258 260186 478494
rect 260422 478258 260464 478494
rect 260144 471494 260464 478258
rect 260144 471258 260186 471494
rect 260422 471258 260464 471494
rect 260144 464494 260464 471258
rect 260144 464258 260186 464494
rect 260422 464258 260464 464494
rect 260144 457494 260464 464258
rect 260144 457258 260186 457494
rect 260422 457258 260464 457494
rect 260144 450494 260464 457258
rect 260144 450258 260186 450494
rect 260422 450258 260464 450494
rect 260144 443494 260464 450258
rect 260144 443258 260186 443494
rect 260422 443258 260464 443494
rect 260144 436494 260464 443258
rect 260144 436258 260186 436494
rect 260422 436258 260464 436494
rect 260144 429494 260464 436258
rect 260144 429258 260186 429494
rect 260422 429258 260464 429494
rect 260144 422494 260464 429258
rect 260144 422258 260186 422494
rect 260422 422258 260464 422494
rect 260144 415494 260464 422258
rect 260144 415258 260186 415494
rect 260422 415258 260464 415494
rect 260144 408494 260464 415258
rect 260144 408258 260186 408494
rect 260422 408258 260464 408494
rect 260144 401494 260464 408258
rect 260144 401258 260186 401494
rect 260422 401258 260464 401494
rect 260144 394494 260464 401258
rect 260144 394258 260186 394494
rect 260422 394258 260464 394494
rect 260144 387494 260464 394258
rect 260144 387258 260186 387494
rect 260422 387258 260464 387494
rect 260144 380494 260464 387258
rect 260144 380258 260186 380494
rect 260422 380258 260464 380494
rect 260144 373494 260464 380258
rect 260144 373258 260186 373494
rect 260422 373258 260464 373494
rect 260144 366494 260464 373258
rect 260144 366258 260186 366494
rect 260422 366258 260464 366494
rect 260144 359494 260464 366258
rect 260144 359258 260186 359494
rect 260422 359258 260464 359494
rect 260144 352494 260464 359258
rect 260144 352258 260186 352494
rect 260422 352258 260464 352494
rect 260144 345494 260464 352258
rect 260144 345258 260186 345494
rect 260422 345258 260464 345494
rect 260144 338494 260464 345258
rect 260144 338258 260186 338494
rect 260422 338258 260464 338494
rect 260144 331494 260464 338258
rect 260144 331258 260186 331494
rect 260422 331258 260464 331494
rect 260144 324494 260464 331258
rect 260144 324258 260186 324494
rect 260422 324258 260464 324494
rect 260144 317494 260464 324258
rect 260144 317258 260186 317494
rect 260422 317258 260464 317494
rect 260144 310494 260464 317258
rect 260144 310258 260186 310494
rect 260422 310258 260464 310494
rect 260144 303494 260464 310258
rect 260144 303258 260186 303494
rect 260422 303258 260464 303494
rect 260144 296494 260464 303258
rect 260144 296258 260186 296494
rect 260422 296258 260464 296494
rect 260144 289494 260464 296258
rect 260144 289258 260186 289494
rect 260422 289258 260464 289494
rect 260144 282494 260464 289258
rect 260144 282258 260186 282494
rect 260422 282258 260464 282494
rect 260144 275494 260464 282258
rect 260144 275258 260186 275494
rect 260422 275258 260464 275494
rect 260144 268494 260464 275258
rect 260144 268258 260186 268494
rect 260422 268258 260464 268494
rect 260144 261494 260464 268258
rect 260144 261258 260186 261494
rect 260422 261258 260464 261494
rect 260144 254494 260464 261258
rect 260144 254258 260186 254494
rect 260422 254258 260464 254494
rect 260144 247494 260464 254258
rect 260144 247258 260186 247494
rect 260422 247258 260464 247494
rect 260144 240494 260464 247258
rect 260144 240258 260186 240494
rect 260422 240258 260464 240494
rect 260144 233494 260464 240258
rect 260144 233258 260186 233494
rect 260422 233258 260464 233494
rect 260144 226494 260464 233258
rect 260144 226258 260186 226494
rect 260422 226258 260464 226494
rect 260144 219494 260464 226258
rect 260144 219258 260186 219494
rect 260422 219258 260464 219494
rect 260144 212494 260464 219258
rect 260144 212258 260186 212494
rect 260422 212258 260464 212494
rect 260144 205494 260464 212258
rect 260144 205258 260186 205494
rect 260422 205258 260464 205494
rect 260144 198494 260464 205258
rect 260144 198258 260186 198494
rect 260422 198258 260464 198494
rect 260144 191494 260464 198258
rect 260144 191258 260186 191494
rect 260422 191258 260464 191494
rect 260144 184494 260464 191258
rect 260144 184258 260186 184494
rect 260422 184258 260464 184494
rect 260144 177494 260464 184258
rect 260144 177258 260186 177494
rect 260422 177258 260464 177494
rect 260144 170494 260464 177258
rect 260144 170258 260186 170494
rect 260422 170258 260464 170494
rect 260144 163494 260464 170258
rect 260144 163258 260186 163494
rect 260422 163258 260464 163494
rect 260144 156494 260464 163258
rect 260144 156258 260186 156494
rect 260422 156258 260464 156494
rect 260144 149494 260464 156258
rect 260144 149258 260186 149494
rect 260422 149258 260464 149494
rect 260144 142494 260464 149258
rect 260144 142258 260186 142494
rect 260422 142258 260464 142494
rect 260144 135494 260464 142258
rect 260144 135258 260186 135494
rect 260422 135258 260464 135494
rect 260144 128494 260464 135258
rect 260144 128258 260186 128494
rect 260422 128258 260464 128494
rect 260144 121494 260464 128258
rect 260144 121258 260186 121494
rect 260422 121258 260464 121494
rect 260144 114494 260464 121258
rect 260144 114258 260186 114494
rect 260422 114258 260464 114494
rect 260144 107494 260464 114258
rect 260144 107258 260186 107494
rect 260422 107258 260464 107494
rect 260144 100494 260464 107258
rect 260144 100258 260186 100494
rect 260422 100258 260464 100494
rect 260144 93494 260464 100258
rect 260144 93258 260186 93494
rect 260422 93258 260464 93494
rect 260144 86494 260464 93258
rect 260144 86258 260186 86494
rect 260422 86258 260464 86494
rect 260144 79494 260464 86258
rect 260144 79258 260186 79494
rect 260422 79258 260464 79494
rect 260144 72494 260464 79258
rect 260144 72258 260186 72494
rect 260422 72258 260464 72494
rect 260144 65494 260464 72258
rect 260144 65258 260186 65494
rect 260422 65258 260464 65494
rect 260144 58494 260464 65258
rect 260144 58258 260186 58494
rect 260422 58258 260464 58494
rect 260144 51494 260464 58258
rect 260144 51258 260186 51494
rect 260422 51258 260464 51494
rect 260144 44494 260464 51258
rect 260144 44258 260186 44494
rect 260422 44258 260464 44494
rect 260144 37494 260464 44258
rect 260144 37258 260186 37494
rect 260422 37258 260464 37494
rect 260144 30494 260464 37258
rect 260144 30258 260186 30494
rect 260422 30258 260464 30494
rect 260144 23494 260464 30258
rect 260144 23258 260186 23494
rect 260422 23258 260464 23494
rect 260144 16494 260464 23258
rect 260144 16258 260186 16494
rect 260422 16258 260464 16494
rect 260144 9494 260464 16258
rect 260144 9258 260186 9494
rect 260422 9258 260464 9494
rect 260144 2494 260464 9258
rect 260144 2258 260186 2494
rect 260422 2258 260464 2494
rect 260144 -746 260464 2258
rect 260144 -982 260186 -746
rect 260422 -982 260464 -746
rect 260144 -1066 260464 -982
rect 260144 -1302 260186 -1066
rect 260422 -1302 260464 -1066
rect 260144 -2294 260464 -1302
rect 261876 706198 262196 706230
rect 261876 705962 261918 706198
rect 262154 705962 262196 706198
rect 261876 705878 262196 705962
rect 261876 705642 261918 705878
rect 262154 705642 262196 705878
rect 261876 696434 262196 705642
rect 261876 696198 261918 696434
rect 262154 696198 262196 696434
rect 261876 689434 262196 696198
rect 261876 689198 261918 689434
rect 262154 689198 262196 689434
rect 261876 682434 262196 689198
rect 261876 682198 261918 682434
rect 262154 682198 262196 682434
rect 261876 675434 262196 682198
rect 261876 675198 261918 675434
rect 262154 675198 262196 675434
rect 261876 668434 262196 675198
rect 261876 668198 261918 668434
rect 262154 668198 262196 668434
rect 261876 661434 262196 668198
rect 261876 661198 261918 661434
rect 262154 661198 262196 661434
rect 261876 654434 262196 661198
rect 261876 654198 261918 654434
rect 262154 654198 262196 654434
rect 261876 647434 262196 654198
rect 261876 647198 261918 647434
rect 262154 647198 262196 647434
rect 261876 640434 262196 647198
rect 261876 640198 261918 640434
rect 262154 640198 262196 640434
rect 261876 633434 262196 640198
rect 261876 633198 261918 633434
rect 262154 633198 262196 633434
rect 261876 626434 262196 633198
rect 261876 626198 261918 626434
rect 262154 626198 262196 626434
rect 261876 619434 262196 626198
rect 261876 619198 261918 619434
rect 262154 619198 262196 619434
rect 261876 612434 262196 619198
rect 261876 612198 261918 612434
rect 262154 612198 262196 612434
rect 261876 605434 262196 612198
rect 261876 605198 261918 605434
rect 262154 605198 262196 605434
rect 261876 598434 262196 605198
rect 261876 598198 261918 598434
rect 262154 598198 262196 598434
rect 261876 591434 262196 598198
rect 261876 591198 261918 591434
rect 262154 591198 262196 591434
rect 261876 584434 262196 591198
rect 261876 584198 261918 584434
rect 262154 584198 262196 584434
rect 261876 577434 262196 584198
rect 261876 577198 261918 577434
rect 262154 577198 262196 577434
rect 261876 570434 262196 577198
rect 261876 570198 261918 570434
rect 262154 570198 262196 570434
rect 261876 563434 262196 570198
rect 261876 563198 261918 563434
rect 262154 563198 262196 563434
rect 261876 556434 262196 563198
rect 261876 556198 261918 556434
rect 262154 556198 262196 556434
rect 261876 549434 262196 556198
rect 261876 549198 261918 549434
rect 262154 549198 262196 549434
rect 261876 542434 262196 549198
rect 261876 542198 261918 542434
rect 262154 542198 262196 542434
rect 261876 535434 262196 542198
rect 261876 535198 261918 535434
rect 262154 535198 262196 535434
rect 261876 528434 262196 535198
rect 261876 528198 261918 528434
rect 262154 528198 262196 528434
rect 261876 521434 262196 528198
rect 261876 521198 261918 521434
rect 262154 521198 262196 521434
rect 261876 514434 262196 521198
rect 261876 514198 261918 514434
rect 262154 514198 262196 514434
rect 261876 507434 262196 514198
rect 261876 507198 261918 507434
rect 262154 507198 262196 507434
rect 261876 500434 262196 507198
rect 261876 500198 261918 500434
rect 262154 500198 262196 500434
rect 261876 493434 262196 500198
rect 261876 493198 261918 493434
rect 262154 493198 262196 493434
rect 261876 486434 262196 493198
rect 261876 486198 261918 486434
rect 262154 486198 262196 486434
rect 261876 479434 262196 486198
rect 261876 479198 261918 479434
rect 262154 479198 262196 479434
rect 261876 472434 262196 479198
rect 261876 472198 261918 472434
rect 262154 472198 262196 472434
rect 261876 465434 262196 472198
rect 261876 465198 261918 465434
rect 262154 465198 262196 465434
rect 261876 458434 262196 465198
rect 261876 458198 261918 458434
rect 262154 458198 262196 458434
rect 261876 451434 262196 458198
rect 261876 451198 261918 451434
rect 262154 451198 262196 451434
rect 261876 444434 262196 451198
rect 261876 444198 261918 444434
rect 262154 444198 262196 444434
rect 261876 437434 262196 444198
rect 261876 437198 261918 437434
rect 262154 437198 262196 437434
rect 261876 430434 262196 437198
rect 261876 430198 261918 430434
rect 262154 430198 262196 430434
rect 261876 423434 262196 430198
rect 261876 423198 261918 423434
rect 262154 423198 262196 423434
rect 261876 416434 262196 423198
rect 261876 416198 261918 416434
rect 262154 416198 262196 416434
rect 261876 409434 262196 416198
rect 261876 409198 261918 409434
rect 262154 409198 262196 409434
rect 261876 402434 262196 409198
rect 261876 402198 261918 402434
rect 262154 402198 262196 402434
rect 261876 395434 262196 402198
rect 261876 395198 261918 395434
rect 262154 395198 262196 395434
rect 261876 388434 262196 395198
rect 261876 388198 261918 388434
rect 262154 388198 262196 388434
rect 261876 381434 262196 388198
rect 261876 381198 261918 381434
rect 262154 381198 262196 381434
rect 261876 374434 262196 381198
rect 261876 374198 261918 374434
rect 262154 374198 262196 374434
rect 261876 367434 262196 374198
rect 261876 367198 261918 367434
rect 262154 367198 262196 367434
rect 261876 360434 262196 367198
rect 261876 360198 261918 360434
rect 262154 360198 262196 360434
rect 261876 353434 262196 360198
rect 261876 353198 261918 353434
rect 262154 353198 262196 353434
rect 261876 346434 262196 353198
rect 261876 346198 261918 346434
rect 262154 346198 262196 346434
rect 261876 339434 262196 346198
rect 261876 339198 261918 339434
rect 262154 339198 262196 339434
rect 261876 332434 262196 339198
rect 261876 332198 261918 332434
rect 262154 332198 262196 332434
rect 261876 325434 262196 332198
rect 261876 325198 261918 325434
rect 262154 325198 262196 325434
rect 261876 318434 262196 325198
rect 261876 318198 261918 318434
rect 262154 318198 262196 318434
rect 261876 311434 262196 318198
rect 261876 311198 261918 311434
rect 262154 311198 262196 311434
rect 261876 304434 262196 311198
rect 261876 304198 261918 304434
rect 262154 304198 262196 304434
rect 261876 297434 262196 304198
rect 261876 297198 261918 297434
rect 262154 297198 262196 297434
rect 261876 290434 262196 297198
rect 261876 290198 261918 290434
rect 262154 290198 262196 290434
rect 261876 283434 262196 290198
rect 261876 283198 261918 283434
rect 262154 283198 262196 283434
rect 261876 276434 262196 283198
rect 261876 276198 261918 276434
rect 262154 276198 262196 276434
rect 261876 269434 262196 276198
rect 261876 269198 261918 269434
rect 262154 269198 262196 269434
rect 261876 262434 262196 269198
rect 261876 262198 261918 262434
rect 262154 262198 262196 262434
rect 261876 255434 262196 262198
rect 261876 255198 261918 255434
rect 262154 255198 262196 255434
rect 261876 248434 262196 255198
rect 261876 248198 261918 248434
rect 262154 248198 262196 248434
rect 261876 241434 262196 248198
rect 261876 241198 261918 241434
rect 262154 241198 262196 241434
rect 261876 234434 262196 241198
rect 261876 234198 261918 234434
rect 262154 234198 262196 234434
rect 261876 227434 262196 234198
rect 261876 227198 261918 227434
rect 262154 227198 262196 227434
rect 261876 220434 262196 227198
rect 261876 220198 261918 220434
rect 262154 220198 262196 220434
rect 261876 213434 262196 220198
rect 261876 213198 261918 213434
rect 262154 213198 262196 213434
rect 261876 206434 262196 213198
rect 261876 206198 261918 206434
rect 262154 206198 262196 206434
rect 261876 199434 262196 206198
rect 261876 199198 261918 199434
rect 262154 199198 262196 199434
rect 261876 192434 262196 199198
rect 261876 192198 261918 192434
rect 262154 192198 262196 192434
rect 261876 185434 262196 192198
rect 261876 185198 261918 185434
rect 262154 185198 262196 185434
rect 261876 178434 262196 185198
rect 261876 178198 261918 178434
rect 262154 178198 262196 178434
rect 261876 171434 262196 178198
rect 261876 171198 261918 171434
rect 262154 171198 262196 171434
rect 261876 164434 262196 171198
rect 261876 164198 261918 164434
rect 262154 164198 262196 164434
rect 261876 157434 262196 164198
rect 261876 157198 261918 157434
rect 262154 157198 262196 157434
rect 261876 150434 262196 157198
rect 261876 150198 261918 150434
rect 262154 150198 262196 150434
rect 261876 143434 262196 150198
rect 261876 143198 261918 143434
rect 262154 143198 262196 143434
rect 261876 136434 262196 143198
rect 261876 136198 261918 136434
rect 262154 136198 262196 136434
rect 261876 129434 262196 136198
rect 261876 129198 261918 129434
rect 262154 129198 262196 129434
rect 261876 122434 262196 129198
rect 261876 122198 261918 122434
rect 262154 122198 262196 122434
rect 261876 115434 262196 122198
rect 261876 115198 261918 115434
rect 262154 115198 262196 115434
rect 261876 108434 262196 115198
rect 261876 108198 261918 108434
rect 262154 108198 262196 108434
rect 261876 101434 262196 108198
rect 261876 101198 261918 101434
rect 262154 101198 262196 101434
rect 261876 94434 262196 101198
rect 261876 94198 261918 94434
rect 262154 94198 262196 94434
rect 261876 87434 262196 94198
rect 261876 87198 261918 87434
rect 262154 87198 262196 87434
rect 261876 80434 262196 87198
rect 261876 80198 261918 80434
rect 262154 80198 262196 80434
rect 261876 73434 262196 80198
rect 261876 73198 261918 73434
rect 262154 73198 262196 73434
rect 261876 66434 262196 73198
rect 261876 66198 261918 66434
rect 262154 66198 262196 66434
rect 261876 59434 262196 66198
rect 261876 59198 261918 59434
rect 262154 59198 262196 59434
rect 261876 52434 262196 59198
rect 261876 52198 261918 52434
rect 262154 52198 262196 52434
rect 261876 45434 262196 52198
rect 261876 45198 261918 45434
rect 262154 45198 262196 45434
rect 261876 38434 262196 45198
rect 261876 38198 261918 38434
rect 262154 38198 262196 38434
rect 261876 31434 262196 38198
rect 261876 31198 261918 31434
rect 262154 31198 262196 31434
rect 261876 24434 262196 31198
rect 261876 24198 261918 24434
rect 262154 24198 262196 24434
rect 261876 17434 262196 24198
rect 261876 17198 261918 17434
rect 262154 17198 262196 17434
rect 261876 10434 262196 17198
rect 261876 10198 261918 10434
rect 262154 10198 262196 10434
rect 261876 3434 262196 10198
rect 261876 3198 261918 3434
rect 262154 3198 262196 3434
rect 261876 -1706 262196 3198
rect 261876 -1942 261918 -1706
rect 262154 -1942 262196 -1706
rect 261876 -2026 262196 -1942
rect 261876 -2262 261918 -2026
rect 262154 -2262 262196 -2026
rect 261876 -2294 262196 -2262
rect 267144 705238 267464 706230
rect 267144 705002 267186 705238
rect 267422 705002 267464 705238
rect 267144 704918 267464 705002
rect 267144 704682 267186 704918
rect 267422 704682 267464 704918
rect 267144 695494 267464 704682
rect 267144 695258 267186 695494
rect 267422 695258 267464 695494
rect 267144 688494 267464 695258
rect 267144 688258 267186 688494
rect 267422 688258 267464 688494
rect 267144 681494 267464 688258
rect 267144 681258 267186 681494
rect 267422 681258 267464 681494
rect 267144 674494 267464 681258
rect 267144 674258 267186 674494
rect 267422 674258 267464 674494
rect 267144 667494 267464 674258
rect 267144 667258 267186 667494
rect 267422 667258 267464 667494
rect 267144 660494 267464 667258
rect 267144 660258 267186 660494
rect 267422 660258 267464 660494
rect 267144 653494 267464 660258
rect 267144 653258 267186 653494
rect 267422 653258 267464 653494
rect 267144 646494 267464 653258
rect 267144 646258 267186 646494
rect 267422 646258 267464 646494
rect 267144 639494 267464 646258
rect 267144 639258 267186 639494
rect 267422 639258 267464 639494
rect 267144 632494 267464 639258
rect 267144 632258 267186 632494
rect 267422 632258 267464 632494
rect 267144 625494 267464 632258
rect 267144 625258 267186 625494
rect 267422 625258 267464 625494
rect 267144 618494 267464 625258
rect 267144 618258 267186 618494
rect 267422 618258 267464 618494
rect 267144 611494 267464 618258
rect 267144 611258 267186 611494
rect 267422 611258 267464 611494
rect 267144 604494 267464 611258
rect 267144 604258 267186 604494
rect 267422 604258 267464 604494
rect 267144 597494 267464 604258
rect 267144 597258 267186 597494
rect 267422 597258 267464 597494
rect 267144 590494 267464 597258
rect 267144 590258 267186 590494
rect 267422 590258 267464 590494
rect 267144 583494 267464 590258
rect 267144 583258 267186 583494
rect 267422 583258 267464 583494
rect 267144 576494 267464 583258
rect 267144 576258 267186 576494
rect 267422 576258 267464 576494
rect 267144 569494 267464 576258
rect 267144 569258 267186 569494
rect 267422 569258 267464 569494
rect 267144 562494 267464 569258
rect 267144 562258 267186 562494
rect 267422 562258 267464 562494
rect 267144 555494 267464 562258
rect 267144 555258 267186 555494
rect 267422 555258 267464 555494
rect 267144 548494 267464 555258
rect 267144 548258 267186 548494
rect 267422 548258 267464 548494
rect 267144 541494 267464 548258
rect 267144 541258 267186 541494
rect 267422 541258 267464 541494
rect 267144 534494 267464 541258
rect 267144 534258 267186 534494
rect 267422 534258 267464 534494
rect 267144 527494 267464 534258
rect 267144 527258 267186 527494
rect 267422 527258 267464 527494
rect 267144 520494 267464 527258
rect 267144 520258 267186 520494
rect 267422 520258 267464 520494
rect 267144 513494 267464 520258
rect 267144 513258 267186 513494
rect 267422 513258 267464 513494
rect 267144 506494 267464 513258
rect 267144 506258 267186 506494
rect 267422 506258 267464 506494
rect 267144 499494 267464 506258
rect 267144 499258 267186 499494
rect 267422 499258 267464 499494
rect 267144 492494 267464 499258
rect 267144 492258 267186 492494
rect 267422 492258 267464 492494
rect 267144 485494 267464 492258
rect 267144 485258 267186 485494
rect 267422 485258 267464 485494
rect 267144 478494 267464 485258
rect 267144 478258 267186 478494
rect 267422 478258 267464 478494
rect 267144 471494 267464 478258
rect 267144 471258 267186 471494
rect 267422 471258 267464 471494
rect 267144 464494 267464 471258
rect 267144 464258 267186 464494
rect 267422 464258 267464 464494
rect 267144 457494 267464 464258
rect 267144 457258 267186 457494
rect 267422 457258 267464 457494
rect 267144 450494 267464 457258
rect 267144 450258 267186 450494
rect 267422 450258 267464 450494
rect 267144 443494 267464 450258
rect 267144 443258 267186 443494
rect 267422 443258 267464 443494
rect 267144 436494 267464 443258
rect 267144 436258 267186 436494
rect 267422 436258 267464 436494
rect 267144 429494 267464 436258
rect 267144 429258 267186 429494
rect 267422 429258 267464 429494
rect 267144 422494 267464 429258
rect 267144 422258 267186 422494
rect 267422 422258 267464 422494
rect 267144 415494 267464 422258
rect 267144 415258 267186 415494
rect 267422 415258 267464 415494
rect 267144 408494 267464 415258
rect 267144 408258 267186 408494
rect 267422 408258 267464 408494
rect 267144 401494 267464 408258
rect 267144 401258 267186 401494
rect 267422 401258 267464 401494
rect 267144 394494 267464 401258
rect 267144 394258 267186 394494
rect 267422 394258 267464 394494
rect 267144 387494 267464 394258
rect 267144 387258 267186 387494
rect 267422 387258 267464 387494
rect 267144 380494 267464 387258
rect 267144 380258 267186 380494
rect 267422 380258 267464 380494
rect 267144 373494 267464 380258
rect 267144 373258 267186 373494
rect 267422 373258 267464 373494
rect 267144 366494 267464 373258
rect 267144 366258 267186 366494
rect 267422 366258 267464 366494
rect 267144 359494 267464 366258
rect 267144 359258 267186 359494
rect 267422 359258 267464 359494
rect 267144 352494 267464 359258
rect 267144 352258 267186 352494
rect 267422 352258 267464 352494
rect 267144 345494 267464 352258
rect 267144 345258 267186 345494
rect 267422 345258 267464 345494
rect 267144 338494 267464 345258
rect 267144 338258 267186 338494
rect 267422 338258 267464 338494
rect 267144 331494 267464 338258
rect 267144 331258 267186 331494
rect 267422 331258 267464 331494
rect 267144 324494 267464 331258
rect 267144 324258 267186 324494
rect 267422 324258 267464 324494
rect 267144 317494 267464 324258
rect 267144 317258 267186 317494
rect 267422 317258 267464 317494
rect 267144 310494 267464 317258
rect 267144 310258 267186 310494
rect 267422 310258 267464 310494
rect 267144 303494 267464 310258
rect 267144 303258 267186 303494
rect 267422 303258 267464 303494
rect 267144 296494 267464 303258
rect 267144 296258 267186 296494
rect 267422 296258 267464 296494
rect 267144 289494 267464 296258
rect 267144 289258 267186 289494
rect 267422 289258 267464 289494
rect 267144 282494 267464 289258
rect 267144 282258 267186 282494
rect 267422 282258 267464 282494
rect 267144 275494 267464 282258
rect 267144 275258 267186 275494
rect 267422 275258 267464 275494
rect 267144 268494 267464 275258
rect 267144 268258 267186 268494
rect 267422 268258 267464 268494
rect 267144 261494 267464 268258
rect 267144 261258 267186 261494
rect 267422 261258 267464 261494
rect 267144 254494 267464 261258
rect 267144 254258 267186 254494
rect 267422 254258 267464 254494
rect 267144 247494 267464 254258
rect 267144 247258 267186 247494
rect 267422 247258 267464 247494
rect 267144 240494 267464 247258
rect 267144 240258 267186 240494
rect 267422 240258 267464 240494
rect 267144 233494 267464 240258
rect 267144 233258 267186 233494
rect 267422 233258 267464 233494
rect 267144 226494 267464 233258
rect 267144 226258 267186 226494
rect 267422 226258 267464 226494
rect 267144 219494 267464 226258
rect 267144 219258 267186 219494
rect 267422 219258 267464 219494
rect 267144 212494 267464 219258
rect 267144 212258 267186 212494
rect 267422 212258 267464 212494
rect 267144 205494 267464 212258
rect 267144 205258 267186 205494
rect 267422 205258 267464 205494
rect 267144 198494 267464 205258
rect 267144 198258 267186 198494
rect 267422 198258 267464 198494
rect 267144 191494 267464 198258
rect 267144 191258 267186 191494
rect 267422 191258 267464 191494
rect 267144 184494 267464 191258
rect 267144 184258 267186 184494
rect 267422 184258 267464 184494
rect 267144 177494 267464 184258
rect 267144 177258 267186 177494
rect 267422 177258 267464 177494
rect 267144 170494 267464 177258
rect 267144 170258 267186 170494
rect 267422 170258 267464 170494
rect 267144 163494 267464 170258
rect 267144 163258 267186 163494
rect 267422 163258 267464 163494
rect 267144 156494 267464 163258
rect 267144 156258 267186 156494
rect 267422 156258 267464 156494
rect 267144 149494 267464 156258
rect 267144 149258 267186 149494
rect 267422 149258 267464 149494
rect 267144 142494 267464 149258
rect 267144 142258 267186 142494
rect 267422 142258 267464 142494
rect 267144 135494 267464 142258
rect 267144 135258 267186 135494
rect 267422 135258 267464 135494
rect 267144 128494 267464 135258
rect 267144 128258 267186 128494
rect 267422 128258 267464 128494
rect 267144 121494 267464 128258
rect 267144 121258 267186 121494
rect 267422 121258 267464 121494
rect 267144 114494 267464 121258
rect 267144 114258 267186 114494
rect 267422 114258 267464 114494
rect 267144 107494 267464 114258
rect 267144 107258 267186 107494
rect 267422 107258 267464 107494
rect 267144 100494 267464 107258
rect 267144 100258 267186 100494
rect 267422 100258 267464 100494
rect 267144 93494 267464 100258
rect 267144 93258 267186 93494
rect 267422 93258 267464 93494
rect 267144 86494 267464 93258
rect 267144 86258 267186 86494
rect 267422 86258 267464 86494
rect 267144 79494 267464 86258
rect 267144 79258 267186 79494
rect 267422 79258 267464 79494
rect 267144 72494 267464 79258
rect 267144 72258 267186 72494
rect 267422 72258 267464 72494
rect 267144 65494 267464 72258
rect 267144 65258 267186 65494
rect 267422 65258 267464 65494
rect 267144 58494 267464 65258
rect 267144 58258 267186 58494
rect 267422 58258 267464 58494
rect 267144 51494 267464 58258
rect 267144 51258 267186 51494
rect 267422 51258 267464 51494
rect 267144 44494 267464 51258
rect 267144 44258 267186 44494
rect 267422 44258 267464 44494
rect 267144 37494 267464 44258
rect 267144 37258 267186 37494
rect 267422 37258 267464 37494
rect 267144 30494 267464 37258
rect 267144 30258 267186 30494
rect 267422 30258 267464 30494
rect 267144 23494 267464 30258
rect 267144 23258 267186 23494
rect 267422 23258 267464 23494
rect 267144 16494 267464 23258
rect 267144 16258 267186 16494
rect 267422 16258 267464 16494
rect 267144 9494 267464 16258
rect 267144 9258 267186 9494
rect 267422 9258 267464 9494
rect 267144 2494 267464 9258
rect 267144 2258 267186 2494
rect 267422 2258 267464 2494
rect 267144 -746 267464 2258
rect 267144 -982 267186 -746
rect 267422 -982 267464 -746
rect 267144 -1066 267464 -982
rect 267144 -1302 267186 -1066
rect 267422 -1302 267464 -1066
rect 267144 -2294 267464 -1302
rect 268876 706198 269196 706230
rect 268876 705962 268918 706198
rect 269154 705962 269196 706198
rect 268876 705878 269196 705962
rect 268876 705642 268918 705878
rect 269154 705642 269196 705878
rect 268876 696434 269196 705642
rect 268876 696198 268918 696434
rect 269154 696198 269196 696434
rect 268876 689434 269196 696198
rect 268876 689198 268918 689434
rect 269154 689198 269196 689434
rect 268876 682434 269196 689198
rect 268876 682198 268918 682434
rect 269154 682198 269196 682434
rect 268876 675434 269196 682198
rect 268876 675198 268918 675434
rect 269154 675198 269196 675434
rect 268876 668434 269196 675198
rect 268876 668198 268918 668434
rect 269154 668198 269196 668434
rect 268876 661434 269196 668198
rect 268876 661198 268918 661434
rect 269154 661198 269196 661434
rect 268876 654434 269196 661198
rect 268876 654198 268918 654434
rect 269154 654198 269196 654434
rect 268876 647434 269196 654198
rect 268876 647198 268918 647434
rect 269154 647198 269196 647434
rect 268876 640434 269196 647198
rect 268876 640198 268918 640434
rect 269154 640198 269196 640434
rect 268876 633434 269196 640198
rect 268876 633198 268918 633434
rect 269154 633198 269196 633434
rect 268876 626434 269196 633198
rect 268876 626198 268918 626434
rect 269154 626198 269196 626434
rect 268876 619434 269196 626198
rect 268876 619198 268918 619434
rect 269154 619198 269196 619434
rect 268876 612434 269196 619198
rect 268876 612198 268918 612434
rect 269154 612198 269196 612434
rect 268876 605434 269196 612198
rect 268876 605198 268918 605434
rect 269154 605198 269196 605434
rect 268876 598434 269196 605198
rect 268876 598198 268918 598434
rect 269154 598198 269196 598434
rect 268876 591434 269196 598198
rect 268876 591198 268918 591434
rect 269154 591198 269196 591434
rect 268876 584434 269196 591198
rect 268876 584198 268918 584434
rect 269154 584198 269196 584434
rect 268876 577434 269196 584198
rect 268876 577198 268918 577434
rect 269154 577198 269196 577434
rect 268876 570434 269196 577198
rect 268876 570198 268918 570434
rect 269154 570198 269196 570434
rect 268876 563434 269196 570198
rect 268876 563198 268918 563434
rect 269154 563198 269196 563434
rect 268876 556434 269196 563198
rect 268876 556198 268918 556434
rect 269154 556198 269196 556434
rect 268876 549434 269196 556198
rect 268876 549198 268918 549434
rect 269154 549198 269196 549434
rect 268876 542434 269196 549198
rect 268876 542198 268918 542434
rect 269154 542198 269196 542434
rect 268876 535434 269196 542198
rect 268876 535198 268918 535434
rect 269154 535198 269196 535434
rect 268876 528434 269196 535198
rect 268876 528198 268918 528434
rect 269154 528198 269196 528434
rect 268876 521434 269196 528198
rect 268876 521198 268918 521434
rect 269154 521198 269196 521434
rect 268876 514434 269196 521198
rect 268876 514198 268918 514434
rect 269154 514198 269196 514434
rect 268876 507434 269196 514198
rect 268876 507198 268918 507434
rect 269154 507198 269196 507434
rect 268876 500434 269196 507198
rect 268876 500198 268918 500434
rect 269154 500198 269196 500434
rect 268876 493434 269196 500198
rect 268876 493198 268918 493434
rect 269154 493198 269196 493434
rect 268876 486434 269196 493198
rect 268876 486198 268918 486434
rect 269154 486198 269196 486434
rect 268876 479434 269196 486198
rect 268876 479198 268918 479434
rect 269154 479198 269196 479434
rect 268876 472434 269196 479198
rect 268876 472198 268918 472434
rect 269154 472198 269196 472434
rect 268876 465434 269196 472198
rect 268876 465198 268918 465434
rect 269154 465198 269196 465434
rect 268876 458434 269196 465198
rect 268876 458198 268918 458434
rect 269154 458198 269196 458434
rect 268876 451434 269196 458198
rect 268876 451198 268918 451434
rect 269154 451198 269196 451434
rect 268876 444434 269196 451198
rect 268876 444198 268918 444434
rect 269154 444198 269196 444434
rect 268876 437434 269196 444198
rect 268876 437198 268918 437434
rect 269154 437198 269196 437434
rect 268876 430434 269196 437198
rect 268876 430198 268918 430434
rect 269154 430198 269196 430434
rect 268876 423434 269196 430198
rect 268876 423198 268918 423434
rect 269154 423198 269196 423434
rect 268876 416434 269196 423198
rect 268876 416198 268918 416434
rect 269154 416198 269196 416434
rect 268876 409434 269196 416198
rect 268876 409198 268918 409434
rect 269154 409198 269196 409434
rect 268876 402434 269196 409198
rect 268876 402198 268918 402434
rect 269154 402198 269196 402434
rect 268876 395434 269196 402198
rect 268876 395198 268918 395434
rect 269154 395198 269196 395434
rect 268876 388434 269196 395198
rect 268876 388198 268918 388434
rect 269154 388198 269196 388434
rect 268876 381434 269196 388198
rect 268876 381198 268918 381434
rect 269154 381198 269196 381434
rect 268876 374434 269196 381198
rect 268876 374198 268918 374434
rect 269154 374198 269196 374434
rect 268876 367434 269196 374198
rect 268876 367198 268918 367434
rect 269154 367198 269196 367434
rect 268876 360434 269196 367198
rect 268876 360198 268918 360434
rect 269154 360198 269196 360434
rect 268876 353434 269196 360198
rect 268876 353198 268918 353434
rect 269154 353198 269196 353434
rect 268876 346434 269196 353198
rect 268876 346198 268918 346434
rect 269154 346198 269196 346434
rect 268876 339434 269196 346198
rect 268876 339198 268918 339434
rect 269154 339198 269196 339434
rect 268876 332434 269196 339198
rect 268876 332198 268918 332434
rect 269154 332198 269196 332434
rect 268876 325434 269196 332198
rect 268876 325198 268918 325434
rect 269154 325198 269196 325434
rect 268876 318434 269196 325198
rect 268876 318198 268918 318434
rect 269154 318198 269196 318434
rect 268876 311434 269196 318198
rect 268876 311198 268918 311434
rect 269154 311198 269196 311434
rect 268876 304434 269196 311198
rect 268876 304198 268918 304434
rect 269154 304198 269196 304434
rect 268876 297434 269196 304198
rect 268876 297198 268918 297434
rect 269154 297198 269196 297434
rect 268876 290434 269196 297198
rect 268876 290198 268918 290434
rect 269154 290198 269196 290434
rect 268876 283434 269196 290198
rect 268876 283198 268918 283434
rect 269154 283198 269196 283434
rect 268876 276434 269196 283198
rect 268876 276198 268918 276434
rect 269154 276198 269196 276434
rect 268876 269434 269196 276198
rect 268876 269198 268918 269434
rect 269154 269198 269196 269434
rect 268876 262434 269196 269198
rect 268876 262198 268918 262434
rect 269154 262198 269196 262434
rect 268876 255434 269196 262198
rect 268876 255198 268918 255434
rect 269154 255198 269196 255434
rect 268876 248434 269196 255198
rect 268876 248198 268918 248434
rect 269154 248198 269196 248434
rect 268876 241434 269196 248198
rect 268876 241198 268918 241434
rect 269154 241198 269196 241434
rect 268876 234434 269196 241198
rect 268876 234198 268918 234434
rect 269154 234198 269196 234434
rect 268876 227434 269196 234198
rect 268876 227198 268918 227434
rect 269154 227198 269196 227434
rect 268876 220434 269196 227198
rect 268876 220198 268918 220434
rect 269154 220198 269196 220434
rect 268876 213434 269196 220198
rect 268876 213198 268918 213434
rect 269154 213198 269196 213434
rect 268876 206434 269196 213198
rect 268876 206198 268918 206434
rect 269154 206198 269196 206434
rect 268876 199434 269196 206198
rect 268876 199198 268918 199434
rect 269154 199198 269196 199434
rect 268876 192434 269196 199198
rect 268876 192198 268918 192434
rect 269154 192198 269196 192434
rect 268876 185434 269196 192198
rect 268876 185198 268918 185434
rect 269154 185198 269196 185434
rect 268876 178434 269196 185198
rect 268876 178198 268918 178434
rect 269154 178198 269196 178434
rect 268876 171434 269196 178198
rect 268876 171198 268918 171434
rect 269154 171198 269196 171434
rect 268876 164434 269196 171198
rect 268876 164198 268918 164434
rect 269154 164198 269196 164434
rect 268876 157434 269196 164198
rect 268876 157198 268918 157434
rect 269154 157198 269196 157434
rect 268876 150434 269196 157198
rect 268876 150198 268918 150434
rect 269154 150198 269196 150434
rect 268876 143434 269196 150198
rect 268876 143198 268918 143434
rect 269154 143198 269196 143434
rect 268876 136434 269196 143198
rect 268876 136198 268918 136434
rect 269154 136198 269196 136434
rect 268876 129434 269196 136198
rect 268876 129198 268918 129434
rect 269154 129198 269196 129434
rect 268876 122434 269196 129198
rect 268876 122198 268918 122434
rect 269154 122198 269196 122434
rect 268876 115434 269196 122198
rect 268876 115198 268918 115434
rect 269154 115198 269196 115434
rect 268876 108434 269196 115198
rect 268876 108198 268918 108434
rect 269154 108198 269196 108434
rect 268876 101434 269196 108198
rect 268876 101198 268918 101434
rect 269154 101198 269196 101434
rect 268876 94434 269196 101198
rect 268876 94198 268918 94434
rect 269154 94198 269196 94434
rect 268876 87434 269196 94198
rect 268876 87198 268918 87434
rect 269154 87198 269196 87434
rect 268876 80434 269196 87198
rect 268876 80198 268918 80434
rect 269154 80198 269196 80434
rect 268876 73434 269196 80198
rect 268876 73198 268918 73434
rect 269154 73198 269196 73434
rect 268876 66434 269196 73198
rect 268876 66198 268918 66434
rect 269154 66198 269196 66434
rect 268876 59434 269196 66198
rect 268876 59198 268918 59434
rect 269154 59198 269196 59434
rect 268876 52434 269196 59198
rect 268876 52198 268918 52434
rect 269154 52198 269196 52434
rect 268876 45434 269196 52198
rect 268876 45198 268918 45434
rect 269154 45198 269196 45434
rect 268876 38434 269196 45198
rect 268876 38198 268918 38434
rect 269154 38198 269196 38434
rect 268876 31434 269196 38198
rect 268876 31198 268918 31434
rect 269154 31198 269196 31434
rect 268876 24434 269196 31198
rect 268876 24198 268918 24434
rect 269154 24198 269196 24434
rect 268876 17434 269196 24198
rect 268876 17198 268918 17434
rect 269154 17198 269196 17434
rect 268876 10434 269196 17198
rect 268876 10198 268918 10434
rect 269154 10198 269196 10434
rect 268876 3434 269196 10198
rect 268876 3198 268918 3434
rect 269154 3198 269196 3434
rect 268876 -1706 269196 3198
rect 268876 -1942 268918 -1706
rect 269154 -1942 269196 -1706
rect 268876 -2026 269196 -1942
rect 268876 -2262 268918 -2026
rect 269154 -2262 269196 -2026
rect 268876 -2294 269196 -2262
rect 274144 705238 274464 706230
rect 274144 705002 274186 705238
rect 274422 705002 274464 705238
rect 274144 704918 274464 705002
rect 274144 704682 274186 704918
rect 274422 704682 274464 704918
rect 274144 695494 274464 704682
rect 274144 695258 274186 695494
rect 274422 695258 274464 695494
rect 274144 688494 274464 695258
rect 274144 688258 274186 688494
rect 274422 688258 274464 688494
rect 274144 681494 274464 688258
rect 274144 681258 274186 681494
rect 274422 681258 274464 681494
rect 274144 674494 274464 681258
rect 274144 674258 274186 674494
rect 274422 674258 274464 674494
rect 274144 667494 274464 674258
rect 274144 667258 274186 667494
rect 274422 667258 274464 667494
rect 274144 660494 274464 667258
rect 274144 660258 274186 660494
rect 274422 660258 274464 660494
rect 274144 653494 274464 660258
rect 274144 653258 274186 653494
rect 274422 653258 274464 653494
rect 274144 646494 274464 653258
rect 274144 646258 274186 646494
rect 274422 646258 274464 646494
rect 274144 639494 274464 646258
rect 274144 639258 274186 639494
rect 274422 639258 274464 639494
rect 274144 632494 274464 639258
rect 274144 632258 274186 632494
rect 274422 632258 274464 632494
rect 274144 625494 274464 632258
rect 274144 625258 274186 625494
rect 274422 625258 274464 625494
rect 274144 618494 274464 625258
rect 274144 618258 274186 618494
rect 274422 618258 274464 618494
rect 274144 611494 274464 618258
rect 274144 611258 274186 611494
rect 274422 611258 274464 611494
rect 274144 604494 274464 611258
rect 274144 604258 274186 604494
rect 274422 604258 274464 604494
rect 274144 597494 274464 604258
rect 274144 597258 274186 597494
rect 274422 597258 274464 597494
rect 274144 590494 274464 597258
rect 274144 590258 274186 590494
rect 274422 590258 274464 590494
rect 274144 583494 274464 590258
rect 274144 583258 274186 583494
rect 274422 583258 274464 583494
rect 274144 576494 274464 583258
rect 274144 576258 274186 576494
rect 274422 576258 274464 576494
rect 274144 569494 274464 576258
rect 274144 569258 274186 569494
rect 274422 569258 274464 569494
rect 274144 562494 274464 569258
rect 274144 562258 274186 562494
rect 274422 562258 274464 562494
rect 274144 555494 274464 562258
rect 274144 555258 274186 555494
rect 274422 555258 274464 555494
rect 274144 548494 274464 555258
rect 274144 548258 274186 548494
rect 274422 548258 274464 548494
rect 274144 541494 274464 548258
rect 274144 541258 274186 541494
rect 274422 541258 274464 541494
rect 274144 534494 274464 541258
rect 274144 534258 274186 534494
rect 274422 534258 274464 534494
rect 274144 527494 274464 534258
rect 274144 527258 274186 527494
rect 274422 527258 274464 527494
rect 274144 520494 274464 527258
rect 274144 520258 274186 520494
rect 274422 520258 274464 520494
rect 274144 513494 274464 520258
rect 274144 513258 274186 513494
rect 274422 513258 274464 513494
rect 274144 506494 274464 513258
rect 274144 506258 274186 506494
rect 274422 506258 274464 506494
rect 274144 499494 274464 506258
rect 274144 499258 274186 499494
rect 274422 499258 274464 499494
rect 274144 492494 274464 499258
rect 274144 492258 274186 492494
rect 274422 492258 274464 492494
rect 274144 485494 274464 492258
rect 274144 485258 274186 485494
rect 274422 485258 274464 485494
rect 274144 478494 274464 485258
rect 274144 478258 274186 478494
rect 274422 478258 274464 478494
rect 274144 471494 274464 478258
rect 274144 471258 274186 471494
rect 274422 471258 274464 471494
rect 274144 464494 274464 471258
rect 274144 464258 274186 464494
rect 274422 464258 274464 464494
rect 274144 457494 274464 464258
rect 274144 457258 274186 457494
rect 274422 457258 274464 457494
rect 274144 450494 274464 457258
rect 274144 450258 274186 450494
rect 274422 450258 274464 450494
rect 274144 443494 274464 450258
rect 274144 443258 274186 443494
rect 274422 443258 274464 443494
rect 274144 436494 274464 443258
rect 274144 436258 274186 436494
rect 274422 436258 274464 436494
rect 274144 429494 274464 436258
rect 274144 429258 274186 429494
rect 274422 429258 274464 429494
rect 274144 422494 274464 429258
rect 274144 422258 274186 422494
rect 274422 422258 274464 422494
rect 274144 415494 274464 422258
rect 274144 415258 274186 415494
rect 274422 415258 274464 415494
rect 274144 408494 274464 415258
rect 274144 408258 274186 408494
rect 274422 408258 274464 408494
rect 274144 401494 274464 408258
rect 274144 401258 274186 401494
rect 274422 401258 274464 401494
rect 274144 394494 274464 401258
rect 274144 394258 274186 394494
rect 274422 394258 274464 394494
rect 274144 387494 274464 394258
rect 274144 387258 274186 387494
rect 274422 387258 274464 387494
rect 274144 380494 274464 387258
rect 274144 380258 274186 380494
rect 274422 380258 274464 380494
rect 274144 373494 274464 380258
rect 274144 373258 274186 373494
rect 274422 373258 274464 373494
rect 274144 366494 274464 373258
rect 274144 366258 274186 366494
rect 274422 366258 274464 366494
rect 274144 359494 274464 366258
rect 274144 359258 274186 359494
rect 274422 359258 274464 359494
rect 274144 352494 274464 359258
rect 274144 352258 274186 352494
rect 274422 352258 274464 352494
rect 274144 345494 274464 352258
rect 274144 345258 274186 345494
rect 274422 345258 274464 345494
rect 274144 338494 274464 345258
rect 274144 338258 274186 338494
rect 274422 338258 274464 338494
rect 274144 331494 274464 338258
rect 274144 331258 274186 331494
rect 274422 331258 274464 331494
rect 274144 324494 274464 331258
rect 274144 324258 274186 324494
rect 274422 324258 274464 324494
rect 274144 317494 274464 324258
rect 274144 317258 274186 317494
rect 274422 317258 274464 317494
rect 274144 310494 274464 317258
rect 274144 310258 274186 310494
rect 274422 310258 274464 310494
rect 274144 303494 274464 310258
rect 274144 303258 274186 303494
rect 274422 303258 274464 303494
rect 274144 296494 274464 303258
rect 274144 296258 274186 296494
rect 274422 296258 274464 296494
rect 274144 289494 274464 296258
rect 274144 289258 274186 289494
rect 274422 289258 274464 289494
rect 274144 282494 274464 289258
rect 274144 282258 274186 282494
rect 274422 282258 274464 282494
rect 274144 275494 274464 282258
rect 274144 275258 274186 275494
rect 274422 275258 274464 275494
rect 274144 268494 274464 275258
rect 274144 268258 274186 268494
rect 274422 268258 274464 268494
rect 274144 261494 274464 268258
rect 274144 261258 274186 261494
rect 274422 261258 274464 261494
rect 274144 254494 274464 261258
rect 274144 254258 274186 254494
rect 274422 254258 274464 254494
rect 274144 247494 274464 254258
rect 274144 247258 274186 247494
rect 274422 247258 274464 247494
rect 274144 240494 274464 247258
rect 274144 240258 274186 240494
rect 274422 240258 274464 240494
rect 274144 233494 274464 240258
rect 274144 233258 274186 233494
rect 274422 233258 274464 233494
rect 274144 226494 274464 233258
rect 274144 226258 274186 226494
rect 274422 226258 274464 226494
rect 274144 219494 274464 226258
rect 274144 219258 274186 219494
rect 274422 219258 274464 219494
rect 274144 212494 274464 219258
rect 274144 212258 274186 212494
rect 274422 212258 274464 212494
rect 274144 205494 274464 212258
rect 274144 205258 274186 205494
rect 274422 205258 274464 205494
rect 274144 198494 274464 205258
rect 274144 198258 274186 198494
rect 274422 198258 274464 198494
rect 274144 191494 274464 198258
rect 274144 191258 274186 191494
rect 274422 191258 274464 191494
rect 274144 184494 274464 191258
rect 274144 184258 274186 184494
rect 274422 184258 274464 184494
rect 274144 177494 274464 184258
rect 274144 177258 274186 177494
rect 274422 177258 274464 177494
rect 274144 170494 274464 177258
rect 274144 170258 274186 170494
rect 274422 170258 274464 170494
rect 274144 163494 274464 170258
rect 274144 163258 274186 163494
rect 274422 163258 274464 163494
rect 274144 156494 274464 163258
rect 274144 156258 274186 156494
rect 274422 156258 274464 156494
rect 274144 149494 274464 156258
rect 274144 149258 274186 149494
rect 274422 149258 274464 149494
rect 274144 142494 274464 149258
rect 274144 142258 274186 142494
rect 274422 142258 274464 142494
rect 274144 135494 274464 142258
rect 274144 135258 274186 135494
rect 274422 135258 274464 135494
rect 274144 128494 274464 135258
rect 274144 128258 274186 128494
rect 274422 128258 274464 128494
rect 274144 121494 274464 128258
rect 274144 121258 274186 121494
rect 274422 121258 274464 121494
rect 274144 114494 274464 121258
rect 274144 114258 274186 114494
rect 274422 114258 274464 114494
rect 274144 107494 274464 114258
rect 274144 107258 274186 107494
rect 274422 107258 274464 107494
rect 274144 100494 274464 107258
rect 274144 100258 274186 100494
rect 274422 100258 274464 100494
rect 274144 93494 274464 100258
rect 274144 93258 274186 93494
rect 274422 93258 274464 93494
rect 274144 86494 274464 93258
rect 274144 86258 274186 86494
rect 274422 86258 274464 86494
rect 274144 79494 274464 86258
rect 274144 79258 274186 79494
rect 274422 79258 274464 79494
rect 274144 72494 274464 79258
rect 274144 72258 274186 72494
rect 274422 72258 274464 72494
rect 274144 65494 274464 72258
rect 274144 65258 274186 65494
rect 274422 65258 274464 65494
rect 274144 58494 274464 65258
rect 274144 58258 274186 58494
rect 274422 58258 274464 58494
rect 274144 51494 274464 58258
rect 274144 51258 274186 51494
rect 274422 51258 274464 51494
rect 274144 44494 274464 51258
rect 274144 44258 274186 44494
rect 274422 44258 274464 44494
rect 274144 37494 274464 44258
rect 274144 37258 274186 37494
rect 274422 37258 274464 37494
rect 274144 30494 274464 37258
rect 274144 30258 274186 30494
rect 274422 30258 274464 30494
rect 274144 23494 274464 30258
rect 274144 23258 274186 23494
rect 274422 23258 274464 23494
rect 274144 16494 274464 23258
rect 274144 16258 274186 16494
rect 274422 16258 274464 16494
rect 274144 9494 274464 16258
rect 274144 9258 274186 9494
rect 274422 9258 274464 9494
rect 274144 2494 274464 9258
rect 274144 2258 274186 2494
rect 274422 2258 274464 2494
rect 274144 -746 274464 2258
rect 274144 -982 274186 -746
rect 274422 -982 274464 -746
rect 274144 -1066 274464 -982
rect 274144 -1302 274186 -1066
rect 274422 -1302 274464 -1066
rect 274144 -2294 274464 -1302
rect 275876 706198 276196 706230
rect 275876 705962 275918 706198
rect 276154 705962 276196 706198
rect 275876 705878 276196 705962
rect 275876 705642 275918 705878
rect 276154 705642 276196 705878
rect 275876 696434 276196 705642
rect 275876 696198 275918 696434
rect 276154 696198 276196 696434
rect 275876 689434 276196 696198
rect 275876 689198 275918 689434
rect 276154 689198 276196 689434
rect 275876 682434 276196 689198
rect 275876 682198 275918 682434
rect 276154 682198 276196 682434
rect 275876 675434 276196 682198
rect 275876 675198 275918 675434
rect 276154 675198 276196 675434
rect 275876 668434 276196 675198
rect 275876 668198 275918 668434
rect 276154 668198 276196 668434
rect 275876 661434 276196 668198
rect 275876 661198 275918 661434
rect 276154 661198 276196 661434
rect 275876 654434 276196 661198
rect 275876 654198 275918 654434
rect 276154 654198 276196 654434
rect 275876 647434 276196 654198
rect 275876 647198 275918 647434
rect 276154 647198 276196 647434
rect 275876 640434 276196 647198
rect 275876 640198 275918 640434
rect 276154 640198 276196 640434
rect 275876 633434 276196 640198
rect 275876 633198 275918 633434
rect 276154 633198 276196 633434
rect 275876 626434 276196 633198
rect 275876 626198 275918 626434
rect 276154 626198 276196 626434
rect 275876 619434 276196 626198
rect 275876 619198 275918 619434
rect 276154 619198 276196 619434
rect 275876 612434 276196 619198
rect 275876 612198 275918 612434
rect 276154 612198 276196 612434
rect 275876 605434 276196 612198
rect 275876 605198 275918 605434
rect 276154 605198 276196 605434
rect 275876 598434 276196 605198
rect 275876 598198 275918 598434
rect 276154 598198 276196 598434
rect 275876 591434 276196 598198
rect 275876 591198 275918 591434
rect 276154 591198 276196 591434
rect 275876 584434 276196 591198
rect 275876 584198 275918 584434
rect 276154 584198 276196 584434
rect 275876 577434 276196 584198
rect 275876 577198 275918 577434
rect 276154 577198 276196 577434
rect 275876 570434 276196 577198
rect 275876 570198 275918 570434
rect 276154 570198 276196 570434
rect 275876 563434 276196 570198
rect 275876 563198 275918 563434
rect 276154 563198 276196 563434
rect 275876 556434 276196 563198
rect 275876 556198 275918 556434
rect 276154 556198 276196 556434
rect 275876 549434 276196 556198
rect 275876 549198 275918 549434
rect 276154 549198 276196 549434
rect 275876 542434 276196 549198
rect 275876 542198 275918 542434
rect 276154 542198 276196 542434
rect 275876 535434 276196 542198
rect 275876 535198 275918 535434
rect 276154 535198 276196 535434
rect 275876 528434 276196 535198
rect 275876 528198 275918 528434
rect 276154 528198 276196 528434
rect 275876 521434 276196 528198
rect 275876 521198 275918 521434
rect 276154 521198 276196 521434
rect 275876 514434 276196 521198
rect 275876 514198 275918 514434
rect 276154 514198 276196 514434
rect 275876 507434 276196 514198
rect 275876 507198 275918 507434
rect 276154 507198 276196 507434
rect 275876 500434 276196 507198
rect 275876 500198 275918 500434
rect 276154 500198 276196 500434
rect 275876 493434 276196 500198
rect 275876 493198 275918 493434
rect 276154 493198 276196 493434
rect 275876 486434 276196 493198
rect 275876 486198 275918 486434
rect 276154 486198 276196 486434
rect 275876 479434 276196 486198
rect 275876 479198 275918 479434
rect 276154 479198 276196 479434
rect 275876 472434 276196 479198
rect 275876 472198 275918 472434
rect 276154 472198 276196 472434
rect 275876 465434 276196 472198
rect 275876 465198 275918 465434
rect 276154 465198 276196 465434
rect 275876 458434 276196 465198
rect 275876 458198 275918 458434
rect 276154 458198 276196 458434
rect 275876 451434 276196 458198
rect 275876 451198 275918 451434
rect 276154 451198 276196 451434
rect 275876 444434 276196 451198
rect 275876 444198 275918 444434
rect 276154 444198 276196 444434
rect 275876 437434 276196 444198
rect 275876 437198 275918 437434
rect 276154 437198 276196 437434
rect 275876 430434 276196 437198
rect 275876 430198 275918 430434
rect 276154 430198 276196 430434
rect 275876 423434 276196 430198
rect 275876 423198 275918 423434
rect 276154 423198 276196 423434
rect 275876 416434 276196 423198
rect 275876 416198 275918 416434
rect 276154 416198 276196 416434
rect 275876 409434 276196 416198
rect 275876 409198 275918 409434
rect 276154 409198 276196 409434
rect 275876 402434 276196 409198
rect 275876 402198 275918 402434
rect 276154 402198 276196 402434
rect 275876 395434 276196 402198
rect 275876 395198 275918 395434
rect 276154 395198 276196 395434
rect 275876 388434 276196 395198
rect 275876 388198 275918 388434
rect 276154 388198 276196 388434
rect 275876 381434 276196 388198
rect 275876 381198 275918 381434
rect 276154 381198 276196 381434
rect 275876 374434 276196 381198
rect 275876 374198 275918 374434
rect 276154 374198 276196 374434
rect 275876 367434 276196 374198
rect 275876 367198 275918 367434
rect 276154 367198 276196 367434
rect 275876 360434 276196 367198
rect 275876 360198 275918 360434
rect 276154 360198 276196 360434
rect 275876 353434 276196 360198
rect 275876 353198 275918 353434
rect 276154 353198 276196 353434
rect 275876 346434 276196 353198
rect 275876 346198 275918 346434
rect 276154 346198 276196 346434
rect 275876 339434 276196 346198
rect 275876 339198 275918 339434
rect 276154 339198 276196 339434
rect 275876 332434 276196 339198
rect 275876 332198 275918 332434
rect 276154 332198 276196 332434
rect 275876 325434 276196 332198
rect 275876 325198 275918 325434
rect 276154 325198 276196 325434
rect 275876 318434 276196 325198
rect 275876 318198 275918 318434
rect 276154 318198 276196 318434
rect 275876 311434 276196 318198
rect 275876 311198 275918 311434
rect 276154 311198 276196 311434
rect 275876 304434 276196 311198
rect 275876 304198 275918 304434
rect 276154 304198 276196 304434
rect 275876 297434 276196 304198
rect 275876 297198 275918 297434
rect 276154 297198 276196 297434
rect 275876 290434 276196 297198
rect 275876 290198 275918 290434
rect 276154 290198 276196 290434
rect 275876 283434 276196 290198
rect 275876 283198 275918 283434
rect 276154 283198 276196 283434
rect 275876 276434 276196 283198
rect 275876 276198 275918 276434
rect 276154 276198 276196 276434
rect 275876 269434 276196 276198
rect 275876 269198 275918 269434
rect 276154 269198 276196 269434
rect 275876 262434 276196 269198
rect 275876 262198 275918 262434
rect 276154 262198 276196 262434
rect 275876 255434 276196 262198
rect 275876 255198 275918 255434
rect 276154 255198 276196 255434
rect 275876 248434 276196 255198
rect 275876 248198 275918 248434
rect 276154 248198 276196 248434
rect 275876 241434 276196 248198
rect 275876 241198 275918 241434
rect 276154 241198 276196 241434
rect 275876 234434 276196 241198
rect 275876 234198 275918 234434
rect 276154 234198 276196 234434
rect 275876 227434 276196 234198
rect 275876 227198 275918 227434
rect 276154 227198 276196 227434
rect 275876 220434 276196 227198
rect 275876 220198 275918 220434
rect 276154 220198 276196 220434
rect 275876 213434 276196 220198
rect 275876 213198 275918 213434
rect 276154 213198 276196 213434
rect 275876 206434 276196 213198
rect 275876 206198 275918 206434
rect 276154 206198 276196 206434
rect 275876 199434 276196 206198
rect 275876 199198 275918 199434
rect 276154 199198 276196 199434
rect 275876 192434 276196 199198
rect 275876 192198 275918 192434
rect 276154 192198 276196 192434
rect 275876 185434 276196 192198
rect 275876 185198 275918 185434
rect 276154 185198 276196 185434
rect 275876 178434 276196 185198
rect 275876 178198 275918 178434
rect 276154 178198 276196 178434
rect 275876 171434 276196 178198
rect 275876 171198 275918 171434
rect 276154 171198 276196 171434
rect 275876 164434 276196 171198
rect 275876 164198 275918 164434
rect 276154 164198 276196 164434
rect 275876 157434 276196 164198
rect 275876 157198 275918 157434
rect 276154 157198 276196 157434
rect 275876 150434 276196 157198
rect 275876 150198 275918 150434
rect 276154 150198 276196 150434
rect 275876 143434 276196 150198
rect 275876 143198 275918 143434
rect 276154 143198 276196 143434
rect 275876 136434 276196 143198
rect 275876 136198 275918 136434
rect 276154 136198 276196 136434
rect 275876 129434 276196 136198
rect 275876 129198 275918 129434
rect 276154 129198 276196 129434
rect 275876 122434 276196 129198
rect 275876 122198 275918 122434
rect 276154 122198 276196 122434
rect 275876 115434 276196 122198
rect 275876 115198 275918 115434
rect 276154 115198 276196 115434
rect 275876 108434 276196 115198
rect 275876 108198 275918 108434
rect 276154 108198 276196 108434
rect 275876 101434 276196 108198
rect 275876 101198 275918 101434
rect 276154 101198 276196 101434
rect 275876 94434 276196 101198
rect 275876 94198 275918 94434
rect 276154 94198 276196 94434
rect 275876 87434 276196 94198
rect 275876 87198 275918 87434
rect 276154 87198 276196 87434
rect 275876 80434 276196 87198
rect 275876 80198 275918 80434
rect 276154 80198 276196 80434
rect 275876 73434 276196 80198
rect 275876 73198 275918 73434
rect 276154 73198 276196 73434
rect 275876 66434 276196 73198
rect 275876 66198 275918 66434
rect 276154 66198 276196 66434
rect 275876 59434 276196 66198
rect 275876 59198 275918 59434
rect 276154 59198 276196 59434
rect 275876 52434 276196 59198
rect 275876 52198 275918 52434
rect 276154 52198 276196 52434
rect 275876 45434 276196 52198
rect 275876 45198 275918 45434
rect 276154 45198 276196 45434
rect 275876 38434 276196 45198
rect 275876 38198 275918 38434
rect 276154 38198 276196 38434
rect 275876 31434 276196 38198
rect 275876 31198 275918 31434
rect 276154 31198 276196 31434
rect 275876 24434 276196 31198
rect 275876 24198 275918 24434
rect 276154 24198 276196 24434
rect 275876 17434 276196 24198
rect 275876 17198 275918 17434
rect 276154 17198 276196 17434
rect 275876 10434 276196 17198
rect 275876 10198 275918 10434
rect 276154 10198 276196 10434
rect 275876 3434 276196 10198
rect 275876 3198 275918 3434
rect 276154 3198 276196 3434
rect 275876 -1706 276196 3198
rect 275876 -1942 275918 -1706
rect 276154 -1942 276196 -1706
rect 275876 -2026 276196 -1942
rect 275876 -2262 275918 -2026
rect 276154 -2262 276196 -2026
rect 275876 -2294 276196 -2262
rect 281144 705238 281464 706230
rect 281144 705002 281186 705238
rect 281422 705002 281464 705238
rect 281144 704918 281464 705002
rect 281144 704682 281186 704918
rect 281422 704682 281464 704918
rect 281144 695494 281464 704682
rect 281144 695258 281186 695494
rect 281422 695258 281464 695494
rect 281144 688494 281464 695258
rect 281144 688258 281186 688494
rect 281422 688258 281464 688494
rect 281144 681494 281464 688258
rect 281144 681258 281186 681494
rect 281422 681258 281464 681494
rect 281144 674494 281464 681258
rect 281144 674258 281186 674494
rect 281422 674258 281464 674494
rect 281144 667494 281464 674258
rect 281144 667258 281186 667494
rect 281422 667258 281464 667494
rect 281144 660494 281464 667258
rect 281144 660258 281186 660494
rect 281422 660258 281464 660494
rect 281144 653494 281464 660258
rect 281144 653258 281186 653494
rect 281422 653258 281464 653494
rect 281144 646494 281464 653258
rect 281144 646258 281186 646494
rect 281422 646258 281464 646494
rect 281144 639494 281464 646258
rect 281144 639258 281186 639494
rect 281422 639258 281464 639494
rect 281144 632494 281464 639258
rect 281144 632258 281186 632494
rect 281422 632258 281464 632494
rect 281144 625494 281464 632258
rect 281144 625258 281186 625494
rect 281422 625258 281464 625494
rect 281144 618494 281464 625258
rect 281144 618258 281186 618494
rect 281422 618258 281464 618494
rect 281144 611494 281464 618258
rect 281144 611258 281186 611494
rect 281422 611258 281464 611494
rect 281144 604494 281464 611258
rect 281144 604258 281186 604494
rect 281422 604258 281464 604494
rect 281144 597494 281464 604258
rect 281144 597258 281186 597494
rect 281422 597258 281464 597494
rect 281144 590494 281464 597258
rect 281144 590258 281186 590494
rect 281422 590258 281464 590494
rect 281144 583494 281464 590258
rect 281144 583258 281186 583494
rect 281422 583258 281464 583494
rect 281144 576494 281464 583258
rect 281144 576258 281186 576494
rect 281422 576258 281464 576494
rect 281144 569494 281464 576258
rect 281144 569258 281186 569494
rect 281422 569258 281464 569494
rect 281144 562494 281464 569258
rect 281144 562258 281186 562494
rect 281422 562258 281464 562494
rect 281144 555494 281464 562258
rect 281144 555258 281186 555494
rect 281422 555258 281464 555494
rect 281144 548494 281464 555258
rect 281144 548258 281186 548494
rect 281422 548258 281464 548494
rect 281144 541494 281464 548258
rect 281144 541258 281186 541494
rect 281422 541258 281464 541494
rect 281144 534494 281464 541258
rect 281144 534258 281186 534494
rect 281422 534258 281464 534494
rect 281144 527494 281464 534258
rect 281144 527258 281186 527494
rect 281422 527258 281464 527494
rect 281144 520494 281464 527258
rect 281144 520258 281186 520494
rect 281422 520258 281464 520494
rect 281144 513494 281464 520258
rect 281144 513258 281186 513494
rect 281422 513258 281464 513494
rect 281144 506494 281464 513258
rect 281144 506258 281186 506494
rect 281422 506258 281464 506494
rect 281144 499494 281464 506258
rect 281144 499258 281186 499494
rect 281422 499258 281464 499494
rect 281144 492494 281464 499258
rect 281144 492258 281186 492494
rect 281422 492258 281464 492494
rect 281144 485494 281464 492258
rect 281144 485258 281186 485494
rect 281422 485258 281464 485494
rect 281144 478494 281464 485258
rect 281144 478258 281186 478494
rect 281422 478258 281464 478494
rect 281144 471494 281464 478258
rect 281144 471258 281186 471494
rect 281422 471258 281464 471494
rect 281144 464494 281464 471258
rect 281144 464258 281186 464494
rect 281422 464258 281464 464494
rect 281144 457494 281464 464258
rect 281144 457258 281186 457494
rect 281422 457258 281464 457494
rect 281144 450494 281464 457258
rect 281144 450258 281186 450494
rect 281422 450258 281464 450494
rect 281144 443494 281464 450258
rect 281144 443258 281186 443494
rect 281422 443258 281464 443494
rect 281144 436494 281464 443258
rect 281144 436258 281186 436494
rect 281422 436258 281464 436494
rect 281144 429494 281464 436258
rect 281144 429258 281186 429494
rect 281422 429258 281464 429494
rect 281144 422494 281464 429258
rect 281144 422258 281186 422494
rect 281422 422258 281464 422494
rect 281144 415494 281464 422258
rect 281144 415258 281186 415494
rect 281422 415258 281464 415494
rect 281144 408494 281464 415258
rect 281144 408258 281186 408494
rect 281422 408258 281464 408494
rect 281144 401494 281464 408258
rect 281144 401258 281186 401494
rect 281422 401258 281464 401494
rect 281144 394494 281464 401258
rect 281144 394258 281186 394494
rect 281422 394258 281464 394494
rect 281144 387494 281464 394258
rect 281144 387258 281186 387494
rect 281422 387258 281464 387494
rect 281144 380494 281464 387258
rect 281144 380258 281186 380494
rect 281422 380258 281464 380494
rect 281144 373494 281464 380258
rect 281144 373258 281186 373494
rect 281422 373258 281464 373494
rect 281144 366494 281464 373258
rect 281144 366258 281186 366494
rect 281422 366258 281464 366494
rect 281144 359494 281464 366258
rect 281144 359258 281186 359494
rect 281422 359258 281464 359494
rect 281144 352494 281464 359258
rect 281144 352258 281186 352494
rect 281422 352258 281464 352494
rect 281144 345494 281464 352258
rect 281144 345258 281186 345494
rect 281422 345258 281464 345494
rect 281144 338494 281464 345258
rect 281144 338258 281186 338494
rect 281422 338258 281464 338494
rect 281144 331494 281464 338258
rect 281144 331258 281186 331494
rect 281422 331258 281464 331494
rect 281144 324494 281464 331258
rect 281144 324258 281186 324494
rect 281422 324258 281464 324494
rect 281144 317494 281464 324258
rect 281144 317258 281186 317494
rect 281422 317258 281464 317494
rect 281144 310494 281464 317258
rect 281144 310258 281186 310494
rect 281422 310258 281464 310494
rect 281144 303494 281464 310258
rect 281144 303258 281186 303494
rect 281422 303258 281464 303494
rect 281144 296494 281464 303258
rect 281144 296258 281186 296494
rect 281422 296258 281464 296494
rect 281144 289494 281464 296258
rect 281144 289258 281186 289494
rect 281422 289258 281464 289494
rect 281144 282494 281464 289258
rect 281144 282258 281186 282494
rect 281422 282258 281464 282494
rect 281144 275494 281464 282258
rect 281144 275258 281186 275494
rect 281422 275258 281464 275494
rect 281144 268494 281464 275258
rect 281144 268258 281186 268494
rect 281422 268258 281464 268494
rect 281144 261494 281464 268258
rect 281144 261258 281186 261494
rect 281422 261258 281464 261494
rect 281144 254494 281464 261258
rect 281144 254258 281186 254494
rect 281422 254258 281464 254494
rect 281144 247494 281464 254258
rect 281144 247258 281186 247494
rect 281422 247258 281464 247494
rect 281144 240494 281464 247258
rect 281144 240258 281186 240494
rect 281422 240258 281464 240494
rect 281144 233494 281464 240258
rect 281144 233258 281186 233494
rect 281422 233258 281464 233494
rect 281144 226494 281464 233258
rect 281144 226258 281186 226494
rect 281422 226258 281464 226494
rect 281144 219494 281464 226258
rect 281144 219258 281186 219494
rect 281422 219258 281464 219494
rect 281144 212494 281464 219258
rect 281144 212258 281186 212494
rect 281422 212258 281464 212494
rect 281144 205494 281464 212258
rect 281144 205258 281186 205494
rect 281422 205258 281464 205494
rect 281144 198494 281464 205258
rect 281144 198258 281186 198494
rect 281422 198258 281464 198494
rect 281144 191494 281464 198258
rect 281144 191258 281186 191494
rect 281422 191258 281464 191494
rect 281144 184494 281464 191258
rect 281144 184258 281186 184494
rect 281422 184258 281464 184494
rect 281144 177494 281464 184258
rect 281144 177258 281186 177494
rect 281422 177258 281464 177494
rect 281144 170494 281464 177258
rect 281144 170258 281186 170494
rect 281422 170258 281464 170494
rect 281144 163494 281464 170258
rect 281144 163258 281186 163494
rect 281422 163258 281464 163494
rect 281144 156494 281464 163258
rect 281144 156258 281186 156494
rect 281422 156258 281464 156494
rect 281144 149494 281464 156258
rect 281144 149258 281186 149494
rect 281422 149258 281464 149494
rect 281144 142494 281464 149258
rect 281144 142258 281186 142494
rect 281422 142258 281464 142494
rect 281144 135494 281464 142258
rect 281144 135258 281186 135494
rect 281422 135258 281464 135494
rect 281144 128494 281464 135258
rect 281144 128258 281186 128494
rect 281422 128258 281464 128494
rect 281144 121494 281464 128258
rect 281144 121258 281186 121494
rect 281422 121258 281464 121494
rect 281144 114494 281464 121258
rect 281144 114258 281186 114494
rect 281422 114258 281464 114494
rect 281144 107494 281464 114258
rect 281144 107258 281186 107494
rect 281422 107258 281464 107494
rect 281144 100494 281464 107258
rect 281144 100258 281186 100494
rect 281422 100258 281464 100494
rect 281144 93494 281464 100258
rect 281144 93258 281186 93494
rect 281422 93258 281464 93494
rect 281144 86494 281464 93258
rect 281144 86258 281186 86494
rect 281422 86258 281464 86494
rect 281144 79494 281464 86258
rect 281144 79258 281186 79494
rect 281422 79258 281464 79494
rect 281144 72494 281464 79258
rect 281144 72258 281186 72494
rect 281422 72258 281464 72494
rect 281144 65494 281464 72258
rect 281144 65258 281186 65494
rect 281422 65258 281464 65494
rect 281144 58494 281464 65258
rect 281144 58258 281186 58494
rect 281422 58258 281464 58494
rect 281144 51494 281464 58258
rect 281144 51258 281186 51494
rect 281422 51258 281464 51494
rect 281144 44494 281464 51258
rect 281144 44258 281186 44494
rect 281422 44258 281464 44494
rect 281144 37494 281464 44258
rect 281144 37258 281186 37494
rect 281422 37258 281464 37494
rect 281144 30494 281464 37258
rect 281144 30258 281186 30494
rect 281422 30258 281464 30494
rect 281144 23494 281464 30258
rect 281144 23258 281186 23494
rect 281422 23258 281464 23494
rect 281144 16494 281464 23258
rect 281144 16258 281186 16494
rect 281422 16258 281464 16494
rect 281144 9494 281464 16258
rect 281144 9258 281186 9494
rect 281422 9258 281464 9494
rect 281144 2494 281464 9258
rect 281144 2258 281186 2494
rect 281422 2258 281464 2494
rect 281144 -746 281464 2258
rect 281144 -982 281186 -746
rect 281422 -982 281464 -746
rect 281144 -1066 281464 -982
rect 281144 -1302 281186 -1066
rect 281422 -1302 281464 -1066
rect 281144 -2294 281464 -1302
rect 282876 706198 283196 706230
rect 282876 705962 282918 706198
rect 283154 705962 283196 706198
rect 282876 705878 283196 705962
rect 282876 705642 282918 705878
rect 283154 705642 283196 705878
rect 282876 696434 283196 705642
rect 282876 696198 282918 696434
rect 283154 696198 283196 696434
rect 282876 689434 283196 696198
rect 282876 689198 282918 689434
rect 283154 689198 283196 689434
rect 282876 682434 283196 689198
rect 282876 682198 282918 682434
rect 283154 682198 283196 682434
rect 282876 675434 283196 682198
rect 282876 675198 282918 675434
rect 283154 675198 283196 675434
rect 282876 668434 283196 675198
rect 282876 668198 282918 668434
rect 283154 668198 283196 668434
rect 282876 661434 283196 668198
rect 282876 661198 282918 661434
rect 283154 661198 283196 661434
rect 282876 654434 283196 661198
rect 282876 654198 282918 654434
rect 283154 654198 283196 654434
rect 282876 647434 283196 654198
rect 282876 647198 282918 647434
rect 283154 647198 283196 647434
rect 282876 640434 283196 647198
rect 282876 640198 282918 640434
rect 283154 640198 283196 640434
rect 282876 633434 283196 640198
rect 282876 633198 282918 633434
rect 283154 633198 283196 633434
rect 282876 626434 283196 633198
rect 282876 626198 282918 626434
rect 283154 626198 283196 626434
rect 282876 619434 283196 626198
rect 282876 619198 282918 619434
rect 283154 619198 283196 619434
rect 282876 612434 283196 619198
rect 282876 612198 282918 612434
rect 283154 612198 283196 612434
rect 282876 605434 283196 612198
rect 282876 605198 282918 605434
rect 283154 605198 283196 605434
rect 282876 598434 283196 605198
rect 282876 598198 282918 598434
rect 283154 598198 283196 598434
rect 282876 591434 283196 598198
rect 282876 591198 282918 591434
rect 283154 591198 283196 591434
rect 282876 584434 283196 591198
rect 282876 584198 282918 584434
rect 283154 584198 283196 584434
rect 282876 577434 283196 584198
rect 282876 577198 282918 577434
rect 283154 577198 283196 577434
rect 282876 570434 283196 577198
rect 282876 570198 282918 570434
rect 283154 570198 283196 570434
rect 282876 563434 283196 570198
rect 282876 563198 282918 563434
rect 283154 563198 283196 563434
rect 282876 556434 283196 563198
rect 282876 556198 282918 556434
rect 283154 556198 283196 556434
rect 282876 549434 283196 556198
rect 282876 549198 282918 549434
rect 283154 549198 283196 549434
rect 282876 542434 283196 549198
rect 282876 542198 282918 542434
rect 283154 542198 283196 542434
rect 282876 535434 283196 542198
rect 282876 535198 282918 535434
rect 283154 535198 283196 535434
rect 282876 528434 283196 535198
rect 282876 528198 282918 528434
rect 283154 528198 283196 528434
rect 282876 521434 283196 528198
rect 282876 521198 282918 521434
rect 283154 521198 283196 521434
rect 282876 514434 283196 521198
rect 282876 514198 282918 514434
rect 283154 514198 283196 514434
rect 282876 507434 283196 514198
rect 282876 507198 282918 507434
rect 283154 507198 283196 507434
rect 282876 500434 283196 507198
rect 282876 500198 282918 500434
rect 283154 500198 283196 500434
rect 282876 493434 283196 500198
rect 282876 493198 282918 493434
rect 283154 493198 283196 493434
rect 282876 486434 283196 493198
rect 282876 486198 282918 486434
rect 283154 486198 283196 486434
rect 282876 479434 283196 486198
rect 282876 479198 282918 479434
rect 283154 479198 283196 479434
rect 282876 472434 283196 479198
rect 282876 472198 282918 472434
rect 283154 472198 283196 472434
rect 282876 465434 283196 472198
rect 282876 465198 282918 465434
rect 283154 465198 283196 465434
rect 282876 458434 283196 465198
rect 282876 458198 282918 458434
rect 283154 458198 283196 458434
rect 282876 451434 283196 458198
rect 282876 451198 282918 451434
rect 283154 451198 283196 451434
rect 282876 444434 283196 451198
rect 282876 444198 282918 444434
rect 283154 444198 283196 444434
rect 282876 437434 283196 444198
rect 282876 437198 282918 437434
rect 283154 437198 283196 437434
rect 282876 430434 283196 437198
rect 282876 430198 282918 430434
rect 283154 430198 283196 430434
rect 282876 423434 283196 430198
rect 282876 423198 282918 423434
rect 283154 423198 283196 423434
rect 282876 416434 283196 423198
rect 282876 416198 282918 416434
rect 283154 416198 283196 416434
rect 282876 409434 283196 416198
rect 282876 409198 282918 409434
rect 283154 409198 283196 409434
rect 282876 402434 283196 409198
rect 282876 402198 282918 402434
rect 283154 402198 283196 402434
rect 282876 395434 283196 402198
rect 282876 395198 282918 395434
rect 283154 395198 283196 395434
rect 282876 388434 283196 395198
rect 282876 388198 282918 388434
rect 283154 388198 283196 388434
rect 282876 381434 283196 388198
rect 282876 381198 282918 381434
rect 283154 381198 283196 381434
rect 282876 374434 283196 381198
rect 282876 374198 282918 374434
rect 283154 374198 283196 374434
rect 282876 367434 283196 374198
rect 282876 367198 282918 367434
rect 283154 367198 283196 367434
rect 282876 360434 283196 367198
rect 282876 360198 282918 360434
rect 283154 360198 283196 360434
rect 282876 353434 283196 360198
rect 282876 353198 282918 353434
rect 283154 353198 283196 353434
rect 282876 346434 283196 353198
rect 282876 346198 282918 346434
rect 283154 346198 283196 346434
rect 282876 339434 283196 346198
rect 282876 339198 282918 339434
rect 283154 339198 283196 339434
rect 282876 332434 283196 339198
rect 282876 332198 282918 332434
rect 283154 332198 283196 332434
rect 282876 325434 283196 332198
rect 282876 325198 282918 325434
rect 283154 325198 283196 325434
rect 282876 318434 283196 325198
rect 282876 318198 282918 318434
rect 283154 318198 283196 318434
rect 282876 311434 283196 318198
rect 282876 311198 282918 311434
rect 283154 311198 283196 311434
rect 282876 304434 283196 311198
rect 282876 304198 282918 304434
rect 283154 304198 283196 304434
rect 282876 297434 283196 304198
rect 282876 297198 282918 297434
rect 283154 297198 283196 297434
rect 282876 290434 283196 297198
rect 282876 290198 282918 290434
rect 283154 290198 283196 290434
rect 282876 283434 283196 290198
rect 282876 283198 282918 283434
rect 283154 283198 283196 283434
rect 282876 276434 283196 283198
rect 282876 276198 282918 276434
rect 283154 276198 283196 276434
rect 282876 269434 283196 276198
rect 282876 269198 282918 269434
rect 283154 269198 283196 269434
rect 282876 262434 283196 269198
rect 282876 262198 282918 262434
rect 283154 262198 283196 262434
rect 282876 255434 283196 262198
rect 282876 255198 282918 255434
rect 283154 255198 283196 255434
rect 282876 248434 283196 255198
rect 282876 248198 282918 248434
rect 283154 248198 283196 248434
rect 282876 241434 283196 248198
rect 282876 241198 282918 241434
rect 283154 241198 283196 241434
rect 282876 234434 283196 241198
rect 282876 234198 282918 234434
rect 283154 234198 283196 234434
rect 282876 227434 283196 234198
rect 282876 227198 282918 227434
rect 283154 227198 283196 227434
rect 282876 220434 283196 227198
rect 282876 220198 282918 220434
rect 283154 220198 283196 220434
rect 282876 213434 283196 220198
rect 282876 213198 282918 213434
rect 283154 213198 283196 213434
rect 282876 206434 283196 213198
rect 282876 206198 282918 206434
rect 283154 206198 283196 206434
rect 282876 199434 283196 206198
rect 282876 199198 282918 199434
rect 283154 199198 283196 199434
rect 282876 192434 283196 199198
rect 282876 192198 282918 192434
rect 283154 192198 283196 192434
rect 282876 185434 283196 192198
rect 282876 185198 282918 185434
rect 283154 185198 283196 185434
rect 282876 178434 283196 185198
rect 282876 178198 282918 178434
rect 283154 178198 283196 178434
rect 282876 171434 283196 178198
rect 282876 171198 282918 171434
rect 283154 171198 283196 171434
rect 282876 164434 283196 171198
rect 282876 164198 282918 164434
rect 283154 164198 283196 164434
rect 282876 157434 283196 164198
rect 282876 157198 282918 157434
rect 283154 157198 283196 157434
rect 282876 150434 283196 157198
rect 282876 150198 282918 150434
rect 283154 150198 283196 150434
rect 282876 143434 283196 150198
rect 282876 143198 282918 143434
rect 283154 143198 283196 143434
rect 282876 136434 283196 143198
rect 282876 136198 282918 136434
rect 283154 136198 283196 136434
rect 282876 129434 283196 136198
rect 282876 129198 282918 129434
rect 283154 129198 283196 129434
rect 282876 122434 283196 129198
rect 282876 122198 282918 122434
rect 283154 122198 283196 122434
rect 282876 115434 283196 122198
rect 282876 115198 282918 115434
rect 283154 115198 283196 115434
rect 282876 108434 283196 115198
rect 282876 108198 282918 108434
rect 283154 108198 283196 108434
rect 282876 101434 283196 108198
rect 282876 101198 282918 101434
rect 283154 101198 283196 101434
rect 282876 94434 283196 101198
rect 282876 94198 282918 94434
rect 283154 94198 283196 94434
rect 282876 87434 283196 94198
rect 282876 87198 282918 87434
rect 283154 87198 283196 87434
rect 282876 80434 283196 87198
rect 282876 80198 282918 80434
rect 283154 80198 283196 80434
rect 282876 73434 283196 80198
rect 282876 73198 282918 73434
rect 283154 73198 283196 73434
rect 282876 66434 283196 73198
rect 282876 66198 282918 66434
rect 283154 66198 283196 66434
rect 282876 59434 283196 66198
rect 282876 59198 282918 59434
rect 283154 59198 283196 59434
rect 282876 52434 283196 59198
rect 282876 52198 282918 52434
rect 283154 52198 283196 52434
rect 282876 45434 283196 52198
rect 282876 45198 282918 45434
rect 283154 45198 283196 45434
rect 282876 38434 283196 45198
rect 282876 38198 282918 38434
rect 283154 38198 283196 38434
rect 282876 31434 283196 38198
rect 282876 31198 282918 31434
rect 283154 31198 283196 31434
rect 282876 24434 283196 31198
rect 282876 24198 282918 24434
rect 283154 24198 283196 24434
rect 282876 17434 283196 24198
rect 282876 17198 282918 17434
rect 283154 17198 283196 17434
rect 282876 10434 283196 17198
rect 282876 10198 282918 10434
rect 283154 10198 283196 10434
rect 282876 3434 283196 10198
rect 282876 3198 282918 3434
rect 283154 3198 283196 3434
rect 282876 -1706 283196 3198
rect 282876 -1942 282918 -1706
rect 283154 -1942 283196 -1706
rect 282876 -2026 283196 -1942
rect 282876 -2262 282918 -2026
rect 283154 -2262 283196 -2026
rect 282876 -2294 283196 -2262
rect 288144 705238 288464 706230
rect 288144 705002 288186 705238
rect 288422 705002 288464 705238
rect 288144 704918 288464 705002
rect 288144 704682 288186 704918
rect 288422 704682 288464 704918
rect 288144 695494 288464 704682
rect 288144 695258 288186 695494
rect 288422 695258 288464 695494
rect 288144 688494 288464 695258
rect 288144 688258 288186 688494
rect 288422 688258 288464 688494
rect 288144 681494 288464 688258
rect 288144 681258 288186 681494
rect 288422 681258 288464 681494
rect 288144 674494 288464 681258
rect 288144 674258 288186 674494
rect 288422 674258 288464 674494
rect 288144 667494 288464 674258
rect 288144 667258 288186 667494
rect 288422 667258 288464 667494
rect 288144 660494 288464 667258
rect 288144 660258 288186 660494
rect 288422 660258 288464 660494
rect 288144 653494 288464 660258
rect 288144 653258 288186 653494
rect 288422 653258 288464 653494
rect 288144 646494 288464 653258
rect 288144 646258 288186 646494
rect 288422 646258 288464 646494
rect 288144 639494 288464 646258
rect 288144 639258 288186 639494
rect 288422 639258 288464 639494
rect 288144 632494 288464 639258
rect 288144 632258 288186 632494
rect 288422 632258 288464 632494
rect 288144 625494 288464 632258
rect 288144 625258 288186 625494
rect 288422 625258 288464 625494
rect 288144 618494 288464 625258
rect 288144 618258 288186 618494
rect 288422 618258 288464 618494
rect 288144 611494 288464 618258
rect 288144 611258 288186 611494
rect 288422 611258 288464 611494
rect 288144 604494 288464 611258
rect 288144 604258 288186 604494
rect 288422 604258 288464 604494
rect 288144 597494 288464 604258
rect 288144 597258 288186 597494
rect 288422 597258 288464 597494
rect 288144 590494 288464 597258
rect 288144 590258 288186 590494
rect 288422 590258 288464 590494
rect 288144 583494 288464 590258
rect 288144 583258 288186 583494
rect 288422 583258 288464 583494
rect 288144 576494 288464 583258
rect 288144 576258 288186 576494
rect 288422 576258 288464 576494
rect 288144 569494 288464 576258
rect 288144 569258 288186 569494
rect 288422 569258 288464 569494
rect 288144 562494 288464 569258
rect 288144 562258 288186 562494
rect 288422 562258 288464 562494
rect 288144 555494 288464 562258
rect 288144 555258 288186 555494
rect 288422 555258 288464 555494
rect 288144 548494 288464 555258
rect 288144 548258 288186 548494
rect 288422 548258 288464 548494
rect 288144 541494 288464 548258
rect 288144 541258 288186 541494
rect 288422 541258 288464 541494
rect 288144 534494 288464 541258
rect 288144 534258 288186 534494
rect 288422 534258 288464 534494
rect 288144 527494 288464 534258
rect 288144 527258 288186 527494
rect 288422 527258 288464 527494
rect 288144 520494 288464 527258
rect 288144 520258 288186 520494
rect 288422 520258 288464 520494
rect 288144 513494 288464 520258
rect 288144 513258 288186 513494
rect 288422 513258 288464 513494
rect 288144 506494 288464 513258
rect 288144 506258 288186 506494
rect 288422 506258 288464 506494
rect 288144 499494 288464 506258
rect 288144 499258 288186 499494
rect 288422 499258 288464 499494
rect 288144 492494 288464 499258
rect 288144 492258 288186 492494
rect 288422 492258 288464 492494
rect 288144 485494 288464 492258
rect 288144 485258 288186 485494
rect 288422 485258 288464 485494
rect 288144 478494 288464 485258
rect 288144 478258 288186 478494
rect 288422 478258 288464 478494
rect 288144 471494 288464 478258
rect 288144 471258 288186 471494
rect 288422 471258 288464 471494
rect 288144 464494 288464 471258
rect 288144 464258 288186 464494
rect 288422 464258 288464 464494
rect 288144 457494 288464 464258
rect 288144 457258 288186 457494
rect 288422 457258 288464 457494
rect 288144 450494 288464 457258
rect 288144 450258 288186 450494
rect 288422 450258 288464 450494
rect 288144 443494 288464 450258
rect 288144 443258 288186 443494
rect 288422 443258 288464 443494
rect 288144 436494 288464 443258
rect 288144 436258 288186 436494
rect 288422 436258 288464 436494
rect 288144 429494 288464 436258
rect 288144 429258 288186 429494
rect 288422 429258 288464 429494
rect 288144 422494 288464 429258
rect 288144 422258 288186 422494
rect 288422 422258 288464 422494
rect 288144 415494 288464 422258
rect 288144 415258 288186 415494
rect 288422 415258 288464 415494
rect 288144 408494 288464 415258
rect 288144 408258 288186 408494
rect 288422 408258 288464 408494
rect 288144 401494 288464 408258
rect 288144 401258 288186 401494
rect 288422 401258 288464 401494
rect 288144 394494 288464 401258
rect 288144 394258 288186 394494
rect 288422 394258 288464 394494
rect 288144 387494 288464 394258
rect 288144 387258 288186 387494
rect 288422 387258 288464 387494
rect 288144 380494 288464 387258
rect 288144 380258 288186 380494
rect 288422 380258 288464 380494
rect 288144 373494 288464 380258
rect 288144 373258 288186 373494
rect 288422 373258 288464 373494
rect 288144 366494 288464 373258
rect 288144 366258 288186 366494
rect 288422 366258 288464 366494
rect 288144 359494 288464 366258
rect 288144 359258 288186 359494
rect 288422 359258 288464 359494
rect 288144 352494 288464 359258
rect 288144 352258 288186 352494
rect 288422 352258 288464 352494
rect 288144 345494 288464 352258
rect 288144 345258 288186 345494
rect 288422 345258 288464 345494
rect 288144 338494 288464 345258
rect 288144 338258 288186 338494
rect 288422 338258 288464 338494
rect 288144 331494 288464 338258
rect 288144 331258 288186 331494
rect 288422 331258 288464 331494
rect 288144 324494 288464 331258
rect 288144 324258 288186 324494
rect 288422 324258 288464 324494
rect 288144 317494 288464 324258
rect 288144 317258 288186 317494
rect 288422 317258 288464 317494
rect 288144 310494 288464 317258
rect 288144 310258 288186 310494
rect 288422 310258 288464 310494
rect 288144 303494 288464 310258
rect 288144 303258 288186 303494
rect 288422 303258 288464 303494
rect 288144 296494 288464 303258
rect 288144 296258 288186 296494
rect 288422 296258 288464 296494
rect 288144 289494 288464 296258
rect 288144 289258 288186 289494
rect 288422 289258 288464 289494
rect 288144 282494 288464 289258
rect 288144 282258 288186 282494
rect 288422 282258 288464 282494
rect 288144 275494 288464 282258
rect 288144 275258 288186 275494
rect 288422 275258 288464 275494
rect 288144 268494 288464 275258
rect 288144 268258 288186 268494
rect 288422 268258 288464 268494
rect 288144 261494 288464 268258
rect 288144 261258 288186 261494
rect 288422 261258 288464 261494
rect 288144 254494 288464 261258
rect 288144 254258 288186 254494
rect 288422 254258 288464 254494
rect 288144 247494 288464 254258
rect 288144 247258 288186 247494
rect 288422 247258 288464 247494
rect 288144 240494 288464 247258
rect 288144 240258 288186 240494
rect 288422 240258 288464 240494
rect 288144 233494 288464 240258
rect 288144 233258 288186 233494
rect 288422 233258 288464 233494
rect 288144 226494 288464 233258
rect 288144 226258 288186 226494
rect 288422 226258 288464 226494
rect 288144 219494 288464 226258
rect 288144 219258 288186 219494
rect 288422 219258 288464 219494
rect 288144 212494 288464 219258
rect 288144 212258 288186 212494
rect 288422 212258 288464 212494
rect 288144 205494 288464 212258
rect 288144 205258 288186 205494
rect 288422 205258 288464 205494
rect 288144 198494 288464 205258
rect 288144 198258 288186 198494
rect 288422 198258 288464 198494
rect 288144 191494 288464 198258
rect 288144 191258 288186 191494
rect 288422 191258 288464 191494
rect 288144 184494 288464 191258
rect 288144 184258 288186 184494
rect 288422 184258 288464 184494
rect 288144 177494 288464 184258
rect 288144 177258 288186 177494
rect 288422 177258 288464 177494
rect 288144 170494 288464 177258
rect 288144 170258 288186 170494
rect 288422 170258 288464 170494
rect 288144 163494 288464 170258
rect 288144 163258 288186 163494
rect 288422 163258 288464 163494
rect 288144 156494 288464 163258
rect 288144 156258 288186 156494
rect 288422 156258 288464 156494
rect 288144 149494 288464 156258
rect 288144 149258 288186 149494
rect 288422 149258 288464 149494
rect 288144 142494 288464 149258
rect 288144 142258 288186 142494
rect 288422 142258 288464 142494
rect 288144 135494 288464 142258
rect 288144 135258 288186 135494
rect 288422 135258 288464 135494
rect 288144 128494 288464 135258
rect 288144 128258 288186 128494
rect 288422 128258 288464 128494
rect 288144 121494 288464 128258
rect 288144 121258 288186 121494
rect 288422 121258 288464 121494
rect 288144 114494 288464 121258
rect 288144 114258 288186 114494
rect 288422 114258 288464 114494
rect 288144 107494 288464 114258
rect 288144 107258 288186 107494
rect 288422 107258 288464 107494
rect 288144 100494 288464 107258
rect 288144 100258 288186 100494
rect 288422 100258 288464 100494
rect 288144 93494 288464 100258
rect 288144 93258 288186 93494
rect 288422 93258 288464 93494
rect 288144 86494 288464 93258
rect 288144 86258 288186 86494
rect 288422 86258 288464 86494
rect 288144 79494 288464 86258
rect 288144 79258 288186 79494
rect 288422 79258 288464 79494
rect 288144 72494 288464 79258
rect 288144 72258 288186 72494
rect 288422 72258 288464 72494
rect 288144 65494 288464 72258
rect 288144 65258 288186 65494
rect 288422 65258 288464 65494
rect 288144 58494 288464 65258
rect 288144 58258 288186 58494
rect 288422 58258 288464 58494
rect 288144 51494 288464 58258
rect 288144 51258 288186 51494
rect 288422 51258 288464 51494
rect 288144 44494 288464 51258
rect 288144 44258 288186 44494
rect 288422 44258 288464 44494
rect 288144 37494 288464 44258
rect 288144 37258 288186 37494
rect 288422 37258 288464 37494
rect 288144 30494 288464 37258
rect 288144 30258 288186 30494
rect 288422 30258 288464 30494
rect 288144 23494 288464 30258
rect 288144 23258 288186 23494
rect 288422 23258 288464 23494
rect 288144 16494 288464 23258
rect 288144 16258 288186 16494
rect 288422 16258 288464 16494
rect 288144 9494 288464 16258
rect 288144 9258 288186 9494
rect 288422 9258 288464 9494
rect 288144 2494 288464 9258
rect 288144 2258 288186 2494
rect 288422 2258 288464 2494
rect 288144 -746 288464 2258
rect 288144 -982 288186 -746
rect 288422 -982 288464 -746
rect 288144 -1066 288464 -982
rect 288144 -1302 288186 -1066
rect 288422 -1302 288464 -1066
rect 288144 -2294 288464 -1302
rect 289876 706198 290196 706230
rect 289876 705962 289918 706198
rect 290154 705962 290196 706198
rect 289876 705878 290196 705962
rect 289876 705642 289918 705878
rect 290154 705642 290196 705878
rect 289876 696434 290196 705642
rect 289876 696198 289918 696434
rect 290154 696198 290196 696434
rect 289876 689434 290196 696198
rect 289876 689198 289918 689434
rect 290154 689198 290196 689434
rect 289876 682434 290196 689198
rect 289876 682198 289918 682434
rect 290154 682198 290196 682434
rect 289876 675434 290196 682198
rect 289876 675198 289918 675434
rect 290154 675198 290196 675434
rect 289876 668434 290196 675198
rect 289876 668198 289918 668434
rect 290154 668198 290196 668434
rect 289876 661434 290196 668198
rect 289876 661198 289918 661434
rect 290154 661198 290196 661434
rect 289876 654434 290196 661198
rect 289876 654198 289918 654434
rect 290154 654198 290196 654434
rect 289876 647434 290196 654198
rect 289876 647198 289918 647434
rect 290154 647198 290196 647434
rect 289876 640434 290196 647198
rect 289876 640198 289918 640434
rect 290154 640198 290196 640434
rect 289876 633434 290196 640198
rect 289876 633198 289918 633434
rect 290154 633198 290196 633434
rect 289876 626434 290196 633198
rect 289876 626198 289918 626434
rect 290154 626198 290196 626434
rect 289876 619434 290196 626198
rect 289876 619198 289918 619434
rect 290154 619198 290196 619434
rect 289876 612434 290196 619198
rect 289876 612198 289918 612434
rect 290154 612198 290196 612434
rect 289876 605434 290196 612198
rect 289876 605198 289918 605434
rect 290154 605198 290196 605434
rect 289876 598434 290196 605198
rect 289876 598198 289918 598434
rect 290154 598198 290196 598434
rect 289876 591434 290196 598198
rect 289876 591198 289918 591434
rect 290154 591198 290196 591434
rect 289876 584434 290196 591198
rect 289876 584198 289918 584434
rect 290154 584198 290196 584434
rect 289876 577434 290196 584198
rect 289876 577198 289918 577434
rect 290154 577198 290196 577434
rect 289876 570434 290196 577198
rect 289876 570198 289918 570434
rect 290154 570198 290196 570434
rect 289876 563434 290196 570198
rect 289876 563198 289918 563434
rect 290154 563198 290196 563434
rect 289876 556434 290196 563198
rect 289876 556198 289918 556434
rect 290154 556198 290196 556434
rect 289876 549434 290196 556198
rect 289876 549198 289918 549434
rect 290154 549198 290196 549434
rect 289876 542434 290196 549198
rect 289876 542198 289918 542434
rect 290154 542198 290196 542434
rect 289876 535434 290196 542198
rect 289876 535198 289918 535434
rect 290154 535198 290196 535434
rect 289876 528434 290196 535198
rect 289876 528198 289918 528434
rect 290154 528198 290196 528434
rect 289876 521434 290196 528198
rect 289876 521198 289918 521434
rect 290154 521198 290196 521434
rect 289876 514434 290196 521198
rect 289876 514198 289918 514434
rect 290154 514198 290196 514434
rect 289876 507434 290196 514198
rect 289876 507198 289918 507434
rect 290154 507198 290196 507434
rect 289876 500434 290196 507198
rect 289876 500198 289918 500434
rect 290154 500198 290196 500434
rect 289876 493434 290196 500198
rect 289876 493198 289918 493434
rect 290154 493198 290196 493434
rect 289876 486434 290196 493198
rect 289876 486198 289918 486434
rect 290154 486198 290196 486434
rect 289876 479434 290196 486198
rect 289876 479198 289918 479434
rect 290154 479198 290196 479434
rect 289876 472434 290196 479198
rect 289876 472198 289918 472434
rect 290154 472198 290196 472434
rect 289876 465434 290196 472198
rect 289876 465198 289918 465434
rect 290154 465198 290196 465434
rect 289876 458434 290196 465198
rect 289876 458198 289918 458434
rect 290154 458198 290196 458434
rect 289876 451434 290196 458198
rect 289876 451198 289918 451434
rect 290154 451198 290196 451434
rect 289876 444434 290196 451198
rect 289876 444198 289918 444434
rect 290154 444198 290196 444434
rect 289876 437434 290196 444198
rect 289876 437198 289918 437434
rect 290154 437198 290196 437434
rect 289876 430434 290196 437198
rect 289876 430198 289918 430434
rect 290154 430198 290196 430434
rect 289876 423434 290196 430198
rect 289876 423198 289918 423434
rect 290154 423198 290196 423434
rect 289876 416434 290196 423198
rect 289876 416198 289918 416434
rect 290154 416198 290196 416434
rect 289876 409434 290196 416198
rect 289876 409198 289918 409434
rect 290154 409198 290196 409434
rect 289876 402434 290196 409198
rect 289876 402198 289918 402434
rect 290154 402198 290196 402434
rect 289876 395434 290196 402198
rect 289876 395198 289918 395434
rect 290154 395198 290196 395434
rect 289876 388434 290196 395198
rect 289876 388198 289918 388434
rect 290154 388198 290196 388434
rect 289876 381434 290196 388198
rect 289876 381198 289918 381434
rect 290154 381198 290196 381434
rect 289876 374434 290196 381198
rect 289876 374198 289918 374434
rect 290154 374198 290196 374434
rect 289876 367434 290196 374198
rect 295144 705238 295464 706230
rect 295144 705002 295186 705238
rect 295422 705002 295464 705238
rect 295144 704918 295464 705002
rect 295144 704682 295186 704918
rect 295422 704682 295464 704918
rect 295144 695494 295464 704682
rect 295144 695258 295186 695494
rect 295422 695258 295464 695494
rect 295144 688494 295464 695258
rect 295144 688258 295186 688494
rect 295422 688258 295464 688494
rect 295144 681494 295464 688258
rect 295144 681258 295186 681494
rect 295422 681258 295464 681494
rect 295144 674494 295464 681258
rect 295144 674258 295186 674494
rect 295422 674258 295464 674494
rect 295144 667494 295464 674258
rect 295144 667258 295186 667494
rect 295422 667258 295464 667494
rect 295144 660494 295464 667258
rect 295144 660258 295186 660494
rect 295422 660258 295464 660494
rect 295144 653494 295464 660258
rect 295144 653258 295186 653494
rect 295422 653258 295464 653494
rect 295144 646494 295464 653258
rect 295144 646258 295186 646494
rect 295422 646258 295464 646494
rect 295144 639494 295464 646258
rect 295144 639258 295186 639494
rect 295422 639258 295464 639494
rect 295144 632494 295464 639258
rect 295144 632258 295186 632494
rect 295422 632258 295464 632494
rect 295144 625494 295464 632258
rect 295144 625258 295186 625494
rect 295422 625258 295464 625494
rect 295144 618494 295464 625258
rect 295144 618258 295186 618494
rect 295422 618258 295464 618494
rect 295144 611494 295464 618258
rect 295144 611258 295186 611494
rect 295422 611258 295464 611494
rect 295144 604494 295464 611258
rect 295144 604258 295186 604494
rect 295422 604258 295464 604494
rect 295144 597494 295464 604258
rect 295144 597258 295186 597494
rect 295422 597258 295464 597494
rect 295144 590494 295464 597258
rect 295144 590258 295186 590494
rect 295422 590258 295464 590494
rect 295144 583494 295464 590258
rect 295144 583258 295186 583494
rect 295422 583258 295464 583494
rect 295144 576494 295464 583258
rect 295144 576258 295186 576494
rect 295422 576258 295464 576494
rect 295144 569494 295464 576258
rect 295144 569258 295186 569494
rect 295422 569258 295464 569494
rect 295144 562494 295464 569258
rect 295144 562258 295186 562494
rect 295422 562258 295464 562494
rect 295144 555494 295464 562258
rect 295144 555258 295186 555494
rect 295422 555258 295464 555494
rect 295144 548494 295464 555258
rect 295144 548258 295186 548494
rect 295422 548258 295464 548494
rect 295144 541494 295464 548258
rect 295144 541258 295186 541494
rect 295422 541258 295464 541494
rect 295144 534494 295464 541258
rect 295144 534258 295186 534494
rect 295422 534258 295464 534494
rect 295144 527494 295464 534258
rect 295144 527258 295186 527494
rect 295422 527258 295464 527494
rect 295144 520494 295464 527258
rect 295144 520258 295186 520494
rect 295422 520258 295464 520494
rect 295144 513494 295464 520258
rect 295144 513258 295186 513494
rect 295422 513258 295464 513494
rect 295144 506494 295464 513258
rect 295144 506258 295186 506494
rect 295422 506258 295464 506494
rect 295144 499494 295464 506258
rect 295144 499258 295186 499494
rect 295422 499258 295464 499494
rect 295144 492494 295464 499258
rect 295144 492258 295186 492494
rect 295422 492258 295464 492494
rect 295144 485494 295464 492258
rect 295144 485258 295186 485494
rect 295422 485258 295464 485494
rect 295144 478494 295464 485258
rect 295144 478258 295186 478494
rect 295422 478258 295464 478494
rect 295144 471494 295464 478258
rect 295144 471258 295186 471494
rect 295422 471258 295464 471494
rect 295144 464494 295464 471258
rect 295144 464258 295186 464494
rect 295422 464258 295464 464494
rect 295144 457494 295464 464258
rect 295144 457258 295186 457494
rect 295422 457258 295464 457494
rect 295144 450494 295464 457258
rect 295144 450258 295186 450494
rect 295422 450258 295464 450494
rect 295144 443494 295464 450258
rect 295144 443258 295186 443494
rect 295422 443258 295464 443494
rect 295144 436494 295464 443258
rect 295144 436258 295186 436494
rect 295422 436258 295464 436494
rect 295144 429494 295464 436258
rect 295144 429258 295186 429494
rect 295422 429258 295464 429494
rect 295144 422494 295464 429258
rect 295144 422258 295186 422494
rect 295422 422258 295464 422494
rect 295144 415494 295464 422258
rect 295144 415258 295186 415494
rect 295422 415258 295464 415494
rect 295144 408494 295464 415258
rect 295144 408258 295186 408494
rect 295422 408258 295464 408494
rect 295144 401494 295464 408258
rect 295144 401258 295186 401494
rect 295422 401258 295464 401494
rect 295144 394494 295464 401258
rect 295144 394258 295186 394494
rect 295422 394258 295464 394494
rect 295144 387494 295464 394258
rect 295144 387258 295186 387494
rect 295422 387258 295464 387494
rect 295144 380494 295464 387258
rect 295144 380258 295186 380494
rect 295422 380258 295464 380494
rect 295144 373494 295464 380258
rect 295144 373258 295186 373494
rect 295422 373258 295464 373494
rect 295144 368380 295464 373258
rect 296876 706198 297196 706230
rect 296876 705962 296918 706198
rect 297154 705962 297196 706198
rect 296876 705878 297196 705962
rect 296876 705642 296918 705878
rect 297154 705642 297196 705878
rect 296876 696434 297196 705642
rect 296876 696198 296918 696434
rect 297154 696198 297196 696434
rect 296876 689434 297196 696198
rect 296876 689198 296918 689434
rect 297154 689198 297196 689434
rect 296876 682434 297196 689198
rect 296876 682198 296918 682434
rect 297154 682198 297196 682434
rect 296876 675434 297196 682198
rect 296876 675198 296918 675434
rect 297154 675198 297196 675434
rect 296876 668434 297196 675198
rect 296876 668198 296918 668434
rect 297154 668198 297196 668434
rect 296876 661434 297196 668198
rect 296876 661198 296918 661434
rect 297154 661198 297196 661434
rect 296876 654434 297196 661198
rect 296876 654198 296918 654434
rect 297154 654198 297196 654434
rect 296876 647434 297196 654198
rect 296876 647198 296918 647434
rect 297154 647198 297196 647434
rect 296876 640434 297196 647198
rect 296876 640198 296918 640434
rect 297154 640198 297196 640434
rect 296876 633434 297196 640198
rect 296876 633198 296918 633434
rect 297154 633198 297196 633434
rect 296876 626434 297196 633198
rect 296876 626198 296918 626434
rect 297154 626198 297196 626434
rect 296876 619434 297196 626198
rect 296876 619198 296918 619434
rect 297154 619198 297196 619434
rect 296876 612434 297196 619198
rect 296876 612198 296918 612434
rect 297154 612198 297196 612434
rect 296876 605434 297196 612198
rect 296876 605198 296918 605434
rect 297154 605198 297196 605434
rect 296876 598434 297196 605198
rect 296876 598198 296918 598434
rect 297154 598198 297196 598434
rect 296876 591434 297196 598198
rect 296876 591198 296918 591434
rect 297154 591198 297196 591434
rect 296876 584434 297196 591198
rect 296876 584198 296918 584434
rect 297154 584198 297196 584434
rect 296876 577434 297196 584198
rect 296876 577198 296918 577434
rect 297154 577198 297196 577434
rect 296876 570434 297196 577198
rect 296876 570198 296918 570434
rect 297154 570198 297196 570434
rect 296876 563434 297196 570198
rect 296876 563198 296918 563434
rect 297154 563198 297196 563434
rect 296876 556434 297196 563198
rect 296876 556198 296918 556434
rect 297154 556198 297196 556434
rect 296876 549434 297196 556198
rect 296876 549198 296918 549434
rect 297154 549198 297196 549434
rect 296876 542434 297196 549198
rect 296876 542198 296918 542434
rect 297154 542198 297196 542434
rect 296876 535434 297196 542198
rect 296876 535198 296918 535434
rect 297154 535198 297196 535434
rect 296876 528434 297196 535198
rect 296876 528198 296918 528434
rect 297154 528198 297196 528434
rect 296876 521434 297196 528198
rect 296876 521198 296918 521434
rect 297154 521198 297196 521434
rect 296876 514434 297196 521198
rect 296876 514198 296918 514434
rect 297154 514198 297196 514434
rect 296876 507434 297196 514198
rect 296876 507198 296918 507434
rect 297154 507198 297196 507434
rect 296876 500434 297196 507198
rect 296876 500198 296918 500434
rect 297154 500198 297196 500434
rect 296876 493434 297196 500198
rect 296876 493198 296918 493434
rect 297154 493198 297196 493434
rect 296876 486434 297196 493198
rect 296876 486198 296918 486434
rect 297154 486198 297196 486434
rect 296876 479434 297196 486198
rect 296876 479198 296918 479434
rect 297154 479198 297196 479434
rect 296876 472434 297196 479198
rect 296876 472198 296918 472434
rect 297154 472198 297196 472434
rect 296876 465434 297196 472198
rect 296876 465198 296918 465434
rect 297154 465198 297196 465434
rect 296876 458434 297196 465198
rect 296876 458198 296918 458434
rect 297154 458198 297196 458434
rect 296876 451434 297196 458198
rect 296876 451198 296918 451434
rect 297154 451198 297196 451434
rect 296876 444434 297196 451198
rect 296876 444198 296918 444434
rect 297154 444198 297196 444434
rect 296876 437434 297196 444198
rect 296876 437198 296918 437434
rect 297154 437198 297196 437434
rect 296876 430434 297196 437198
rect 296876 430198 296918 430434
rect 297154 430198 297196 430434
rect 296876 423434 297196 430198
rect 296876 423198 296918 423434
rect 297154 423198 297196 423434
rect 296876 416434 297196 423198
rect 296876 416198 296918 416434
rect 297154 416198 297196 416434
rect 296876 409434 297196 416198
rect 296876 409198 296918 409434
rect 297154 409198 297196 409434
rect 296876 402434 297196 409198
rect 296876 402198 296918 402434
rect 297154 402198 297196 402434
rect 296876 395434 297196 402198
rect 296876 395198 296918 395434
rect 297154 395198 297196 395434
rect 296876 388434 297196 395198
rect 296876 388198 296918 388434
rect 297154 388198 297196 388434
rect 296876 381434 297196 388198
rect 296876 381198 296918 381434
rect 297154 381198 297196 381434
rect 296876 374434 297196 381198
rect 296876 374198 296918 374434
rect 297154 374198 297196 374434
rect 296876 368380 297196 374198
rect 302144 705238 302464 706230
rect 302144 705002 302186 705238
rect 302422 705002 302464 705238
rect 302144 704918 302464 705002
rect 302144 704682 302186 704918
rect 302422 704682 302464 704918
rect 302144 695494 302464 704682
rect 302144 695258 302186 695494
rect 302422 695258 302464 695494
rect 302144 688494 302464 695258
rect 302144 688258 302186 688494
rect 302422 688258 302464 688494
rect 302144 681494 302464 688258
rect 302144 681258 302186 681494
rect 302422 681258 302464 681494
rect 302144 674494 302464 681258
rect 302144 674258 302186 674494
rect 302422 674258 302464 674494
rect 302144 667494 302464 674258
rect 302144 667258 302186 667494
rect 302422 667258 302464 667494
rect 302144 660494 302464 667258
rect 302144 660258 302186 660494
rect 302422 660258 302464 660494
rect 302144 653494 302464 660258
rect 302144 653258 302186 653494
rect 302422 653258 302464 653494
rect 302144 646494 302464 653258
rect 302144 646258 302186 646494
rect 302422 646258 302464 646494
rect 302144 639494 302464 646258
rect 302144 639258 302186 639494
rect 302422 639258 302464 639494
rect 302144 632494 302464 639258
rect 302144 632258 302186 632494
rect 302422 632258 302464 632494
rect 302144 625494 302464 632258
rect 302144 625258 302186 625494
rect 302422 625258 302464 625494
rect 302144 618494 302464 625258
rect 302144 618258 302186 618494
rect 302422 618258 302464 618494
rect 302144 611494 302464 618258
rect 302144 611258 302186 611494
rect 302422 611258 302464 611494
rect 302144 604494 302464 611258
rect 302144 604258 302186 604494
rect 302422 604258 302464 604494
rect 302144 597494 302464 604258
rect 302144 597258 302186 597494
rect 302422 597258 302464 597494
rect 302144 590494 302464 597258
rect 302144 590258 302186 590494
rect 302422 590258 302464 590494
rect 302144 583494 302464 590258
rect 302144 583258 302186 583494
rect 302422 583258 302464 583494
rect 302144 576494 302464 583258
rect 302144 576258 302186 576494
rect 302422 576258 302464 576494
rect 302144 569494 302464 576258
rect 302144 569258 302186 569494
rect 302422 569258 302464 569494
rect 302144 562494 302464 569258
rect 302144 562258 302186 562494
rect 302422 562258 302464 562494
rect 302144 555494 302464 562258
rect 302144 555258 302186 555494
rect 302422 555258 302464 555494
rect 302144 548494 302464 555258
rect 302144 548258 302186 548494
rect 302422 548258 302464 548494
rect 302144 541494 302464 548258
rect 302144 541258 302186 541494
rect 302422 541258 302464 541494
rect 302144 534494 302464 541258
rect 302144 534258 302186 534494
rect 302422 534258 302464 534494
rect 302144 527494 302464 534258
rect 302144 527258 302186 527494
rect 302422 527258 302464 527494
rect 302144 520494 302464 527258
rect 302144 520258 302186 520494
rect 302422 520258 302464 520494
rect 302144 513494 302464 520258
rect 302144 513258 302186 513494
rect 302422 513258 302464 513494
rect 302144 506494 302464 513258
rect 302144 506258 302186 506494
rect 302422 506258 302464 506494
rect 302144 499494 302464 506258
rect 302144 499258 302186 499494
rect 302422 499258 302464 499494
rect 302144 492494 302464 499258
rect 302144 492258 302186 492494
rect 302422 492258 302464 492494
rect 302144 485494 302464 492258
rect 302144 485258 302186 485494
rect 302422 485258 302464 485494
rect 302144 478494 302464 485258
rect 302144 478258 302186 478494
rect 302422 478258 302464 478494
rect 302144 471494 302464 478258
rect 302144 471258 302186 471494
rect 302422 471258 302464 471494
rect 302144 464494 302464 471258
rect 302144 464258 302186 464494
rect 302422 464258 302464 464494
rect 302144 457494 302464 464258
rect 302144 457258 302186 457494
rect 302422 457258 302464 457494
rect 302144 450494 302464 457258
rect 302144 450258 302186 450494
rect 302422 450258 302464 450494
rect 302144 443494 302464 450258
rect 302144 443258 302186 443494
rect 302422 443258 302464 443494
rect 302144 436494 302464 443258
rect 302144 436258 302186 436494
rect 302422 436258 302464 436494
rect 302144 429494 302464 436258
rect 302144 429258 302186 429494
rect 302422 429258 302464 429494
rect 302144 422494 302464 429258
rect 302144 422258 302186 422494
rect 302422 422258 302464 422494
rect 302144 415494 302464 422258
rect 302144 415258 302186 415494
rect 302422 415258 302464 415494
rect 302144 408494 302464 415258
rect 302144 408258 302186 408494
rect 302422 408258 302464 408494
rect 302144 401494 302464 408258
rect 302144 401258 302186 401494
rect 302422 401258 302464 401494
rect 302144 394494 302464 401258
rect 302144 394258 302186 394494
rect 302422 394258 302464 394494
rect 302144 387494 302464 394258
rect 302144 387258 302186 387494
rect 302422 387258 302464 387494
rect 302144 380494 302464 387258
rect 302144 380258 302186 380494
rect 302422 380258 302464 380494
rect 302144 373494 302464 380258
rect 302144 373258 302186 373494
rect 302422 373258 302464 373494
rect 302144 368380 302464 373258
rect 303876 706198 304196 706230
rect 303876 705962 303918 706198
rect 304154 705962 304196 706198
rect 303876 705878 304196 705962
rect 303876 705642 303918 705878
rect 304154 705642 304196 705878
rect 303876 696434 304196 705642
rect 303876 696198 303918 696434
rect 304154 696198 304196 696434
rect 303876 689434 304196 696198
rect 303876 689198 303918 689434
rect 304154 689198 304196 689434
rect 303876 682434 304196 689198
rect 303876 682198 303918 682434
rect 304154 682198 304196 682434
rect 303876 675434 304196 682198
rect 303876 675198 303918 675434
rect 304154 675198 304196 675434
rect 303876 668434 304196 675198
rect 303876 668198 303918 668434
rect 304154 668198 304196 668434
rect 303876 661434 304196 668198
rect 303876 661198 303918 661434
rect 304154 661198 304196 661434
rect 303876 654434 304196 661198
rect 303876 654198 303918 654434
rect 304154 654198 304196 654434
rect 303876 647434 304196 654198
rect 303876 647198 303918 647434
rect 304154 647198 304196 647434
rect 303876 640434 304196 647198
rect 303876 640198 303918 640434
rect 304154 640198 304196 640434
rect 303876 633434 304196 640198
rect 303876 633198 303918 633434
rect 304154 633198 304196 633434
rect 303876 626434 304196 633198
rect 303876 626198 303918 626434
rect 304154 626198 304196 626434
rect 303876 619434 304196 626198
rect 303876 619198 303918 619434
rect 304154 619198 304196 619434
rect 303876 612434 304196 619198
rect 303876 612198 303918 612434
rect 304154 612198 304196 612434
rect 303876 605434 304196 612198
rect 303876 605198 303918 605434
rect 304154 605198 304196 605434
rect 303876 598434 304196 605198
rect 303876 598198 303918 598434
rect 304154 598198 304196 598434
rect 303876 591434 304196 598198
rect 303876 591198 303918 591434
rect 304154 591198 304196 591434
rect 303876 584434 304196 591198
rect 303876 584198 303918 584434
rect 304154 584198 304196 584434
rect 303876 577434 304196 584198
rect 303876 577198 303918 577434
rect 304154 577198 304196 577434
rect 303876 570434 304196 577198
rect 303876 570198 303918 570434
rect 304154 570198 304196 570434
rect 303876 563434 304196 570198
rect 303876 563198 303918 563434
rect 304154 563198 304196 563434
rect 303876 556434 304196 563198
rect 303876 556198 303918 556434
rect 304154 556198 304196 556434
rect 303876 549434 304196 556198
rect 303876 549198 303918 549434
rect 304154 549198 304196 549434
rect 303876 542434 304196 549198
rect 303876 542198 303918 542434
rect 304154 542198 304196 542434
rect 303876 535434 304196 542198
rect 303876 535198 303918 535434
rect 304154 535198 304196 535434
rect 303876 528434 304196 535198
rect 303876 528198 303918 528434
rect 304154 528198 304196 528434
rect 303876 521434 304196 528198
rect 303876 521198 303918 521434
rect 304154 521198 304196 521434
rect 303876 514434 304196 521198
rect 303876 514198 303918 514434
rect 304154 514198 304196 514434
rect 303876 507434 304196 514198
rect 303876 507198 303918 507434
rect 304154 507198 304196 507434
rect 303876 500434 304196 507198
rect 303876 500198 303918 500434
rect 304154 500198 304196 500434
rect 303876 493434 304196 500198
rect 303876 493198 303918 493434
rect 304154 493198 304196 493434
rect 303876 486434 304196 493198
rect 303876 486198 303918 486434
rect 304154 486198 304196 486434
rect 303876 479434 304196 486198
rect 303876 479198 303918 479434
rect 304154 479198 304196 479434
rect 303876 472434 304196 479198
rect 303876 472198 303918 472434
rect 304154 472198 304196 472434
rect 303876 465434 304196 472198
rect 303876 465198 303918 465434
rect 304154 465198 304196 465434
rect 303876 458434 304196 465198
rect 303876 458198 303918 458434
rect 304154 458198 304196 458434
rect 303876 451434 304196 458198
rect 303876 451198 303918 451434
rect 304154 451198 304196 451434
rect 303876 444434 304196 451198
rect 303876 444198 303918 444434
rect 304154 444198 304196 444434
rect 303876 437434 304196 444198
rect 303876 437198 303918 437434
rect 304154 437198 304196 437434
rect 303876 430434 304196 437198
rect 303876 430198 303918 430434
rect 304154 430198 304196 430434
rect 303876 423434 304196 430198
rect 303876 423198 303918 423434
rect 304154 423198 304196 423434
rect 303876 416434 304196 423198
rect 303876 416198 303918 416434
rect 304154 416198 304196 416434
rect 303876 409434 304196 416198
rect 303876 409198 303918 409434
rect 304154 409198 304196 409434
rect 303876 402434 304196 409198
rect 303876 402198 303918 402434
rect 304154 402198 304196 402434
rect 303876 395434 304196 402198
rect 303876 395198 303918 395434
rect 304154 395198 304196 395434
rect 303876 388434 304196 395198
rect 303876 388198 303918 388434
rect 304154 388198 304196 388434
rect 303876 381434 304196 388198
rect 303876 381198 303918 381434
rect 304154 381198 304196 381434
rect 303876 374434 304196 381198
rect 303876 374198 303918 374434
rect 304154 374198 304196 374434
rect 303876 368380 304196 374198
rect 309144 705238 309464 706230
rect 309144 705002 309186 705238
rect 309422 705002 309464 705238
rect 309144 704918 309464 705002
rect 309144 704682 309186 704918
rect 309422 704682 309464 704918
rect 309144 695494 309464 704682
rect 309144 695258 309186 695494
rect 309422 695258 309464 695494
rect 309144 688494 309464 695258
rect 309144 688258 309186 688494
rect 309422 688258 309464 688494
rect 309144 681494 309464 688258
rect 309144 681258 309186 681494
rect 309422 681258 309464 681494
rect 309144 674494 309464 681258
rect 309144 674258 309186 674494
rect 309422 674258 309464 674494
rect 309144 667494 309464 674258
rect 309144 667258 309186 667494
rect 309422 667258 309464 667494
rect 309144 660494 309464 667258
rect 309144 660258 309186 660494
rect 309422 660258 309464 660494
rect 309144 653494 309464 660258
rect 309144 653258 309186 653494
rect 309422 653258 309464 653494
rect 309144 646494 309464 653258
rect 309144 646258 309186 646494
rect 309422 646258 309464 646494
rect 309144 639494 309464 646258
rect 309144 639258 309186 639494
rect 309422 639258 309464 639494
rect 309144 632494 309464 639258
rect 309144 632258 309186 632494
rect 309422 632258 309464 632494
rect 309144 625494 309464 632258
rect 309144 625258 309186 625494
rect 309422 625258 309464 625494
rect 309144 618494 309464 625258
rect 309144 618258 309186 618494
rect 309422 618258 309464 618494
rect 309144 611494 309464 618258
rect 309144 611258 309186 611494
rect 309422 611258 309464 611494
rect 309144 604494 309464 611258
rect 309144 604258 309186 604494
rect 309422 604258 309464 604494
rect 309144 597494 309464 604258
rect 309144 597258 309186 597494
rect 309422 597258 309464 597494
rect 309144 590494 309464 597258
rect 309144 590258 309186 590494
rect 309422 590258 309464 590494
rect 309144 583494 309464 590258
rect 309144 583258 309186 583494
rect 309422 583258 309464 583494
rect 309144 576494 309464 583258
rect 309144 576258 309186 576494
rect 309422 576258 309464 576494
rect 309144 569494 309464 576258
rect 309144 569258 309186 569494
rect 309422 569258 309464 569494
rect 309144 562494 309464 569258
rect 309144 562258 309186 562494
rect 309422 562258 309464 562494
rect 309144 555494 309464 562258
rect 309144 555258 309186 555494
rect 309422 555258 309464 555494
rect 309144 548494 309464 555258
rect 309144 548258 309186 548494
rect 309422 548258 309464 548494
rect 309144 541494 309464 548258
rect 309144 541258 309186 541494
rect 309422 541258 309464 541494
rect 309144 534494 309464 541258
rect 309144 534258 309186 534494
rect 309422 534258 309464 534494
rect 309144 527494 309464 534258
rect 309144 527258 309186 527494
rect 309422 527258 309464 527494
rect 309144 520494 309464 527258
rect 309144 520258 309186 520494
rect 309422 520258 309464 520494
rect 309144 513494 309464 520258
rect 309144 513258 309186 513494
rect 309422 513258 309464 513494
rect 309144 506494 309464 513258
rect 309144 506258 309186 506494
rect 309422 506258 309464 506494
rect 309144 499494 309464 506258
rect 309144 499258 309186 499494
rect 309422 499258 309464 499494
rect 309144 492494 309464 499258
rect 309144 492258 309186 492494
rect 309422 492258 309464 492494
rect 309144 485494 309464 492258
rect 309144 485258 309186 485494
rect 309422 485258 309464 485494
rect 309144 478494 309464 485258
rect 309144 478258 309186 478494
rect 309422 478258 309464 478494
rect 309144 471494 309464 478258
rect 309144 471258 309186 471494
rect 309422 471258 309464 471494
rect 309144 464494 309464 471258
rect 309144 464258 309186 464494
rect 309422 464258 309464 464494
rect 309144 457494 309464 464258
rect 309144 457258 309186 457494
rect 309422 457258 309464 457494
rect 309144 450494 309464 457258
rect 309144 450258 309186 450494
rect 309422 450258 309464 450494
rect 309144 443494 309464 450258
rect 309144 443258 309186 443494
rect 309422 443258 309464 443494
rect 309144 436494 309464 443258
rect 309144 436258 309186 436494
rect 309422 436258 309464 436494
rect 309144 429494 309464 436258
rect 309144 429258 309186 429494
rect 309422 429258 309464 429494
rect 309144 422494 309464 429258
rect 309144 422258 309186 422494
rect 309422 422258 309464 422494
rect 309144 415494 309464 422258
rect 309144 415258 309186 415494
rect 309422 415258 309464 415494
rect 309144 408494 309464 415258
rect 309144 408258 309186 408494
rect 309422 408258 309464 408494
rect 309144 401494 309464 408258
rect 309144 401258 309186 401494
rect 309422 401258 309464 401494
rect 309144 394494 309464 401258
rect 309144 394258 309186 394494
rect 309422 394258 309464 394494
rect 309144 387494 309464 394258
rect 309144 387258 309186 387494
rect 309422 387258 309464 387494
rect 309144 380494 309464 387258
rect 309144 380258 309186 380494
rect 309422 380258 309464 380494
rect 309144 373494 309464 380258
rect 309144 373258 309186 373494
rect 309422 373258 309464 373494
rect 289876 367198 289918 367434
rect 290154 367198 290196 367434
rect 289876 360434 290196 367198
rect 309144 366494 309464 373258
rect 309144 366258 309186 366494
rect 309422 366258 309464 366494
rect 289876 360198 289918 360434
rect 290154 360198 290196 360434
rect 289876 353434 290196 360198
rect 289876 353198 289918 353434
rect 290154 353198 290196 353434
rect 289876 346434 290196 353198
rect 289876 346198 289918 346434
rect 290154 346198 290196 346434
rect 289876 339434 290196 346198
rect 289876 339198 289918 339434
rect 290154 339198 290196 339434
rect 289876 332434 290196 339198
rect 289876 332198 289918 332434
rect 290154 332198 290196 332434
rect 289876 325434 290196 332198
rect 289876 325198 289918 325434
rect 290154 325198 290196 325434
rect 289876 318434 290196 325198
rect 289876 318198 289918 318434
rect 290154 318198 290196 318434
rect 289876 311434 290196 318198
rect 289876 311198 289918 311434
rect 290154 311198 290196 311434
rect 289876 304434 290196 311198
rect 289876 304198 289918 304434
rect 290154 304198 290196 304434
rect 289876 297434 290196 304198
rect 289876 297198 289918 297434
rect 290154 297198 290196 297434
rect 289876 290434 290196 297198
rect 289876 290198 289918 290434
rect 290154 290198 290196 290434
rect 289876 283434 290196 290198
rect 289876 283198 289918 283434
rect 290154 283198 290196 283434
rect 289876 276434 290196 283198
rect 289876 276198 289918 276434
rect 290154 276198 290196 276434
rect 289876 269434 290196 276198
rect 289876 269198 289918 269434
rect 290154 269198 290196 269434
rect 289876 262434 290196 269198
rect 289876 262198 289918 262434
rect 290154 262198 290196 262434
rect 289876 255434 290196 262198
rect 289876 255198 289918 255434
rect 290154 255198 290196 255434
rect 289876 248434 290196 255198
rect 289876 248198 289918 248434
rect 290154 248198 290196 248434
rect 289876 241434 290196 248198
rect 289876 241198 289918 241434
rect 290154 241198 290196 241434
rect 289876 234434 290196 241198
rect 289876 234198 289918 234434
rect 290154 234198 290196 234434
rect 289876 227434 290196 234198
rect 289876 227198 289918 227434
rect 290154 227198 290196 227434
rect 289876 220434 290196 227198
rect 289876 220198 289918 220434
rect 290154 220198 290196 220434
rect 289876 213434 290196 220198
rect 289876 213198 289918 213434
rect 290154 213198 290196 213434
rect 289876 206434 290196 213198
rect 289876 206198 289918 206434
rect 290154 206198 290196 206434
rect 289876 199434 290196 206198
rect 295144 359494 295464 363976
rect 295144 359258 295186 359494
rect 295422 359258 295464 359494
rect 295144 352494 295464 359258
rect 295144 352258 295186 352494
rect 295422 352258 295464 352494
rect 295144 345494 295464 352258
rect 295144 345258 295186 345494
rect 295422 345258 295464 345494
rect 295144 338494 295464 345258
rect 295144 338258 295186 338494
rect 295422 338258 295464 338494
rect 295144 331494 295464 338258
rect 295144 331258 295186 331494
rect 295422 331258 295464 331494
rect 295144 324494 295464 331258
rect 295144 324258 295186 324494
rect 295422 324258 295464 324494
rect 295144 317494 295464 324258
rect 295144 317258 295186 317494
rect 295422 317258 295464 317494
rect 295144 310494 295464 317258
rect 295144 310258 295186 310494
rect 295422 310258 295464 310494
rect 295144 303494 295464 310258
rect 295144 303258 295186 303494
rect 295422 303258 295464 303494
rect 295144 296494 295464 303258
rect 295144 296258 295186 296494
rect 295422 296258 295464 296494
rect 295144 289494 295464 296258
rect 295144 289258 295186 289494
rect 295422 289258 295464 289494
rect 295144 282494 295464 289258
rect 295144 282258 295186 282494
rect 295422 282258 295464 282494
rect 295144 275494 295464 282258
rect 295144 275258 295186 275494
rect 295422 275258 295464 275494
rect 295144 268494 295464 275258
rect 295144 268258 295186 268494
rect 295422 268258 295464 268494
rect 295144 261494 295464 268258
rect 295144 261258 295186 261494
rect 295422 261258 295464 261494
rect 295144 254494 295464 261258
rect 295144 254258 295186 254494
rect 295422 254258 295464 254494
rect 295144 247494 295464 254258
rect 295144 247258 295186 247494
rect 295422 247258 295464 247494
rect 295144 240494 295464 247258
rect 295144 240258 295186 240494
rect 295422 240258 295464 240494
rect 295144 233494 295464 240258
rect 295144 233258 295186 233494
rect 295422 233258 295464 233494
rect 295144 226494 295464 233258
rect 295144 226258 295186 226494
rect 295422 226258 295464 226494
rect 295144 219494 295464 226258
rect 295144 219258 295186 219494
rect 295422 219258 295464 219494
rect 295144 212494 295464 219258
rect 295144 212258 295186 212494
rect 295422 212258 295464 212494
rect 295144 205494 295464 212258
rect 295144 205258 295186 205494
rect 295422 205258 295464 205494
rect 295144 200380 295464 205258
rect 296876 360434 297196 363976
rect 296876 360198 296918 360434
rect 297154 360198 297196 360434
rect 296876 353434 297196 360198
rect 296876 353198 296918 353434
rect 297154 353198 297196 353434
rect 296876 346434 297196 353198
rect 296876 346198 296918 346434
rect 297154 346198 297196 346434
rect 296876 339434 297196 346198
rect 296876 339198 296918 339434
rect 297154 339198 297196 339434
rect 296876 332434 297196 339198
rect 296876 332198 296918 332434
rect 297154 332198 297196 332434
rect 296876 325434 297196 332198
rect 296876 325198 296918 325434
rect 297154 325198 297196 325434
rect 296876 318434 297196 325198
rect 296876 318198 296918 318434
rect 297154 318198 297196 318434
rect 296876 311434 297196 318198
rect 296876 311198 296918 311434
rect 297154 311198 297196 311434
rect 296876 304434 297196 311198
rect 296876 304198 296918 304434
rect 297154 304198 297196 304434
rect 296876 297434 297196 304198
rect 296876 297198 296918 297434
rect 297154 297198 297196 297434
rect 296876 290434 297196 297198
rect 296876 290198 296918 290434
rect 297154 290198 297196 290434
rect 296876 283434 297196 290198
rect 296876 283198 296918 283434
rect 297154 283198 297196 283434
rect 296876 276434 297196 283198
rect 296876 276198 296918 276434
rect 297154 276198 297196 276434
rect 296876 269434 297196 276198
rect 296876 269198 296918 269434
rect 297154 269198 297196 269434
rect 296876 262434 297196 269198
rect 296876 262198 296918 262434
rect 297154 262198 297196 262434
rect 296876 255434 297196 262198
rect 296876 255198 296918 255434
rect 297154 255198 297196 255434
rect 296876 248434 297196 255198
rect 296876 248198 296918 248434
rect 297154 248198 297196 248434
rect 296876 241434 297196 248198
rect 296876 241198 296918 241434
rect 297154 241198 297196 241434
rect 296876 234434 297196 241198
rect 296876 234198 296918 234434
rect 297154 234198 297196 234434
rect 296876 227434 297196 234198
rect 296876 227198 296918 227434
rect 297154 227198 297196 227434
rect 296876 220434 297196 227198
rect 296876 220198 296918 220434
rect 297154 220198 297196 220434
rect 296876 213434 297196 220198
rect 296876 213198 296918 213434
rect 297154 213198 297196 213434
rect 296876 206434 297196 213198
rect 296876 206198 296918 206434
rect 297154 206198 297196 206434
rect 296876 200380 297196 206198
rect 302144 359494 302464 363976
rect 302144 359258 302186 359494
rect 302422 359258 302464 359494
rect 302144 352494 302464 359258
rect 302144 352258 302186 352494
rect 302422 352258 302464 352494
rect 302144 345494 302464 352258
rect 302144 345258 302186 345494
rect 302422 345258 302464 345494
rect 302144 338494 302464 345258
rect 302144 338258 302186 338494
rect 302422 338258 302464 338494
rect 302144 331494 302464 338258
rect 302144 331258 302186 331494
rect 302422 331258 302464 331494
rect 302144 324494 302464 331258
rect 302144 324258 302186 324494
rect 302422 324258 302464 324494
rect 302144 317494 302464 324258
rect 302144 317258 302186 317494
rect 302422 317258 302464 317494
rect 302144 310494 302464 317258
rect 302144 310258 302186 310494
rect 302422 310258 302464 310494
rect 302144 303494 302464 310258
rect 302144 303258 302186 303494
rect 302422 303258 302464 303494
rect 302144 296494 302464 303258
rect 302144 296258 302186 296494
rect 302422 296258 302464 296494
rect 302144 289494 302464 296258
rect 302144 289258 302186 289494
rect 302422 289258 302464 289494
rect 302144 282494 302464 289258
rect 302144 282258 302186 282494
rect 302422 282258 302464 282494
rect 302144 275494 302464 282258
rect 302144 275258 302186 275494
rect 302422 275258 302464 275494
rect 302144 268494 302464 275258
rect 302144 268258 302186 268494
rect 302422 268258 302464 268494
rect 302144 261494 302464 268258
rect 302144 261258 302186 261494
rect 302422 261258 302464 261494
rect 302144 254494 302464 261258
rect 302144 254258 302186 254494
rect 302422 254258 302464 254494
rect 302144 247494 302464 254258
rect 302144 247258 302186 247494
rect 302422 247258 302464 247494
rect 302144 240494 302464 247258
rect 302144 240258 302186 240494
rect 302422 240258 302464 240494
rect 302144 233494 302464 240258
rect 302144 233258 302186 233494
rect 302422 233258 302464 233494
rect 302144 226494 302464 233258
rect 302144 226258 302186 226494
rect 302422 226258 302464 226494
rect 302144 219494 302464 226258
rect 302144 219258 302186 219494
rect 302422 219258 302464 219494
rect 302144 212494 302464 219258
rect 302144 212258 302186 212494
rect 302422 212258 302464 212494
rect 302144 205494 302464 212258
rect 302144 205258 302186 205494
rect 302422 205258 302464 205494
rect 302144 200380 302464 205258
rect 303876 360434 304196 363976
rect 303876 360198 303918 360434
rect 304154 360198 304196 360434
rect 303876 353434 304196 360198
rect 303876 353198 303918 353434
rect 304154 353198 304196 353434
rect 303876 346434 304196 353198
rect 303876 346198 303918 346434
rect 304154 346198 304196 346434
rect 303876 339434 304196 346198
rect 303876 339198 303918 339434
rect 304154 339198 304196 339434
rect 303876 332434 304196 339198
rect 303876 332198 303918 332434
rect 304154 332198 304196 332434
rect 303876 325434 304196 332198
rect 303876 325198 303918 325434
rect 304154 325198 304196 325434
rect 303876 318434 304196 325198
rect 303876 318198 303918 318434
rect 304154 318198 304196 318434
rect 303876 311434 304196 318198
rect 303876 311198 303918 311434
rect 304154 311198 304196 311434
rect 303876 304434 304196 311198
rect 303876 304198 303918 304434
rect 304154 304198 304196 304434
rect 303876 297434 304196 304198
rect 303876 297198 303918 297434
rect 304154 297198 304196 297434
rect 303876 290434 304196 297198
rect 303876 290198 303918 290434
rect 304154 290198 304196 290434
rect 303876 283434 304196 290198
rect 303876 283198 303918 283434
rect 304154 283198 304196 283434
rect 303876 276434 304196 283198
rect 303876 276198 303918 276434
rect 304154 276198 304196 276434
rect 303876 269434 304196 276198
rect 303876 269198 303918 269434
rect 304154 269198 304196 269434
rect 303876 262434 304196 269198
rect 303876 262198 303918 262434
rect 304154 262198 304196 262434
rect 303876 255434 304196 262198
rect 303876 255198 303918 255434
rect 304154 255198 304196 255434
rect 303876 248434 304196 255198
rect 303876 248198 303918 248434
rect 304154 248198 304196 248434
rect 303876 241434 304196 248198
rect 303876 241198 303918 241434
rect 304154 241198 304196 241434
rect 303876 234434 304196 241198
rect 303876 234198 303918 234434
rect 304154 234198 304196 234434
rect 303876 227434 304196 234198
rect 303876 227198 303918 227434
rect 304154 227198 304196 227434
rect 303876 220434 304196 227198
rect 303876 220198 303918 220434
rect 304154 220198 304196 220434
rect 303876 213434 304196 220198
rect 303876 213198 303918 213434
rect 304154 213198 304196 213434
rect 303876 206434 304196 213198
rect 303876 206198 303918 206434
rect 304154 206198 304196 206434
rect 303876 200380 304196 206198
rect 309144 359494 309464 366258
rect 309144 359258 309186 359494
rect 309422 359258 309464 359494
rect 309144 352494 309464 359258
rect 309144 352258 309186 352494
rect 309422 352258 309464 352494
rect 309144 345494 309464 352258
rect 309144 345258 309186 345494
rect 309422 345258 309464 345494
rect 309144 338494 309464 345258
rect 309144 338258 309186 338494
rect 309422 338258 309464 338494
rect 309144 331494 309464 338258
rect 309144 331258 309186 331494
rect 309422 331258 309464 331494
rect 309144 324494 309464 331258
rect 309144 324258 309186 324494
rect 309422 324258 309464 324494
rect 309144 317494 309464 324258
rect 309144 317258 309186 317494
rect 309422 317258 309464 317494
rect 309144 310494 309464 317258
rect 309144 310258 309186 310494
rect 309422 310258 309464 310494
rect 309144 303494 309464 310258
rect 309144 303258 309186 303494
rect 309422 303258 309464 303494
rect 309144 296494 309464 303258
rect 309144 296258 309186 296494
rect 309422 296258 309464 296494
rect 309144 289494 309464 296258
rect 309144 289258 309186 289494
rect 309422 289258 309464 289494
rect 309144 282494 309464 289258
rect 309144 282258 309186 282494
rect 309422 282258 309464 282494
rect 309144 275494 309464 282258
rect 309144 275258 309186 275494
rect 309422 275258 309464 275494
rect 309144 268494 309464 275258
rect 309144 268258 309186 268494
rect 309422 268258 309464 268494
rect 309144 261494 309464 268258
rect 309144 261258 309186 261494
rect 309422 261258 309464 261494
rect 309144 254494 309464 261258
rect 309144 254258 309186 254494
rect 309422 254258 309464 254494
rect 309144 247494 309464 254258
rect 309144 247258 309186 247494
rect 309422 247258 309464 247494
rect 309144 240494 309464 247258
rect 309144 240258 309186 240494
rect 309422 240258 309464 240494
rect 309144 233494 309464 240258
rect 309144 233258 309186 233494
rect 309422 233258 309464 233494
rect 309144 226494 309464 233258
rect 309144 226258 309186 226494
rect 309422 226258 309464 226494
rect 309144 219494 309464 226258
rect 309144 219258 309186 219494
rect 309422 219258 309464 219494
rect 309144 212494 309464 219258
rect 309144 212258 309186 212494
rect 309422 212258 309464 212494
rect 309144 205494 309464 212258
rect 309144 205258 309186 205494
rect 309422 205258 309464 205494
rect 289876 199198 289918 199434
rect 290154 199198 290196 199434
rect 289876 192434 290196 199198
rect 309144 198494 309464 205258
rect 309144 198258 309186 198494
rect 309422 198258 309464 198494
rect 289876 192198 289918 192434
rect 290154 192198 290196 192434
rect 289876 185434 290196 192198
rect 289876 185198 289918 185434
rect 290154 185198 290196 185434
rect 289876 178434 290196 185198
rect 289876 178198 289918 178434
rect 290154 178198 290196 178434
rect 289876 171434 290196 178198
rect 289876 171198 289918 171434
rect 290154 171198 290196 171434
rect 289876 164434 290196 171198
rect 289876 164198 289918 164434
rect 290154 164198 290196 164434
rect 289876 157434 290196 164198
rect 289876 157198 289918 157434
rect 290154 157198 290196 157434
rect 289876 150434 290196 157198
rect 289876 150198 289918 150434
rect 290154 150198 290196 150434
rect 289876 143434 290196 150198
rect 289876 143198 289918 143434
rect 290154 143198 290196 143434
rect 289876 136434 290196 143198
rect 289876 136198 289918 136434
rect 290154 136198 290196 136434
rect 289876 129434 290196 136198
rect 289876 129198 289918 129434
rect 290154 129198 290196 129434
rect 289876 122434 290196 129198
rect 289876 122198 289918 122434
rect 290154 122198 290196 122434
rect 289876 115434 290196 122198
rect 289876 115198 289918 115434
rect 290154 115198 290196 115434
rect 289876 108434 290196 115198
rect 289876 108198 289918 108434
rect 290154 108198 290196 108434
rect 289876 101434 290196 108198
rect 289876 101198 289918 101434
rect 290154 101198 290196 101434
rect 289876 94434 290196 101198
rect 289876 94198 289918 94434
rect 290154 94198 290196 94434
rect 289876 87434 290196 94198
rect 289876 87198 289918 87434
rect 290154 87198 290196 87434
rect 289876 80434 290196 87198
rect 289876 80198 289918 80434
rect 290154 80198 290196 80434
rect 289876 73434 290196 80198
rect 289876 73198 289918 73434
rect 290154 73198 290196 73434
rect 289876 66434 290196 73198
rect 289876 66198 289918 66434
rect 290154 66198 290196 66434
rect 289876 59434 290196 66198
rect 289876 59198 289918 59434
rect 290154 59198 290196 59434
rect 289876 52434 290196 59198
rect 289876 52198 289918 52434
rect 290154 52198 290196 52434
rect 289876 45434 290196 52198
rect 289876 45198 289918 45434
rect 290154 45198 290196 45434
rect 289876 38434 290196 45198
rect 289876 38198 289918 38434
rect 290154 38198 290196 38434
rect 289876 31434 290196 38198
rect 289876 31198 289918 31434
rect 290154 31198 290196 31434
rect 289876 24434 290196 31198
rect 289876 24198 289918 24434
rect 290154 24198 290196 24434
rect 289876 17434 290196 24198
rect 289876 17198 289918 17434
rect 290154 17198 290196 17434
rect 289876 10434 290196 17198
rect 289876 10198 289918 10434
rect 290154 10198 290196 10434
rect 289876 3434 290196 10198
rect 289876 3198 289918 3434
rect 290154 3198 290196 3434
rect 289876 -1706 290196 3198
rect 289876 -1942 289918 -1706
rect 290154 -1942 290196 -1706
rect 289876 -2026 290196 -1942
rect 289876 -2262 289918 -2026
rect 290154 -2262 290196 -2026
rect 289876 -2294 290196 -2262
rect 295144 191494 295464 195976
rect 295144 191258 295186 191494
rect 295422 191258 295464 191494
rect 295144 184494 295464 191258
rect 295144 184258 295186 184494
rect 295422 184258 295464 184494
rect 295144 177494 295464 184258
rect 295144 177258 295186 177494
rect 295422 177258 295464 177494
rect 295144 170494 295464 177258
rect 295144 170258 295186 170494
rect 295422 170258 295464 170494
rect 295144 163494 295464 170258
rect 295144 163258 295186 163494
rect 295422 163258 295464 163494
rect 295144 156494 295464 163258
rect 295144 156258 295186 156494
rect 295422 156258 295464 156494
rect 295144 149494 295464 156258
rect 295144 149258 295186 149494
rect 295422 149258 295464 149494
rect 295144 142494 295464 149258
rect 295144 142258 295186 142494
rect 295422 142258 295464 142494
rect 295144 135494 295464 142258
rect 295144 135258 295186 135494
rect 295422 135258 295464 135494
rect 295144 128494 295464 135258
rect 295144 128258 295186 128494
rect 295422 128258 295464 128494
rect 295144 121494 295464 128258
rect 295144 121258 295186 121494
rect 295422 121258 295464 121494
rect 295144 114494 295464 121258
rect 295144 114258 295186 114494
rect 295422 114258 295464 114494
rect 295144 107494 295464 114258
rect 295144 107258 295186 107494
rect 295422 107258 295464 107494
rect 295144 100494 295464 107258
rect 295144 100258 295186 100494
rect 295422 100258 295464 100494
rect 295144 93494 295464 100258
rect 295144 93258 295186 93494
rect 295422 93258 295464 93494
rect 295144 86494 295464 93258
rect 295144 86258 295186 86494
rect 295422 86258 295464 86494
rect 295144 79494 295464 86258
rect 295144 79258 295186 79494
rect 295422 79258 295464 79494
rect 295144 72494 295464 79258
rect 295144 72258 295186 72494
rect 295422 72258 295464 72494
rect 295144 65494 295464 72258
rect 295144 65258 295186 65494
rect 295422 65258 295464 65494
rect 295144 58494 295464 65258
rect 295144 58258 295186 58494
rect 295422 58258 295464 58494
rect 295144 51494 295464 58258
rect 295144 51258 295186 51494
rect 295422 51258 295464 51494
rect 295144 44494 295464 51258
rect 295144 44258 295186 44494
rect 295422 44258 295464 44494
rect 295144 37494 295464 44258
rect 295144 37258 295186 37494
rect 295422 37258 295464 37494
rect 295144 30494 295464 37258
rect 295144 30258 295186 30494
rect 295422 30258 295464 30494
rect 295144 23494 295464 30258
rect 295144 23258 295186 23494
rect 295422 23258 295464 23494
rect 295144 16494 295464 23258
rect 295144 16258 295186 16494
rect 295422 16258 295464 16494
rect 295144 9494 295464 16258
rect 295144 9258 295186 9494
rect 295422 9258 295464 9494
rect 295144 2494 295464 9258
rect 295144 2258 295186 2494
rect 295422 2258 295464 2494
rect 295144 -746 295464 2258
rect 295144 -982 295186 -746
rect 295422 -982 295464 -746
rect 295144 -1066 295464 -982
rect 295144 -1302 295186 -1066
rect 295422 -1302 295464 -1066
rect 295144 -2294 295464 -1302
rect 296876 192434 297196 195976
rect 296876 192198 296918 192434
rect 297154 192198 297196 192434
rect 296876 185434 297196 192198
rect 296876 185198 296918 185434
rect 297154 185198 297196 185434
rect 296876 178434 297196 185198
rect 296876 178198 296918 178434
rect 297154 178198 297196 178434
rect 296876 171434 297196 178198
rect 296876 171198 296918 171434
rect 297154 171198 297196 171434
rect 296876 164434 297196 171198
rect 296876 164198 296918 164434
rect 297154 164198 297196 164434
rect 296876 157434 297196 164198
rect 296876 157198 296918 157434
rect 297154 157198 297196 157434
rect 296876 150434 297196 157198
rect 296876 150198 296918 150434
rect 297154 150198 297196 150434
rect 296876 143434 297196 150198
rect 296876 143198 296918 143434
rect 297154 143198 297196 143434
rect 296876 136434 297196 143198
rect 296876 136198 296918 136434
rect 297154 136198 297196 136434
rect 296876 129434 297196 136198
rect 296876 129198 296918 129434
rect 297154 129198 297196 129434
rect 296876 122434 297196 129198
rect 296876 122198 296918 122434
rect 297154 122198 297196 122434
rect 296876 115434 297196 122198
rect 296876 115198 296918 115434
rect 297154 115198 297196 115434
rect 296876 108434 297196 115198
rect 296876 108198 296918 108434
rect 297154 108198 297196 108434
rect 296876 101434 297196 108198
rect 296876 101198 296918 101434
rect 297154 101198 297196 101434
rect 296876 94434 297196 101198
rect 296876 94198 296918 94434
rect 297154 94198 297196 94434
rect 296876 87434 297196 94198
rect 296876 87198 296918 87434
rect 297154 87198 297196 87434
rect 296876 80434 297196 87198
rect 296876 80198 296918 80434
rect 297154 80198 297196 80434
rect 296876 73434 297196 80198
rect 296876 73198 296918 73434
rect 297154 73198 297196 73434
rect 296876 66434 297196 73198
rect 296876 66198 296918 66434
rect 297154 66198 297196 66434
rect 296876 59434 297196 66198
rect 296876 59198 296918 59434
rect 297154 59198 297196 59434
rect 296876 52434 297196 59198
rect 296876 52198 296918 52434
rect 297154 52198 297196 52434
rect 296876 45434 297196 52198
rect 296876 45198 296918 45434
rect 297154 45198 297196 45434
rect 296876 38434 297196 45198
rect 296876 38198 296918 38434
rect 297154 38198 297196 38434
rect 296876 31434 297196 38198
rect 296876 31198 296918 31434
rect 297154 31198 297196 31434
rect 296876 24434 297196 31198
rect 296876 24198 296918 24434
rect 297154 24198 297196 24434
rect 296876 17434 297196 24198
rect 296876 17198 296918 17434
rect 297154 17198 297196 17434
rect 296876 10434 297196 17198
rect 296876 10198 296918 10434
rect 297154 10198 297196 10434
rect 296876 3434 297196 10198
rect 296876 3198 296918 3434
rect 297154 3198 297196 3434
rect 296876 -1706 297196 3198
rect 296876 -1942 296918 -1706
rect 297154 -1942 297196 -1706
rect 296876 -2026 297196 -1942
rect 296876 -2262 296918 -2026
rect 297154 -2262 297196 -2026
rect 296876 -2294 297196 -2262
rect 302144 191494 302464 195976
rect 302144 191258 302186 191494
rect 302422 191258 302464 191494
rect 302144 184494 302464 191258
rect 302144 184258 302186 184494
rect 302422 184258 302464 184494
rect 302144 177494 302464 184258
rect 302144 177258 302186 177494
rect 302422 177258 302464 177494
rect 302144 170494 302464 177258
rect 302144 170258 302186 170494
rect 302422 170258 302464 170494
rect 302144 163494 302464 170258
rect 302144 163258 302186 163494
rect 302422 163258 302464 163494
rect 302144 156494 302464 163258
rect 302144 156258 302186 156494
rect 302422 156258 302464 156494
rect 302144 149494 302464 156258
rect 302144 149258 302186 149494
rect 302422 149258 302464 149494
rect 302144 142494 302464 149258
rect 302144 142258 302186 142494
rect 302422 142258 302464 142494
rect 302144 135494 302464 142258
rect 302144 135258 302186 135494
rect 302422 135258 302464 135494
rect 302144 128494 302464 135258
rect 302144 128258 302186 128494
rect 302422 128258 302464 128494
rect 302144 121494 302464 128258
rect 302144 121258 302186 121494
rect 302422 121258 302464 121494
rect 302144 114494 302464 121258
rect 302144 114258 302186 114494
rect 302422 114258 302464 114494
rect 302144 107494 302464 114258
rect 302144 107258 302186 107494
rect 302422 107258 302464 107494
rect 302144 100494 302464 107258
rect 302144 100258 302186 100494
rect 302422 100258 302464 100494
rect 302144 93494 302464 100258
rect 302144 93258 302186 93494
rect 302422 93258 302464 93494
rect 302144 86494 302464 93258
rect 302144 86258 302186 86494
rect 302422 86258 302464 86494
rect 302144 79494 302464 86258
rect 302144 79258 302186 79494
rect 302422 79258 302464 79494
rect 302144 72494 302464 79258
rect 302144 72258 302186 72494
rect 302422 72258 302464 72494
rect 302144 65494 302464 72258
rect 302144 65258 302186 65494
rect 302422 65258 302464 65494
rect 302144 58494 302464 65258
rect 302144 58258 302186 58494
rect 302422 58258 302464 58494
rect 302144 51494 302464 58258
rect 302144 51258 302186 51494
rect 302422 51258 302464 51494
rect 302144 44494 302464 51258
rect 302144 44258 302186 44494
rect 302422 44258 302464 44494
rect 302144 37494 302464 44258
rect 302144 37258 302186 37494
rect 302422 37258 302464 37494
rect 302144 30494 302464 37258
rect 302144 30258 302186 30494
rect 302422 30258 302464 30494
rect 302144 23494 302464 30258
rect 302144 23258 302186 23494
rect 302422 23258 302464 23494
rect 302144 16494 302464 23258
rect 302144 16258 302186 16494
rect 302422 16258 302464 16494
rect 302144 9494 302464 16258
rect 302144 9258 302186 9494
rect 302422 9258 302464 9494
rect 302144 2494 302464 9258
rect 302144 2258 302186 2494
rect 302422 2258 302464 2494
rect 302144 -746 302464 2258
rect 302144 -982 302186 -746
rect 302422 -982 302464 -746
rect 302144 -1066 302464 -982
rect 302144 -1302 302186 -1066
rect 302422 -1302 302464 -1066
rect 302144 -2294 302464 -1302
rect 303876 192434 304196 195976
rect 303876 192198 303918 192434
rect 304154 192198 304196 192434
rect 303876 185434 304196 192198
rect 303876 185198 303918 185434
rect 304154 185198 304196 185434
rect 303876 178434 304196 185198
rect 303876 178198 303918 178434
rect 304154 178198 304196 178434
rect 303876 171434 304196 178198
rect 303876 171198 303918 171434
rect 304154 171198 304196 171434
rect 303876 164434 304196 171198
rect 303876 164198 303918 164434
rect 304154 164198 304196 164434
rect 303876 157434 304196 164198
rect 303876 157198 303918 157434
rect 304154 157198 304196 157434
rect 303876 150434 304196 157198
rect 303876 150198 303918 150434
rect 304154 150198 304196 150434
rect 303876 143434 304196 150198
rect 303876 143198 303918 143434
rect 304154 143198 304196 143434
rect 303876 136434 304196 143198
rect 303876 136198 303918 136434
rect 304154 136198 304196 136434
rect 303876 129434 304196 136198
rect 303876 129198 303918 129434
rect 304154 129198 304196 129434
rect 303876 122434 304196 129198
rect 303876 122198 303918 122434
rect 304154 122198 304196 122434
rect 303876 115434 304196 122198
rect 303876 115198 303918 115434
rect 304154 115198 304196 115434
rect 303876 108434 304196 115198
rect 303876 108198 303918 108434
rect 304154 108198 304196 108434
rect 303876 101434 304196 108198
rect 303876 101198 303918 101434
rect 304154 101198 304196 101434
rect 303876 94434 304196 101198
rect 303876 94198 303918 94434
rect 304154 94198 304196 94434
rect 303876 87434 304196 94198
rect 303876 87198 303918 87434
rect 304154 87198 304196 87434
rect 303876 80434 304196 87198
rect 303876 80198 303918 80434
rect 304154 80198 304196 80434
rect 303876 73434 304196 80198
rect 303876 73198 303918 73434
rect 304154 73198 304196 73434
rect 303876 66434 304196 73198
rect 303876 66198 303918 66434
rect 304154 66198 304196 66434
rect 303876 59434 304196 66198
rect 303876 59198 303918 59434
rect 304154 59198 304196 59434
rect 303876 52434 304196 59198
rect 303876 52198 303918 52434
rect 304154 52198 304196 52434
rect 303876 45434 304196 52198
rect 303876 45198 303918 45434
rect 304154 45198 304196 45434
rect 303876 38434 304196 45198
rect 303876 38198 303918 38434
rect 304154 38198 304196 38434
rect 303876 31434 304196 38198
rect 303876 31198 303918 31434
rect 304154 31198 304196 31434
rect 303876 24434 304196 31198
rect 303876 24198 303918 24434
rect 304154 24198 304196 24434
rect 303876 17434 304196 24198
rect 303876 17198 303918 17434
rect 304154 17198 304196 17434
rect 303876 10434 304196 17198
rect 303876 10198 303918 10434
rect 304154 10198 304196 10434
rect 303876 3434 304196 10198
rect 303876 3198 303918 3434
rect 304154 3198 304196 3434
rect 303876 -1706 304196 3198
rect 303876 -1942 303918 -1706
rect 304154 -1942 304196 -1706
rect 303876 -2026 304196 -1942
rect 303876 -2262 303918 -2026
rect 304154 -2262 304196 -2026
rect 303876 -2294 304196 -2262
rect 309144 191494 309464 198258
rect 309144 191258 309186 191494
rect 309422 191258 309464 191494
rect 309144 184494 309464 191258
rect 309144 184258 309186 184494
rect 309422 184258 309464 184494
rect 309144 177494 309464 184258
rect 309144 177258 309186 177494
rect 309422 177258 309464 177494
rect 309144 170494 309464 177258
rect 309144 170258 309186 170494
rect 309422 170258 309464 170494
rect 309144 163494 309464 170258
rect 309144 163258 309186 163494
rect 309422 163258 309464 163494
rect 309144 156494 309464 163258
rect 309144 156258 309186 156494
rect 309422 156258 309464 156494
rect 309144 149494 309464 156258
rect 309144 149258 309186 149494
rect 309422 149258 309464 149494
rect 309144 142494 309464 149258
rect 309144 142258 309186 142494
rect 309422 142258 309464 142494
rect 309144 135494 309464 142258
rect 309144 135258 309186 135494
rect 309422 135258 309464 135494
rect 309144 128494 309464 135258
rect 309144 128258 309186 128494
rect 309422 128258 309464 128494
rect 309144 121494 309464 128258
rect 309144 121258 309186 121494
rect 309422 121258 309464 121494
rect 309144 114494 309464 121258
rect 309144 114258 309186 114494
rect 309422 114258 309464 114494
rect 309144 107494 309464 114258
rect 309144 107258 309186 107494
rect 309422 107258 309464 107494
rect 309144 100494 309464 107258
rect 309144 100258 309186 100494
rect 309422 100258 309464 100494
rect 309144 93494 309464 100258
rect 309144 93258 309186 93494
rect 309422 93258 309464 93494
rect 309144 86494 309464 93258
rect 309144 86258 309186 86494
rect 309422 86258 309464 86494
rect 309144 79494 309464 86258
rect 309144 79258 309186 79494
rect 309422 79258 309464 79494
rect 309144 72494 309464 79258
rect 309144 72258 309186 72494
rect 309422 72258 309464 72494
rect 309144 65494 309464 72258
rect 309144 65258 309186 65494
rect 309422 65258 309464 65494
rect 309144 58494 309464 65258
rect 309144 58258 309186 58494
rect 309422 58258 309464 58494
rect 309144 51494 309464 58258
rect 309144 51258 309186 51494
rect 309422 51258 309464 51494
rect 309144 44494 309464 51258
rect 309144 44258 309186 44494
rect 309422 44258 309464 44494
rect 309144 37494 309464 44258
rect 309144 37258 309186 37494
rect 309422 37258 309464 37494
rect 309144 30494 309464 37258
rect 309144 30258 309186 30494
rect 309422 30258 309464 30494
rect 309144 23494 309464 30258
rect 309144 23258 309186 23494
rect 309422 23258 309464 23494
rect 309144 16494 309464 23258
rect 309144 16258 309186 16494
rect 309422 16258 309464 16494
rect 309144 9494 309464 16258
rect 309144 9258 309186 9494
rect 309422 9258 309464 9494
rect 309144 2494 309464 9258
rect 309144 2258 309186 2494
rect 309422 2258 309464 2494
rect 309144 -746 309464 2258
rect 309144 -982 309186 -746
rect 309422 -982 309464 -746
rect 309144 -1066 309464 -982
rect 309144 -1302 309186 -1066
rect 309422 -1302 309464 -1066
rect 309144 -2294 309464 -1302
rect 310876 706198 311196 706230
rect 310876 705962 310918 706198
rect 311154 705962 311196 706198
rect 310876 705878 311196 705962
rect 310876 705642 310918 705878
rect 311154 705642 311196 705878
rect 310876 696434 311196 705642
rect 310876 696198 310918 696434
rect 311154 696198 311196 696434
rect 310876 689434 311196 696198
rect 310876 689198 310918 689434
rect 311154 689198 311196 689434
rect 310876 682434 311196 689198
rect 310876 682198 310918 682434
rect 311154 682198 311196 682434
rect 310876 675434 311196 682198
rect 310876 675198 310918 675434
rect 311154 675198 311196 675434
rect 310876 668434 311196 675198
rect 310876 668198 310918 668434
rect 311154 668198 311196 668434
rect 310876 661434 311196 668198
rect 310876 661198 310918 661434
rect 311154 661198 311196 661434
rect 310876 654434 311196 661198
rect 310876 654198 310918 654434
rect 311154 654198 311196 654434
rect 310876 647434 311196 654198
rect 310876 647198 310918 647434
rect 311154 647198 311196 647434
rect 310876 640434 311196 647198
rect 310876 640198 310918 640434
rect 311154 640198 311196 640434
rect 310876 633434 311196 640198
rect 310876 633198 310918 633434
rect 311154 633198 311196 633434
rect 310876 626434 311196 633198
rect 310876 626198 310918 626434
rect 311154 626198 311196 626434
rect 310876 619434 311196 626198
rect 310876 619198 310918 619434
rect 311154 619198 311196 619434
rect 310876 612434 311196 619198
rect 310876 612198 310918 612434
rect 311154 612198 311196 612434
rect 310876 605434 311196 612198
rect 310876 605198 310918 605434
rect 311154 605198 311196 605434
rect 310876 598434 311196 605198
rect 310876 598198 310918 598434
rect 311154 598198 311196 598434
rect 310876 591434 311196 598198
rect 310876 591198 310918 591434
rect 311154 591198 311196 591434
rect 310876 584434 311196 591198
rect 310876 584198 310918 584434
rect 311154 584198 311196 584434
rect 310876 577434 311196 584198
rect 310876 577198 310918 577434
rect 311154 577198 311196 577434
rect 310876 570434 311196 577198
rect 310876 570198 310918 570434
rect 311154 570198 311196 570434
rect 310876 563434 311196 570198
rect 310876 563198 310918 563434
rect 311154 563198 311196 563434
rect 310876 556434 311196 563198
rect 310876 556198 310918 556434
rect 311154 556198 311196 556434
rect 310876 549434 311196 556198
rect 310876 549198 310918 549434
rect 311154 549198 311196 549434
rect 310876 542434 311196 549198
rect 310876 542198 310918 542434
rect 311154 542198 311196 542434
rect 310876 535434 311196 542198
rect 310876 535198 310918 535434
rect 311154 535198 311196 535434
rect 310876 528434 311196 535198
rect 310876 528198 310918 528434
rect 311154 528198 311196 528434
rect 310876 521434 311196 528198
rect 310876 521198 310918 521434
rect 311154 521198 311196 521434
rect 310876 514434 311196 521198
rect 310876 514198 310918 514434
rect 311154 514198 311196 514434
rect 310876 507434 311196 514198
rect 310876 507198 310918 507434
rect 311154 507198 311196 507434
rect 310876 500434 311196 507198
rect 310876 500198 310918 500434
rect 311154 500198 311196 500434
rect 310876 493434 311196 500198
rect 310876 493198 310918 493434
rect 311154 493198 311196 493434
rect 310876 486434 311196 493198
rect 310876 486198 310918 486434
rect 311154 486198 311196 486434
rect 310876 479434 311196 486198
rect 310876 479198 310918 479434
rect 311154 479198 311196 479434
rect 310876 472434 311196 479198
rect 310876 472198 310918 472434
rect 311154 472198 311196 472434
rect 310876 465434 311196 472198
rect 310876 465198 310918 465434
rect 311154 465198 311196 465434
rect 310876 458434 311196 465198
rect 310876 458198 310918 458434
rect 311154 458198 311196 458434
rect 310876 451434 311196 458198
rect 310876 451198 310918 451434
rect 311154 451198 311196 451434
rect 310876 444434 311196 451198
rect 310876 444198 310918 444434
rect 311154 444198 311196 444434
rect 310876 437434 311196 444198
rect 310876 437198 310918 437434
rect 311154 437198 311196 437434
rect 310876 430434 311196 437198
rect 310876 430198 310918 430434
rect 311154 430198 311196 430434
rect 310876 423434 311196 430198
rect 310876 423198 310918 423434
rect 311154 423198 311196 423434
rect 310876 416434 311196 423198
rect 310876 416198 310918 416434
rect 311154 416198 311196 416434
rect 310876 409434 311196 416198
rect 310876 409198 310918 409434
rect 311154 409198 311196 409434
rect 310876 402434 311196 409198
rect 310876 402198 310918 402434
rect 311154 402198 311196 402434
rect 310876 395434 311196 402198
rect 310876 395198 310918 395434
rect 311154 395198 311196 395434
rect 310876 388434 311196 395198
rect 310876 388198 310918 388434
rect 311154 388198 311196 388434
rect 310876 381434 311196 388198
rect 310876 381198 310918 381434
rect 311154 381198 311196 381434
rect 310876 374434 311196 381198
rect 310876 374198 310918 374434
rect 311154 374198 311196 374434
rect 310876 367434 311196 374198
rect 310876 367198 310918 367434
rect 311154 367198 311196 367434
rect 310876 360434 311196 367198
rect 310876 360198 310918 360434
rect 311154 360198 311196 360434
rect 310876 353434 311196 360198
rect 310876 353198 310918 353434
rect 311154 353198 311196 353434
rect 310876 346434 311196 353198
rect 310876 346198 310918 346434
rect 311154 346198 311196 346434
rect 310876 339434 311196 346198
rect 310876 339198 310918 339434
rect 311154 339198 311196 339434
rect 310876 332434 311196 339198
rect 310876 332198 310918 332434
rect 311154 332198 311196 332434
rect 310876 325434 311196 332198
rect 310876 325198 310918 325434
rect 311154 325198 311196 325434
rect 310876 318434 311196 325198
rect 310876 318198 310918 318434
rect 311154 318198 311196 318434
rect 310876 311434 311196 318198
rect 310876 311198 310918 311434
rect 311154 311198 311196 311434
rect 310876 304434 311196 311198
rect 310876 304198 310918 304434
rect 311154 304198 311196 304434
rect 310876 297434 311196 304198
rect 310876 297198 310918 297434
rect 311154 297198 311196 297434
rect 310876 290434 311196 297198
rect 310876 290198 310918 290434
rect 311154 290198 311196 290434
rect 310876 283434 311196 290198
rect 310876 283198 310918 283434
rect 311154 283198 311196 283434
rect 310876 276434 311196 283198
rect 310876 276198 310918 276434
rect 311154 276198 311196 276434
rect 310876 269434 311196 276198
rect 310876 269198 310918 269434
rect 311154 269198 311196 269434
rect 310876 262434 311196 269198
rect 310876 262198 310918 262434
rect 311154 262198 311196 262434
rect 310876 255434 311196 262198
rect 310876 255198 310918 255434
rect 311154 255198 311196 255434
rect 310876 248434 311196 255198
rect 310876 248198 310918 248434
rect 311154 248198 311196 248434
rect 310876 241434 311196 248198
rect 310876 241198 310918 241434
rect 311154 241198 311196 241434
rect 310876 234434 311196 241198
rect 310876 234198 310918 234434
rect 311154 234198 311196 234434
rect 310876 227434 311196 234198
rect 310876 227198 310918 227434
rect 311154 227198 311196 227434
rect 310876 220434 311196 227198
rect 310876 220198 310918 220434
rect 311154 220198 311196 220434
rect 310876 213434 311196 220198
rect 310876 213198 310918 213434
rect 311154 213198 311196 213434
rect 310876 206434 311196 213198
rect 310876 206198 310918 206434
rect 311154 206198 311196 206434
rect 310876 199434 311196 206198
rect 310876 199198 310918 199434
rect 311154 199198 311196 199434
rect 310876 192434 311196 199198
rect 310876 192198 310918 192434
rect 311154 192198 311196 192434
rect 310876 185434 311196 192198
rect 310876 185198 310918 185434
rect 311154 185198 311196 185434
rect 310876 178434 311196 185198
rect 310876 178198 310918 178434
rect 311154 178198 311196 178434
rect 310876 171434 311196 178198
rect 310876 171198 310918 171434
rect 311154 171198 311196 171434
rect 310876 164434 311196 171198
rect 310876 164198 310918 164434
rect 311154 164198 311196 164434
rect 310876 157434 311196 164198
rect 310876 157198 310918 157434
rect 311154 157198 311196 157434
rect 310876 150434 311196 157198
rect 310876 150198 310918 150434
rect 311154 150198 311196 150434
rect 310876 143434 311196 150198
rect 310876 143198 310918 143434
rect 311154 143198 311196 143434
rect 310876 136434 311196 143198
rect 310876 136198 310918 136434
rect 311154 136198 311196 136434
rect 310876 129434 311196 136198
rect 310876 129198 310918 129434
rect 311154 129198 311196 129434
rect 310876 122434 311196 129198
rect 310876 122198 310918 122434
rect 311154 122198 311196 122434
rect 310876 115434 311196 122198
rect 310876 115198 310918 115434
rect 311154 115198 311196 115434
rect 310876 108434 311196 115198
rect 310876 108198 310918 108434
rect 311154 108198 311196 108434
rect 310876 101434 311196 108198
rect 310876 101198 310918 101434
rect 311154 101198 311196 101434
rect 310876 94434 311196 101198
rect 310876 94198 310918 94434
rect 311154 94198 311196 94434
rect 310876 87434 311196 94198
rect 310876 87198 310918 87434
rect 311154 87198 311196 87434
rect 310876 80434 311196 87198
rect 310876 80198 310918 80434
rect 311154 80198 311196 80434
rect 310876 73434 311196 80198
rect 310876 73198 310918 73434
rect 311154 73198 311196 73434
rect 310876 66434 311196 73198
rect 310876 66198 310918 66434
rect 311154 66198 311196 66434
rect 310876 59434 311196 66198
rect 310876 59198 310918 59434
rect 311154 59198 311196 59434
rect 310876 52434 311196 59198
rect 310876 52198 310918 52434
rect 311154 52198 311196 52434
rect 310876 45434 311196 52198
rect 310876 45198 310918 45434
rect 311154 45198 311196 45434
rect 310876 38434 311196 45198
rect 310876 38198 310918 38434
rect 311154 38198 311196 38434
rect 310876 31434 311196 38198
rect 310876 31198 310918 31434
rect 311154 31198 311196 31434
rect 310876 24434 311196 31198
rect 310876 24198 310918 24434
rect 311154 24198 311196 24434
rect 310876 17434 311196 24198
rect 310876 17198 310918 17434
rect 311154 17198 311196 17434
rect 310876 10434 311196 17198
rect 310876 10198 310918 10434
rect 311154 10198 311196 10434
rect 310876 3434 311196 10198
rect 310876 3198 310918 3434
rect 311154 3198 311196 3434
rect 310876 -1706 311196 3198
rect 310876 -1942 310918 -1706
rect 311154 -1942 311196 -1706
rect 310876 -2026 311196 -1942
rect 310876 -2262 310918 -2026
rect 311154 -2262 311196 -2026
rect 310876 -2294 311196 -2262
rect 316144 705238 316464 706230
rect 316144 705002 316186 705238
rect 316422 705002 316464 705238
rect 316144 704918 316464 705002
rect 316144 704682 316186 704918
rect 316422 704682 316464 704918
rect 316144 695494 316464 704682
rect 316144 695258 316186 695494
rect 316422 695258 316464 695494
rect 316144 688494 316464 695258
rect 316144 688258 316186 688494
rect 316422 688258 316464 688494
rect 316144 681494 316464 688258
rect 316144 681258 316186 681494
rect 316422 681258 316464 681494
rect 316144 674494 316464 681258
rect 316144 674258 316186 674494
rect 316422 674258 316464 674494
rect 316144 667494 316464 674258
rect 316144 667258 316186 667494
rect 316422 667258 316464 667494
rect 316144 660494 316464 667258
rect 316144 660258 316186 660494
rect 316422 660258 316464 660494
rect 316144 653494 316464 660258
rect 316144 653258 316186 653494
rect 316422 653258 316464 653494
rect 316144 646494 316464 653258
rect 316144 646258 316186 646494
rect 316422 646258 316464 646494
rect 316144 639494 316464 646258
rect 316144 639258 316186 639494
rect 316422 639258 316464 639494
rect 316144 632494 316464 639258
rect 316144 632258 316186 632494
rect 316422 632258 316464 632494
rect 316144 625494 316464 632258
rect 316144 625258 316186 625494
rect 316422 625258 316464 625494
rect 316144 618494 316464 625258
rect 316144 618258 316186 618494
rect 316422 618258 316464 618494
rect 316144 611494 316464 618258
rect 316144 611258 316186 611494
rect 316422 611258 316464 611494
rect 316144 604494 316464 611258
rect 316144 604258 316186 604494
rect 316422 604258 316464 604494
rect 316144 597494 316464 604258
rect 316144 597258 316186 597494
rect 316422 597258 316464 597494
rect 316144 590494 316464 597258
rect 316144 590258 316186 590494
rect 316422 590258 316464 590494
rect 316144 583494 316464 590258
rect 316144 583258 316186 583494
rect 316422 583258 316464 583494
rect 316144 576494 316464 583258
rect 316144 576258 316186 576494
rect 316422 576258 316464 576494
rect 316144 569494 316464 576258
rect 316144 569258 316186 569494
rect 316422 569258 316464 569494
rect 316144 562494 316464 569258
rect 316144 562258 316186 562494
rect 316422 562258 316464 562494
rect 316144 555494 316464 562258
rect 316144 555258 316186 555494
rect 316422 555258 316464 555494
rect 316144 548494 316464 555258
rect 316144 548258 316186 548494
rect 316422 548258 316464 548494
rect 316144 541494 316464 548258
rect 316144 541258 316186 541494
rect 316422 541258 316464 541494
rect 316144 534494 316464 541258
rect 316144 534258 316186 534494
rect 316422 534258 316464 534494
rect 316144 527494 316464 534258
rect 316144 527258 316186 527494
rect 316422 527258 316464 527494
rect 316144 520494 316464 527258
rect 316144 520258 316186 520494
rect 316422 520258 316464 520494
rect 316144 513494 316464 520258
rect 316144 513258 316186 513494
rect 316422 513258 316464 513494
rect 316144 506494 316464 513258
rect 316144 506258 316186 506494
rect 316422 506258 316464 506494
rect 316144 499494 316464 506258
rect 316144 499258 316186 499494
rect 316422 499258 316464 499494
rect 316144 492494 316464 499258
rect 316144 492258 316186 492494
rect 316422 492258 316464 492494
rect 316144 485494 316464 492258
rect 316144 485258 316186 485494
rect 316422 485258 316464 485494
rect 316144 478494 316464 485258
rect 316144 478258 316186 478494
rect 316422 478258 316464 478494
rect 316144 471494 316464 478258
rect 316144 471258 316186 471494
rect 316422 471258 316464 471494
rect 316144 464494 316464 471258
rect 316144 464258 316186 464494
rect 316422 464258 316464 464494
rect 316144 457494 316464 464258
rect 316144 457258 316186 457494
rect 316422 457258 316464 457494
rect 316144 450494 316464 457258
rect 316144 450258 316186 450494
rect 316422 450258 316464 450494
rect 316144 443494 316464 450258
rect 316144 443258 316186 443494
rect 316422 443258 316464 443494
rect 316144 436494 316464 443258
rect 316144 436258 316186 436494
rect 316422 436258 316464 436494
rect 316144 429494 316464 436258
rect 316144 429258 316186 429494
rect 316422 429258 316464 429494
rect 316144 422494 316464 429258
rect 316144 422258 316186 422494
rect 316422 422258 316464 422494
rect 316144 415494 316464 422258
rect 316144 415258 316186 415494
rect 316422 415258 316464 415494
rect 316144 408494 316464 415258
rect 316144 408258 316186 408494
rect 316422 408258 316464 408494
rect 316144 401494 316464 408258
rect 316144 401258 316186 401494
rect 316422 401258 316464 401494
rect 316144 394494 316464 401258
rect 316144 394258 316186 394494
rect 316422 394258 316464 394494
rect 316144 387494 316464 394258
rect 316144 387258 316186 387494
rect 316422 387258 316464 387494
rect 316144 380494 316464 387258
rect 316144 380258 316186 380494
rect 316422 380258 316464 380494
rect 316144 373494 316464 380258
rect 316144 373258 316186 373494
rect 316422 373258 316464 373494
rect 316144 366494 316464 373258
rect 316144 366258 316186 366494
rect 316422 366258 316464 366494
rect 316144 359494 316464 366258
rect 316144 359258 316186 359494
rect 316422 359258 316464 359494
rect 316144 352494 316464 359258
rect 316144 352258 316186 352494
rect 316422 352258 316464 352494
rect 316144 345494 316464 352258
rect 316144 345258 316186 345494
rect 316422 345258 316464 345494
rect 316144 338494 316464 345258
rect 316144 338258 316186 338494
rect 316422 338258 316464 338494
rect 316144 331494 316464 338258
rect 316144 331258 316186 331494
rect 316422 331258 316464 331494
rect 316144 324494 316464 331258
rect 316144 324258 316186 324494
rect 316422 324258 316464 324494
rect 316144 317494 316464 324258
rect 316144 317258 316186 317494
rect 316422 317258 316464 317494
rect 316144 310494 316464 317258
rect 316144 310258 316186 310494
rect 316422 310258 316464 310494
rect 316144 303494 316464 310258
rect 316144 303258 316186 303494
rect 316422 303258 316464 303494
rect 316144 296494 316464 303258
rect 316144 296258 316186 296494
rect 316422 296258 316464 296494
rect 316144 289494 316464 296258
rect 316144 289258 316186 289494
rect 316422 289258 316464 289494
rect 316144 282494 316464 289258
rect 316144 282258 316186 282494
rect 316422 282258 316464 282494
rect 316144 275494 316464 282258
rect 316144 275258 316186 275494
rect 316422 275258 316464 275494
rect 316144 268494 316464 275258
rect 316144 268258 316186 268494
rect 316422 268258 316464 268494
rect 316144 261494 316464 268258
rect 316144 261258 316186 261494
rect 316422 261258 316464 261494
rect 316144 254494 316464 261258
rect 316144 254258 316186 254494
rect 316422 254258 316464 254494
rect 316144 247494 316464 254258
rect 316144 247258 316186 247494
rect 316422 247258 316464 247494
rect 316144 240494 316464 247258
rect 316144 240258 316186 240494
rect 316422 240258 316464 240494
rect 316144 233494 316464 240258
rect 316144 233258 316186 233494
rect 316422 233258 316464 233494
rect 316144 226494 316464 233258
rect 316144 226258 316186 226494
rect 316422 226258 316464 226494
rect 316144 219494 316464 226258
rect 316144 219258 316186 219494
rect 316422 219258 316464 219494
rect 316144 212494 316464 219258
rect 316144 212258 316186 212494
rect 316422 212258 316464 212494
rect 316144 205494 316464 212258
rect 316144 205258 316186 205494
rect 316422 205258 316464 205494
rect 316144 198494 316464 205258
rect 316144 198258 316186 198494
rect 316422 198258 316464 198494
rect 316144 191494 316464 198258
rect 316144 191258 316186 191494
rect 316422 191258 316464 191494
rect 316144 184494 316464 191258
rect 316144 184258 316186 184494
rect 316422 184258 316464 184494
rect 316144 177494 316464 184258
rect 316144 177258 316186 177494
rect 316422 177258 316464 177494
rect 316144 170494 316464 177258
rect 316144 170258 316186 170494
rect 316422 170258 316464 170494
rect 316144 163494 316464 170258
rect 316144 163258 316186 163494
rect 316422 163258 316464 163494
rect 316144 156494 316464 163258
rect 316144 156258 316186 156494
rect 316422 156258 316464 156494
rect 316144 149494 316464 156258
rect 316144 149258 316186 149494
rect 316422 149258 316464 149494
rect 316144 142494 316464 149258
rect 316144 142258 316186 142494
rect 316422 142258 316464 142494
rect 316144 135494 316464 142258
rect 316144 135258 316186 135494
rect 316422 135258 316464 135494
rect 316144 128494 316464 135258
rect 316144 128258 316186 128494
rect 316422 128258 316464 128494
rect 316144 121494 316464 128258
rect 316144 121258 316186 121494
rect 316422 121258 316464 121494
rect 316144 114494 316464 121258
rect 316144 114258 316186 114494
rect 316422 114258 316464 114494
rect 316144 107494 316464 114258
rect 316144 107258 316186 107494
rect 316422 107258 316464 107494
rect 316144 100494 316464 107258
rect 316144 100258 316186 100494
rect 316422 100258 316464 100494
rect 316144 93494 316464 100258
rect 316144 93258 316186 93494
rect 316422 93258 316464 93494
rect 316144 86494 316464 93258
rect 316144 86258 316186 86494
rect 316422 86258 316464 86494
rect 316144 79494 316464 86258
rect 316144 79258 316186 79494
rect 316422 79258 316464 79494
rect 316144 72494 316464 79258
rect 316144 72258 316186 72494
rect 316422 72258 316464 72494
rect 316144 65494 316464 72258
rect 316144 65258 316186 65494
rect 316422 65258 316464 65494
rect 316144 58494 316464 65258
rect 316144 58258 316186 58494
rect 316422 58258 316464 58494
rect 316144 51494 316464 58258
rect 316144 51258 316186 51494
rect 316422 51258 316464 51494
rect 316144 44494 316464 51258
rect 316144 44258 316186 44494
rect 316422 44258 316464 44494
rect 316144 37494 316464 44258
rect 316144 37258 316186 37494
rect 316422 37258 316464 37494
rect 316144 30494 316464 37258
rect 316144 30258 316186 30494
rect 316422 30258 316464 30494
rect 316144 23494 316464 30258
rect 316144 23258 316186 23494
rect 316422 23258 316464 23494
rect 316144 16494 316464 23258
rect 316144 16258 316186 16494
rect 316422 16258 316464 16494
rect 316144 9494 316464 16258
rect 316144 9258 316186 9494
rect 316422 9258 316464 9494
rect 316144 2494 316464 9258
rect 316144 2258 316186 2494
rect 316422 2258 316464 2494
rect 316144 -746 316464 2258
rect 316144 -982 316186 -746
rect 316422 -982 316464 -746
rect 316144 -1066 316464 -982
rect 316144 -1302 316186 -1066
rect 316422 -1302 316464 -1066
rect 316144 -2294 316464 -1302
rect 317876 706198 318196 706230
rect 317876 705962 317918 706198
rect 318154 705962 318196 706198
rect 317876 705878 318196 705962
rect 317876 705642 317918 705878
rect 318154 705642 318196 705878
rect 317876 696434 318196 705642
rect 317876 696198 317918 696434
rect 318154 696198 318196 696434
rect 317876 689434 318196 696198
rect 317876 689198 317918 689434
rect 318154 689198 318196 689434
rect 317876 682434 318196 689198
rect 317876 682198 317918 682434
rect 318154 682198 318196 682434
rect 317876 675434 318196 682198
rect 317876 675198 317918 675434
rect 318154 675198 318196 675434
rect 317876 668434 318196 675198
rect 317876 668198 317918 668434
rect 318154 668198 318196 668434
rect 317876 661434 318196 668198
rect 317876 661198 317918 661434
rect 318154 661198 318196 661434
rect 317876 654434 318196 661198
rect 317876 654198 317918 654434
rect 318154 654198 318196 654434
rect 317876 647434 318196 654198
rect 317876 647198 317918 647434
rect 318154 647198 318196 647434
rect 317876 640434 318196 647198
rect 317876 640198 317918 640434
rect 318154 640198 318196 640434
rect 317876 633434 318196 640198
rect 317876 633198 317918 633434
rect 318154 633198 318196 633434
rect 317876 626434 318196 633198
rect 317876 626198 317918 626434
rect 318154 626198 318196 626434
rect 317876 619434 318196 626198
rect 317876 619198 317918 619434
rect 318154 619198 318196 619434
rect 317876 612434 318196 619198
rect 317876 612198 317918 612434
rect 318154 612198 318196 612434
rect 317876 605434 318196 612198
rect 317876 605198 317918 605434
rect 318154 605198 318196 605434
rect 317876 598434 318196 605198
rect 317876 598198 317918 598434
rect 318154 598198 318196 598434
rect 317876 591434 318196 598198
rect 317876 591198 317918 591434
rect 318154 591198 318196 591434
rect 317876 584434 318196 591198
rect 317876 584198 317918 584434
rect 318154 584198 318196 584434
rect 317876 577434 318196 584198
rect 317876 577198 317918 577434
rect 318154 577198 318196 577434
rect 317876 570434 318196 577198
rect 317876 570198 317918 570434
rect 318154 570198 318196 570434
rect 317876 563434 318196 570198
rect 317876 563198 317918 563434
rect 318154 563198 318196 563434
rect 317876 556434 318196 563198
rect 317876 556198 317918 556434
rect 318154 556198 318196 556434
rect 317876 549434 318196 556198
rect 317876 549198 317918 549434
rect 318154 549198 318196 549434
rect 317876 542434 318196 549198
rect 317876 542198 317918 542434
rect 318154 542198 318196 542434
rect 317876 535434 318196 542198
rect 317876 535198 317918 535434
rect 318154 535198 318196 535434
rect 317876 528434 318196 535198
rect 317876 528198 317918 528434
rect 318154 528198 318196 528434
rect 317876 521434 318196 528198
rect 317876 521198 317918 521434
rect 318154 521198 318196 521434
rect 317876 514434 318196 521198
rect 317876 514198 317918 514434
rect 318154 514198 318196 514434
rect 317876 507434 318196 514198
rect 317876 507198 317918 507434
rect 318154 507198 318196 507434
rect 317876 500434 318196 507198
rect 317876 500198 317918 500434
rect 318154 500198 318196 500434
rect 317876 493434 318196 500198
rect 317876 493198 317918 493434
rect 318154 493198 318196 493434
rect 317876 486434 318196 493198
rect 317876 486198 317918 486434
rect 318154 486198 318196 486434
rect 317876 479434 318196 486198
rect 317876 479198 317918 479434
rect 318154 479198 318196 479434
rect 317876 472434 318196 479198
rect 317876 472198 317918 472434
rect 318154 472198 318196 472434
rect 317876 465434 318196 472198
rect 317876 465198 317918 465434
rect 318154 465198 318196 465434
rect 317876 458434 318196 465198
rect 317876 458198 317918 458434
rect 318154 458198 318196 458434
rect 317876 451434 318196 458198
rect 317876 451198 317918 451434
rect 318154 451198 318196 451434
rect 317876 444434 318196 451198
rect 317876 444198 317918 444434
rect 318154 444198 318196 444434
rect 317876 437434 318196 444198
rect 317876 437198 317918 437434
rect 318154 437198 318196 437434
rect 317876 430434 318196 437198
rect 317876 430198 317918 430434
rect 318154 430198 318196 430434
rect 317876 423434 318196 430198
rect 317876 423198 317918 423434
rect 318154 423198 318196 423434
rect 317876 416434 318196 423198
rect 317876 416198 317918 416434
rect 318154 416198 318196 416434
rect 317876 409434 318196 416198
rect 317876 409198 317918 409434
rect 318154 409198 318196 409434
rect 317876 402434 318196 409198
rect 317876 402198 317918 402434
rect 318154 402198 318196 402434
rect 317876 395434 318196 402198
rect 317876 395198 317918 395434
rect 318154 395198 318196 395434
rect 317876 388434 318196 395198
rect 317876 388198 317918 388434
rect 318154 388198 318196 388434
rect 317876 381434 318196 388198
rect 317876 381198 317918 381434
rect 318154 381198 318196 381434
rect 317876 374434 318196 381198
rect 317876 374198 317918 374434
rect 318154 374198 318196 374434
rect 317876 367434 318196 374198
rect 317876 367198 317918 367434
rect 318154 367198 318196 367434
rect 317876 360434 318196 367198
rect 317876 360198 317918 360434
rect 318154 360198 318196 360434
rect 317876 353434 318196 360198
rect 317876 353198 317918 353434
rect 318154 353198 318196 353434
rect 317876 346434 318196 353198
rect 317876 346198 317918 346434
rect 318154 346198 318196 346434
rect 317876 339434 318196 346198
rect 317876 339198 317918 339434
rect 318154 339198 318196 339434
rect 317876 332434 318196 339198
rect 317876 332198 317918 332434
rect 318154 332198 318196 332434
rect 317876 325434 318196 332198
rect 317876 325198 317918 325434
rect 318154 325198 318196 325434
rect 317876 318434 318196 325198
rect 317876 318198 317918 318434
rect 318154 318198 318196 318434
rect 317876 311434 318196 318198
rect 317876 311198 317918 311434
rect 318154 311198 318196 311434
rect 317876 304434 318196 311198
rect 317876 304198 317918 304434
rect 318154 304198 318196 304434
rect 317876 297434 318196 304198
rect 317876 297198 317918 297434
rect 318154 297198 318196 297434
rect 317876 290434 318196 297198
rect 317876 290198 317918 290434
rect 318154 290198 318196 290434
rect 317876 283434 318196 290198
rect 317876 283198 317918 283434
rect 318154 283198 318196 283434
rect 317876 276434 318196 283198
rect 317876 276198 317918 276434
rect 318154 276198 318196 276434
rect 317876 269434 318196 276198
rect 317876 269198 317918 269434
rect 318154 269198 318196 269434
rect 317876 262434 318196 269198
rect 317876 262198 317918 262434
rect 318154 262198 318196 262434
rect 317876 255434 318196 262198
rect 317876 255198 317918 255434
rect 318154 255198 318196 255434
rect 317876 248434 318196 255198
rect 317876 248198 317918 248434
rect 318154 248198 318196 248434
rect 317876 241434 318196 248198
rect 317876 241198 317918 241434
rect 318154 241198 318196 241434
rect 317876 234434 318196 241198
rect 317876 234198 317918 234434
rect 318154 234198 318196 234434
rect 317876 227434 318196 234198
rect 317876 227198 317918 227434
rect 318154 227198 318196 227434
rect 317876 220434 318196 227198
rect 317876 220198 317918 220434
rect 318154 220198 318196 220434
rect 317876 213434 318196 220198
rect 317876 213198 317918 213434
rect 318154 213198 318196 213434
rect 317876 206434 318196 213198
rect 317876 206198 317918 206434
rect 318154 206198 318196 206434
rect 317876 199434 318196 206198
rect 317876 199198 317918 199434
rect 318154 199198 318196 199434
rect 317876 192434 318196 199198
rect 317876 192198 317918 192434
rect 318154 192198 318196 192434
rect 317876 185434 318196 192198
rect 317876 185198 317918 185434
rect 318154 185198 318196 185434
rect 317876 178434 318196 185198
rect 317876 178198 317918 178434
rect 318154 178198 318196 178434
rect 317876 171434 318196 178198
rect 317876 171198 317918 171434
rect 318154 171198 318196 171434
rect 317876 164434 318196 171198
rect 317876 164198 317918 164434
rect 318154 164198 318196 164434
rect 317876 157434 318196 164198
rect 317876 157198 317918 157434
rect 318154 157198 318196 157434
rect 317876 150434 318196 157198
rect 317876 150198 317918 150434
rect 318154 150198 318196 150434
rect 317876 143434 318196 150198
rect 317876 143198 317918 143434
rect 318154 143198 318196 143434
rect 317876 136434 318196 143198
rect 317876 136198 317918 136434
rect 318154 136198 318196 136434
rect 317876 129434 318196 136198
rect 317876 129198 317918 129434
rect 318154 129198 318196 129434
rect 317876 122434 318196 129198
rect 317876 122198 317918 122434
rect 318154 122198 318196 122434
rect 317876 115434 318196 122198
rect 317876 115198 317918 115434
rect 318154 115198 318196 115434
rect 317876 108434 318196 115198
rect 317876 108198 317918 108434
rect 318154 108198 318196 108434
rect 317876 101434 318196 108198
rect 317876 101198 317918 101434
rect 318154 101198 318196 101434
rect 317876 94434 318196 101198
rect 317876 94198 317918 94434
rect 318154 94198 318196 94434
rect 317876 87434 318196 94198
rect 317876 87198 317918 87434
rect 318154 87198 318196 87434
rect 317876 80434 318196 87198
rect 317876 80198 317918 80434
rect 318154 80198 318196 80434
rect 317876 73434 318196 80198
rect 317876 73198 317918 73434
rect 318154 73198 318196 73434
rect 317876 66434 318196 73198
rect 317876 66198 317918 66434
rect 318154 66198 318196 66434
rect 317876 59434 318196 66198
rect 317876 59198 317918 59434
rect 318154 59198 318196 59434
rect 317876 52434 318196 59198
rect 317876 52198 317918 52434
rect 318154 52198 318196 52434
rect 317876 45434 318196 52198
rect 317876 45198 317918 45434
rect 318154 45198 318196 45434
rect 317876 38434 318196 45198
rect 317876 38198 317918 38434
rect 318154 38198 318196 38434
rect 317876 31434 318196 38198
rect 317876 31198 317918 31434
rect 318154 31198 318196 31434
rect 317876 24434 318196 31198
rect 317876 24198 317918 24434
rect 318154 24198 318196 24434
rect 317876 17434 318196 24198
rect 317876 17198 317918 17434
rect 318154 17198 318196 17434
rect 317876 10434 318196 17198
rect 317876 10198 317918 10434
rect 318154 10198 318196 10434
rect 317876 3434 318196 10198
rect 317876 3198 317918 3434
rect 318154 3198 318196 3434
rect 317876 -1706 318196 3198
rect 317876 -1942 317918 -1706
rect 318154 -1942 318196 -1706
rect 317876 -2026 318196 -1942
rect 317876 -2262 317918 -2026
rect 318154 -2262 318196 -2026
rect 317876 -2294 318196 -2262
rect 323144 705238 323464 706230
rect 323144 705002 323186 705238
rect 323422 705002 323464 705238
rect 323144 704918 323464 705002
rect 323144 704682 323186 704918
rect 323422 704682 323464 704918
rect 323144 695494 323464 704682
rect 323144 695258 323186 695494
rect 323422 695258 323464 695494
rect 323144 688494 323464 695258
rect 323144 688258 323186 688494
rect 323422 688258 323464 688494
rect 323144 681494 323464 688258
rect 323144 681258 323186 681494
rect 323422 681258 323464 681494
rect 323144 674494 323464 681258
rect 323144 674258 323186 674494
rect 323422 674258 323464 674494
rect 323144 667494 323464 674258
rect 323144 667258 323186 667494
rect 323422 667258 323464 667494
rect 323144 660494 323464 667258
rect 323144 660258 323186 660494
rect 323422 660258 323464 660494
rect 323144 653494 323464 660258
rect 323144 653258 323186 653494
rect 323422 653258 323464 653494
rect 323144 646494 323464 653258
rect 323144 646258 323186 646494
rect 323422 646258 323464 646494
rect 323144 639494 323464 646258
rect 323144 639258 323186 639494
rect 323422 639258 323464 639494
rect 323144 632494 323464 639258
rect 323144 632258 323186 632494
rect 323422 632258 323464 632494
rect 323144 625494 323464 632258
rect 323144 625258 323186 625494
rect 323422 625258 323464 625494
rect 323144 618494 323464 625258
rect 323144 618258 323186 618494
rect 323422 618258 323464 618494
rect 323144 611494 323464 618258
rect 323144 611258 323186 611494
rect 323422 611258 323464 611494
rect 323144 604494 323464 611258
rect 323144 604258 323186 604494
rect 323422 604258 323464 604494
rect 323144 597494 323464 604258
rect 323144 597258 323186 597494
rect 323422 597258 323464 597494
rect 323144 590494 323464 597258
rect 323144 590258 323186 590494
rect 323422 590258 323464 590494
rect 323144 583494 323464 590258
rect 323144 583258 323186 583494
rect 323422 583258 323464 583494
rect 323144 576494 323464 583258
rect 323144 576258 323186 576494
rect 323422 576258 323464 576494
rect 323144 569494 323464 576258
rect 323144 569258 323186 569494
rect 323422 569258 323464 569494
rect 323144 562494 323464 569258
rect 323144 562258 323186 562494
rect 323422 562258 323464 562494
rect 323144 555494 323464 562258
rect 323144 555258 323186 555494
rect 323422 555258 323464 555494
rect 323144 548494 323464 555258
rect 323144 548258 323186 548494
rect 323422 548258 323464 548494
rect 323144 541494 323464 548258
rect 323144 541258 323186 541494
rect 323422 541258 323464 541494
rect 323144 534494 323464 541258
rect 323144 534258 323186 534494
rect 323422 534258 323464 534494
rect 323144 527494 323464 534258
rect 323144 527258 323186 527494
rect 323422 527258 323464 527494
rect 323144 520494 323464 527258
rect 323144 520258 323186 520494
rect 323422 520258 323464 520494
rect 323144 513494 323464 520258
rect 323144 513258 323186 513494
rect 323422 513258 323464 513494
rect 323144 506494 323464 513258
rect 323144 506258 323186 506494
rect 323422 506258 323464 506494
rect 323144 499494 323464 506258
rect 323144 499258 323186 499494
rect 323422 499258 323464 499494
rect 323144 492494 323464 499258
rect 323144 492258 323186 492494
rect 323422 492258 323464 492494
rect 323144 485494 323464 492258
rect 323144 485258 323186 485494
rect 323422 485258 323464 485494
rect 323144 478494 323464 485258
rect 323144 478258 323186 478494
rect 323422 478258 323464 478494
rect 323144 471494 323464 478258
rect 323144 471258 323186 471494
rect 323422 471258 323464 471494
rect 323144 464494 323464 471258
rect 323144 464258 323186 464494
rect 323422 464258 323464 464494
rect 323144 457494 323464 464258
rect 323144 457258 323186 457494
rect 323422 457258 323464 457494
rect 323144 450494 323464 457258
rect 323144 450258 323186 450494
rect 323422 450258 323464 450494
rect 323144 443494 323464 450258
rect 323144 443258 323186 443494
rect 323422 443258 323464 443494
rect 323144 436494 323464 443258
rect 323144 436258 323186 436494
rect 323422 436258 323464 436494
rect 323144 429494 323464 436258
rect 323144 429258 323186 429494
rect 323422 429258 323464 429494
rect 323144 422494 323464 429258
rect 323144 422258 323186 422494
rect 323422 422258 323464 422494
rect 323144 415494 323464 422258
rect 323144 415258 323186 415494
rect 323422 415258 323464 415494
rect 323144 408494 323464 415258
rect 323144 408258 323186 408494
rect 323422 408258 323464 408494
rect 323144 401494 323464 408258
rect 323144 401258 323186 401494
rect 323422 401258 323464 401494
rect 323144 394494 323464 401258
rect 323144 394258 323186 394494
rect 323422 394258 323464 394494
rect 323144 387494 323464 394258
rect 323144 387258 323186 387494
rect 323422 387258 323464 387494
rect 323144 380494 323464 387258
rect 323144 380258 323186 380494
rect 323422 380258 323464 380494
rect 323144 373494 323464 380258
rect 323144 373258 323186 373494
rect 323422 373258 323464 373494
rect 323144 366494 323464 373258
rect 323144 366258 323186 366494
rect 323422 366258 323464 366494
rect 323144 359494 323464 366258
rect 323144 359258 323186 359494
rect 323422 359258 323464 359494
rect 323144 352494 323464 359258
rect 323144 352258 323186 352494
rect 323422 352258 323464 352494
rect 323144 345494 323464 352258
rect 323144 345258 323186 345494
rect 323422 345258 323464 345494
rect 323144 338494 323464 345258
rect 323144 338258 323186 338494
rect 323422 338258 323464 338494
rect 323144 331494 323464 338258
rect 323144 331258 323186 331494
rect 323422 331258 323464 331494
rect 323144 324494 323464 331258
rect 323144 324258 323186 324494
rect 323422 324258 323464 324494
rect 323144 317494 323464 324258
rect 323144 317258 323186 317494
rect 323422 317258 323464 317494
rect 323144 310494 323464 317258
rect 323144 310258 323186 310494
rect 323422 310258 323464 310494
rect 323144 303494 323464 310258
rect 323144 303258 323186 303494
rect 323422 303258 323464 303494
rect 323144 296494 323464 303258
rect 323144 296258 323186 296494
rect 323422 296258 323464 296494
rect 323144 289494 323464 296258
rect 323144 289258 323186 289494
rect 323422 289258 323464 289494
rect 323144 282494 323464 289258
rect 323144 282258 323186 282494
rect 323422 282258 323464 282494
rect 323144 275494 323464 282258
rect 323144 275258 323186 275494
rect 323422 275258 323464 275494
rect 323144 268494 323464 275258
rect 323144 268258 323186 268494
rect 323422 268258 323464 268494
rect 323144 261494 323464 268258
rect 323144 261258 323186 261494
rect 323422 261258 323464 261494
rect 323144 254494 323464 261258
rect 323144 254258 323186 254494
rect 323422 254258 323464 254494
rect 323144 247494 323464 254258
rect 323144 247258 323186 247494
rect 323422 247258 323464 247494
rect 323144 240494 323464 247258
rect 323144 240258 323186 240494
rect 323422 240258 323464 240494
rect 323144 233494 323464 240258
rect 323144 233258 323186 233494
rect 323422 233258 323464 233494
rect 323144 226494 323464 233258
rect 323144 226258 323186 226494
rect 323422 226258 323464 226494
rect 323144 219494 323464 226258
rect 323144 219258 323186 219494
rect 323422 219258 323464 219494
rect 323144 212494 323464 219258
rect 323144 212258 323186 212494
rect 323422 212258 323464 212494
rect 323144 205494 323464 212258
rect 323144 205258 323186 205494
rect 323422 205258 323464 205494
rect 323144 198494 323464 205258
rect 323144 198258 323186 198494
rect 323422 198258 323464 198494
rect 323144 191494 323464 198258
rect 323144 191258 323186 191494
rect 323422 191258 323464 191494
rect 323144 184494 323464 191258
rect 323144 184258 323186 184494
rect 323422 184258 323464 184494
rect 323144 177494 323464 184258
rect 323144 177258 323186 177494
rect 323422 177258 323464 177494
rect 323144 170494 323464 177258
rect 323144 170258 323186 170494
rect 323422 170258 323464 170494
rect 323144 163494 323464 170258
rect 323144 163258 323186 163494
rect 323422 163258 323464 163494
rect 323144 156494 323464 163258
rect 323144 156258 323186 156494
rect 323422 156258 323464 156494
rect 323144 149494 323464 156258
rect 323144 149258 323186 149494
rect 323422 149258 323464 149494
rect 323144 142494 323464 149258
rect 323144 142258 323186 142494
rect 323422 142258 323464 142494
rect 323144 135494 323464 142258
rect 323144 135258 323186 135494
rect 323422 135258 323464 135494
rect 323144 128494 323464 135258
rect 323144 128258 323186 128494
rect 323422 128258 323464 128494
rect 323144 121494 323464 128258
rect 323144 121258 323186 121494
rect 323422 121258 323464 121494
rect 323144 114494 323464 121258
rect 323144 114258 323186 114494
rect 323422 114258 323464 114494
rect 323144 107494 323464 114258
rect 323144 107258 323186 107494
rect 323422 107258 323464 107494
rect 323144 100494 323464 107258
rect 323144 100258 323186 100494
rect 323422 100258 323464 100494
rect 323144 93494 323464 100258
rect 323144 93258 323186 93494
rect 323422 93258 323464 93494
rect 323144 86494 323464 93258
rect 323144 86258 323186 86494
rect 323422 86258 323464 86494
rect 323144 79494 323464 86258
rect 323144 79258 323186 79494
rect 323422 79258 323464 79494
rect 323144 72494 323464 79258
rect 323144 72258 323186 72494
rect 323422 72258 323464 72494
rect 323144 65494 323464 72258
rect 323144 65258 323186 65494
rect 323422 65258 323464 65494
rect 323144 58494 323464 65258
rect 323144 58258 323186 58494
rect 323422 58258 323464 58494
rect 323144 51494 323464 58258
rect 323144 51258 323186 51494
rect 323422 51258 323464 51494
rect 323144 44494 323464 51258
rect 323144 44258 323186 44494
rect 323422 44258 323464 44494
rect 323144 37494 323464 44258
rect 323144 37258 323186 37494
rect 323422 37258 323464 37494
rect 323144 30494 323464 37258
rect 323144 30258 323186 30494
rect 323422 30258 323464 30494
rect 323144 23494 323464 30258
rect 323144 23258 323186 23494
rect 323422 23258 323464 23494
rect 323144 16494 323464 23258
rect 323144 16258 323186 16494
rect 323422 16258 323464 16494
rect 323144 9494 323464 16258
rect 323144 9258 323186 9494
rect 323422 9258 323464 9494
rect 323144 2494 323464 9258
rect 323144 2258 323186 2494
rect 323422 2258 323464 2494
rect 323144 -746 323464 2258
rect 323144 -982 323186 -746
rect 323422 -982 323464 -746
rect 323144 -1066 323464 -982
rect 323144 -1302 323186 -1066
rect 323422 -1302 323464 -1066
rect 323144 -2294 323464 -1302
rect 324876 706198 325196 706230
rect 324876 705962 324918 706198
rect 325154 705962 325196 706198
rect 324876 705878 325196 705962
rect 324876 705642 324918 705878
rect 325154 705642 325196 705878
rect 324876 696434 325196 705642
rect 324876 696198 324918 696434
rect 325154 696198 325196 696434
rect 324876 689434 325196 696198
rect 324876 689198 324918 689434
rect 325154 689198 325196 689434
rect 324876 682434 325196 689198
rect 324876 682198 324918 682434
rect 325154 682198 325196 682434
rect 324876 675434 325196 682198
rect 324876 675198 324918 675434
rect 325154 675198 325196 675434
rect 324876 668434 325196 675198
rect 324876 668198 324918 668434
rect 325154 668198 325196 668434
rect 324876 661434 325196 668198
rect 324876 661198 324918 661434
rect 325154 661198 325196 661434
rect 324876 654434 325196 661198
rect 324876 654198 324918 654434
rect 325154 654198 325196 654434
rect 324876 647434 325196 654198
rect 324876 647198 324918 647434
rect 325154 647198 325196 647434
rect 324876 640434 325196 647198
rect 324876 640198 324918 640434
rect 325154 640198 325196 640434
rect 324876 633434 325196 640198
rect 324876 633198 324918 633434
rect 325154 633198 325196 633434
rect 324876 626434 325196 633198
rect 324876 626198 324918 626434
rect 325154 626198 325196 626434
rect 324876 619434 325196 626198
rect 324876 619198 324918 619434
rect 325154 619198 325196 619434
rect 324876 612434 325196 619198
rect 324876 612198 324918 612434
rect 325154 612198 325196 612434
rect 324876 605434 325196 612198
rect 324876 605198 324918 605434
rect 325154 605198 325196 605434
rect 324876 598434 325196 605198
rect 324876 598198 324918 598434
rect 325154 598198 325196 598434
rect 324876 591434 325196 598198
rect 324876 591198 324918 591434
rect 325154 591198 325196 591434
rect 324876 584434 325196 591198
rect 324876 584198 324918 584434
rect 325154 584198 325196 584434
rect 324876 577434 325196 584198
rect 324876 577198 324918 577434
rect 325154 577198 325196 577434
rect 324876 570434 325196 577198
rect 324876 570198 324918 570434
rect 325154 570198 325196 570434
rect 324876 563434 325196 570198
rect 324876 563198 324918 563434
rect 325154 563198 325196 563434
rect 324876 556434 325196 563198
rect 324876 556198 324918 556434
rect 325154 556198 325196 556434
rect 324876 549434 325196 556198
rect 324876 549198 324918 549434
rect 325154 549198 325196 549434
rect 324876 542434 325196 549198
rect 324876 542198 324918 542434
rect 325154 542198 325196 542434
rect 324876 535434 325196 542198
rect 324876 535198 324918 535434
rect 325154 535198 325196 535434
rect 324876 528434 325196 535198
rect 324876 528198 324918 528434
rect 325154 528198 325196 528434
rect 324876 521434 325196 528198
rect 324876 521198 324918 521434
rect 325154 521198 325196 521434
rect 324876 514434 325196 521198
rect 324876 514198 324918 514434
rect 325154 514198 325196 514434
rect 324876 507434 325196 514198
rect 324876 507198 324918 507434
rect 325154 507198 325196 507434
rect 324876 500434 325196 507198
rect 324876 500198 324918 500434
rect 325154 500198 325196 500434
rect 324876 493434 325196 500198
rect 324876 493198 324918 493434
rect 325154 493198 325196 493434
rect 324876 486434 325196 493198
rect 324876 486198 324918 486434
rect 325154 486198 325196 486434
rect 324876 479434 325196 486198
rect 324876 479198 324918 479434
rect 325154 479198 325196 479434
rect 324876 472434 325196 479198
rect 324876 472198 324918 472434
rect 325154 472198 325196 472434
rect 324876 465434 325196 472198
rect 324876 465198 324918 465434
rect 325154 465198 325196 465434
rect 324876 458434 325196 465198
rect 324876 458198 324918 458434
rect 325154 458198 325196 458434
rect 324876 451434 325196 458198
rect 324876 451198 324918 451434
rect 325154 451198 325196 451434
rect 324876 444434 325196 451198
rect 324876 444198 324918 444434
rect 325154 444198 325196 444434
rect 324876 437434 325196 444198
rect 324876 437198 324918 437434
rect 325154 437198 325196 437434
rect 324876 430434 325196 437198
rect 324876 430198 324918 430434
rect 325154 430198 325196 430434
rect 324876 423434 325196 430198
rect 324876 423198 324918 423434
rect 325154 423198 325196 423434
rect 324876 416434 325196 423198
rect 324876 416198 324918 416434
rect 325154 416198 325196 416434
rect 324876 409434 325196 416198
rect 324876 409198 324918 409434
rect 325154 409198 325196 409434
rect 324876 402434 325196 409198
rect 324876 402198 324918 402434
rect 325154 402198 325196 402434
rect 324876 395434 325196 402198
rect 324876 395198 324918 395434
rect 325154 395198 325196 395434
rect 324876 388434 325196 395198
rect 324876 388198 324918 388434
rect 325154 388198 325196 388434
rect 324876 381434 325196 388198
rect 324876 381198 324918 381434
rect 325154 381198 325196 381434
rect 324876 374434 325196 381198
rect 324876 374198 324918 374434
rect 325154 374198 325196 374434
rect 324876 367434 325196 374198
rect 324876 367198 324918 367434
rect 325154 367198 325196 367434
rect 324876 360434 325196 367198
rect 324876 360198 324918 360434
rect 325154 360198 325196 360434
rect 324876 353434 325196 360198
rect 324876 353198 324918 353434
rect 325154 353198 325196 353434
rect 324876 346434 325196 353198
rect 324876 346198 324918 346434
rect 325154 346198 325196 346434
rect 324876 339434 325196 346198
rect 324876 339198 324918 339434
rect 325154 339198 325196 339434
rect 324876 332434 325196 339198
rect 324876 332198 324918 332434
rect 325154 332198 325196 332434
rect 324876 325434 325196 332198
rect 324876 325198 324918 325434
rect 325154 325198 325196 325434
rect 324876 318434 325196 325198
rect 324876 318198 324918 318434
rect 325154 318198 325196 318434
rect 324876 311434 325196 318198
rect 324876 311198 324918 311434
rect 325154 311198 325196 311434
rect 324876 304434 325196 311198
rect 324876 304198 324918 304434
rect 325154 304198 325196 304434
rect 324876 297434 325196 304198
rect 324876 297198 324918 297434
rect 325154 297198 325196 297434
rect 324876 290434 325196 297198
rect 324876 290198 324918 290434
rect 325154 290198 325196 290434
rect 324876 283434 325196 290198
rect 324876 283198 324918 283434
rect 325154 283198 325196 283434
rect 324876 276434 325196 283198
rect 324876 276198 324918 276434
rect 325154 276198 325196 276434
rect 324876 269434 325196 276198
rect 324876 269198 324918 269434
rect 325154 269198 325196 269434
rect 324876 262434 325196 269198
rect 324876 262198 324918 262434
rect 325154 262198 325196 262434
rect 324876 255434 325196 262198
rect 324876 255198 324918 255434
rect 325154 255198 325196 255434
rect 324876 248434 325196 255198
rect 324876 248198 324918 248434
rect 325154 248198 325196 248434
rect 324876 241434 325196 248198
rect 324876 241198 324918 241434
rect 325154 241198 325196 241434
rect 324876 234434 325196 241198
rect 324876 234198 324918 234434
rect 325154 234198 325196 234434
rect 324876 227434 325196 234198
rect 324876 227198 324918 227434
rect 325154 227198 325196 227434
rect 324876 220434 325196 227198
rect 324876 220198 324918 220434
rect 325154 220198 325196 220434
rect 324876 213434 325196 220198
rect 324876 213198 324918 213434
rect 325154 213198 325196 213434
rect 324876 206434 325196 213198
rect 324876 206198 324918 206434
rect 325154 206198 325196 206434
rect 324876 199434 325196 206198
rect 324876 199198 324918 199434
rect 325154 199198 325196 199434
rect 324876 192434 325196 199198
rect 324876 192198 324918 192434
rect 325154 192198 325196 192434
rect 324876 185434 325196 192198
rect 324876 185198 324918 185434
rect 325154 185198 325196 185434
rect 324876 178434 325196 185198
rect 324876 178198 324918 178434
rect 325154 178198 325196 178434
rect 324876 171434 325196 178198
rect 324876 171198 324918 171434
rect 325154 171198 325196 171434
rect 324876 164434 325196 171198
rect 324876 164198 324918 164434
rect 325154 164198 325196 164434
rect 324876 157434 325196 164198
rect 324876 157198 324918 157434
rect 325154 157198 325196 157434
rect 324876 150434 325196 157198
rect 324876 150198 324918 150434
rect 325154 150198 325196 150434
rect 324876 143434 325196 150198
rect 324876 143198 324918 143434
rect 325154 143198 325196 143434
rect 324876 136434 325196 143198
rect 324876 136198 324918 136434
rect 325154 136198 325196 136434
rect 324876 129434 325196 136198
rect 324876 129198 324918 129434
rect 325154 129198 325196 129434
rect 324876 122434 325196 129198
rect 324876 122198 324918 122434
rect 325154 122198 325196 122434
rect 324876 115434 325196 122198
rect 324876 115198 324918 115434
rect 325154 115198 325196 115434
rect 324876 108434 325196 115198
rect 324876 108198 324918 108434
rect 325154 108198 325196 108434
rect 324876 101434 325196 108198
rect 324876 101198 324918 101434
rect 325154 101198 325196 101434
rect 324876 94434 325196 101198
rect 324876 94198 324918 94434
rect 325154 94198 325196 94434
rect 324876 87434 325196 94198
rect 324876 87198 324918 87434
rect 325154 87198 325196 87434
rect 324876 80434 325196 87198
rect 324876 80198 324918 80434
rect 325154 80198 325196 80434
rect 324876 73434 325196 80198
rect 324876 73198 324918 73434
rect 325154 73198 325196 73434
rect 324876 66434 325196 73198
rect 324876 66198 324918 66434
rect 325154 66198 325196 66434
rect 324876 59434 325196 66198
rect 324876 59198 324918 59434
rect 325154 59198 325196 59434
rect 324876 52434 325196 59198
rect 324876 52198 324918 52434
rect 325154 52198 325196 52434
rect 324876 45434 325196 52198
rect 324876 45198 324918 45434
rect 325154 45198 325196 45434
rect 324876 38434 325196 45198
rect 324876 38198 324918 38434
rect 325154 38198 325196 38434
rect 324876 31434 325196 38198
rect 324876 31198 324918 31434
rect 325154 31198 325196 31434
rect 324876 24434 325196 31198
rect 324876 24198 324918 24434
rect 325154 24198 325196 24434
rect 324876 17434 325196 24198
rect 324876 17198 324918 17434
rect 325154 17198 325196 17434
rect 324876 10434 325196 17198
rect 324876 10198 324918 10434
rect 325154 10198 325196 10434
rect 324876 3434 325196 10198
rect 324876 3198 324918 3434
rect 325154 3198 325196 3434
rect 324876 -1706 325196 3198
rect 324876 -1942 324918 -1706
rect 325154 -1942 325196 -1706
rect 324876 -2026 325196 -1942
rect 324876 -2262 324918 -2026
rect 325154 -2262 325196 -2026
rect 324876 -2294 325196 -2262
rect 330144 705238 330464 706230
rect 330144 705002 330186 705238
rect 330422 705002 330464 705238
rect 330144 704918 330464 705002
rect 330144 704682 330186 704918
rect 330422 704682 330464 704918
rect 330144 695494 330464 704682
rect 330144 695258 330186 695494
rect 330422 695258 330464 695494
rect 330144 688494 330464 695258
rect 330144 688258 330186 688494
rect 330422 688258 330464 688494
rect 330144 681494 330464 688258
rect 330144 681258 330186 681494
rect 330422 681258 330464 681494
rect 330144 674494 330464 681258
rect 330144 674258 330186 674494
rect 330422 674258 330464 674494
rect 330144 667494 330464 674258
rect 330144 667258 330186 667494
rect 330422 667258 330464 667494
rect 330144 660494 330464 667258
rect 330144 660258 330186 660494
rect 330422 660258 330464 660494
rect 330144 653494 330464 660258
rect 330144 653258 330186 653494
rect 330422 653258 330464 653494
rect 330144 646494 330464 653258
rect 330144 646258 330186 646494
rect 330422 646258 330464 646494
rect 330144 639494 330464 646258
rect 330144 639258 330186 639494
rect 330422 639258 330464 639494
rect 330144 632494 330464 639258
rect 330144 632258 330186 632494
rect 330422 632258 330464 632494
rect 330144 625494 330464 632258
rect 330144 625258 330186 625494
rect 330422 625258 330464 625494
rect 330144 618494 330464 625258
rect 330144 618258 330186 618494
rect 330422 618258 330464 618494
rect 330144 611494 330464 618258
rect 330144 611258 330186 611494
rect 330422 611258 330464 611494
rect 330144 604494 330464 611258
rect 330144 604258 330186 604494
rect 330422 604258 330464 604494
rect 330144 597494 330464 604258
rect 330144 597258 330186 597494
rect 330422 597258 330464 597494
rect 330144 590494 330464 597258
rect 330144 590258 330186 590494
rect 330422 590258 330464 590494
rect 330144 583494 330464 590258
rect 330144 583258 330186 583494
rect 330422 583258 330464 583494
rect 330144 576494 330464 583258
rect 330144 576258 330186 576494
rect 330422 576258 330464 576494
rect 330144 569494 330464 576258
rect 330144 569258 330186 569494
rect 330422 569258 330464 569494
rect 330144 562494 330464 569258
rect 330144 562258 330186 562494
rect 330422 562258 330464 562494
rect 330144 555494 330464 562258
rect 330144 555258 330186 555494
rect 330422 555258 330464 555494
rect 330144 548494 330464 555258
rect 330144 548258 330186 548494
rect 330422 548258 330464 548494
rect 330144 541494 330464 548258
rect 330144 541258 330186 541494
rect 330422 541258 330464 541494
rect 330144 534494 330464 541258
rect 330144 534258 330186 534494
rect 330422 534258 330464 534494
rect 330144 527494 330464 534258
rect 330144 527258 330186 527494
rect 330422 527258 330464 527494
rect 330144 520494 330464 527258
rect 330144 520258 330186 520494
rect 330422 520258 330464 520494
rect 330144 513494 330464 520258
rect 330144 513258 330186 513494
rect 330422 513258 330464 513494
rect 330144 506494 330464 513258
rect 330144 506258 330186 506494
rect 330422 506258 330464 506494
rect 330144 499494 330464 506258
rect 330144 499258 330186 499494
rect 330422 499258 330464 499494
rect 330144 492494 330464 499258
rect 330144 492258 330186 492494
rect 330422 492258 330464 492494
rect 330144 485494 330464 492258
rect 330144 485258 330186 485494
rect 330422 485258 330464 485494
rect 330144 478494 330464 485258
rect 330144 478258 330186 478494
rect 330422 478258 330464 478494
rect 330144 471494 330464 478258
rect 330144 471258 330186 471494
rect 330422 471258 330464 471494
rect 330144 464494 330464 471258
rect 330144 464258 330186 464494
rect 330422 464258 330464 464494
rect 330144 457494 330464 464258
rect 330144 457258 330186 457494
rect 330422 457258 330464 457494
rect 330144 450494 330464 457258
rect 330144 450258 330186 450494
rect 330422 450258 330464 450494
rect 330144 443494 330464 450258
rect 330144 443258 330186 443494
rect 330422 443258 330464 443494
rect 330144 436494 330464 443258
rect 330144 436258 330186 436494
rect 330422 436258 330464 436494
rect 330144 429494 330464 436258
rect 330144 429258 330186 429494
rect 330422 429258 330464 429494
rect 330144 422494 330464 429258
rect 330144 422258 330186 422494
rect 330422 422258 330464 422494
rect 330144 415494 330464 422258
rect 330144 415258 330186 415494
rect 330422 415258 330464 415494
rect 330144 408494 330464 415258
rect 330144 408258 330186 408494
rect 330422 408258 330464 408494
rect 330144 401494 330464 408258
rect 330144 401258 330186 401494
rect 330422 401258 330464 401494
rect 330144 394494 330464 401258
rect 330144 394258 330186 394494
rect 330422 394258 330464 394494
rect 330144 387494 330464 394258
rect 330144 387258 330186 387494
rect 330422 387258 330464 387494
rect 330144 380494 330464 387258
rect 330144 380258 330186 380494
rect 330422 380258 330464 380494
rect 330144 373494 330464 380258
rect 330144 373258 330186 373494
rect 330422 373258 330464 373494
rect 330144 366494 330464 373258
rect 330144 366258 330186 366494
rect 330422 366258 330464 366494
rect 330144 359494 330464 366258
rect 330144 359258 330186 359494
rect 330422 359258 330464 359494
rect 330144 352494 330464 359258
rect 330144 352258 330186 352494
rect 330422 352258 330464 352494
rect 330144 345494 330464 352258
rect 330144 345258 330186 345494
rect 330422 345258 330464 345494
rect 330144 338494 330464 345258
rect 330144 338258 330186 338494
rect 330422 338258 330464 338494
rect 330144 331494 330464 338258
rect 330144 331258 330186 331494
rect 330422 331258 330464 331494
rect 330144 324494 330464 331258
rect 330144 324258 330186 324494
rect 330422 324258 330464 324494
rect 330144 317494 330464 324258
rect 330144 317258 330186 317494
rect 330422 317258 330464 317494
rect 330144 310494 330464 317258
rect 330144 310258 330186 310494
rect 330422 310258 330464 310494
rect 330144 303494 330464 310258
rect 330144 303258 330186 303494
rect 330422 303258 330464 303494
rect 330144 296494 330464 303258
rect 330144 296258 330186 296494
rect 330422 296258 330464 296494
rect 330144 289494 330464 296258
rect 330144 289258 330186 289494
rect 330422 289258 330464 289494
rect 330144 282494 330464 289258
rect 330144 282258 330186 282494
rect 330422 282258 330464 282494
rect 330144 275494 330464 282258
rect 330144 275258 330186 275494
rect 330422 275258 330464 275494
rect 330144 268494 330464 275258
rect 330144 268258 330186 268494
rect 330422 268258 330464 268494
rect 330144 261494 330464 268258
rect 330144 261258 330186 261494
rect 330422 261258 330464 261494
rect 330144 254494 330464 261258
rect 330144 254258 330186 254494
rect 330422 254258 330464 254494
rect 330144 247494 330464 254258
rect 330144 247258 330186 247494
rect 330422 247258 330464 247494
rect 330144 240494 330464 247258
rect 330144 240258 330186 240494
rect 330422 240258 330464 240494
rect 330144 233494 330464 240258
rect 330144 233258 330186 233494
rect 330422 233258 330464 233494
rect 330144 226494 330464 233258
rect 330144 226258 330186 226494
rect 330422 226258 330464 226494
rect 330144 219494 330464 226258
rect 330144 219258 330186 219494
rect 330422 219258 330464 219494
rect 330144 212494 330464 219258
rect 330144 212258 330186 212494
rect 330422 212258 330464 212494
rect 330144 205494 330464 212258
rect 330144 205258 330186 205494
rect 330422 205258 330464 205494
rect 330144 198494 330464 205258
rect 330144 198258 330186 198494
rect 330422 198258 330464 198494
rect 330144 191494 330464 198258
rect 330144 191258 330186 191494
rect 330422 191258 330464 191494
rect 330144 184494 330464 191258
rect 330144 184258 330186 184494
rect 330422 184258 330464 184494
rect 330144 177494 330464 184258
rect 330144 177258 330186 177494
rect 330422 177258 330464 177494
rect 330144 170494 330464 177258
rect 330144 170258 330186 170494
rect 330422 170258 330464 170494
rect 330144 163494 330464 170258
rect 330144 163258 330186 163494
rect 330422 163258 330464 163494
rect 330144 156494 330464 163258
rect 330144 156258 330186 156494
rect 330422 156258 330464 156494
rect 330144 149494 330464 156258
rect 330144 149258 330186 149494
rect 330422 149258 330464 149494
rect 330144 142494 330464 149258
rect 330144 142258 330186 142494
rect 330422 142258 330464 142494
rect 330144 135494 330464 142258
rect 330144 135258 330186 135494
rect 330422 135258 330464 135494
rect 330144 128494 330464 135258
rect 330144 128258 330186 128494
rect 330422 128258 330464 128494
rect 330144 121494 330464 128258
rect 330144 121258 330186 121494
rect 330422 121258 330464 121494
rect 330144 114494 330464 121258
rect 330144 114258 330186 114494
rect 330422 114258 330464 114494
rect 330144 107494 330464 114258
rect 330144 107258 330186 107494
rect 330422 107258 330464 107494
rect 330144 100494 330464 107258
rect 330144 100258 330186 100494
rect 330422 100258 330464 100494
rect 330144 93494 330464 100258
rect 330144 93258 330186 93494
rect 330422 93258 330464 93494
rect 330144 86494 330464 93258
rect 330144 86258 330186 86494
rect 330422 86258 330464 86494
rect 330144 79494 330464 86258
rect 330144 79258 330186 79494
rect 330422 79258 330464 79494
rect 330144 72494 330464 79258
rect 330144 72258 330186 72494
rect 330422 72258 330464 72494
rect 330144 65494 330464 72258
rect 330144 65258 330186 65494
rect 330422 65258 330464 65494
rect 330144 58494 330464 65258
rect 330144 58258 330186 58494
rect 330422 58258 330464 58494
rect 330144 51494 330464 58258
rect 330144 51258 330186 51494
rect 330422 51258 330464 51494
rect 330144 44494 330464 51258
rect 330144 44258 330186 44494
rect 330422 44258 330464 44494
rect 330144 37494 330464 44258
rect 330144 37258 330186 37494
rect 330422 37258 330464 37494
rect 330144 30494 330464 37258
rect 330144 30258 330186 30494
rect 330422 30258 330464 30494
rect 330144 23494 330464 30258
rect 330144 23258 330186 23494
rect 330422 23258 330464 23494
rect 330144 16494 330464 23258
rect 330144 16258 330186 16494
rect 330422 16258 330464 16494
rect 330144 9494 330464 16258
rect 330144 9258 330186 9494
rect 330422 9258 330464 9494
rect 330144 2494 330464 9258
rect 330144 2258 330186 2494
rect 330422 2258 330464 2494
rect 330144 -746 330464 2258
rect 330144 -982 330186 -746
rect 330422 -982 330464 -746
rect 330144 -1066 330464 -982
rect 330144 -1302 330186 -1066
rect 330422 -1302 330464 -1066
rect 330144 -2294 330464 -1302
rect 331876 706198 332196 706230
rect 331876 705962 331918 706198
rect 332154 705962 332196 706198
rect 331876 705878 332196 705962
rect 331876 705642 331918 705878
rect 332154 705642 332196 705878
rect 331876 696434 332196 705642
rect 331876 696198 331918 696434
rect 332154 696198 332196 696434
rect 331876 689434 332196 696198
rect 331876 689198 331918 689434
rect 332154 689198 332196 689434
rect 331876 682434 332196 689198
rect 331876 682198 331918 682434
rect 332154 682198 332196 682434
rect 331876 675434 332196 682198
rect 331876 675198 331918 675434
rect 332154 675198 332196 675434
rect 331876 668434 332196 675198
rect 331876 668198 331918 668434
rect 332154 668198 332196 668434
rect 331876 661434 332196 668198
rect 331876 661198 331918 661434
rect 332154 661198 332196 661434
rect 331876 654434 332196 661198
rect 331876 654198 331918 654434
rect 332154 654198 332196 654434
rect 331876 647434 332196 654198
rect 331876 647198 331918 647434
rect 332154 647198 332196 647434
rect 331876 640434 332196 647198
rect 331876 640198 331918 640434
rect 332154 640198 332196 640434
rect 331876 633434 332196 640198
rect 331876 633198 331918 633434
rect 332154 633198 332196 633434
rect 331876 626434 332196 633198
rect 331876 626198 331918 626434
rect 332154 626198 332196 626434
rect 331876 619434 332196 626198
rect 331876 619198 331918 619434
rect 332154 619198 332196 619434
rect 331876 612434 332196 619198
rect 331876 612198 331918 612434
rect 332154 612198 332196 612434
rect 331876 605434 332196 612198
rect 331876 605198 331918 605434
rect 332154 605198 332196 605434
rect 331876 598434 332196 605198
rect 331876 598198 331918 598434
rect 332154 598198 332196 598434
rect 331876 591434 332196 598198
rect 331876 591198 331918 591434
rect 332154 591198 332196 591434
rect 331876 584434 332196 591198
rect 331876 584198 331918 584434
rect 332154 584198 332196 584434
rect 331876 577434 332196 584198
rect 331876 577198 331918 577434
rect 332154 577198 332196 577434
rect 331876 570434 332196 577198
rect 331876 570198 331918 570434
rect 332154 570198 332196 570434
rect 331876 563434 332196 570198
rect 331876 563198 331918 563434
rect 332154 563198 332196 563434
rect 331876 556434 332196 563198
rect 331876 556198 331918 556434
rect 332154 556198 332196 556434
rect 331876 549434 332196 556198
rect 331876 549198 331918 549434
rect 332154 549198 332196 549434
rect 331876 542434 332196 549198
rect 331876 542198 331918 542434
rect 332154 542198 332196 542434
rect 331876 535434 332196 542198
rect 331876 535198 331918 535434
rect 332154 535198 332196 535434
rect 331876 528434 332196 535198
rect 331876 528198 331918 528434
rect 332154 528198 332196 528434
rect 331876 521434 332196 528198
rect 331876 521198 331918 521434
rect 332154 521198 332196 521434
rect 331876 514434 332196 521198
rect 331876 514198 331918 514434
rect 332154 514198 332196 514434
rect 331876 507434 332196 514198
rect 331876 507198 331918 507434
rect 332154 507198 332196 507434
rect 331876 500434 332196 507198
rect 331876 500198 331918 500434
rect 332154 500198 332196 500434
rect 331876 493434 332196 500198
rect 331876 493198 331918 493434
rect 332154 493198 332196 493434
rect 331876 486434 332196 493198
rect 331876 486198 331918 486434
rect 332154 486198 332196 486434
rect 331876 479434 332196 486198
rect 331876 479198 331918 479434
rect 332154 479198 332196 479434
rect 331876 472434 332196 479198
rect 331876 472198 331918 472434
rect 332154 472198 332196 472434
rect 331876 465434 332196 472198
rect 331876 465198 331918 465434
rect 332154 465198 332196 465434
rect 331876 458434 332196 465198
rect 331876 458198 331918 458434
rect 332154 458198 332196 458434
rect 331876 451434 332196 458198
rect 331876 451198 331918 451434
rect 332154 451198 332196 451434
rect 331876 444434 332196 451198
rect 331876 444198 331918 444434
rect 332154 444198 332196 444434
rect 331876 437434 332196 444198
rect 331876 437198 331918 437434
rect 332154 437198 332196 437434
rect 331876 430434 332196 437198
rect 331876 430198 331918 430434
rect 332154 430198 332196 430434
rect 331876 423434 332196 430198
rect 331876 423198 331918 423434
rect 332154 423198 332196 423434
rect 331876 416434 332196 423198
rect 331876 416198 331918 416434
rect 332154 416198 332196 416434
rect 331876 409434 332196 416198
rect 331876 409198 331918 409434
rect 332154 409198 332196 409434
rect 331876 402434 332196 409198
rect 331876 402198 331918 402434
rect 332154 402198 332196 402434
rect 331876 395434 332196 402198
rect 331876 395198 331918 395434
rect 332154 395198 332196 395434
rect 331876 388434 332196 395198
rect 331876 388198 331918 388434
rect 332154 388198 332196 388434
rect 331876 381434 332196 388198
rect 331876 381198 331918 381434
rect 332154 381198 332196 381434
rect 331876 374434 332196 381198
rect 331876 374198 331918 374434
rect 332154 374198 332196 374434
rect 331876 367434 332196 374198
rect 331876 367198 331918 367434
rect 332154 367198 332196 367434
rect 331876 360434 332196 367198
rect 331876 360198 331918 360434
rect 332154 360198 332196 360434
rect 331876 353434 332196 360198
rect 331876 353198 331918 353434
rect 332154 353198 332196 353434
rect 331876 346434 332196 353198
rect 331876 346198 331918 346434
rect 332154 346198 332196 346434
rect 331876 339434 332196 346198
rect 331876 339198 331918 339434
rect 332154 339198 332196 339434
rect 331876 332434 332196 339198
rect 331876 332198 331918 332434
rect 332154 332198 332196 332434
rect 331876 325434 332196 332198
rect 331876 325198 331918 325434
rect 332154 325198 332196 325434
rect 331876 318434 332196 325198
rect 331876 318198 331918 318434
rect 332154 318198 332196 318434
rect 331876 311434 332196 318198
rect 331876 311198 331918 311434
rect 332154 311198 332196 311434
rect 331876 304434 332196 311198
rect 331876 304198 331918 304434
rect 332154 304198 332196 304434
rect 331876 297434 332196 304198
rect 331876 297198 331918 297434
rect 332154 297198 332196 297434
rect 331876 290434 332196 297198
rect 331876 290198 331918 290434
rect 332154 290198 332196 290434
rect 331876 283434 332196 290198
rect 331876 283198 331918 283434
rect 332154 283198 332196 283434
rect 331876 276434 332196 283198
rect 331876 276198 331918 276434
rect 332154 276198 332196 276434
rect 331876 269434 332196 276198
rect 331876 269198 331918 269434
rect 332154 269198 332196 269434
rect 331876 262434 332196 269198
rect 331876 262198 331918 262434
rect 332154 262198 332196 262434
rect 331876 255434 332196 262198
rect 331876 255198 331918 255434
rect 332154 255198 332196 255434
rect 331876 248434 332196 255198
rect 331876 248198 331918 248434
rect 332154 248198 332196 248434
rect 331876 241434 332196 248198
rect 331876 241198 331918 241434
rect 332154 241198 332196 241434
rect 331876 234434 332196 241198
rect 331876 234198 331918 234434
rect 332154 234198 332196 234434
rect 331876 227434 332196 234198
rect 331876 227198 331918 227434
rect 332154 227198 332196 227434
rect 331876 220434 332196 227198
rect 331876 220198 331918 220434
rect 332154 220198 332196 220434
rect 331876 213434 332196 220198
rect 331876 213198 331918 213434
rect 332154 213198 332196 213434
rect 331876 206434 332196 213198
rect 331876 206198 331918 206434
rect 332154 206198 332196 206434
rect 331876 199434 332196 206198
rect 331876 199198 331918 199434
rect 332154 199198 332196 199434
rect 331876 192434 332196 199198
rect 331876 192198 331918 192434
rect 332154 192198 332196 192434
rect 331876 185434 332196 192198
rect 331876 185198 331918 185434
rect 332154 185198 332196 185434
rect 331876 178434 332196 185198
rect 331876 178198 331918 178434
rect 332154 178198 332196 178434
rect 331876 171434 332196 178198
rect 331876 171198 331918 171434
rect 332154 171198 332196 171434
rect 331876 164434 332196 171198
rect 331876 164198 331918 164434
rect 332154 164198 332196 164434
rect 331876 157434 332196 164198
rect 331876 157198 331918 157434
rect 332154 157198 332196 157434
rect 331876 150434 332196 157198
rect 331876 150198 331918 150434
rect 332154 150198 332196 150434
rect 331876 143434 332196 150198
rect 331876 143198 331918 143434
rect 332154 143198 332196 143434
rect 331876 136434 332196 143198
rect 331876 136198 331918 136434
rect 332154 136198 332196 136434
rect 331876 129434 332196 136198
rect 331876 129198 331918 129434
rect 332154 129198 332196 129434
rect 331876 122434 332196 129198
rect 331876 122198 331918 122434
rect 332154 122198 332196 122434
rect 331876 115434 332196 122198
rect 331876 115198 331918 115434
rect 332154 115198 332196 115434
rect 331876 108434 332196 115198
rect 331876 108198 331918 108434
rect 332154 108198 332196 108434
rect 331876 101434 332196 108198
rect 331876 101198 331918 101434
rect 332154 101198 332196 101434
rect 331876 94434 332196 101198
rect 331876 94198 331918 94434
rect 332154 94198 332196 94434
rect 331876 87434 332196 94198
rect 331876 87198 331918 87434
rect 332154 87198 332196 87434
rect 331876 80434 332196 87198
rect 331876 80198 331918 80434
rect 332154 80198 332196 80434
rect 331876 73434 332196 80198
rect 331876 73198 331918 73434
rect 332154 73198 332196 73434
rect 331876 66434 332196 73198
rect 331876 66198 331918 66434
rect 332154 66198 332196 66434
rect 331876 59434 332196 66198
rect 331876 59198 331918 59434
rect 332154 59198 332196 59434
rect 331876 52434 332196 59198
rect 331876 52198 331918 52434
rect 332154 52198 332196 52434
rect 331876 45434 332196 52198
rect 331876 45198 331918 45434
rect 332154 45198 332196 45434
rect 331876 38434 332196 45198
rect 331876 38198 331918 38434
rect 332154 38198 332196 38434
rect 331876 31434 332196 38198
rect 331876 31198 331918 31434
rect 332154 31198 332196 31434
rect 331876 24434 332196 31198
rect 331876 24198 331918 24434
rect 332154 24198 332196 24434
rect 331876 17434 332196 24198
rect 331876 17198 331918 17434
rect 332154 17198 332196 17434
rect 331876 10434 332196 17198
rect 331876 10198 331918 10434
rect 332154 10198 332196 10434
rect 331876 3434 332196 10198
rect 331876 3198 331918 3434
rect 332154 3198 332196 3434
rect 331876 -1706 332196 3198
rect 331876 -1942 331918 -1706
rect 332154 -1942 332196 -1706
rect 331876 -2026 332196 -1942
rect 331876 -2262 331918 -2026
rect 332154 -2262 332196 -2026
rect 331876 -2294 332196 -2262
rect 337144 705238 337464 706230
rect 337144 705002 337186 705238
rect 337422 705002 337464 705238
rect 337144 704918 337464 705002
rect 337144 704682 337186 704918
rect 337422 704682 337464 704918
rect 337144 695494 337464 704682
rect 337144 695258 337186 695494
rect 337422 695258 337464 695494
rect 337144 688494 337464 695258
rect 337144 688258 337186 688494
rect 337422 688258 337464 688494
rect 337144 681494 337464 688258
rect 337144 681258 337186 681494
rect 337422 681258 337464 681494
rect 337144 674494 337464 681258
rect 337144 674258 337186 674494
rect 337422 674258 337464 674494
rect 337144 667494 337464 674258
rect 337144 667258 337186 667494
rect 337422 667258 337464 667494
rect 337144 660494 337464 667258
rect 337144 660258 337186 660494
rect 337422 660258 337464 660494
rect 337144 653494 337464 660258
rect 337144 653258 337186 653494
rect 337422 653258 337464 653494
rect 337144 646494 337464 653258
rect 337144 646258 337186 646494
rect 337422 646258 337464 646494
rect 337144 639494 337464 646258
rect 337144 639258 337186 639494
rect 337422 639258 337464 639494
rect 337144 632494 337464 639258
rect 337144 632258 337186 632494
rect 337422 632258 337464 632494
rect 337144 625494 337464 632258
rect 337144 625258 337186 625494
rect 337422 625258 337464 625494
rect 337144 618494 337464 625258
rect 337144 618258 337186 618494
rect 337422 618258 337464 618494
rect 337144 611494 337464 618258
rect 337144 611258 337186 611494
rect 337422 611258 337464 611494
rect 337144 604494 337464 611258
rect 337144 604258 337186 604494
rect 337422 604258 337464 604494
rect 337144 597494 337464 604258
rect 337144 597258 337186 597494
rect 337422 597258 337464 597494
rect 337144 590494 337464 597258
rect 337144 590258 337186 590494
rect 337422 590258 337464 590494
rect 337144 583494 337464 590258
rect 337144 583258 337186 583494
rect 337422 583258 337464 583494
rect 337144 576494 337464 583258
rect 337144 576258 337186 576494
rect 337422 576258 337464 576494
rect 337144 569494 337464 576258
rect 337144 569258 337186 569494
rect 337422 569258 337464 569494
rect 337144 562494 337464 569258
rect 337144 562258 337186 562494
rect 337422 562258 337464 562494
rect 337144 555494 337464 562258
rect 337144 555258 337186 555494
rect 337422 555258 337464 555494
rect 337144 548494 337464 555258
rect 337144 548258 337186 548494
rect 337422 548258 337464 548494
rect 337144 541494 337464 548258
rect 337144 541258 337186 541494
rect 337422 541258 337464 541494
rect 337144 534494 337464 541258
rect 337144 534258 337186 534494
rect 337422 534258 337464 534494
rect 337144 527494 337464 534258
rect 337144 527258 337186 527494
rect 337422 527258 337464 527494
rect 337144 520494 337464 527258
rect 337144 520258 337186 520494
rect 337422 520258 337464 520494
rect 337144 513494 337464 520258
rect 337144 513258 337186 513494
rect 337422 513258 337464 513494
rect 337144 506494 337464 513258
rect 337144 506258 337186 506494
rect 337422 506258 337464 506494
rect 337144 499494 337464 506258
rect 337144 499258 337186 499494
rect 337422 499258 337464 499494
rect 337144 492494 337464 499258
rect 337144 492258 337186 492494
rect 337422 492258 337464 492494
rect 337144 485494 337464 492258
rect 337144 485258 337186 485494
rect 337422 485258 337464 485494
rect 337144 478494 337464 485258
rect 337144 478258 337186 478494
rect 337422 478258 337464 478494
rect 337144 471494 337464 478258
rect 337144 471258 337186 471494
rect 337422 471258 337464 471494
rect 337144 464494 337464 471258
rect 337144 464258 337186 464494
rect 337422 464258 337464 464494
rect 337144 457494 337464 464258
rect 337144 457258 337186 457494
rect 337422 457258 337464 457494
rect 337144 450494 337464 457258
rect 337144 450258 337186 450494
rect 337422 450258 337464 450494
rect 337144 443494 337464 450258
rect 337144 443258 337186 443494
rect 337422 443258 337464 443494
rect 337144 436494 337464 443258
rect 337144 436258 337186 436494
rect 337422 436258 337464 436494
rect 337144 429494 337464 436258
rect 337144 429258 337186 429494
rect 337422 429258 337464 429494
rect 337144 422494 337464 429258
rect 337144 422258 337186 422494
rect 337422 422258 337464 422494
rect 337144 415494 337464 422258
rect 337144 415258 337186 415494
rect 337422 415258 337464 415494
rect 337144 408494 337464 415258
rect 337144 408258 337186 408494
rect 337422 408258 337464 408494
rect 337144 401494 337464 408258
rect 337144 401258 337186 401494
rect 337422 401258 337464 401494
rect 337144 394494 337464 401258
rect 337144 394258 337186 394494
rect 337422 394258 337464 394494
rect 337144 387494 337464 394258
rect 337144 387258 337186 387494
rect 337422 387258 337464 387494
rect 337144 380494 337464 387258
rect 337144 380258 337186 380494
rect 337422 380258 337464 380494
rect 337144 373494 337464 380258
rect 337144 373258 337186 373494
rect 337422 373258 337464 373494
rect 337144 366494 337464 373258
rect 337144 366258 337186 366494
rect 337422 366258 337464 366494
rect 337144 359494 337464 366258
rect 337144 359258 337186 359494
rect 337422 359258 337464 359494
rect 337144 352494 337464 359258
rect 337144 352258 337186 352494
rect 337422 352258 337464 352494
rect 337144 345494 337464 352258
rect 337144 345258 337186 345494
rect 337422 345258 337464 345494
rect 337144 338494 337464 345258
rect 337144 338258 337186 338494
rect 337422 338258 337464 338494
rect 337144 331494 337464 338258
rect 337144 331258 337186 331494
rect 337422 331258 337464 331494
rect 337144 324494 337464 331258
rect 337144 324258 337186 324494
rect 337422 324258 337464 324494
rect 337144 317494 337464 324258
rect 337144 317258 337186 317494
rect 337422 317258 337464 317494
rect 337144 310494 337464 317258
rect 337144 310258 337186 310494
rect 337422 310258 337464 310494
rect 337144 303494 337464 310258
rect 337144 303258 337186 303494
rect 337422 303258 337464 303494
rect 337144 296494 337464 303258
rect 337144 296258 337186 296494
rect 337422 296258 337464 296494
rect 337144 289494 337464 296258
rect 337144 289258 337186 289494
rect 337422 289258 337464 289494
rect 337144 282494 337464 289258
rect 337144 282258 337186 282494
rect 337422 282258 337464 282494
rect 337144 275494 337464 282258
rect 337144 275258 337186 275494
rect 337422 275258 337464 275494
rect 337144 268494 337464 275258
rect 337144 268258 337186 268494
rect 337422 268258 337464 268494
rect 337144 261494 337464 268258
rect 337144 261258 337186 261494
rect 337422 261258 337464 261494
rect 337144 254494 337464 261258
rect 337144 254258 337186 254494
rect 337422 254258 337464 254494
rect 337144 247494 337464 254258
rect 337144 247258 337186 247494
rect 337422 247258 337464 247494
rect 337144 240494 337464 247258
rect 337144 240258 337186 240494
rect 337422 240258 337464 240494
rect 337144 233494 337464 240258
rect 337144 233258 337186 233494
rect 337422 233258 337464 233494
rect 337144 226494 337464 233258
rect 337144 226258 337186 226494
rect 337422 226258 337464 226494
rect 337144 219494 337464 226258
rect 337144 219258 337186 219494
rect 337422 219258 337464 219494
rect 337144 212494 337464 219258
rect 337144 212258 337186 212494
rect 337422 212258 337464 212494
rect 337144 205494 337464 212258
rect 337144 205258 337186 205494
rect 337422 205258 337464 205494
rect 337144 198494 337464 205258
rect 337144 198258 337186 198494
rect 337422 198258 337464 198494
rect 337144 191494 337464 198258
rect 337144 191258 337186 191494
rect 337422 191258 337464 191494
rect 337144 184494 337464 191258
rect 337144 184258 337186 184494
rect 337422 184258 337464 184494
rect 337144 177494 337464 184258
rect 337144 177258 337186 177494
rect 337422 177258 337464 177494
rect 337144 170494 337464 177258
rect 337144 170258 337186 170494
rect 337422 170258 337464 170494
rect 337144 163494 337464 170258
rect 337144 163258 337186 163494
rect 337422 163258 337464 163494
rect 337144 156494 337464 163258
rect 337144 156258 337186 156494
rect 337422 156258 337464 156494
rect 337144 149494 337464 156258
rect 337144 149258 337186 149494
rect 337422 149258 337464 149494
rect 337144 142494 337464 149258
rect 337144 142258 337186 142494
rect 337422 142258 337464 142494
rect 337144 135494 337464 142258
rect 337144 135258 337186 135494
rect 337422 135258 337464 135494
rect 337144 128494 337464 135258
rect 337144 128258 337186 128494
rect 337422 128258 337464 128494
rect 337144 121494 337464 128258
rect 337144 121258 337186 121494
rect 337422 121258 337464 121494
rect 337144 114494 337464 121258
rect 337144 114258 337186 114494
rect 337422 114258 337464 114494
rect 337144 107494 337464 114258
rect 337144 107258 337186 107494
rect 337422 107258 337464 107494
rect 337144 100494 337464 107258
rect 337144 100258 337186 100494
rect 337422 100258 337464 100494
rect 337144 93494 337464 100258
rect 337144 93258 337186 93494
rect 337422 93258 337464 93494
rect 337144 86494 337464 93258
rect 337144 86258 337186 86494
rect 337422 86258 337464 86494
rect 337144 79494 337464 86258
rect 337144 79258 337186 79494
rect 337422 79258 337464 79494
rect 337144 72494 337464 79258
rect 337144 72258 337186 72494
rect 337422 72258 337464 72494
rect 337144 65494 337464 72258
rect 337144 65258 337186 65494
rect 337422 65258 337464 65494
rect 337144 58494 337464 65258
rect 337144 58258 337186 58494
rect 337422 58258 337464 58494
rect 337144 51494 337464 58258
rect 337144 51258 337186 51494
rect 337422 51258 337464 51494
rect 337144 44494 337464 51258
rect 337144 44258 337186 44494
rect 337422 44258 337464 44494
rect 337144 37494 337464 44258
rect 337144 37258 337186 37494
rect 337422 37258 337464 37494
rect 337144 30494 337464 37258
rect 337144 30258 337186 30494
rect 337422 30258 337464 30494
rect 337144 23494 337464 30258
rect 337144 23258 337186 23494
rect 337422 23258 337464 23494
rect 337144 16494 337464 23258
rect 337144 16258 337186 16494
rect 337422 16258 337464 16494
rect 337144 9494 337464 16258
rect 337144 9258 337186 9494
rect 337422 9258 337464 9494
rect 337144 2494 337464 9258
rect 337144 2258 337186 2494
rect 337422 2258 337464 2494
rect 337144 -746 337464 2258
rect 337144 -982 337186 -746
rect 337422 -982 337464 -746
rect 337144 -1066 337464 -982
rect 337144 -1302 337186 -1066
rect 337422 -1302 337464 -1066
rect 337144 -2294 337464 -1302
rect 338876 706198 339196 706230
rect 338876 705962 338918 706198
rect 339154 705962 339196 706198
rect 338876 705878 339196 705962
rect 338876 705642 338918 705878
rect 339154 705642 339196 705878
rect 338876 696434 339196 705642
rect 338876 696198 338918 696434
rect 339154 696198 339196 696434
rect 338876 689434 339196 696198
rect 338876 689198 338918 689434
rect 339154 689198 339196 689434
rect 338876 682434 339196 689198
rect 338876 682198 338918 682434
rect 339154 682198 339196 682434
rect 338876 675434 339196 682198
rect 338876 675198 338918 675434
rect 339154 675198 339196 675434
rect 338876 668434 339196 675198
rect 338876 668198 338918 668434
rect 339154 668198 339196 668434
rect 338876 661434 339196 668198
rect 338876 661198 338918 661434
rect 339154 661198 339196 661434
rect 338876 654434 339196 661198
rect 338876 654198 338918 654434
rect 339154 654198 339196 654434
rect 338876 647434 339196 654198
rect 338876 647198 338918 647434
rect 339154 647198 339196 647434
rect 338876 640434 339196 647198
rect 338876 640198 338918 640434
rect 339154 640198 339196 640434
rect 338876 633434 339196 640198
rect 338876 633198 338918 633434
rect 339154 633198 339196 633434
rect 338876 626434 339196 633198
rect 338876 626198 338918 626434
rect 339154 626198 339196 626434
rect 338876 619434 339196 626198
rect 338876 619198 338918 619434
rect 339154 619198 339196 619434
rect 338876 612434 339196 619198
rect 338876 612198 338918 612434
rect 339154 612198 339196 612434
rect 338876 605434 339196 612198
rect 338876 605198 338918 605434
rect 339154 605198 339196 605434
rect 338876 598434 339196 605198
rect 338876 598198 338918 598434
rect 339154 598198 339196 598434
rect 338876 591434 339196 598198
rect 338876 591198 338918 591434
rect 339154 591198 339196 591434
rect 338876 584434 339196 591198
rect 338876 584198 338918 584434
rect 339154 584198 339196 584434
rect 338876 577434 339196 584198
rect 338876 577198 338918 577434
rect 339154 577198 339196 577434
rect 338876 570434 339196 577198
rect 338876 570198 338918 570434
rect 339154 570198 339196 570434
rect 338876 563434 339196 570198
rect 338876 563198 338918 563434
rect 339154 563198 339196 563434
rect 338876 556434 339196 563198
rect 338876 556198 338918 556434
rect 339154 556198 339196 556434
rect 338876 549434 339196 556198
rect 338876 549198 338918 549434
rect 339154 549198 339196 549434
rect 338876 542434 339196 549198
rect 338876 542198 338918 542434
rect 339154 542198 339196 542434
rect 338876 535434 339196 542198
rect 338876 535198 338918 535434
rect 339154 535198 339196 535434
rect 338876 528434 339196 535198
rect 338876 528198 338918 528434
rect 339154 528198 339196 528434
rect 338876 521434 339196 528198
rect 338876 521198 338918 521434
rect 339154 521198 339196 521434
rect 338876 514434 339196 521198
rect 338876 514198 338918 514434
rect 339154 514198 339196 514434
rect 338876 507434 339196 514198
rect 338876 507198 338918 507434
rect 339154 507198 339196 507434
rect 338876 500434 339196 507198
rect 338876 500198 338918 500434
rect 339154 500198 339196 500434
rect 338876 493434 339196 500198
rect 338876 493198 338918 493434
rect 339154 493198 339196 493434
rect 338876 486434 339196 493198
rect 338876 486198 338918 486434
rect 339154 486198 339196 486434
rect 338876 479434 339196 486198
rect 338876 479198 338918 479434
rect 339154 479198 339196 479434
rect 338876 472434 339196 479198
rect 338876 472198 338918 472434
rect 339154 472198 339196 472434
rect 338876 465434 339196 472198
rect 338876 465198 338918 465434
rect 339154 465198 339196 465434
rect 338876 458434 339196 465198
rect 338876 458198 338918 458434
rect 339154 458198 339196 458434
rect 338876 451434 339196 458198
rect 338876 451198 338918 451434
rect 339154 451198 339196 451434
rect 338876 444434 339196 451198
rect 338876 444198 338918 444434
rect 339154 444198 339196 444434
rect 338876 437434 339196 444198
rect 338876 437198 338918 437434
rect 339154 437198 339196 437434
rect 338876 430434 339196 437198
rect 338876 430198 338918 430434
rect 339154 430198 339196 430434
rect 338876 423434 339196 430198
rect 338876 423198 338918 423434
rect 339154 423198 339196 423434
rect 338876 416434 339196 423198
rect 338876 416198 338918 416434
rect 339154 416198 339196 416434
rect 338876 409434 339196 416198
rect 338876 409198 338918 409434
rect 339154 409198 339196 409434
rect 338876 402434 339196 409198
rect 338876 402198 338918 402434
rect 339154 402198 339196 402434
rect 338876 395434 339196 402198
rect 338876 395198 338918 395434
rect 339154 395198 339196 395434
rect 338876 388434 339196 395198
rect 338876 388198 338918 388434
rect 339154 388198 339196 388434
rect 338876 381434 339196 388198
rect 338876 381198 338918 381434
rect 339154 381198 339196 381434
rect 338876 374434 339196 381198
rect 338876 374198 338918 374434
rect 339154 374198 339196 374434
rect 338876 367434 339196 374198
rect 338876 367198 338918 367434
rect 339154 367198 339196 367434
rect 338876 360434 339196 367198
rect 338876 360198 338918 360434
rect 339154 360198 339196 360434
rect 338876 353434 339196 360198
rect 338876 353198 338918 353434
rect 339154 353198 339196 353434
rect 338876 346434 339196 353198
rect 338876 346198 338918 346434
rect 339154 346198 339196 346434
rect 338876 339434 339196 346198
rect 338876 339198 338918 339434
rect 339154 339198 339196 339434
rect 338876 332434 339196 339198
rect 338876 332198 338918 332434
rect 339154 332198 339196 332434
rect 338876 325434 339196 332198
rect 338876 325198 338918 325434
rect 339154 325198 339196 325434
rect 338876 318434 339196 325198
rect 338876 318198 338918 318434
rect 339154 318198 339196 318434
rect 338876 311434 339196 318198
rect 338876 311198 338918 311434
rect 339154 311198 339196 311434
rect 338876 304434 339196 311198
rect 338876 304198 338918 304434
rect 339154 304198 339196 304434
rect 338876 297434 339196 304198
rect 338876 297198 338918 297434
rect 339154 297198 339196 297434
rect 338876 290434 339196 297198
rect 338876 290198 338918 290434
rect 339154 290198 339196 290434
rect 338876 283434 339196 290198
rect 338876 283198 338918 283434
rect 339154 283198 339196 283434
rect 338876 276434 339196 283198
rect 338876 276198 338918 276434
rect 339154 276198 339196 276434
rect 338876 269434 339196 276198
rect 338876 269198 338918 269434
rect 339154 269198 339196 269434
rect 338876 262434 339196 269198
rect 338876 262198 338918 262434
rect 339154 262198 339196 262434
rect 338876 255434 339196 262198
rect 338876 255198 338918 255434
rect 339154 255198 339196 255434
rect 338876 248434 339196 255198
rect 338876 248198 338918 248434
rect 339154 248198 339196 248434
rect 338876 241434 339196 248198
rect 338876 241198 338918 241434
rect 339154 241198 339196 241434
rect 338876 234434 339196 241198
rect 338876 234198 338918 234434
rect 339154 234198 339196 234434
rect 338876 227434 339196 234198
rect 338876 227198 338918 227434
rect 339154 227198 339196 227434
rect 338876 220434 339196 227198
rect 338876 220198 338918 220434
rect 339154 220198 339196 220434
rect 338876 213434 339196 220198
rect 338876 213198 338918 213434
rect 339154 213198 339196 213434
rect 338876 206434 339196 213198
rect 338876 206198 338918 206434
rect 339154 206198 339196 206434
rect 338876 199434 339196 206198
rect 338876 199198 338918 199434
rect 339154 199198 339196 199434
rect 338876 192434 339196 199198
rect 338876 192198 338918 192434
rect 339154 192198 339196 192434
rect 338876 185434 339196 192198
rect 338876 185198 338918 185434
rect 339154 185198 339196 185434
rect 338876 178434 339196 185198
rect 338876 178198 338918 178434
rect 339154 178198 339196 178434
rect 338876 171434 339196 178198
rect 338876 171198 338918 171434
rect 339154 171198 339196 171434
rect 338876 164434 339196 171198
rect 338876 164198 338918 164434
rect 339154 164198 339196 164434
rect 338876 157434 339196 164198
rect 338876 157198 338918 157434
rect 339154 157198 339196 157434
rect 338876 150434 339196 157198
rect 338876 150198 338918 150434
rect 339154 150198 339196 150434
rect 338876 143434 339196 150198
rect 338876 143198 338918 143434
rect 339154 143198 339196 143434
rect 338876 136434 339196 143198
rect 338876 136198 338918 136434
rect 339154 136198 339196 136434
rect 338876 129434 339196 136198
rect 338876 129198 338918 129434
rect 339154 129198 339196 129434
rect 338876 122434 339196 129198
rect 338876 122198 338918 122434
rect 339154 122198 339196 122434
rect 338876 115434 339196 122198
rect 338876 115198 338918 115434
rect 339154 115198 339196 115434
rect 338876 108434 339196 115198
rect 338876 108198 338918 108434
rect 339154 108198 339196 108434
rect 338876 101434 339196 108198
rect 338876 101198 338918 101434
rect 339154 101198 339196 101434
rect 338876 94434 339196 101198
rect 338876 94198 338918 94434
rect 339154 94198 339196 94434
rect 338876 87434 339196 94198
rect 338876 87198 338918 87434
rect 339154 87198 339196 87434
rect 338876 80434 339196 87198
rect 338876 80198 338918 80434
rect 339154 80198 339196 80434
rect 338876 73434 339196 80198
rect 338876 73198 338918 73434
rect 339154 73198 339196 73434
rect 338876 66434 339196 73198
rect 338876 66198 338918 66434
rect 339154 66198 339196 66434
rect 338876 59434 339196 66198
rect 338876 59198 338918 59434
rect 339154 59198 339196 59434
rect 338876 52434 339196 59198
rect 338876 52198 338918 52434
rect 339154 52198 339196 52434
rect 338876 45434 339196 52198
rect 338876 45198 338918 45434
rect 339154 45198 339196 45434
rect 338876 38434 339196 45198
rect 338876 38198 338918 38434
rect 339154 38198 339196 38434
rect 338876 31434 339196 38198
rect 338876 31198 338918 31434
rect 339154 31198 339196 31434
rect 338876 24434 339196 31198
rect 338876 24198 338918 24434
rect 339154 24198 339196 24434
rect 338876 17434 339196 24198
rect 338876 17198 338918 17434
rect 339154 17198 339196 17434
rect 338876 10434 339196 17198
rect 338876 10198 338918 10434
rect 339154 10198 339196 10434
rect 338876 3434 339196 10198
rect 338876 3198 338918 3434
rect 339154 3198 339196 3434
rect 338876 -1706 339196 3198
rect 338876 -1942 338918 -1706
rect 339154 -1942 339196 -1706
rect 338876 -2026 339196 -1942
rect 338876 -2262 338918 -2026
rect 339154 -2262 339196 -2026
rect 338876 -2294 339196 -2262
rect 344144 705238 344464 706230
rect 344144 705002 344186 705238
rect 344422 705002 344464 705238
rect 344144 704918 344464 705002
rect 344144 704682 344186 704918
rect 344422 704682 344464 704918
rect 344144 695494 344464 704682
rect 344144 695258 344186 695494
rect 344422 695258 344464 695494
rect 344144 688494 344464 695258
rect 344144 688258 344186 688494
rect 344422 688258 344464 688494
rect 344144 681494 344464 688258
rect 344144 681258 344186 681494
rect 344422 681258 344464 681494
rect 344144 674494 344464 681258
rect 344144 674258 344186 674494
rect 344422 674258 344464 674494
rect 344144 667494 344464 674258
rect 344144 667258 344186 667494
rect 344422 667258 344464 667494
rect 344144 660494 344464 667258
rect 344144 660258 344186 660494
rect 344422 660258 344464 660494
rect 344144 653494 344464 660258
rect 344144 653258 344186 653494
rect 344422 653258 344464 653494
rect 344144 646494 344464 653258
rect 344144 646258 344186 646494
rect 344422 646258 344464 646494
rect 344144 639494 344464 646258
rect 344144 639258 344186 639494
rect 344422 639258 344464 639494
rect 344144 632494 344464 639258
rect 344144 632258 344186 632494
rect 344422 632258 344464 632494
rect 344144 625494 344464 632258
rect 344144 625258 344186 625494
rect 344422 625258 344464 625494
rect 344144 618494 344464 625258
rect 344144 618258 344186 618494
rect 344422 618258 344464 618494
rect 344144 611494 344464 618258
rect 344144 611258 344186 611494
rect 344422 611258 344464 611494
rect 344144 604494 344464 611258
rect 344144 604258 344186 604494
rect 344422 604258 344464 604494
rect 344144 597494 344464 604258
rect 344144 597258 344186 597494
rect 344422 597258 344464 597494
rect 344144 590494 344464 597258
rect 344144 590258 344186 590494
rect 344422 590258 344464 590494
rect 344144 583494 344464 590258
rect 344144 583258 344186 583494
rect 344422 583258 344464 583494
rect 344144 576494 344464 583258
rect 344144 576258 344186 576494
rect 344422 576258 344464 576494
rect 344144 569494 344464 576258
rect 344144 569258 344186 569494
rect 344422 569258 344464 569494
rect 344144 562494 344464 569258
rect 344144 562258 344186 562494
rect 344422 562258 344464 562494
rect 344144 555494 344464 562258
rect 344144 555258 344186 555494
rect 344422 555258 344464 555494
rect 344144 548494 344464 555258
rect 344144 548258 344186 548494
rect 344422 548258 344464 548494
rect 344144 541494 344464 548258
rect 344144 541258 344186 541494
rect 344422 541258 344464 541494
rect 344144 534494 344464 541258
rect 344144 534258 344186 534494
rect 344422 534258 344464 534494
rect 344144 527494 344464 534258
rect 344144 527258 344186 527494
rect 344422 527258 344464 527494
rect 344144 520494 344464 527258
rect 344144 520258 344186 520494
rect 344422 520258 344464 520494
rect 344144 513494 344464 520258
rect 344144 513258 344186 513494
rect 344422 513258 344464 513494
rect 344144 506494 344464 513258
rect 344144 506258 344186 506494
rect 344422 506258 344464 506494
rect 344144 499494 344464 506258
rect 344144 499258 344186 499494
rect 344422 499258 344464 499494
rect 344144 492494 344464 499258
rect 344144 492258 344186 492494
rect 344422 492258 344464 492494
rect 344144 485494 344464 492258
rect 344144 485258 344186 485494
rect 344422 485258 344464 485494
rect 344144 478494 344464 485258
rect 344144 478258 344186 478494
rect 344422 478258 344464 478494
rect 344144 471494 344464 478258
rect 344144 471258 344186 471494
rect 344422 471258 344464 471494
rect 344144 464494 344464 471258
rect 344144 464258 344186 464494
rect 344422 464258 344464 464494
rect 344144 457494 344464 464258
rect 344144 457258 344186 457494
rect 344422 457258 344464 457494
rect 344144 450494 344464 457258
rect 344144 450258 344186 450494
rect 344422 450258 344464 450494
rect 344144 443494 344464 450258
rect 344144 443258 344186 443494
rect 344422 443258 344464 443494
rect 344144 436494 344464 443258
rect 344144 436258 344186 436494
rect 344422 436258 344464 436494
rect 344144 429494 344464 436258
rect 344144 429258 344186 429494
rect 344422 429258 344464 429494
rect 344144 422494 344464 429258
rect 344144 422258 344186 422494
rect 344422 422258 344464 422494
rect 344144 415494 344464 422258
rect 344144 415258 344186 415494
rect 344422 415258 344464 415494
rect 344144 408494 344464 415258
rect 344144 408258 344186 408494
rect 344422 408258 344464 408494
rect 344144 401494 344464 408258
rect 344144 401258 344186 401494
rect 344422 401258 344464 401494
rect 344144 394494 344464 401258
rect 344144 394258 344186 394494
rect 344422 394258 344464 394494
rect 344144 387494 344464 394258
rect 344144 387258 344186 387494
rect 344422 387258 344464 387494
rect 344144 380494 344464 387258
rect 344144 380258 344186 380494
rect 344422 380258 344464 380494
rect 344144 373494 344464 380258
rect 344144 373258 344186 373494
rect 344422 373258 344464 373494
rect 344144 366494 344464 373258
rect 344144 366258 344186 366494
rect 344422 366258 344464 366494
rect 344144 359494 344464 366258
rect 344144 359258 344186 359494
rect 344422 359258 344464 359494
rect 344144 352494 344464 359258
rect 344144 352258 344186 352494
rect 344422 352258 344464 352494
rect 344144 345494 344464 352258
rect 344144 345258 344186 345494
rect 344422 345258 344464 345494
rect 344144 338494 344464 345258
rect 344144 338258 344186 338494
rect 344422 338258 344464 338494
rect 344144 331494 344464 338258
rect 344144 331258 344186 331494
rect 344422 331258 344464 331494
rect 344144 324494 344464 331258
rect 344144 324258 344186 324494
rect 344422 324258 344464 324494
rect 344144 317494 344464 324258
rect 344144 317258 344186 317494
rect 344422 317258 344464 317494
rect 344144 310494 344464 317258
rect 344144 310258 344186 310494
rect 344422 310258 344464 310494
rect 344144 303494 344464 310258
rect 344144 303258 344186 303494
rect 344422 303258 344464 303494
rect 344144 296494 344464 303258
rect 344144 296258 344186 296494
rect 344422 296258 344464 296494
rect 344144 289494 344464 296258
rect 344144 289258 344186 289494
rect 344422 289258 344464 289494
rect 344144 282494 344464 289258
rect 344144 282258 344186 282494
rect 344422 282258 344464 282494
rect 344144 275494 344464 282258
rect 344144 275258 344186 275494
rect 344422 275258 344464 275494
rect 344144 268494 344464 275258
rect 344144 268258 344186 268494
rect 344422 268258 344464 268494
rect 344144 261494 344464 268258
rect 344144 261258 344186 261494
rect 344422 261258 344464 261494
rect 344144 254494 344464 261258
rect 344144 254258 344186 254494
rect 344422 254258 344464 254494
rect 344144 247494 344464 254258
rect 344144 247258 344186 247494
rect 344422 247258 344464 247494
rect 344144 240494 344464 247258
rect 344144 240258 344186 240494
rect 344422 240258 344464 240494
rect 344144 233494 344464 240258
rect 344144 233258 344186 233494
rect 344422 233258 344464 233494
rect 344144 226494 344464 233258
rect 344144 226258 344186 226494
rect 344422 226258 344464 226494
rect 344144 219494 344464 226258
rect 344144 219258 344186 219494
rect 344422 219258 344464 219494
rect 344144 212494 344464 219258
rect 344144 212258 344186 212494
rect 344422 212258 344464 212494
rect 344144 205494 344464 212258
rect 344144 205258 344186 205494
rect 344422 205258 344464 205494
rect 344144 198494 344464 205258
rect 344144 198258 344186 198494
rect 344422 198258 344464 198494
rect 344144 191494 344464 198258
rect 344144 191258 344186 191494
rect 344422 191258 344464 191494
rect 344144 184494 344464 191258
rect 344144 184258 344186 184494
rect 344422 184258 344464 184494
rect 344144 177494 344464 184258
rect 344144 177258 344186 177494
rect 344422 177258 344464 177494
rect 344144 170494 344464 177258
rect 344144 170258 344186 170494
rect 344422 170258 344464 170494
rect 344144 163494 344464 170258
rect 344144 163258 344186 163494
rect 344422 163258 344464 163494
rect 344144 156494 344464 163258
rect 344144 156258 344186 156494
rect 344422 156258 344464 156494
rect 344144 149494 344464 156258
rect 344144 149258 344186 149494
rect 344422 149258 344464 149494
rect 344144 142494 344464 149258
rect 344144 142258 344186 142494
rect 344422 142258 344464 142494
rect 344144 135494 344464 142258
rect 344144 135258 344186 135494
rect 344422 135258 344464 135494
rect 344144 128494 344464 135258
rect 344144 128258 344186 128494
rect 344422 128258 344464 128494
rect 344144 121494 344464 128258
rect 344144 121258 344186 121494
rect 344422 121258 344464 121494
rect 344144 114494 344464 121258
rect 344144 114258 344186 114494
rect 344422 114258 344464 114494
rect 344144 107494 344464 114258
rect 344144 107258 344186 107494
rect 344422 107258 344464 107494
rect 344144 100494 344464 107258
rect 344144 100258 344186 100494
rect 344422 100258 344464 100494
rect 344144 93494 344464 100258
rect 344144 93258 344186 93494
rect 344422 93258 344464 93494
rect 344144 86494 344464 93258
rect 344144 86258 344186 86494
rect 344422 86258 344464 86494
rect 344144 79494 344464 86258
rect 344144 79258 344186 79494
rect 344422 79258 344464 79494
rect 344144 72494 344464 79258
rect 344144 72258 344186 72494
rect 344422 72258 344464 72494
rect 344144 65494 344464 72258
rect 344144 65258 344186 65494
rect 344422 65258 344464 65494
rect 344144 58494 344464 65258
rect 344144 58258 344186 58494
rect 344422 58258 344464 58494
rect 344144 51494 344464 58258
rect 344144 51258 344186 51494
rect 344422 51258 344464 51494
rect 344144 44494 344464 51258
rect 344144 44258 344186 44494
rect 344422 44258 344464 44494
rect 344144 37494 344464 44258
rect 344144 37258 344186 37494
rect 344422 37258 344464 37494
rect 344144 30494 344464 37258
rect 344144 30258 344186 30494
rect 344422 30258 344464 30494
rect 344144 23494 344464 30258
rect 344144 23258 344186 23494
rect 344422 23258 344464 23494
rect 344144 16494 344464 23258
rect 344144 16258 344186 16494
rect 344422 16258 344464 16494
rect 344144 9494 344464 16258
rect 344144 9258 344186 9494
rect 344422 9258 344464 9494
rect 344144 2494 344464 9258
rect 344144 2258 344186 2494
rect 344422 2258 344464 2494
rect 344144 -746 344464 2258
rect 344144 -982 344186 -746
rect 344422 -982 344464 -746
rect 344144 -1066 344464 -982
rect 344144 -1302 344186 -1066
rect 344422 -1302 344464 -1066
rect 344144 -2294 344464 -1302
rect 345876 706198 346196 706230
rect 345876 705962 345918 706198
rect 346154 705962 346196 706198
rect 345876 705878 346196 705962
rect 345876 705642 345918 705878
rect 346154 705642 346196 705878
rect 345876 696434 346196 705642
rect 345876 696198 345918 696434
rect 346154 696198 346196 696434
rect 345876 689434 346196 696198
rect 345876 689198 345918 689434
rect 346154 689198 346196 689434
rect 345876 682434 346196 689198
rect 345876 682198 345918 682434
rect 346154 682198 346196 682434
rect 345876 675434 346196 682198
rect 345876 675198 345918 675434
rect 346154 675198 346196 675434
rect 345876 668434 346196 675198
rect 345876 668198 345918 668434
rect 346154 668198 346196 668434
rect 345876 661434 346196 668198
rect 345876 661198 345918 661434
rect 346154 661198 346196 661434
rect 345876 654434 346196 661198
rect 345876 654198 345918 654434
rect 346154 654198 346196 654434
rect 345876 647434 346196 654198
rect 345876 647198 345918 647434
rect 346154 647198 346196 647434
rect 345876 640434 346196 647198
rect 345876 640198 345918 640434
rect 346154 640198 346196 640434
rect 345876 633434 346196 640198
rect 345876 633198 345918 633434
rect 346154 633198 346196 633434
rect 345876 626434 346196 633198
rect 345876 626198 345918 626434
rect 346154 626198 346196 626434
rect 345876 619434 346196 626198
rect 345876 619198 345918 619434
rect 346154 619198 346196 619434
rect 345876 612434 346196 619198
rect 345876 612198 345918 612434
rect 346154 612198 346196 612434
rect 345876 605434 346196 612198
rect 345876 605198 345918 605434
rect 346154 605198 346196 605434
rect 345876 598434 346196 605198
rect 345876 598198 345918 598434
rect 346154 598198 346196 598434
rect 345876 591434 346196 598198
rect 345876 591198 345918 591434
rect 346154 591198 346196 591434
rect 345876 584434 346196 591198
rect 345876 584198 345918 584434
rect 346154 584198 346196 584434
rect 345876 577434 346196 584198
rect 345876 577198 345918 577434
rect 346154 577198 346196 577434
rect 345876 570434 346196 577198
rect 345876 570198 345918 570434
rect 346154 570198 346196 570434
rect 345876 563434 346196 570198
rect 345876 563198 345918 563434
rect 346154 563198 346196 563434
rect 345876 556434 346196 563198
rect 345876 556198 345918 556434
rect 346154 556198 346196 556434
rect 345876 549434 346196 556198
rect 345876 549198 345918 549434
rect 346154 549198 346196 549434
rect 345876 542434 346196 549198
rect 345876 542198 345918 542434
rect 346154 542198 346196 542434
rect 345876 535434 346196 542198
rect 345876 535198 345918 535434
rect 346154 535198 346196 535434
rect 345876 528434 346196 535198
rect 345876 528198 345918 528434
rect 346154 528198 346196 528434
rect 345876 521434 346196 528198
rect 345876 521198 345918 521434
rect 346154 521198 346196 521434
rect 345876 514434 346196 521198
rect 345876 514198 345918 514434
rect 346154 514198 346196 514434
rect 345876 507434 346196 514198
rect 345876 507198 345918 507434
rect 346154 507198 346196 507434
rect 345876 500434 346196 507198
rect 345876 500198 345918 500434
rect 346154 500198 346196 500434
rect 345876 493434 346196 500198
rect 345876 493198 345918 493434
rect 346154 493198 346196 493434
rect 345876 486434 346196 493198
rect 345876 486198 345918 486434
rect 346154 486198 346196 486434
rect 345876 479434 346196 486198
rect 345876 479198 345918 479434
rect 346154 479198 346196 479434
rect 345876 472434 346196 479198
rect 345876 472198 345918 472434
rect 346154 472198 346196 472434
rect 345876 465434 346196 472198
rect 345876 465198 345918 465434
rect 346154 465198 346196 465434
rect 345876 458434 346196 465198
rect 345876 458198 345918 458434
rect 346154 458198 346196 458434
rect 345876 451434 346196 458198
rect 345876 451198 345918 451434
rect 346154 451198 346196 451434
rect 345876 444434 346196 451198
rect 345876 444198 345918 444434
rect 346154 444198 346196 444434
rect 345876 437434 346196 444198
rect 345876 437198 345918 437434
rect 346154 437198 346196 437434
rect 345876 430434 346196 437198
rect 345876 430198 345918 430434
rect 346154 430198 346196 430434
rect 345876 423434 346196 430198
rect 345876 423198 345918 423434
rect 346154 423198 346196 423434
rect 345876 416434 346196 423198
rect 345876 416198 345918 416434
rect 346154 416198 346196 416434
rect 345876 409434 346196 416198
rect 345876 409198 345918 409434
rect 346154 409198 346196 409434
rect 345876 402434 346196 409198
rect 345876 402198 345918 402434
rect 346154 402198 346196 402434
rect 345876 395434 346196 402198
rect 345876 395198 345918 395434
rect 346154 395198 346196 395434
rect 345876 388434 346196 395198
rect 345876 388198 345918 388434
rect 346154 388198 346196 388434
rect 345876 381434 346196 388198
rect 345876 381198 345918 381434
rect 346154 381198 346196 381434
rect 345876 374434 346196 381198
rect 345876 374198 345918 374434
rect 346154 374198 346196 374434
rect 345876 367434 346196 374198
rect 345876 367198 345918 367434
rect 346154 367198 346196 367434
rect 345876 360434 346196 367198
rect 345876 360198 345918 360434
rect 346154 360198 346196 360434
rect 345876 353434 346196 360198
rect 345876 353198 345918 353434
rect 346154 353198 346196 353434
rect 345876 346434 346196 353198
rect 345876 346198 345918 346434
rect 346154 346198 346196 346434
rect 345876 339434 346196 346198
rect 345876 339198 345918 339434
rect 346154 339198 346196 339434
rect 345876 332434 346196 339198
rect 345876 332198 345918 332434
rect 346154 332198 346196 332434
rect 345876 325434 346196 332198
rect 345876 325198 345918 325434
rect 346154 325198 346196 325434
rect 345876 318434 346196 325198
rect 345876 318198 345918 318434
rect 346154 318198 346196 318434
rect 345876 311434 346196 318198
rect 345876 311198 345918 311434
rect 346154 311198 346196 311434
rect 345876 304434 346196 311198
rect 345876 304198 345918 304434
rect 346154 304198 346196 304434
rect 345876 297434 346196 304198
rect 345876 297198 345918 297434
rect 346154 297198 346196 297434
rect 345876 290434 346196 297198
rect 345876 290198 345918 290434
rect 346154 290198 346196 290434
rect 345876 283434 346196 290198
rect 345876 283198 345918 283434
rect 346154 283198 346196 283434
rect 345876 276434 346196 283198
rect 345876 276198 345918 276434
rect 346154 276198 346196 276434
rect 345876 269434 346196 276198
rect 345876 269198 345918 269434
rect 346154 269198 346196 269434
rect 345876 262434 346196 269198
rect 345876 262198 345918 262434
rect 346154 262198 346196 262434
rect 345876 255434 346196 262198
rect 345876 255198 345918 255434
rect 346154 255198 346196 255434
rect 345876 248434 346196 255198
rect 345876 248198 345918 248434
rect 346154 248198 346196 248434
rect 345876 241434 346196 248198
rect 345876 241198 345918 241434
rect 346154 241198 346196 241434
rect 345876 234434 346196 241198
rect 345876 234198 345918 234434
rect 346154 234198 346196 234434
rect 345876 227434 346196 234198
rect 345876 227198 345918 227434
rect 346154 227198 346196 227434
rect 345876 220434 346196 227198
rect 345876 220198 345918 220434
rect 346154 220198 346196 220434
rect 345876 213434 346196 220198
rect 345876 213198 345918 213434
rect 346154 213198 346196 213434
rect 345876 206434 346196 213198
rect 345876 206198 345918 206434
rect 346154 206198 346196 206434
rect 345876 199434 346196 206198
rect 345876 199198 345918 199434
rect 346154 199198 346196 199434
rect 345876 192434 346196 199198
rect 345876 192198 345918 192434
rect 346154 192198 346196 192434
rect 345876 185434 346196 192198
rect 345876 185198 345918 185434
rect 346154 185198 346196 185434
rect 345876 178434 346196 185198
rect 345876 178198 345918 178434
rect 346154 178198 346196 178434
rect 345876 171434 346196 178198
rect 345876 171198 345918 171434
rect 346154 171198 346196 171434
rect 345876 164434 346196 171198
rect 345876 164198 345918 164434
rect 346154 164198 346196 164434
rect 345876 157434 346196 164198
rect 345876 157198 345918 157434
rect 346154 157198 346196 157434
rect 345876 150434 346196 157198
rect 345876 150198 345918 150434
rect 346154 150198 346196 150434
rect 345876 143434 346196 150198
rect 345876 143198 345918 143434
rect 346154 143198 346196 143434
rect 345876 136434 346196 143198
rect 345876 136198 345918 136434
rect 346154 136198 346196 136434
rect 345876 129434 346196 136198
rect 345876 129198 345918 129434
rect 346154 129198 346196 129434
rect 345876 122434 346196 129198
rect 345876 122198 345918 122434
rect 346154 122198 346196 122434
rect 345876 115434 346196 122198
rect 345876 115198 345918 115434
rect 346154 115198 346196 115434
rect 345876 108434 346196 115198
rect 345876 108198 345918 108434
rect 346154 108198 346196 108434
rect 345876 101434 346196 108198
rect 345876 101198 345918 101434
rect 346154 101198 346196 101434
rect 345876 94434 346196 101198
rect 345876 94198 345918 94434
rect 346154 94198 346196 94434
rect 345876 87434 346196 94198
rect 345876 87198 345918 87434
rect 346154 87198 346196 87434
rect 345876 80434 346196 87198
rect 345876 80198 345918 80434
rect 346154 80198 346196 80434
rect 345876 73434 346196 80198
rect 345876 73198 345918 73434
rect 346154 73198 346196 73434
rect 345876 66434 346196 73198
rect 345876 66198 345918 66434
rect 346154 66198 346196 66434
rect 345876 59434 346196 66198
rect 345876 59198 345918 59434
rect 346154 59198 346196 59434
rect 345876 52434 346196 59198
rect 345876 52198 345918 52434
rect 346154 52198 346196 52434
rect 345876 45434 346196 52198
rect 345876 45198 345918 45434
rect 346154 45198 346196 45434
rect 345876 38434 346196 45198
rect 345876 38198 345918 38434
rect 346154 38198 346196 38434
rect 345876 31434 346196 38198
rect 345876 31198 345918 31434
rect 346154 31198 346196 31434
rect 345876 24434 346196 31198
rect 345876 24198 345918 24434
rect 346154 24198 346196 24434
rect 345876 17434 346196 24198
rect 345876 17198 345918 17434
rect 346154 17198 346196 17434
rect 345876 10434 346196 17198
rect 345876 10198 345918 10434
rect 346154 10198 346196 10434
rect 345876 3434 346196 10198
rect 345876 3198 345918 3434
rect 346154 3198 346196 3434
rect 345876 -1706 346196 3198
rect 345876 -1942 345918 -1706
rect 346154 -1942 346196 -1706
rect 345876 -2026 346196 -1942
rect 345876 -2262 345918 -2026
rect 346154 -2262 346196 -2026
rect 345876 -2294 346196 -2262
rect 351144 705238 351464 706230
rect 351144 705002 351186 705238
rect 351422 705002 351464 705238
rect 351144 704918 351464 705002
rect 351144 704682 351186 704918
rect 351422 704682 351464 704918
rect 351144 695494 351464 704682
rect 351144 695258 351186 695494
rect 351422 695258 351464 695494
rect 351144 688494 351464 695258
rect 351144 688258 351186 688494
rect 351422 688258 351464 688494
rect 351144 681494 351464 688258
rect 351144 681258 351186 681494
rect 351422 681258 351464 681494
rect 351144 674494 351464 681258
rect 351144 674258 351186 674494
rect 351422 674258 351464 674494
rect 351144 667494 351464 674258
rect 351144 667258 351186 667494
rect 351422 667258 351464 667494
rect 351144 660494 351464 667258
rect 351144 660258 351186 660494
rect 351422 660258 351464 660494
rect 351144 653494 351464 660258
rect 351144 653258 351186 653494
rect 351422 653258 351464 653494
rect 351144 646494 351464 653258
rect 351144 646258 351186 646494
rect 351422 646258 351464 646494
rect 351144 639494 351464 646258
rect 351144 639258 351186 639494
rect 351422 639258 351464 639494
rect 351144 632494 351464 639258
rect 351144 632258 351186 632494
rect 351422 632258 351464 632494
rect 351144 625494 351464 632258
rect 351144 625258 351186 625494
rect 351422 625258 351464 625494
rect 351144 618494 351464 625258
rect 351144 618258 351186 618494
rect 351422 618258 351464 618494
rect 351144 611494 351464 618258
rect 351144 611258 351186 611494
rect 351422 611258 351464 611494
rect 351144 604494 351464 611258
rect 351144 604258 351186 604494
rect 351422 604258 351464 604494
rect 351144 597494 351464 604258
rect 351144 597258 351186 597494
rect 351422 597258 351464 597494
rect 351144 590494 351464 597258
rect 351144 590258 351186 590494
rect 351422 590258 351464 590494
rect 351144 583494 351464 590258
rect 351144 583258 351186 583494
rect 351422 583258 351464 583494
rect 351144 576494 351464 583258
rect 351144 576258 351186 576494
rect 351422 576258 351464 576494
rect 351144 569494 351464 576258
rect 351144 569258 351186 569494
rect 351422 569258 351464 569494
rect 351144 562494 351464 569258
rect 351144 562258 351186 562494
rect 351422 562258 351464 562494
rect 351144 555494 351464 562258
rect 351144 555258 351186 555494
rect 351422 555258 351464 555494
rect 351144 548494 351464 555258
rect 351144 548258 351186 548494
rect 351422 548258 351464 548494
rect 351144 541494 351464 548258
rect 351144 541258 351186 541494
rect 351422 541258 351464 541494
rect 351144 534494 351464 541258
rect 351144 534258 351186 534494
rect 351422 534258 351464 534494
rect 351144 527494 351464 534258
rect 351144 527258 351186 527494
rect 351422 527258 351464 527494
rect 351144 520494 351464 527258
rect 351144 520258 351186 520494
rect 351422 520258 351464 520494
rect 351144 513494 351464 520258
rect 351144 513258 351186 513494
rect 351422 513258 351464 513494
rect 351144 506494 351464 513258
rect 351144 506258 351186 506494
rect 351422 506258 351464 506494
rect 351144 499494 351464 506258
rect 351144 499258 351186 499494
rect 351422 499258 351464 499494
rect 351144 492494 351464 499258
rect 351144 492258 351186 492494
rect 351422 492258 351464 492494
rect 351144 485494 351464 492258
rect 351144 485258 351186 485494
rect 351422 485258 351464 485494
rect 351144 478494 351464 485258
rect 351144 478258 351186 478494
rect 351422 478258 351464 478494
rect 351144 471494 351464 478258
rect 351144 471258 351186 471494
rect 351422 471258 351464 471494
rect 351144 464494 351464 471258
rect 351144 464258 351186 464494
rect 351422 464258 351464 464494
rect 351144 457494 351464 464258
rect 351144 457258 351186 457494
rect 351422 457258 351464 457494
rect 351144 450494 351464 457258
rect 351144 450258 351186 450494
rect 351422 450258 351464 450494
rect 351144 443494 351464 450258
rect 351144 443258 351186 443494
rect 351422 443258 351464 443494
rect 351144 436494 351464 443258
rect 351144 436258 351186 436494
rect 351422 436258 351464 436494
rect 351144 429494 351464 436258
rect 351144 429258 351186 429494
rect 351422 429258 351464 429494
rect 351144 422494 351464 429258
rect 351144 422258 351186 422494
rect 351422 422258 351464 422494
rect 351144 415494 351464 422258
rect 351144 415258 351186 415494
rect 351422 415258 351464 415494
rect 351144 408494 351464 415258
rect 351144 408258 351186 408494
rect 351422 408258 351464 408494
rect 351144 401494 351464 408258
rect 351144 401258 351186 401494
rect 351422 401258 351464 401494
rect 351144 394494 351464 401258
rect 351144 394258 351186 394494
rect 351422 394258 351464 394494
rect 351144 387494 351464 394258
rect 351144 387258 351186 387494
rect 351422 387258 351464 387494
rect 351144 380494 351464 387258
rect 351144 380258 351186 380494
rect 351422 380258 351464 380494
rect 351144 373494 351464 380258
rect 351144 373258 351186 373494
rect 351422 373258 351464 373494
rect 351144 366494 351464 373258
rect 351144 366258 351186 366494
rect 351422 366258 351464 366494
rect 351144 359494 351464 366258
rect 351144 359258 351186 359494
rect 351422 359258 351464 359494
rect 351144 352494 351464 359258
rect 351144 352258 351186 352494
rect 351422 352258 351464 352494
rect 351144 345494 351464 352258
rect 351144 345258 351186 345494
rect 351422 345258 351464 345494
rect 351144 338494 351464 345258
rect 351144 338258 351186 338494
rect 351422 338258 351464 338494
rect 351144 331494 351464 338258
rect 351144 331258 351186 331494
rect 351422 331258 351464 331494
rect 351144 324494 351464 331258
rect 351144 324258 351186 324494
rect 351422 324258 351464 324494
rect 351144 317494 351464 324258
rect 351144 317258 351186 317494
rect 351422 317258 351464 317494
rect 351144 310494 351464 317258
rect 351144 310258 351186 310494
rect 351422 310258 351464 310494
rect 351144 303494 351464 310258
rect 351144 303258 351186 303494
rect 351422 303258 351464 303494
rect 351144 296494 351464 303258
rect 351144 296258 351186 296494
rect 351422 296258 351464 296494
rect 351144 289494 351464 296258
rect 351144 289258 351186 289494
rect 351422 289258 351464 289494
rect 351144 282494 351464 289258
rect 351144 282258 351186 282494
rect 351422 282258 351464 282494
rect 351144 275494 351464 282258
rect 351144 275258 351186 275494
rect 351422 275258 351464 275494
rect 351144 268494 351464 275258
rect 351144 268258 351186 268494
rect 351422 268258 351464 268494
rect 351144 261494 351464 268258
rect 351144 261258 351186 261494
rect 351422 261258 351464 261494
rect 351144 254494 351464 261258
rect 351144 254258 351186 254494
rect 351422 254258 351464 254494
rect 351144 247494 351464 254258
rect 351144 247258 351186 247494
rect 351422 247258 351464 247494
rect 351144 240494 351464 247258
rect 351144 240258 351186 240494
rect 351422 240258 351464 240494
rect 351144 233494 351464 240258
rect 351144 233258 351186 233494
rect 351422 233258 351464 233494
rect 351144 226494 351464 233258
rect 351144 226258 351186 226494
rect 351422 226258 351464 226494
rect 351144 219494 351464 226258
rect 351144 219258 351186 219494
rect 351422 219258 351464 219494
rect 351144 212494 351464 219258
rect 351144 212258 351186 212494
rect 351422 212258 351464 212494
rect 351144 205494 351464 212258
rect 351144 205258 351186 205494
rect 351422 205258 351464 205494
rect 351144 198494 351464 205258
rect 351144 198258 351186 198494
rect 351422 198258 351464 198494
rect 351144 191494 351464 198258
rect 351144 191258 351186 191494
rect 351422 191258 351464 191494
rect 351144 184494 351464 191258
rect 351144 184258 351186 184494
rect 351422 184258 351464 184494
rect 351144 177494 351464 184258
rect 351144 177258 351186 177494
rect 351422 177258 351464 177494
rect 351144 170494 351464 177258
rect 351144 170258 351186 170494
rect 351422 170258 351464 170494
rect 351144 163494 351464 170258
rect 351144 163258 351186 163494
rect 351422 163258 351464 163494
rect 351144 156494 351464 163258
rect 351144 156258 351186 156494
rect 351422 156258 351464 156494
rect 351144 149494 351464 156258
rect 351144 149258 351186 149494
rect 351422 149258 351464 149494
rect 351144 142494 351464 149258
rect 351144 142258 351186 142494
rect 351422 142258 351464 142494
rect 351144 135494 351464 142258
rect 351144 135258 351186 135494
rect 351422 135258 351464 135494
rect 351144 128494 351464 135258
rect 351144 128258 351186 128494
rect 351422 128258 351464 128494
rect 351144 121494 351464 128258
rect 351144 121258 351186 121494
rect 351422 121258 351464 121494
rect 351144 114494 351464 121258
rect 351144 114258 351186 114494
rect 351422 114258 351464 114494
rect 351144 107494 351464 114258
rect 351144 107258 351186 107494
rect 351422 107258 351464 107494
rect 351144 100494 351464 107258
rect 351144 100258 351186 100494
rect 351422 100258 351464 100494
rect 351144 93494 351464 100258
rect 351144 93258 351186 93494
rect 351422 93258 351464 93494
rect 351144 86494 351464 93258
rect 351144 86258 351186 86494
rect 351422 86258 351464 86494
rect 351144 79494 351464 86258
rect 351144 79258 351186 79494
rect 351422 79258 351464 79494
rect 351144 72494 351464 79258
rect 351144 72258 351186 72494
rect 351422 72258 351464 72494
rect 351144 65494 351464 72258
rect 351144 65258 351186 65494
rect 351422 65258 351464 65494
rect 351144 58494 351464 65258
rect 351144 58258 351186 58494
rect 351422 58258 351464 58494
rect 351144 51494 351464 58258
rect 351144 51258 351186 51494
rect 351422 51258 351464 51494
rect 351144 44494 351464 51258
rect 351144 44258 351186 44494
rect 351422 44258 351464 44494
rect 351144 37494 351464 44258
rect 351144 37258 351186 37494
rect 351422 37258 351464 37494
rect 351144 30494 351464 37258
rect 351144 30258 351186 30494
rect 351422 30258 351464 30494
rect 351144 23494 351464 30258
rect 351144 23258 351186 23494
rect 351422 23258 351464 23494
rect 351144 16494 351464 23258
rect 351144 16258 351186 16494
rect 351422 16258 351464 16494
rect 351144 9494 351464 16258
rect 351144 9258 351186 9494
rect 351422 9258 351464 9494
rect 351144 2494 351464 9258
rect 351144 2258 351186 2494
rect 351422 2258 351464 2494
rect 351144 -746 351464 2258
rect 351144 -982 351186 -746
rect 351422 -982 351464 -746
rect 351144 -1066 351464 -982
rect 351144 -1302 351186 -1066
rect 351422 -1302 351464 -1066
rect 351144 -2294 351464 -1302
rect 352876 706198 353196 706230
rect 352876 705962 352918 706198
rect 353154 705962 353196 706198
rect 352876 705878 353196 705962
rect 352876 705642 352918 705878
rect 353154 705642 353196 705878
rect 352876 696434 353196 705642
rect 352876 696198 352918 696434
rect 353154 696198 353196 696434
rect 352876 689434 353196 696198
rect 352876 689198 352918 689434
rect 353154 689198 353196 689434
rect 352876 682434 353196 689198
rect 352876 682198 352918 682434
rect 353154 682198 353196 682434
rect 352876 675434 353196 682198
rect 352876 675198 352918 675434
rect 353154 675198 353196 675434
rect 352876 668434 353196 675198
rect 352876 668198 352918 668434
rect 353154 668198 353196 668434
rect 352876 661434 353196 668198
rect 352876 661198 352918 661434
rect 353154 661198 353196 661434
rect 352876 654434 353196 661198
rect 352876 654198 352918 654434
rect 353154 654198 353196 654434
rect 352876 647434 353196 654198
rect 352876 647198 352918 647434
rect 353154 647198 353196 647434
rect 352876 640434 353196 647198
rect 352876 640198 352918 640434
rect 353154 640198 353196 640434
rect 352876 633434 353196 640198
rect 352876 633198 352918 633434
rect 353154 633198 353196 633434
rect 352876 626434 353196 633198
rect 352876 626198 352918 626434
rect 353154 626198 353196 626434
rect 352876 619434 353196 626198
rect 352876 619198 352918 619434
rect 353154 619198 353196 619434
rect 352876 612434 353196 619198
rect 352876 612198 352918 612434
rect 353154 612198 353196 612434
rect 352876 605434 353196 612198
rect 352876 605198 352918 605434
rect 353154 605198 353196 605434
rect 352876 598434 353196 605198
rect 352876 598198 352918 598434
rect 353154 598198 353196 598434
rect 352876 591434 353196 598198
rect 352876 591198 352918 591434
rect 353154 591198 353196 591434
rect 352876 584434 353196 591198
rect 352876 584198 352918 584434
rect 353154 584198 353196 584434
rect 352876 577434 353196 584198
rect 352876 577198 352918 577434
rect 353154 577198 353196 577434
rect 352876 570434 353196 577198
rect 352876 570198 352918 570434
rect 353154 570198 353196 570434
rect 352876 563434 353196 570198
rect 352876 563198 352918 563434
rect 353154 563198 353196 563434
rect 352876 556434 353196 563198
rect 352876 556198 352918 556434
rect 353154 556198 353196 556434
rect 352876 549434 353196 556198
rect 352876 549198 352918 549434
rect 353154 549198 353196 549434
rect 352876 542434 353196 549198
rect 352876 542198 352918 542434
rect 353154 542198 353196 542434
rect 352876 535434 353196 542198
rect 352876 535198 352918 535434
rect 353154 535198 353196 535434
rect 352876 528434 353196 535198
rect 352876 528198 352918 528434
rect 353154 528198 353196 528434
rect 352876 521434 353196 528198
rect 352876 521198 352918 521434
rect 353154 521198 353196 521434
rect 352876 514434 353196 521198
rect 352876 514198 352918 514434
rect 353154 514198 353196 514434
rect 352876 507434 353196 514198
rect 352876 507198 352918 507434
rect 353154 507198 353196 507434
rect 352876 500434 353196 507198
rect 352876 500198 352918 500434
rect 353154 500198 353196 500434
rect 352876 493434 353196 500198
rect 352876 493198 352918 493434
rect 353154 493198 353196 493434
rect 352876 486434 353196 493198
rect 352876 486198 352918 486434
rect 353154 486198 353196 486434
rect 352876 479434 353196 486198
rect 352876 479198 352918 479434
rect 353154 479198 353196 479434
rect 352876 472434 353196 479198
rect 352876 472198 352918 472434
rect 353154 472198 353196 472434
rect 352876 465434 353196 472198
rect 352876 465198 352918 465434
rect 353154 465198 353196 465434
rect 352876 458434 353196 465198
rect 352876 458198 352918 458434
rect 353154 458198 353196 458434
rect 352876 451434 353196 458198
rect 352876 451198 352918 451434
rect 353154 451198 353196 451434
rect 352876 444434 353196 451198
rect 352876 444198 352918 444434
rect 353154 444198 353196 444434
rect 352876 437434 353196 444198
rect 352876 437198 352918 437434
rect 353154 437198 353196 437434
rect 352876 430434 353196 437198
rect 352876 430198 352918 430434
rect 353154 430198 353196 430434
rect 352876 423434 353196 430198
rect 352876 423198 352918 423434
rect 353154 423198 353196 423434
rect 352876 416434 353196 423198
rect 352876 416198 352918 416434
rect 353154 416198 353196 416434
rect 352876 409434 353196 416198
rect 352876 409198 352918 409434
rect 353154 409198 353196 409434
rect 352876 402434 353196 409198
rect 352876 402198 352918 402434
rect 353154 402198 353196 402434
rect 352876 395434 353196 402198
rect 352876 395198 352918 395434
rect 353154 395198 353196 395434
rect 352876 388434 353196 395198
rect 352876 388198 352918 388434
rect 353154 388198 353196 388434
rect 352876 381434 353196 388198
rect 352876 381198 352918 381434
rect 353154 381198 353196 381434
rect 352876 374434 353196 381198
rect 352876 374198 352918 374434
rect 353154 374198 353196 374434
rect 352876 367434 353196 374198
rect 352876 367198 352918 367434
rect 353154 367198 353196 367434
rect 352876 360434 353196 367198
rect 352876 360198 352918 360434
rect 353154 360198 353196 360434
rect 352876 353434 353196 360198
rect 352876 353198 352918 353434
rect 353154 353198 353196 353434
rect 352876 346434 353196 353198
rect 352876 346198 352918 346434
rect 353154 346198 353196 346434
rect 352876 339434 353196 346198
rect 352876 339198 352918 339434
rect 353154 339198 353196 339434
rect 352876 332434 353196 339198
rect 352876 332198 352918 332434
rect 353154 332198 353196 332434
rect 352876 325434 353196 332198
rect 352876 325198 352918 325434
rect 353154 325198 353196 325434
rect 352876 318434 353196 325198
rect 352876 318198 352918 318434
rect 353154 318198 353196 318434
rect 352876 311434 353196 318198
rect 352876 311198 352918 311434
rect 353154 311198 353196 311434
rect 352876 304434 353196 311198
rect 352876 304198 352918 304434
rect 353154 304198 353196 304434
rect 352876 297434 353196 304198
rect 352876 297198 352918 297434
rect 353154 297198 353196 297434
rect 352876 290434 353196 297198
rect 352876 290198 352918 290434
rect 353154 290198 353196 290434
rect 352876 283434 353196 290198
rect 352876 283198 352918 283434
rect 353154 283198 353196 283434
rect 352876 276434 353196 283198
rect 352876 276198 352918 276434
rect 353154 276198 353196 276434
rect 352876 269434 353196 276198
rect 352876 269198 352918 269434
rect 353154 269198 353196 269434
rect 352876 262434 353196 269198
rect 352876 262198 352918 262434
rect 353154 262198 353196 262434
rect 352876 255434 353196 262198
rect 352876 255198 352918 255434
rect 353154 255198 353196 255434
rect 352876 248434 353196 255198
rect 352876 248198 352918 248434
rect 353154 248198 353196 248434
rect 352876 241434 353196 248198
rect 352876 241198 352918 241434
rect 353154 241198 353196 241434
rect 352876 234434 353196 241198
rect 352876 234198 352918 234434
rect 353154 234198 353196 234434
rect 352876 227434 353196 234198
rect 352876 227198 352918 227434
rect 353154 227198 353196 227434
rect 352876 220434 353196 227198
rect 352876 220198 352918 220434
rect 353154 220198 353196 220434
rect 352876 213434 353196 220198
rect 352876 213198 352918 213434
rect 353154 213198 353196 213434
rect 352876 206434 353196 213198
rect 352876 206198 352918 206434
rect 353154 206198 353196 206434
rect 352876 199434 353196 206198
rect 352876 199198 352918 199434
rect 353154 199198 353196 199434
rect 352876 192434 353196 199198
rect 352876 192198 352918 192434
rect 353154 192198 353196 192434
rect 352876 185434 353196 192198
rect 352876 185198 352918 185434
rect 353154 185198 353196 185434
rect 352876 178434 353196 185198
rect 352876 178198 352918 178434
rect 353154 178198 353196 178434
rect 352876 171434 353196 178198
rect 352876 171198 352918 171434
rect 353154 171198 353196 171434
rect 352876 164434 353196 171198
rect 352876 164198 352918 164434
rect 353154 164198 353196 164434
rect 352876 157434 353196 164198
rect 352876 157198 352918 157434
rect 353154 157198 353196 157434
rect 352876 150434 353196 157198
rect 352876 150198 352918 150434
rect 353154 150198 353196 150434
rect 352876 143434 353196 150198
rect 352876 143198 352918 143434
rect 353154 143198 353196 143434
rect 352876 136434 353196 143198
rect 352876 136198 352918 136434
rect 353154 136198 353196 136434
rect 352876 129434 353196 136198
rect 352876 129198 352918 129434
rect 353154 129198 353196 129434
rect 352876 122434 353196 129198
rect 352876 122198 352918 122434
rect 353154 122198 353196 122434
rect 352876 115434 353196 122198
rect 352876 115198 352918 115434
rect 353154 115198 353196 115434
rect 352876 108434 353196 115198
rect 352876 108198 352918 108434
rect 353154 108198 353196 108434
rect 352876 101434 353196 108198
rect 352876 101198 352918 101434
rect 353154 101198 353196 101434
rect 352876 94434 353196 101198
rect 352876 94198 352918 94434
rect 353154 94198 353196 94434
rect 352876 87434 353196 94198
rect 352876 87198 352918 87434
rect 353154 87198 353196 87434
rect 352876 80434 353196 87198
rect 352876 80198 352918 80434
rect 353154 80198 353196 80434
rect 352876 73434 353196 80198
rect 352876 73198 352918 73434
rect 353154 73198 353196 73434
rect 352876 66434 353196 73198
rect 352876 66198 352918 66434
rect 353154 66198 353196 66434
rect 352876 59434 353196 66198
rect 352876 59198 352918 59434
rect 353154 59198 353196 59434
rect 352876 52434 353196 59198
rect 352876 52198 352918 52434
rect 353154 52198 353196 52434
rect 352876 45434 353196 52198
rect 352876 45198 352918 45434
rect 353154 45198 353196 45434
rect 352876 38434 353196 45198
rect 352876 38198 352918 38434
rect 353154 38198 353196 38434
rect 352876 31434 353196 38198
rect 352876 31198 352918 31434
rect 353154 31198 353196 31434
rect 352876 24434 353196 31198
rect 352876 24198 352918 24434
rect 353154 24198 353196 24434
rect 352876 17434 353196 24198
rect 352876 17198 352918 17434
rect 353154 17198 353196 17434
rect 352876 10434 353196 17198
rect 352876 10198 352918 10434
rect 353154 10198 353196 10434
rect 352876 3434 353196 10198
rect 352876 3198 352918 3434
rect 353154 3198 353196 3434
rect 352876 -1706 353196 3198
rect 352876 -1942 352918 -1706
rect 353154 -1942 353196 -1706
rect 352876 -2026 353196 -1942
rect 352876 -2262 352918 -2026
rect 353154 -2262 353196 -2026
rect 352876 -2294 353196 -2262
rect 358144 705238 358464 706230
rect 358144 705002 358186 705238
rect 358422 705002 358464 705238
rect 358144 704918 358464 705002
rect 358144 704682 358186 704918
rect 358422 704682 358464 704918
rect 358144 695494 358464 704682
rect 358144 695258 358186 695494
rect 358422 695258 358464 695494
rect 358144 688494 358464 695258
rect 358144 688258 358186 688494
rect 358422 688258 358464 688494
rect 358144 681494 358464 688258
rect 358144 681258 358186 681494
rect 358422 681258 358464 681494
rect 358144 674494 358464 681258
rect 358144 674258 358186 674494
rect 358422 674258 358464 674494
rect 358144 667494 358464 674258
rect 358144 667258 358186 667494
rect 358422 667258 358464 667494
rect 358144 660494 358464 667258
rect 358144 660258 358186 660494
rect 358422 660258 358464 660494
rect 358144 653494 358464 660258
rect 358144 653258 358186 653494
rect 358422 653258 358464 653494
rect 358144 646494 358464 653258
rect 358144 646258 358186 646494
rect 358422 646258 358464 646494
rect 358144 639494 358464 646258
rect 358144 639258 358186 639494
rect 358422 639258 358464 639494
rect 358144 632494 358464 639258
rect 358144 632258 358186 632494
rect 358422 632258 358464 632494
rect 358144 625494 358464 632258
rect 358144 625258 358186 625494
rect 358422 625258 358464 625494
rect 358144 618494 358464 625258
rect 358144 618258 358186 618494
rect 358422 618258 358464 618494
rect 358144 611494 358464 618258
rect 358144 611258 358186 611494
rect 358422 611258 358464 611494
rect 358144 604494 358464 611258
rect 358144 604258 358186 604494
rect 358422 604258 358464 604494
rect 358144 597494 358464 604258
rect 358144 597258 358186 597494
rect 358422 597258 358464 597494
rect 358144 590494 358464 597258
rect 358144 590258 358186 590494
rect 358422 590258 358464 590494
rect 358144 583494 358464 590258
rect 358144 583258 358186 583494
rect 358422 583258 358464 583494
rect 358144 576494 358464 583258
rect 358144 576258 358186 576494
rect 358422 576258 358464 576494
rect 358144 569494 358464 576258
rect 358144 569258 358186 569494
rect 358422 569258 358464 569494
rect 358144 562494 358464 569258
rect 358144 562258 358186 562494
rect 358422 562258 358464 562494
rect 358144 555494 358464 562258
rect 358144 555258 358186 555494
rect 358422 555258 358464 555494
rect 358144 548494 358464 555258
rect 358144 548258 358186 548494
rect 358422 548258 358464 548494
rect 358144 541494 358464 548258
rect 358144 541258 358186 541494
rect 358422 541258 358464 541494
rect 358144 534494 358464 541258
rect 358144 534258 358186 534494
rect 358422 534258 358464 534494
rect 358144 527494 358464 534258
rect 358144 527258 358186 527494
rect 358422 527258 358464 527494
rect 358144 520494 358464 527258
rect 358144 520258 358186 520494
rect 358422 520258 358464 520494
rect 358144 513494 358464 520258
rect 358144 513258 358186 513494
rect 358422 513258 358464 513494
rect 358144 506494 358464 513258
rect 358144 506258 358186 506494
rect 358422 506258 358464 506494
rect 358144 499494 358464 506258
rect 358144 499258 358186 499494
rect 358422 499258 358464 499494
rect 358144 492494 358464 499258
rect 358144 492258 358186 492494
rect 358422 492258 358464 492494
rect 358144 485494 358464 492258
rect 358144 485258 358186 485494
rect 358422 485258 358464 485494
rect 358144 478494 358464 485258
rect 358144 478258 358186 478494
rect 358422 478258 358464 478494
rect 358144 471494 358464 478258
rect 358144 471258 358186 471494
rect 358422 471258 358464 471494
rect 358144 464494 358464 471258
rect 358144 464258 358186 464494
rect 358422 464258 358464 464494
rect 358144 457494 358464 464258
rect 358144 457258 358186 457494
rect 358422 457258 358464 457494
rect 358144 450494 358464 457258
rect 358144 450258 358186 450494
rect 358422 450258 358464 450494
rect 358144 443494 358464 450258
rect 358144 443258 358186 443494
rect 358422 443258 358464 443494
rect 358144 436494 358464 443258
rect 358144 436258 358186 436494
rect 358422 436258 358464 436494
rect 358144 429494 358464 436258
rect 358144 429258 358186 429494
rect 358422 429258 358464 429494
rect 358144 422494 358464 429258
rect 358144 422258 358186 422494
rect 358422 422258 358464 422494
rect 358144 415494 358464 422258
rect 358144 415258 358186 415494
rect 358422 415258 358464 415494
rect 358144 408494 358464 415258
rect 358144 408258 358186 408494
rect 358422 408258 358464 408494
rect 358144 401494 358464 408258
rect 358144 401258 358186 401494
rect 358422 401258 358464 401494
rect 358144 394494 358464 401258
rect 358144 394258 358186 394494
rect 358422 394258 358464 394494
rect 358144 387494 358464 394258
rect 358144 387258 358186 387494
rect 358422 387258 358464 387494
rect 358144 380494 358464 387258
rect 358144 380258 358186 380494
rect 358422 380258 358464 380494
rect 358144 373494 358464 380258
rect 358144 373258 358186 373494
rect 358422 373258 358464 373494
rect 358144 366494 358464 373258
rect 358144 366258 358186 366494
rect 358422 366258 358464 366494
rect 358144 359494 358464 366258
rect 358144 359258 358186 359494
rect 358422 359258 358464 359494
rect 358144 352494 358464 359258
rect 358144 352258 358186 352494
rect 358422 352258 358464 352494
rect 358144 345494 358464 352258
rect 358144 345258 358186 345494
rect 358422 345258 358464 345494
rect 358144 338494 358464 345258
rect 358144 338258 358186 338494
rect 358422 338258 358464 338494
rect 358144 331494 358464 338258
rect 358144 331258 358186 331494
rect 358422 331258 358464 331494
rect 358144 324494 358464 331258
rect 358144 324258 358186 324494
rect 358422 324258 358464 324494
rect 358144 317494 358464 324258
rect 358144 317258 358186 317494
rect 358422 317258 358464 317494
rect 358144 310494 358464 317258
rect 358144 310258 358186 310494
rect 358422 310258 358464 310494
rect 358144 303494 358464 310258
rect 358144 303258 358186 303494
rect 358422 303258 358464 303494
rect 358144 296494 358464 303258
rect 358144 296258 358186 296494
rect 358422 296258 358464 296494
rect 358144 289494 358464 296258
rect 358144 289258 358186 289494
rect 358422 289258 358464 289494
rect 358144 282494 358464 289258
rect 358144 282258 358186 282494
rect 358422 282258 358464 282494
rect 358144 275494 358464 282258
rect 358144 275258 358186 275494
rect 358422 275258 358464 275494
rect 358144 268494 358464 275258
rect 358144 268258 358186 268494
rect 358422 268258 358464 268494
rect 358144 261494 358464 268258
rect 358144 261258 358186 261494
rect 358422 261258 358464 261494
rect 358144 254494 358464 261258
rect 358144 254258 358186 254494
rect 358422 254258 358464 254494
rect 358144 247494 358464 254258
rect 358144 247258 358186 247494
rect 358422 247258 358464 247494
rect 358144 240494 358464 247258
rect 358144 240258 358186 240494
rect 358422 240258 358464 240494
rect 358144 233494 358464 240258
rect 358144 233258 358186 233494
rect 358422 233258 358464 233494
rect 358144 226494 358464 233258
rect 358144 226258 358186 226494
rect 358422 226258 358464 226494
rect 358144 219494 358464 226258
rect 358144 219258 358186 219494
rect 358422 219258 358464 219494
rect 358144 212494 358464 219258
rect 358144 212258 358186 212494
rect 358422 212258 358464 212494
rect 358144 205494 358464 212258
rect 358144 205258 358186 205494
rect 358422 205258 358464 205494
rect 358144 198494 358464 205258
rect 358144 198258 358186 198494
rect 358422 198258 358464 198494
rect 358144 191494 358464 198258
rect 358144 191258 358186 191494
rect 358422 191258 358464 191494
rect 358144 184494 358464 191258
rect 358144 184258 358186 184494
rect 358422 184258 358464 184494
rect 358144 177494 358464 184258
rect 358144 177258 358186 177494
rect 358422 177258 358464 177494
rect 358144 170494 358464 177258
rect 358144 170258 358186 170494
rect 358422 170258 358464 170494
rect 358144 163494 358464 170258
rect 358144 163258 358186 163494
rect 358422 163258 358464 163494
rect 358144 156494 358464 163258
rect 358144 156258 358186 156494
rect 358422 156258 358464 156494
rect 358144 149494 358464 156258
rect 358144 149258 358186 149494
rect 358422 149258 358464 149494
rect 358144 142494 358464 149258
rect 358144 142258 358186 142494
rect 358422 142258 358464 142494
rect 358144 135494 358464 142258
rect 358144 135258 358186 135494
rect 358422 135258 358464 135494
rect 358144 128494 358464 135258
rect 358144 128258 358186 128494
rect 358422 128258 358464 128494
rect 358144 121494 358464 128258
rect 358144 121258 358186 121494
rect 358422 121258 358464 121494
rect 358144 114494 358464 121258
rect 358144 114258 358186 114494
rect 358422 114258 358464 114494
rect 358144 107494 358464 114258
rect 358144 107258 358186 107494
rect 358422 107258 358464 107494
rect 358144 100494 358464 107258
rect 358144 100258 358186 100494
rect 358422 100258 358464 100494
rect 358144 93494 358464 100258
rect 358144 93258 358186 93494
rect 358422 93258 358464 93494
rect 358144 86494 358464 93258
rect 358144 86258 358186 86494
rect 358422 86258 358464 86494
rect 358144 79494 358464 86258
rect 358144 79258 358186 79494
rect 358422 79258 358464 79494
rect 358144 72494 358464 79258
rect 358144 72258 358186 72494
rect 358422 72258 358464 72494
rect 358144 65494 358464 72258
rect 358144 65258 358186 65494
rect 358422 65258 358464 65494
rect 358144 58494 358464 65258
rect 358144 58258 358186 58494
rect 358422 58258 358464 58494
rect 358144 51494 358464 58258
rect 358144 51258 358186 51494
rect 358422 51258 358464 51494
rect 358144 44494 358464 51258
rect 358144 44258 358186 44494
rect 358422 44258 358464 44494
rect 358144 37494 358464 44258
rect 358144 37258 358186 37494
rect 358422 37258 358464 37494
rect 358144 30494 358464 37258
rect 358144 30258 358186 30494
rect 358422 30258 358464 30494
rect 358144 23494 358464 30258
rect 358144 23258 358186 23494
rect 358422 23258 358464 23494
rect 358144 16494 358464 23258
rect 358144 16258 358186 16494
rect 358422 16258 358464 16494
rect 358144 9494 358464 16258
rect 358144 9258 358186 9494
rect 358422 9258 358464 9494
rect 358144 2494 358464 9258
rect 358144 2258 358186 2494
rect 358422 2258 358464 2494
rect 358144 -746 358464 2258
rect 358144 -982 358186 -746
rect 358422 -982 358464 -746
rect 358144 -1066 358464 -982
rect 358144 -1302 358186 -1066
rect 358422 -1302 358464 -1066
rect 358144 -2294 358464 -1302
rect 359876 706198 360196 706230
rect 359876 705962 359918 706198
rect 360154 705962 360196 706198
rect 359876 705878 360196 705962
rect 359876 705642 359918 705878
rect 360154 705642 360196 705878
rect 359876 696434 360196 705642
rect 359876 696198 359918 696434
rect 360154 696198 360196 696434
rect 359876 689434 360196 696198
rect 359876 689198 359918 689434
rect 360154 689198 360196 689434
rect 359876 682434 360196 689198
rect 359876 682198 359918 682434
rect 360154 682198 360196 682434
rect 359876 675434 360196 682198
rect 359876 675198 359918 675434
rect 360154 675198 360196 675434
rect 359876 668434 360196 675198
rect 359876 668198 359918 668434
rect 360154 668198 360196 668434
rect 359876 661434 360196 668198
rect 359876 661198 359918 661434
rect 360154 661198 360196 661434
rect 359876 654434 360196 661198
rect 359876 654198 359918 654434
rect 360154 654198 360196 654434
rect 359876 647434 360196 654198
rect 359876 647198 359918 647434
rect 360154 647198 360196 647434
rect 359876 640434 360196 647198
rect 359876 640198 359918 640434
rect 360154 640198 360196 640434
rect 359876 633434 360196 640198
rect 359876 633198 359918 633434
rect 360154 633198 360196 633434
rect 359876 626434 360196 633198
rect 359876 626198 359918 626434
rect 360154 626198 360196 626434
rect 359876 619434 360196 626198
rect 359876 619198 359918 619434
rect 360154 619198 360196 619434
rect 359876 612434 360196 619198
rect 359876 612198 359918 612434
rect 360154 612198 360196 612434
rect 359876 605434 360196 612198
rect 359876 605198 359918 605434
rect 360154 605198 360196 605434
rect 359876 598434 360196 605198
rect 359876 598198 359918 598434
rect 360154 598198 360196 598434
rect 359876 591434 360196 598198
rect 359876 591198 359918 591434
rect 360154 591198 360196 591434
rect 359876 584434 360196 591198
rect 359876 584198 359918 584434
rect 360154 584198 360196 584434
rect 359876 577434 360196 584198
rect 359876 577198 359918 577434
rect 360154 577198 360196 577434
rect 359876 570434 360196 577198
rect 359876 570198 359918 570434
rect 360154 570198 360196 570434
rect 359876 563434 360196 570198
rect 359876 563198 359918 563434
rect 360154 563198 360196 563434
rect 359876 556434 360196 563198
rect 359876 556198 359918 556434
rect 360154 556198 360196 556434
rect 359876 549434 360196 556198
rect 359876 549198 359918 549434
rect 360154 549198 360196 549434
rect 359876 542434 360196 549198
rect 359876 542198 359918 542434
rect 360154 542198 360196 542434
rect 359876 535434 360196 542198
rect 359876 535198 359918 535434
rect 360154 535198 360196 535434
rect 359876 528434 360196 535198
rect 359876 528198 359918 528434
rect 360154 528198 360196 528434
rect 359876 521434 360196 528198
rect 359876 521198 359918 521434
rect 360154 521198 360196 521434
rect 359876 514434 360196 521198
rect 359876 514198 359918 514434
rect 360154 514198 360196 514434
rect 359876 507434 360196 514198
rect 359876 507198 359918 507434
rect 360154 507198 360196 507434
rect 359876 500434 360196 507198
rect 359876 500198 359918 500434
rect 360154 500198 360196 500434
rect 359876 493434 360196 500198
rect 359876 493198 359918 493434
rect 360154 493198 360196 493434
rect 359876 486434 360196 493198
rect 359876 486198 359918 486434
rect 360154 486198 360196 486434
rect 359876 479434 360196 486198
rect 359876 479198 359918 479434
rect 360154 479198 360196 479434
rect 359876 472434 360196 479198
rect 359876 472198 359918 472434
rect 360154 472198 360196 472434
rect 359876 465434 360196 472198
rect 359876 465198 359918 465434
rect 360154 465198 360196 465434
rect 359876 458434 360196 465198
rect 359876 458198 359918 458434
rect 360154 458198 360196 458434
rect 359876 451434 360196 458198
rect 359876 451198 359918 451434
rect 360154 451198 360196 451434
rect 359876 444434 360196 451198
rect 359876 444198 359918 444434
rect 360154 444198 360196 444434
rect 359876 437434 360196 444198
rect 359876 437198 359918 437434
rect 360154 437198 360196 437434
rect 359876 430434 360196 437198
rect 359876 430198 359918 430434
rect 360154 430198 360196 430434
rect 359876 423434 360196 430198
rect 359876 423198 359918 423434
rect 360154 423198 360196 423434
rect 359876 416434 360196 423198
rect 359876 416198 359918 416434
rect 360154 416198 360196 416434
rect 359876 409434 360196 416198
rect 359876 409198 359918 409434
rect 360154 409198 360196 409434
rect 359876 402434 360196 409198
rect 359876 402198 359918 402434
rect 360154 402198 360196 402434
rect 359876 395434 360196 402198
rect 359876 395198 359918 395434
rect 360154 395198 360196 395434
rect 359876 388434 360196 395198
rect 359876 388198 359918 388434
rect 360154 388198 360196 388434
rect 359876 381434 360196 388198
rect 359876 381198 359918 381434
rect 360154 381198 360196 381434
rect 359876 374434 360196 381198
rect 359876 374198 359918 374434
rect 360154 374198 360196 374434
rect 359876 367434 360196 374198
rect 359876 367198 359918 367434
rect 360154 367198 360196 367434
rect 359876 360434 360196 367198
rect 359876 360198 359918 360434
rect 360154 360198 360196 360434
rect 359876 353434 360196 360198
rect 359876 353198 359918 353434
rect 360154 353198 360196 353434
rect 359876 346434 360196 353198
rect 359876 346198 359918 346434
rect 360154 346198 360196 346434
rect 359876 339434 360196 346198
rect 359876 339198 359918 339434
rect 360154 339198 360196 339434
rect 359876 332434 360196 339198
rect 359876 332198 359918 332434
rect 360154 332198 360196 332434
rect 359876 325434 360196 332198
rect 359876 325198 359918 325434
rect 360154 325198 360196 325434
rect 359876 318434 360196 325198
rect 359876 318198 359918 318434
rect 360154 318198 360196 318434
rect 359876 311434 360196 318198
rect 359876 311198 359918 311434
rect 360154 311198 360196 311434
rect 359876 304434 360196 311198
rect 359876 304198 359918 304434
rect 360154 304198 360196 304434
rect 359876 297434 360196 304198
rect 359876 297198 359918 297434
rect 360154 297198 360196 297434
rect 359876 290434 360196 297198
rect 359876 290198 359918 290434
rect 360154 290198 360196 290434
rect 359876 283434 360196 290198
rect 359876 283198 359918 283434
rect 360154 283198 360196 283434
rect 359876 276434 360196 283198
rect 359876 276198 359918 276434
rect 360154 276198 360196 276434
rect 359876 269434 360196 276198
rect 359876 269198 359918 269434
rect 360154 269198 360196 269434
rect 359876 262434 360196 269198
rect 359876 262198 359918 262434
rect 360154 262198 360196 262434
rect 359876 255434 360196 262198
rect 359876 255198 359918 255434
rect 360154 255198 360196 255434
rect 359876 248434 360196 255198
rect 359876 248198 359918 248434
rect 360154 248198 360196 248434
rect 359876 241434 360196 248198
rect 359876 241198 359918 241434
rect 360154 241198 360196 241434
rect 359876 234434 360196 241198
rect 359876 234198 359918 234434
rect 360154 234198 360196 234434
rect 359876 227434 360196 234198
rect 359876 227198 359918 227434
rect 360154 227198 360196 227434
rect 359876 220434 360196 227198
rect 359876 220198 359918 220434
rect 360154 220198 360196 220434
rect 359876 213434 360196 220198
rect 359876 213198 359918 213434
rect 360154 213198 360196 213434
rect 359876 206434 360196 213198
rect 359876 206198 359918 206434
rect 360154 206198 360196 206434
rect 359876 199434 360196 206198
rect 359876 199198 359918 199434
rect 360154 199198 360196 199434
rect 359876 192434 360196 199198
rect 359876 192198 359918 192434
rect 360154 192198 360196 192434
rect 359876 185434 360196 192198
rect 359876 185198 359918 185434
rect 360154 185198 360196 185434
rect 359876 178434 360196 185198
rect 359876 178198 359918 178434
rect 360154 178198 360196 178434
rect 359876 171434 360196 178198
rect 359876 171198 359918 171434
rect 360154 171198 360196 171434
rect 359876 164434 360196 171198
rect 359876 164198 359918 164434
rect 360154 164198 360196 164434
rect 359876 157434 360196 164198
rect 359876 157198 359918 157434
rect 360154 157198 360196 157434
rect 359876 150434 360196 157198
rect 359876 150198 359918 150434
rect 360154 150198 360196 150434
rect 359876 143434 360196 150198
rect 359876 143198 359918 143434
rect 360154 143198 360196 143434
rect 359876 136434 360196 143198
rect 359876 136198 359918 136434
rect 360154 136198 360196 136434
rect 359876 129434 360196 136198
rect 359876 129198 359918 129434
rect 360154 129198 360196 129434
rect 359876 122434 360196 129198
rect 359876 122198 359918 122434
rect 360154 122198 360196 122434
rect 359876 115434 360196 122198
rect 359876 115198 359918 115434
rect 360154 115198 360196 115434
rect 359876 108434 360196 115198
rect 359876 108198 359918 108434
rect 360154 108198 360196 108434
rect 359876 101434 360196 108198
rect 359876 101198 359918 101434
rect 360154 101198 360196 101434
rect 359876 94434 360196 101198
rect 359876 94198 359918 94434
rect 360154 94198 360196 94434
rect 359876 87434 360196 94198
rect 359876 87198 359918 87434
rect 360154 87198 360196 87434
rect 359876 80434 360196 87198
rect 359876 80198 359918 80434
rect 360154 80198 360196 80434
rect 359876 73434 360196 80198
rect 359876 73198 359918 73434
rect 360154 73198 360196 73434
rect 359876 66434 360196 73198
rect 359876 66198 359918 66434
rect 360154 66198 360196 66434
rect 359876 59434 360196 66198
rect 359876 59198 359918 59434
rect 360154 59198 360196 59434
rect 359876 52434 360196 59198
rect 359876 52198 359918 52434
rect 360154 52198 360196 52434
rect 359876 45434 360196 52198
rect 359876 45198 359918 45434
rect 360154 45198 360196 45434
rect 359876 38434 360196 45198
rect 359876 38198 359918 38434
rect 360154 38198 360196 38434
rect 359876 31434 360196 38198
rect 359876 31198 359918 31434
rect 360154 31198 360196 31434
rect 359876 24434 360196 31198
rect 359876 24198 359918 24434
rect 360154 24198 360196 24434
rect 359876 17434 360196 24198
rect 359876 17198 359918 17434
rect 360154 17198 360196 17434
rect 359876 10434 360196 17198
rect 359876 10198 359918 10434
rect 360154 10198 360196 10434
rect 359876 3434 360196 10198
rect 359876 3198 359918 3434
rect 360154 3198 360196 3434
rect 359876 -1706 360196 3198
rect 359876 -1942 359918 -1706
rect 360154 -1942 360196 -1706
rect 359876 -2026 360196 -1942
rect 359876 -2262 359918 -2026
rect 360154 -2262 360196 -2026
rect 359876 -2294 360196 -2262
rect 365144 705238 365464 706230
rect 365144 705002 365186 705238
rect 365422 705002 365464 705238
rect 365144 704918 365464 705002
rect 365144 704682 365186 704918
rect 365422 704682 365464 704918
rect 365144 695494 365464 704682
rect 365144 695258 365186 695494
rect 365422 695258 365464 695494
rect 365144 688494 365464 695258
rect 365144 688258 365186 688494
rect 365422 688258 365464 688494
rect 365144 681494 365464 688258
rect 365144 681258 365186 681494
rect 365422 681258 365464 681494
rect 365144 674494 365464 681258
rect 365144 674258 365186 674494
rect 365422 674258 365464 674494
rect 365144 667494 365464 674258
rect 365144 667258 365186 667494
rect 365422 667258 365464 667494
rect 365144 660494 365464 667258
rect 365144 660258 365186 660494
rect 365422 660258 365464 660494
rect 365144 653494 365464 660258
rect 365144 653258 365186 653494
rect 365422 653258 365464 653494
rect 365144 646494 365464 653258
rect 365144 646258 365186 646494
rect 365422 646258 365464 646494
rect 365144 639494 365464 646258
rect 365144 639258 365186 639494
rect 365422 639258 365464 639494
rect 365144 632494 365464 639258
rect 365144 632258 365186 632494
rect 365422 632258 365464 632494
rect 365144 625494 365464 632258
rect 365144 625258 365186 625494
rect 365422 625258 365464 625494
rect 365144 618494 365464 625258
rect 365144 618258 365186 618494
rect 365422 618258 365464 618494
rect 365144 611494 365464 618258
rect 365144 611258 365186 611494
rect 365422 611258 365464 611494
rect 365144 604494 365464 611258
rect 365144 604258 365186 604494
rect 365422 604258 365464 604494
rect 365144 597494 365464 604258
rect 365144 597258 365186 597494
rect 365422 597258 365464 597494
rect 365144 590494 365464 597258
rect 365144 590258 365186 590494
rect 365422 590258 365464 590494
rect 365144 583494 365464 590258
rect 365144 583258 365186 583494
rect 365422 583258 365464 583494
rect 365144 576494 365464 583258
rect 365144 576258 365186 576494
rect 365422 576258 365464 576494
rect 365144 569494 365464 576258
rect 365144 569258 365186 569494
rect 365422 569258 365464 569494
rect 365144 562494 365464 569258
rect 365144 562258 365186 562494
rect 365422 562258 365464 562494
rect 365144 555494 365464 562258
rect 365144 555258 365186 555494
rect 365422 555258 365464 555494
rect 365144 548494 365464 555258
rect 365144 548258 365186 548494
rect 365422 548258 365464 548494
rect 365144 541494 365464 548258
rect 365144 541258 365186 541494
rect 365422 541258 365464 541494
rect 365144 534494 365464 541258
rect 365144 534258 365186 534494
rect 365422 534258 365464 534494
rect 365144 527494 365464 534258
rect 365144 527258 365186 527494
rect 365422 527258 365464 527494
rect 365144 520494 365464 527258
rect 365144 520258 365186 520494
rect 365422 520258 365464 520494
rect 365144 513494 365464 520258
rect 365144 513258 365186 513494
rect 365422 513258 365464 513494
rect 365144 506494 365464 513258
rect 365144 506258 365186 506494
rect 365422 506258 365464 506494
rect 365144 499494 365464 506258
rect 365144 499258 365186 499494
rect 365422 499258 365464 499494
rect 365144 492494 365464 499258
rect 365144 492258 365186 492494
rect 365422 492258 365464 492494
rect 365144 485494 365464 492258
rect 365144 485258 365186 485494
rect 365422 485258 365464 485494
rect 365144 478494 365464 485258
rect 365144 478258 365186 478494
rect 365422 478258 365464 478494
rect 365144 471494 365464 478258
rect 365144 471258 365186 471494
rect 365422 471258 365464 471494
rect 365144 464494 365464 471258
rect 365144 464258 365186 464494
rect 365422 464258 365464 464494
rect 365144 457494 365464 464258
rect 365144 457258 365186 457494
rect 365422 457258 365464 457494
rect 365144 450494 365464 457258
rect 365144 450258 365186 450494
rect 365422 450258 365464 450494
rect 365144 443494 365464 450258
rect 365144 443258 365186 443494
rect 365422 443258 365464 443494
rect 365144 436494 365464 443258
rect 365144 436258 365186 436494
rect 365422 436258 365464 436494
rect 365144 429494 365464 436258
rect 365144 429258 365186 429494
rect 365422 429258 365464 429494
rect 365144 422494 365464 429258
rect 365144 422258 365186 422494
rect 365422 422258 365464 422494
rect 365144 415494 365464 422258
rect 365144 415258 365186 415494
rect 365422 415258 365464 415494
rect 365144 408494 365464 415258
rect 365144 408258 365186 408494
rect 365422 408258 365464 408494
rect 365144 401494 365464 408258
rect 365144 401258 365186 401494
rect 365422 401258 365464 401494
rect 365144 394494 365464 401258
rect 365144 394258 365186 394494
rect 365422 394258 365464 394494
rect 365144 387494 365464 394258
rect 365144 387258 365186 387494
rect 365422 387258 365464 387494
rect 365144 380494 365464 387258
rect 365144 380258 365186 380494
rect 365422 380258 365464 380494
rect 365144 373494 365464 380258
rect 365144 373258 365186 373494
rect 365422 373258 365464 373494
rect 365144 366494 365464 373258
rect 365144 366258 365186 366494
rect 365422 366258 365464 366494
rect 365144 359494 365464 366258
rect 365144 359258 365186 359494
rect 365422 359258 365464 359494
rect 365144 352494 365464 359258
rect 365144 352258 365186 352494
rect 365422 352258 365464 352494
rect 365144 345494 365464 352258
rect 365144 345258 365186 345494
rect 365422 345258 365464 345494
rect 365144 338494 365464 345258
rect 365144 338258 365186 338494
rect 365422 338258 365464 338494
rect 365144 331494 365464 338258
rect 365144 331258 365186 331494
rect 365422 331258 365464 331494
rect 365144 324494 365464 331258
rect 365144 324258 365186 324494
rect 365422 324258 365464 324494
rect 365144 317494 365464 324258
rect 365144 317258 365186 317494
rect 365422 317258 365464 317494
rect 365144 310494 365464 317258
rect 365144 310258 365186 310494
rect 365422 310258 365464 310494
rect 365144 303494 365464 310258
rect 365144 303258 365186 303494
rect 365422 303258 365464 303494
rect 365144 296494 365464 303258
rect 365144 296258 365186 296494
rect 365422 296258 365464 296494
rect 365144 289494 365464 296258
rect 365144 289258 365186 289494
rect 365422 289258 365464 289494
rect 365144 282494 365464 289258
rect 365144 282258 365186 282494
rect 365422 282258 365464 282494
rect 365144 275494 365464 282258
rect 365144 275258 365186 275494
rect 365422 275258 365464 275494
rect 365144 268494 365464 275258
rect 365144 268258 365186 268494
rect 365422 268258 365464 268494
rect 365144 261494 365464 268258
rect 365144 261258 365186 261494
rect 365422 261258 365464 261494
rect 365144 254494 365464 261258
rect 365144 254258 365186 254494
rect 365422 254258 365464 254494
rect 365144 247494 365464 254258
rect 365144 247258 365186 247494
rect 365422 247258 365464 247494
rect 365144 240494 365464 247258
rect 365144 240258 365186 240494
rect 365422 240258 365464 240494
rect 365144 233494 365464 240258
rect 365144 233258 365186 233494
rect 365422 233258 365464 233494
rect 365144 226494 365464 233258
rect 365144 226258 365186 226494
rect 365422 226258 365464 226494
rect 365144 219494 365464 226258
rect 365144 219258 365186 219494
rect 365422 219258 365464 219494
rect 365144 212494 365464 219258
rect 365144 212258 365186 212494
rect 365422 212258 365464 212494
rect 365144 205494 365464 212258
rect 365144 205258 365186 205494
rect 365422 205258 365464 205494
rect 365144 198494 365464 205258
rect 365144 198258 365186 198494
rect 365422 198258 365464 198494
rect 365144 191494 365464 198258
rect 365144 191258 365186 191494
rect 365422 191258 365464 191494
rect 365144 184494 365464 191258
rect 365144 184258 365186 184494
rect 365422 184258 365464 184494
rect 365144 177494 365464 184258
rect 365144 177258 365186 177494
rect 365422 177258 365464 177494
rect 365144 170494 365464 177258
rect 365144 170258 365186 170494
rect 365422 170258 365464 170494
rect 365144 163494 365464 170258
rect 365144 163258 365186 163494
rect 365422 163258 365464 163494
rect 365144 156494 365464 163258
rect 365144 156258 365186 156494
rect 365422 156258 365464 156494
rect 365144 149494 365464 156258
rect 365144 149258 365186 149494
rect 365422 149258 365464 149494
rect 365144 142494 365464 149258
rect 365144 142258 365186 142494
rect 365422 142258 365464 142494
rect 365144 135494 365464 142258
rect 365144 135258 365186 135494
rect 365422 135258 365464 135494
rect 365144 128494 365464 135258
rect 365144 128258 365186 128494
rect 365422 128258 365464 128494
rect 365144 121494 365464 128258
rect 365144 121258 365186 121494
rect 365422 121258 365464 121494
rect 365144 114494 365464 121258
rect 365144 114258 365186 114494
rect 365422 114258 365464 114494
rect 365144 107494 365464 114258
rect 365144 107258 365186 107494
rect 365422 107258 365464 107494
rect 365144 100494 365464 107258
rect 365144 100258 365186 100494
rect 365422 100258 365464 100494
rect 365144 93494 365464 100258
rect 365144 93258 365186 93494
rect 365422 93258 365464 93494
rect 365144 86494 365464 93258
rect 365144 86258 365186 86494
rect 365422 86258 365464 86494
rect 365144 79494 365464 86258
rect 365144 79258 365186 79494
rect 365422 79258 365464 79494
rect 365144 72494 365464 79258
rect 365144 72258 365186 72494
rect 365422 72258 365464 72494
rect 365144 65494 365464 72258
rect 365144 65258 365186 65494
rect 365422 65258 365464 65494
rect 365144 58494 365464 65258
rect 365144 58258 365186 58494
rect 365422 58258 365464 58494
rect 365144 51494 365464 58258
rect 365144 51258 365186 51494
rect 365422 51258 365464 51494
rect 365144 44494 365464 51258
rect 365144 44258 365186 44494
rect 365422 44258 365464 44494
rect 365144 37494 365464 44258
rect 365144 37258 365186 37494
rect 365422 37258 365464 37494
rect 365144 30494 365464 37258
rect 365144 30258 365186 30494
rect 365422 30258 365464 30494
rect 365144 23494 365464 30258
rect 365144 23258 365186 23494
rect 365422 23258 365464 23494
rect 365144 16494 365464 23258
rect 365144 16258 365186 16494
rect 365422 16258 365464 16494
rect 365144 9494 365464 16258
rect 365144 9258 365186 9494
rect 365422 9258 365464 9494
rect 365144 2494 365464 9258
rect 365144 2258 365186 2494
rect 365422 2258 365464 2494
rect 365144 -746 365464 2258
rect 365144 -982 365186 -746
rect 365422 -982 365464 -746
rect 365144 -1066 365464 -982
rect 365144 -1302 365186 -1066
rect 365422 -1302 365464 -1066
rect 365144 -2294 365464 -1302
rect 366876 706198 367196 706230
rect 366876 705962 366918 706198
rect 367154 705962 367196 706198
rect 366876 705878 367196 705962
rect 366876 705642 366918 705878
rect 367154 705642 367196 705878
rect 366876 696434 367196 705642
rect 366876 696198 366918 696434
rect 367154 696198 367196 696434
rect 366876 689434 367196 696198
rect 366876 689198 366918 689434
rect 367154 689198 367196 689434
rect 366876 682434 367196 689198
rect 366876 682198 366918 682434
rect 367154 682198 367196 682434
rect 366876 675434 367196 682198
rect 366876 675198 366918 675434
rect 367154 675198 367196 675434
rect 366876 668434 367196 675198
rect 366876 668198 366918 668434
rect 367154 668198 367196 668434
rect 366876 661434 367196 668198
rect 366876 661198 366918 661434
rect 367154 661198 367196 661434
rect 366876 654434 367196 661198
rect 366876 654198 366918 654434
rect 367154 654198 367196 654434
rect 366876 647434 367196 654198
rect 366876 647198 366918 647434
rect 367154 647198 367196 647434
rect 366876 640434 367196 647198
rect 366876 640198 366918 640434
rect 367154 640198 367196 640434
rect 366876 633434 367196 640198
rect 366876 633198 366918 633434
rect 367154 633198 367196 633434
rect 366876 626434 367196 633198
rect 366876 626198 366918 626434
rect 367154 626198 367196 626434
rect 366876 619434 367196 626198
rect 366876 619198 366918 619434
rect 367154 619198 367196 619434
rect 366876 612434 367196 619198
rect 366876 612198 366918 612434
rect 367154 612198 367196 612434
rect 366876 605434 367196 612198
rect 366876 605198 366918 605434
rect 367154 605198 367196 605434
rect 366876 598434 367196 605198
rect 366876 598198 366918 598434
rect 367154 598198 367196 598434
rect 366876 591434 367196 598198
rect 366876 591198 366918 591434
rect 367154 591198 367196 591434
rect 366876 584434 367196 591198
rect 366876 584198 366918 584434
rect 367154 584198 367196 584434
rect 366876 577434 367196 584198
rect 366876 577198 366918 577434
rect 367154 577198 367196 577434
rect 366876 570434 367196 577198
rect 366876 570198 366918 570434
rect 367154 570198 367196 570434
rect 366876 563434 367196 570198
rect 366876 563198 366918 563434
rect 367154 563198 367196 563434
rect 366876 556434 367196 563198
rect 366876 556198 366918 556434
rect 367154 556198 367196 556434
rect 366876 549434 367196 556198
rect 366876 549198 366918 549434
rect 367154 549198 367196 549434
rect 366876 542434 367196 549198
rect 366876 542198 366918 542434
rect 367154 542198 367196 542434
rect 366876 535434 367196 542198
rect 366876 535198 366918 535434
rect 367154 535198 367196 535434
rect 366876 528434 367196 535198
rect 366876 528198 366918 528434
rect 367154 528198 367196 528434
rect 366876 521434 367196 528198
rect 366876 521198 366918 521434
rect 367154 521198 367196 521434
rect 366876 514434 367196 521198
rect 366876 514198 366918 514434
rect 367154 514198 367196 514434
rect 366876 507434 367196 514198
rect 366876 507198 366918 507434
rect 367154 507198 367196 507434
rect 366876 500434 367196 507198
rect 366876 500198 366918 500434
rect 367154 500198 367196 500434
rect 366876 493434 367196 500198
rect 366876 493198 366918 493434
rect 367154 493198 367196 493434
rect 366876 486434 367196 493198
rect 366876 486198 366918 486434
rect 367154 486198 367196 486434
rect 366876 479434 367196 486198
rect 366876 479198 366918 479434
rect 367154 479198 367196 479434
rect 366876 472434 367196 479198
rect 366876 472198 366918 472434
rect 367154 472198 367196 472434
rect 366876 465434 367196 472198
rect 366876 465198 366918 465434
rect 367154 465198 367196 465434
rect 366876 458434 367196 465198
rect 366876 458198 366918 458434
rect 367154 458198 367196 458434
rect 366876 451434 367196 458198
rect 366876 451198 366918 451434
rect 367154 451198 367196 451434
rect 366876 444434 367196 451198
rect 366876 444198 366918 444434
rect 367154 444198 367196 444434
rect 366876 437434 367196 444198
rect 366876 437198 366918 437434
rect 367154 437198 367196 437434
rect 366876 430434 367196 437198
rect 366876 430198 366918 430434
rect 367154 430198 367196 430434
rect 366876 423434 367196 430198
rect 366876 423198 366918 423434
rect 367154 423198 367196 423434
rect 366876 416434 367196 423198
rect 366876 416198 366918 416434
rect 367154 416198 367196 416434
rect 366876 409434 367196 416198
rect 366876 409198 366918 409434
rect 367154 409198 367196 409434
rect 366876 402434 367196 409198
rect 366876 402198 366918 402434
rect 367154 402198 367196 402434
rect 366876 395434 367196 402198
rect 366876 395198 366918 395434
rect 367154 395198 367196 395434
rect 366876 388434 367196 395198
rect 366876 388198 366918 388434
rect 367154 388198 367196 388434
rect 366876 381434 367196 388198
rect 366876 381198 366918 381434
rect 367154 381198 367196 381434
rect 366876 374434 367196 381198
rect 366876 374198 366918 374434
rect 367154 374198 367196 374434
rect 366876 367434 367196 374198
rect 366876 367198 366918 367434
rect 367154 367198 367196 367434
rect 366876 360434 367196 367198
rect 366876 360198 366918 360434
rect 367154 360198 367196 360434
rect 366876 353434 367196 360198
rect 366876 353198 366918 353434
rect 367154 353198 367196 353434
rect 366876 346434 367196 353198
rect 366876 346198 366918 346434
rect 367154 346198 367196 346434
rect 366876 339434 367196 346198
rect 366876 339198 366918 339434
rect 367154 339198 367196 339434
rect 366876 332434 367196 339198
rect 366876 332198 366918 332434
rect 367154 332198 367196 332434
rect 366876 325434 367196 332198
rect 366876 325198 366918 325434
rect 367154 325198 367196 325434
rect 366876 318434 367196 325198
rect 366876 318198 366918 318434
rect 367154 318198 367196 318434
rect 366876 311434 367196 318198
rect 366876 311198 366918 311434
rect 367154 311198 367196 311434
rect 366876 304434 367196 311198
rect 366876 304198 366918 304434
rect 367154 304198 367196 304434
rect 366876 297434 367196 304198
rect 366876 297198 366918 297434
rect 367154 297198 367196 297434
rect 366876 290434 367196 297198
rect 366876 290198 366918 290434
rect 367154 290198 367196 290434
rect 366876 283434 367196 290198
rect 366876 283198 366918 283434
rect 367154 283198 367196 283434
rect 366876 276434 367196 283198
rect 366876 276198 366918 276434
rect 367154 276198 367196 276434
rect 366876 269434 367196 276198
rect 366876 269198 366918 269434
rect 367154 269198 367196 269434
rect 366876 262434 367196 269198
rect 366876 262198 366918 262434
rect 367154 262198 367196 262434
rect 366876 255434 367196 262198
rect 366876 255198 366918 255434
rect 367154 255198 367196 255434
rect 366876 248434 367196 255198
rect 366876 248198 366918 248434
rect 367154 248198 367196 248434
rect 366876 241434 367196 248198
rect 366876 241198 366918 241434
rect 367154 241198 367196 241434
rect 366876 234434 367196 241198
rect 366876 234198 366918 234434
rect 367154 234198 367196 234434
rect 366876 227434 367196 234198
rect 366876 227198 366918 227434
rect 367154 227198 367196 227434
rect 366876 220434 367196 227198
rect 366876 220198 366918 220434
rect 367154 220198 367196 220434
rect 366876 213434 367196 220198
rect 366876 213198 366918 213434
rect 367154 213198 367196 213434
rect 366876 206434 367196 213198
rect 366876 206198 366918 206434
rect 367154 206198 367196 206434
rect 366876 199434 367196 206198
rect 366876 199198 366918 199434
rect 367154 199198 367196 199434
rect 366876 192434 367196 199198
rect 366876 192198 366918 192434
rect 367154 192198 367196 192434
rect 366876 185434 367196 192198
rect 366876 185198 366918 185434
rect 367154 185198 367196 185434
rect 366876 178434 367196 185198
rect 366876 178198 366918 178434
rect 367154 178198 367196 178434
rect 366876 171434 367196 178198
rect 366876 171198 366918 171434
rect 367154 171198 367196 171434
rect 366876 164434 367196 171198
rect 366876 164198 366918 164434
rect 367154 164198 367196 164434
rect 366876 157434 367196 164198
rect 366876 157198 366918 157434
rect 367154 157198 367196 157434
rect 366876 150434 367196 157198
rect 366876 150198 366918 150434
rect 367154 150198 367196 150434
rect 366876 143434 367196 150198
rect 366876 143198 366918 143434
rect 367154 143198 367196 143434
rect 366876 136434 367196 143198
rect 366876 136198 366918 136434
rect 367154 136198 367196 136434
rect 366876 129434 367196 136198
rect 366876 129198 366918 129434
rect 367154 129198 367196 129434
rect 366876 122434 367196 129198
rect 366876 122198 366918 122434
rect 367154 122198 367196 122434
rect 366876 115434 367196 122198
rect 366876 115198 366918 115434
rect 367154 115198 367196 115434
rect 366876 108434 367196 115198
rect 366876 108198 366918 108434
rect 367154 108198 367196 108434
rect 366876 101434 367196 108198
rect 366876 101198 366918 101434
rect 367154 101198 367196 101434
rect 366876 94434 367196 101198
rect 366876 94198 366918 94434
rect 367154 94198 367196 94434
rect 366876 87434 367196 94198
rect 366876 87198 366918 87434
rect 367154 87198 367196 87434
rect 366876 80434 367196 87198
rect 366876 80198 366918 80434
rect 367154 80198 367196 80434
rect 366876 73434 367196 80198
rect 366876 73198 366918 73434
rect 367154 73198 367196 73434
rect 366876 66434 367196 73198
rect 366876 66198 366918 66434
rect 367154 66198 367196 66434
rect 366876 59434 367196 66198
rect 366876 59198 366918 59434
rect 367154 59198 367196 59434
rect 366876 52434 367196 59198
rect 366876 52198 366918 52434
rect 367154 52198 367196 52434
rect 366876 45434 367196 52198
rect 366876 45198 366918 45434
rect 367154 45198 367196 45434
rect 366876 38434 367196 45198
rect 366876 38198 366918 38434
rect 367154 38198 367196 38434
rect 366876 31434 367196 38198
rect 366876 31198 366918 31434
rect 367154 31198 367196 31434
rect 366876 24434 367196 31198
rect 366876 24198 366918 24434
rect 367154 24198 367196 24434
rect 366876 17434 367196 24198
rect 366876 17198 366918 17434
rect 367154 17198 367196 17434
rect 366876 10434 367196 17198
rect 366876 10198 366918 10434
rect 367154 10198 367196 10434
rect 366876 3434 367196 10198
rect 366876 3198 366918 3434
rect 367154 3198 367196 3434
rect 366876 -1706 367196 3198
rect 366876 -1942 366918 -1706
rect 367154 -1942 367196 -1706
rect 366876 -2026 367196 -1942
rect 366876 -2262 366918 -2026
rect 367154 -2262 367196 -2026
rect 366876 -2294 367196 -2262
rect 372144 705238 372464 706230
rect 372144 705002 372186 705238
rect 372422 705002 372464 705238
rect 372144 704918 372464 705002
rect 372144 704682 372186 704918
rect 372422 704682 372464 704918
rect 372144 695494 372464 704682
rect 372144 695258 372186 695494
rect 372422 695258 372464 695494
rect 372144 688494 372464 695258
rect 372144 688258 372186 688494
rect 372422 688258 372464 688494
rect 372144 681494 372464 688258
rect 372144 681258 372186 681494
rect 372422 681258 372464 681494
rect 372144 674494 372464 681258
rect 372144 674258 372186 674494
rect 372422 674258 372464 674494
rect 372144 667494 372464 674258
rect 372144 667258 372186 667494
rect 372422 667258 372464 667494
rect 372144 660494 372464 667258
rect 372144 660258 372186 660494
rect 372422 660258 372464 660494
rect 372144 653494 372464 660258
rect 372144 653258 372186 653494
rect 372422 653258 372464 653494
rect 372144 646494 372464 653258
rect 372144 646258 372186 646494
rect 372422 646258 372464 646494
rect 372144 639494 372464 646258
rect 372144 639258 372186 639494
rect 372422 639258 372464 639494
rect 372144 632494 372464 639258
rect 372144 632258 372186 632494
rect 372422 632258 372464 632494
rect 372144 625494 372464 632258
rect 372144 625258 372186 625494
rect 372422 625258 372464 625494
rect 372144 618494 372464 625258
rect 372144 618258 372186 618494
rect 372422 618258 372464 618494
rect 372144 611494 372464 618258
rect 372144 611258 372186 611494
rect 372422 611258 372464 611494
rect 372144 604494 372464 611258
rect 372144 604258 372186 604494
rect 372422 604258 372464 604494
rect 372144 597494 372464 604258
rect 372144 597258 372186 597494
rect 372422 597258 372464 597494
rect 372144 590494 372464 597258
rect 372144 590258 372186 590494
rect 372422 590258 372464 590494
rect 372144 583494 372464 590258
rect 372144 583258 372186 583494
rect 372422 583258 372464 583494
rect 372144 576494 372464 583258
rect 372144 576258 372186 576494
rect 372422 576258 372464 576494
rect 372144 569494 372464 576258
rect 372144 569258 372186 569494
rect 372422 569258 372464 569494
rect 372144 562494 372464 569258
rect 372144 562258 372186 562494
rect 372422 562258 372464 562494
rect 372144 555494 372464 562258
rect 372144 555258 372186 555494
rect 372422 555258 372464 555494
rect 372144 548494 372464 555258
rect 372144 548258 372186 548494
rect 372422 548258 372464 548494
rect 372144 541494 372464 548258
rect 372144 541258 372186 541494
rect 372422 541258 372464 541494
rect 372144 534494 372464 541258
rect 372144 534258 372186 534494
rect 372422 534258 372464 534494
rect 372144 527494 372464 534258
rect 372144 527258 372186 527494
rect 372422 527258 372464 527494
rect 372144 520494 372464 527258
rect 372144 520258 372186 520494
rect 372422 520258 372464 520494
rect 372144 513494 372464 520258
rect 372144 513258 372186 513494
rect 372422 513258 372464 513494
rect 372144 506494 372464 513258
rect 372144 506258 372186 506494
rect 372422 506258 372464 506494
rect 372144 499494 372464 506258
rect 372144 499258 372186 499494
rect 372422 499258 372464 499494
rect 372144 492494 372464 499258
rect 372144 492258 372186 492494
rect 372422 492258 372464 492494
rect 372144 485494 372464 492258
rect 372144 485258 372186 485494
rect 372422 485258 372464 485494
rect 372144 478494 372464 485258
rect 372144 478258 372186 478494
rect 372422 478258 372464 478494
rect 372144 471494 372464 478258
rect 372144 471258 372186 471494
rect 372422 471258 372464 471494
rect 372144 464494 372464 471258
rect 372144 464258 372186 464494
rect 372422 464258 372464 464494
rect 372144 457494 372464 464258
rect 372144 457258 372186 457494
rect 372422 457258 372464 457494
rect 372144 450494 372464 457258
rect 372144 450258 372186 450494
rect 372422 450258 372464 450494
rect 372144 443494 372464 450258
rect 372144 443258 372186 443494
rect 372422 443258 372464 443494
rect 372144 436494 372464 443258
rect 372144 436258 372186 436494
rect 372422 436258 372464 436494
rect 372144 429494 372464 436258
rect 372144 429258 372186 429494
rect 372422 429258 372464 429494
rect 372144 422494 372464 429258
rect 372144 422258 372186 422494
rect 372422 422258 372464 422494
rect 372144 415494 372464 422258
rect 372144 415258 372186 415494
rect 372422 415258 372464 415494
rect 372144 408494 372464 415258
rect 372144 408258 372186 408494
rect 372422 408258 372464 408494
rect 372144 401494 372464 408258
rect 372144 401258 372186 401494
rect 372422 401258 372464 401494
rect 372144 394494 372464 401258
rect 372144 394258 372186 394494
rect 372422 394258 372464 394494
rect 372144 387494 372464 394258
rect 372144 387258 372186 387494
rect 372422 387258 372464 387494
rect 372144 380494 372464 387258
rect 372144 380258 372186 380494
rect 372422 380258 372464 380494
rect 372144 373494 372464 380258
rect 372144 373258 372186 373494
rect 372422 373258 372464 373494
rect 372144 366494 372464 373258
rect 372144 366258 372186 366494
rect 372422 366258 372464 366494
rect 372144 359494 372464 366258
rect 372144 359258 372186 359494
rect 372422 359258 372464 359494
rect 372144 352494 372464 359258
rect 372144 352258 372186 352494
rect 372422 352258 372464 352494
rect 372144 345494 372464 352258
rect 372144 345258 372186 345494
rect 372422 345258 372464 345494
rect 372144 338494 372464 345258
rect 372144 338258 372186 338494
rect 372422 338258 372464 338494
rect 372144 331494 372464 338258
rect 372144 331258 372186 331494
rect 372422 331258 372464 331494
rect 372144 324494 372464 331258
rect 372144 324258 372186 324494
rect 372422 324258 372464 324494
rect 372144 317494 372464 324258
rect 372144 317258 372186 317494
rect 372422 317258 372464 317494
rect 372144 310494 372464 317258
rect 372144 310258 372186 310494
rect 372422 310258 372464 310494
rect 372144 303494 372464 310258
rect 372144 303258 372186 303494
rect 372422 303258 372464 303494
rect 372144 296494 372464 303258
rect 372144 296258 372186 296494
rect 372422 296258 372464 296494
rect 372144 289494 372464 296258
rect 372144 289258 372186 289494
rect 372422 289258 372464 289494
rect 372144 282494 372464 289258
rect 372144 282258 372186 282494
rect 372422 282258 372464 282494
rect 372144 275494 372464 282258
rect 372144 275258 372186 275494
rect 372422 275258 372464 275494
rect 372144 268494 372464 275258
rect 372144 268258 372186 268494
rect 372422 268258 372464 268494
rect 372144 261494 372464 268258
rect 372144 261258 372186 261494
rect 372422 261258 372464 261494
rect 372144 254494 372464 261258
rect 372144 254258 372186 254494
rect 372422 254258 372464 254494
rect 372144 247494 372464 254258
rect 372144 247258 372186 247494
rect 372422 247258 372464 247494
rect 372144 240494 372464 247258
rect 372144 240258 372186 240494
rect 372422 240258 372464 240494
rect 372144 233494 372464 240258
rect 372144 233258 372186 233494
rect 372422 233258 372464 233494
rect 372144 226494 372464 233258
rect 372144 226258 372186 226494
rect 372422 226258 372464 226494
rect 372144 219494 372464 226258
rect 372144 219258 372186 219494
rect 372422 219258 372464 219494
rect 372144 212494 372464 219258
rect 372144 212258 372186 212494
rect 372422 212258 372464 212494
rect 372144 205494 372464 212258
rect 372144 205258 372186 205494
rect 372422 205258 372464 205494
rect 372144 198494 372464 205258
rect 372144 198258 372186 198494
rect 372422 198258 372464 198494
rect 372144 191494 372464 198258
rect 372144 191258 372186 191494
rect 372422 191258 372464 191494
rect 372144 184494 372464 191258
rect 372144 184258 372186 184494
rect 372422 184258 372464 184494
rect 372144 177494 372464 184258
rect 372144 177258 372186 177494
rect 372422 177258 372464 177494
rect 372144 170494 372464 177258
rect 372144 170258 372186 170494
rect 372422 170258 372464 170494
rect 372144 163494 372464 170258
rect 372144 163258 372186 163494
rect 372422 163258 372464 163494
rect 372144 156494 372464 163258
rect 372144 156258 372186 156494
rect 372422 156258 372464 156494
rect 372144 149494 372464 156258
rect 372144 149258 372186 149494
rect 372422 149258 372464 149494
rect 372144 142494 372464 149258
rect 372144 142258 372186 142494
rect 372422 142258 372464 142494
rect 372144 135494 372464 142258
rect 372144 135258 372186 135494
rect 372422 135258 372464 135494
rect 372144 128494 372464 135258
rect 372144 128258 372186 128494
rect 372422 128258 372464 128494
rect 372144 121494 372464 128258
rect 372144 121258 372186 121494
rect 372422 121258 372464 121494
rect 372144 114494 372464 121258
rect 372144 114258 372186 114494
rect 372422 114258 372464 114494
rect 372144 107494 372464 114258
rect 372144 107258 372186 107494
rect 372422 107258 372464 107494
rect 372144 100494 372464 107258
rect 372144 100258 372186 100494
rect 372422 100258 372464 100494
rect 372144 93494 372464 100258
rect 372144 93258 372186 93494
rect 372422 93258 372464 93494
rect 372144 86494 372464 93258
rect 372144 86258 372186 86494
rect 372422 86258 372464 86494
rect 372144 79494 372464 86258
rect 372144 79258 372186 79494
rect 372422 79258 372464 79494
rect 372144 72494 372464 79258
rect 372144 72258 372186 72494
rect 372422 72258 372464 72494
rect 372144 65494 372464 72258
rect 372144 65258 372186 65494
rect 372422 65258 372464 65494
rect 372144 58494 372464 65258
rect 372144 58258 372186 58494
rect 372422 58258 372464 58494
rect 372144 51494 372464 58258
rect 372144 51258 372186 51494
rect 372422 51258 372464 51494
rect 372144 44494 372464 51258
rect 372144 44258 372186 44494
rect 372422 44258 372464 44494
rect 372144 37494 372464 44258
rect 372144 37258 372186 37494
rect 372422 37258 372464 37494
rect 372144 30494 372464 37258
rect 372144 30258 372186 30494
rect 372422 30258 372464 30494
rect 372144 23494 372464 30258
rect 372144 23258 372186 23494
rect 372422 23258 372464 23494
rect 372144 16494 372464 23258
rect 372144 16258 372186 16494
rect 372422 16258 372464 16494
rect 372144 9494 372464 16258
rect 372144 9258 372186 9494
rect 372422 9258 372464 9494
rect 372144 2494 372464 9258
rect 372144 2258 372186 2494
rect 372422 2258 372464 2494
rect 372144 -746 372464 2258
rect 372144 -982 372186 -746
rect 372422 -982 372464 -746
rect 372144 -1066 372464 -982
rect 372144 -1302 372186 -1066
rect 372422 -1302 372464 -1066
rect 372144 -2294 372464 -1302
rect 373876 706198 374196 706230
rect 373876 705962 373918 706198
rect 374154 705962 374196 706198
rect 373876 705878 374196 705962
rect 373876 705642 373918 705878
rect 374154 705642 374196 705878
rect 373876 696434 374196 705642
rect 373876 696198 373918 696434
rect 374154 696198 374196 696434
rect 373876 689434 374196 696198
rect 373876 689198 373918 689434
rect 374154 689198 374196 689434
rect 373876 682434 374196 689198
rect 373876 682198 373918 682434
rect 374154 682198 374196 682434
rect 373876 675434 374196 682198
rect 373876 675198 373918 675434
rect 374154 675198 374196 675434
rect 373876 668434 374196 675198
rect 373876 668198 373918 668434
rect 374154 668198 374196 668434
rect 373876 661434 374196 668198
rect 373876 661198 373918 661434
rect 374154 661198 374196 661434
rect 373876 654434 374196 661198
rect 373876 654198 373918 654434
rect 374154 654198 374196 654434
rect 373876 647434 374196 654198
rect 373876 647198 373918 647434
rect 374154 647198 374196 647434
rect 373876 640434 374196 647198
rect 373876 640198 373918 640434
rect 374154 640198 374196 640434
rect 373876 633434 374196 640198
rect 373876 633198 373918 633434
rect 374154 633198 374196 633434
rect 373876 626434 374196 633198
rect 373876 626198 373918 626434
rect 374154 626198 374196 626434
rect 373876 619434 374196 626198
rect 373876 619198 373918 619434
rect 374154 619198 374196 619434
rect 373876 612434 374196 619198
rect 373876 612198 373918 612434
rect 374154 612198 374196 612434
rect 373876 605434 374196 612198
rect 373876 605198 373918 605434
rect 374154 605198 374196 605434
rect 373876 598434 374196 605198
rect 373876 598198 373918 598434
rect 374154 598198 374196 598434
rect 373876 591434 374196 598198
rect 373876 591198 373918 591434
rect 374154 591198 374196 591434
rect 373876 584434 374196 591198
rect 373876 584198 373918 584434
rect 374154 584198 374196 584434
rect 373876 577434 374196 584198
rect 373876 577198 373918 577434
rect 374154 577198 374196 577434
rect 373876 570434 374196 577198
rect 373876 570198 373918 570434
rect 374154 570198 374196 570434
rect 373876 563434 374196 570198
rect 373876 563198 373918 563434
rect 374154 563198 374196 563434
rect 373876 556434 374196 563198
rect 373876 556198 373918 556434
rect 374154 556198 374196 556434
rect 373876 549434 374196 556198
rect 373876 549198 373918 549434
rect 374154 549198 374196 549434
rect 373876 542434 374196 549198
rect 373876 542198 373918 542434
rect 374154 542198 374196 542434
rect 373876 535434 374196 542198
rect 373876 535198 373918 535434
rect 374154 535198 374196 535434
rect 373876 528434 374196 535198
rect 373876 528198 373918 528434
rect 374154 528198 374196 528434
rect 373876 521434 374196 528198
rect 373876 521198 373918 521434
rect 374154 521198 374196 521434
rect 373876 514434 374196 521198
rect 373876 514198 373918 514434
rect 374154 514198 374196 514434
rect 373876 507434 374196 514198
rect 373876 507198 373918 507434
rect 374154 507198 374196 507434
rect 373876 500434 374196 507198
rect 373876 500198 373918 500434
rect 374154 500198 374196 500434
rect 373876 493434 374196 500198
rect 373876 493198 373918 493434
rect 374154 493198 374196 493434
rect 373876 486434 374196 493198
rect 373876 486198 373918 486434
rect 374154 486198 374196 486434
rect 373876 479434 374196 486198
rect 373876 479198 373918 479434
rect 374154 479198 374196 479434
rect 373876 472434 374196 479198
rect 373876 472198 373918 472434
rect 374154 472198 374196 472434
rect 373876 465434 374196 472198
rect 373876 465198 373918 465434
rect 374154 465198 374196 465434
rect 373876 458434 374196 465198
rect 373876 458198 373918 458434
rect 374154 458198 374196 458434
rect 373876 451434 374196 458198
rect 373876 451198 373918 451434
rect 374154 451198 374196 451434
rect 373876 444434 374196 451198
rect 373876 444198 373918 444434
rect 374154 444198 374196 444434
rect 373876 437434 374196 444198
rect 373876 437198 373918 437434
rect 374154 437198 374196 437434
rect 373876 430434 374196 437198
rect 373876 430198 373918 430434
rect 374154 430198 374196 430434
rect 373876 423434 374196 430198
rect 373876 423198 373918 423434
rect 374154 423198 374196 423434
rect 373876 416434 374196 423198
rect 373876 416198 373918 416434
rect 374154 416198 374196 416434
rect 373876 409434 374196 416198
rect 373876 409198 373918 409434
rect 374154 409198 374196 409434
rect 373876 402434 374196 409198
rect 373876 402198 373918 402434
rect 374154 402198 374196 402434
rect 373876 395434 374196 402198
rect 373876 395198 373918 395434
rect 374154 395198 374196 395434
rect 373876 388434 374196 395198
rect 373876 388198 373918 388434
rect 374154 388198 374196 388434
rect 373876 381434 374196 388198
rect 373876 381198 373918 381434
rect 374154 381198 374196 381434
rect 373876 374434 374196 381198
rect 373876 374198 373918 374434
rect 374154 374198 374196 374434
rect 373876 367434 374196 374198
rect 373876 367198 373918 367434
rect 374154 367198 374196 367434
rect 373876 360434 374196 367198
rect 373876 360198 373918 360434
rect 374154 360198 374196 360434
rect 373876 353434 374196 360198
rect 373876 353198 373918 353434
rect 374154 353198 374196 353434
rect 373876 346434 374196 353198
rect 373876 346198 373918 346434
rect 374154 346198 374196 346434
rect 373876 339434 374196 346198
rect 373876 339198 373918 339434
rect 374154 339198 374196 339434
rect 373876 332434 374196 339198
rect 373876 332198 373918 332434
rect 374154 332198 374196 332434
rect 373876 325434 374196 332198
rect 373876 325198 373918 325434
rect 374154 325198 374196 325434
rect 373876 318434 374196 325198
rect 373876 318198 373918 318434
rect 374154 318198 374196 318434
rect 373876 311434 374196 318198
rect 373876 311198 373918 311434
rect 374154 311198 374196 311434
rect 373876 304434 374196 311198
rect 373876 304198 373918 304434
rect 374154 304198 374196 304434
rect 373876 297434 374196 304198
rect 373876 297198 373918 297434
rect 374154 297198 374196 297434
rect 373876 290434 374196 297198
rect 373876 290198 373918 290434
rect 374154 290198 374196 290434
rect 373876 283434 374196 290198
rect 373876 283198 373918 283434
rect 374154 283198 374196 283434
rect 373876 276434 374196 283198
rect 373876 276198 373918 276434
rect 374154 276198 374196 276434
rect 373876 269434 374196 276198
rect 373876 269198 373918 269434
rect 374154 269198 374196 269434
rect 373876 262434 374196 269198
rect 373876 262198 373918 262434
rect 374154 262198 374196 262434
rect 373876 255434 374196 262198
rect 373876 255198 373918 255434
rect 374154 255198 374196 255434
rect 373876 248434 374196 255198
rect 373876 248198 373918 248434
rect 374154 248198 374196 248434
rect 373876 241434 374196 248198
rect 373876 241198 373918 241434
rect 374154 241198 374196 241434
rect 373876 234434 374196 241198
rect 373876 234198 373918 234434
rect 374154 234198 374196 234434
rect 373876 227434 374196 234198
rect 373876 227198 373918 227434
rect 374154 227198 374196 227434
rect 373876 220434 374196 227198
rect 373876 220198 373918 220434
rect 374154 220198 374196 220434
rect 373876 213434 374196 220198
rect 373876 213198 373918 213434
rect 374154 213198 374196 213434
rect 373876 206434 374196 213198
rect 373876 206198 373918 206434
rect 374154 206198 374196 206434
rect 373876 199434 374196 206198
rect 373876 199198 373918 199434
rect 374154 199198 374196 199434
rect 373876 192434 374196 199198
rect 373876 192198 373918 192434
rect 374154 192198 374196 192434
rect 373876 185434 374196 192198
rect 373876 185198 373918 185434
rect 374154 185198 374196 185434
rect 373876 178434 374196 185198
rect 373876 178198 373918 178434
rect 374154 178198 374196 178434
rect 373876 171434 374196 178198
rect 373876 171198 373918 171434
rect 374154 171198 374196 171434
rect 373876 164434 374196 171198
rect 373876 164198 373918 164434
rect 374154 164198 374196 164434
rect 373876 157434 374196 164198
rect 373876 157198 373918 157434
rect 374154 157198 374196 157434
rect 373876 150434 374196 157198
rect 373876 150198 373918 150434
rect 374154 150198 374196 150434
rect 373876 143434 374196 150198
rect 373876 143198 373918 143434
rect 374154 143198 374196 143434
rect 373876 136434 374196 143198
rect 373876 136198 373918 136434
rect 374154 136198 374196 136434
rect 373876 129434 374196 136198
rect 373876 129198 373918 129434
rect 374154 129198 374196 129434
rect 373876 122434 374196 129198
rect 373876 122198 373918 122434
rect 374154 122198 374196 122434
rect 373876 115434 374196 122198
rect 373876 115198 373918 115434
rect 374154 115198 374196 115434
rect 373876 108434 374196 115198
rect 373876 108198 373918 108434
rect 374154 108198 374196 108434
rect 373876 101434 374196 108198
rect 373876 101198 373918 101434
rect 374154 101198 374196 101434
rect 373876 94434 374196 101198
rect 373876 94198 373918 94434
rect 374154 94198 374196 94434
rect 373876 87434 374196 94198
rect 373876 87198 373918 87434
rect 374154 87198 374196 87434
rect 373876 80434 374196 87198
rect 373876 80198 373918 80434
rect 374154 80198 374196 80434
rect 373876 73434 374196 80198
rect 373876 73198 373918 73434
rect 374154 73198 374196 73434
rect 373876 66434 374196 73198
rect 373876 66198 373918 66434
rect 374154 66198 374196 66434
rect 373876 59434 374196 66198
rect 373876 59198 373918 59434
rect 374154 59198 374196 59434
rect 373876 52434 374196 59198
rect 373876 52198 373918 52434
rect 374154 52198 374196 52434
rect 373876 45434 374196 52198
rect 373876 45198 373918 45434
rect 374154 45198 374196 45434
rect 373876 38434 374196 45198
rect 373876 38198 373918 38434
rect 374154 38198 374196 38434
rect 373876 31434 374196 38198
rect 373876 31198 373918 31434
rect 374154 31198 374196 31434
rect 373876 24434 374196 31198
rect 373876 24198 373918 24434
rect 374154 24198 374196 24434
rect 373876 17434 374196 24198
rect 373876 17198 373918 17434
rect 374154 17198 374196 17434
rect 373876 10434 374196 17198
rect 373876 10198 373918 10434
rect 374154 10198 374196 10434
rect 373876 3434 374196 10198
rect 373876 3198 373918 3434
rect 374154 3198 374196 3434
rect 373876 -1706 374196 3198
rect 373876 -1942 373918 -1706
rect 374154 -1942 374196 -1706
rect 373876 -2026 374196 -1942
rect 373876 -2262 373918 -2026
rect 374154 -2262 374196 -2026
rect 373876 -2294 374196 -2262
rect 379144 705238 379464 706230
rect 379144 705002 379186 705238
rect 379422 705002 379464 705238
rect 379144 704918 379464 705002
rect 379144 704682 379186 704918
rect 379422 704682 379464 704918
rect 379144 695494 379464 704682
rect 379144 695258 379186 695494
rect 379422 695258 379464 695494
rect 379144 688494 379464 695258
rect 379144 688258 379186 688494
rect 379422 688258 379464 688494
rect 379144 681494 379464 688258
rect 379144 681258 379186 681494
rect 379422 681258 379464 681494
rect 379144 674494 379464 681258
rect 379144 674258 379186 674494
rect 379422 674258 379464 674494
rect 379144 667494 379464 674258
rect 379144 667258 379186 667494
rect 379422 667258 379464 667494
rect 379144 660494 379464 667258
rect 379144 660258 379186 660494
rect 379422 660258 379464 660494
rect 379144 653494 379464 660258
rect 379144 653258 379186 653494
rect 379422 653258 379464 653494
rect 379144 646494 379464 653258
rect 379144 646258 379186 646494
rect 379422 646258 379464 646494
rect 379144 639494 379464 646258
rect 379144 639258 379186 639494
rect 379422 639258 379464 639494
rect 379144 632494 379464 639258
rect 379144 632258 379186 632494
rect 379422 632258 379464 632494
rect 379144 625494 379464 632258
rect 379144 625258 379186 625494
rect 379422 625258 379464 625494
rect 379144 618494 379464 625258
rect 379144 618258 379186 618494
rect 379422 618258 379464 618494
rect 379144 611494 379464 618258
rect 379144 611258 379186 611494
rect 379422 611258 379464 611494
rect 379144 604494 379464 611258
rect 379144 604258 379186 604494
rect 379422 604258 379464 604494
rect 379144 597494 379464 604258
rect 379144 597258 379186 597494
rect 379422 597258 379464 597494
rect 379144 590494 379464 597258
rect 379144 590258 379186 590494
rect 379422 590258 379464 590494
rect 379144 583494 379464 590258
rect 379144 583258 379186 583494
rect 379422 583258 379464 583494
rect 379144 576494 379464 583258
rect 379144 576258 379186 576494
rect 379422 576258 379464 576494
rect 379144 569494 379464 576258
rect 379144 569258 379186 569494
rect 379422 569258 379464 569494
rect 379144 562494 379464 569258
rect 379144 562258 379186 562494
rect 379422 562258 379464 562494
rect 379144 555494 379464 562258
rect 379144 555258 379186 555494
rect 379422 555258 379464 555494
rect 379144 548494 379464 555258
rect 379144 548258 379186 548494
rect 379422 548258 379464 548494
rect 379144 541494 379464 548258
rect 379144 541258 379186 541494
rect 379422 541258 379464 541494
rect 379144 534494 379464 541258
rect 379144 534258 379186 534494
rect 379422 534258 379464 534494
rect 379144 527494 379464 534258
rect 379144 527258 379186 527494
rect 379422 527258 379464 527494
rect 379144 520494 379464 527258
rect 379144 520258 379186 520494
rect 379422 520258 379464 520494
rect 379144 513494 379464 520258
rect 379144 513258 379186 513494
rect 379422 513258 379464 513494
rect 379144 506494 379464 513258
rect 379144 506258 379186 506494
rect 379422 506258 379464 506494
rect 379144 499494 379464 506258
rect 379144 499258 379186 499494
rect 379422 499258 379464 499494
rect 379144 492494 379464 499258
rect 379144 492258 379186 492494
rect 379422 492258 379464 492494
rect 379144 485494 379464 492258
rect 379144 485258 379186 485494
rect 379422 485258 379464 485494
rect 379144 478494 379464 485258
rect 379144 478258 379186 478494
rect 379422 478258 379464 478494
rect 379144 471494 379464 478258
rect 379144 471258 379186 471494
rect 379422 471258 379464 471494
rect 379144 464494 379464 471258
rect 379144 464258 379186 464494
rect 379422 464258 379464 464494
rect 379144 457494 379464 464258
rect 379144 457258 379186 457494
rect 379422 457258 379464 457494
rect 379144 450494 379464 457258
rect 379144 450258 379186 450494
rect 379422 450258 379464 450494
rect 379144 443494 379464 450258
rect 379144 443258 379186 443494
rect 379422 443258 379464 443494
rect 379144 436494 379464 443258
rect 379144 436258 379186 436494
rect 379422 436258 379464 436494
rect 379144 429494 379464 436258
rect 379144 429258 379186 429494
rect 379422 429258 379464 429494
rect 379144 422494 379464 429258
rect 379144 422258 379186 422494
rect 379422 422258 379464 422494
rect 379144 415494 379464 422258
rect 379144 415258 379186 415494
rect 379422 415258 379464 415494
rect 379144 408494 379464 415258
rect 379144 408258 379186 408494
rect 379422 408258 379464 408494
rect 379144 401494 379464 408258
rect 379144 401258 379186 401494
rect 379422 401258 379464 401494
rect 379144 394494 379464 401258
rect 379144 394258 379186 394494
rect 379422 394258 379464 394494
rect 379144 387494 379464 394258
rect 379144 387258 379186 387494
rect 379422 387258 379464 387494
rect 379144 380494 379464 387258
rect 379144 380258 379186 380494
rect 379422 380258 379464 380494
rect 379144 373494 379464 380258
rect 379144 373258 379186 373494
rect 379422 373258 379464 373494
rect 379144 366494 379464 373258
rect 379144 366258 379186 366494
rect 379422 366258 379464 366494
rect 379144 359494 379464 366258
rect 379144 359258 379186 359494
rect 379422 359258 379464 359494
rect 379144 352494 379464 359258
rect 379144 352258 379186 352494
rect 379422 352258 379464 352494
rect 379144 345494 379464 352258
rect 379144 345258 379186 345494
rect 379422 345258 379464 345494
rect 379144 338494 379464 345258
rect 379144 338258 379186 338494
rect 379422 338258 379464 338494
rect 379144 331494 379464 338258
rect 379144 331258 379186 331494
rect 379422 331258 379464 331494
rect 379144 324494 379464 331258
rect 379144 324258 379186 324494
rect 379422 324258 379464 324494
rect 379144 317494 379464 324258
rect 379144 317258 379186 317494
rect 379422 317258 379464 317494
rect 379144 310494 379464 317258
rect 379144 310258 379186 310494
rect 379422 310258 379464 310494
rect 379144 303494 379464 310258
rect 379144 303258 379186 303494
rect 379422 303258 379464 303494
rect 379144 296494 379464 303258
rect 379144 296258 379186 296494
rect 379422 296258 379464 296494
rect 379144 289494 379464 296258
rect 379144 289258 379186 289494
rect 379422 289258 379464 289494
rect 379144 282494 379464 289258
rect 379144 282258 379186 282494
rect 379422 282258 379464 282494
rect 379144 275494 379464 282258
rect 379144 275258 379186 275494
rect 379422 275258 379464 275494
rect 379144 268494 379464 275258
rect 379144 268258 379186 268494
rect 379422 268258 379464 268494
rect 379144 261494 379464 268258
rect 379144 261258 379186 261494
rect 379422 261258 379464 261494
rect 379144 254494 379464 261258
rect 379144 254258 379186 254494
rect 379422 254258 379464 254494
rect 379144 247494 379464 254258
rect 379144 247258 379186 247494
rect 379422 247258 379464 247494
rect 379144 240494 379464 247258
rect 379144 240258 379186 240494
rect 379422 240258 379464 240494
rect 379144 233494 379464 240258
rect 379144 233258 379186 233494
rect 379422 233258 379464 233494
rect 379144 226494 379464 233258
rect 379144 226258 379186 226494
rect 379422 226258 379464 226494
rect 379144 219494 379464 226258
rect 379144 219258 379186 219494
rect 379422 219258 379464 219494
rect 379144 212494 379464 219258
rect 379144 212258 379186 212494
rect 379422 212258 379464 212494
rect 379144 205494 379464 212258
rect 379144 205258 379186 205494
rect 379422 205258 379464 205494
rect 379144 198494 379464 205258
rect 379144 198258 379186 198494
rect 379422 198258 379464 198494
rect 379144 191494 379464 198258
rect 379144 191258 379186 191494
rect 379422 191258 379464 191494
rect 379144 184494 379464 191258
rect 379144 184258 379186 184494
rect 379422 184258 379464 184494
rect 379144 177494 379464 184258
rect 379144 177258 379186 177494
rect 379422 177258 379464 177494
rect 379144 170494 379464 177258
rect 379144 170258 379186 170494
rect 379422 170258 379464 170494
rect 379144 163494 379464 170258
rect 379144 163258 379186 163494
rect 379422 163258 379464 163494
rect 379144 156494 379464 163258
rect 379144 156258 379186 156494
rect 379422 156258 379464 156494
rect 379144 149494 379464 156258
rect 379144 149258 379186 149494
rect 379422 149258 379464 149494
rect 379144 142494 379464 149258
rect 379144 142258 379186 142494
rect 379422 142258 379464 142494
rect 379144 135494 379464 142258
rect 379144 135258 379186 135494
rect 379422 135258 379464 135494
rect 379144 128494 379464 135258
rect 379144 128258 379186 128494
rect 379422 128258 379464 128494
rect 379144 121494 379464 128258
rect 379144 121258 379186 121494
rect 379422 121258 379464 121494
rect 379144 114494 379464 121258
rect 379144 114258 379186 114494
rect 379422 114258 379464 114494
rect 379144 107494 379464 114258
rect 379144 107258 379186 107494
rect 379422 107258 379464 107494
rect 379144 100494 379464 107258
rect 379144 100258 379186 100494
rect 379422 100258 379464 100494
rect 379144 93494 379464 100258
rect 379144 93258 379186 93494
rect 379422 93258 379464 93494
rect 379144 86494 379464 93258
rect 379144 86258 379186 86494
rect 379422 86258 379464 86494
rect 379144 79494 379464 86258
rect 379144 79258 379186 79494
rect 379422 79258 379464 79494
rect 379144 72494 379464 79258
rect 379144 72258 379186 72494
rect 379422 72258 379464 72494
rect 379144 65494 379464 72258
rect 379144 65258 379186 65494
rect 379422 65258 379464 65494
rect 379144 58494 379464 65258
rect 379144 58258 379186 58494
rect 379422 58258 379464 58494
rect 379144 51494 379464 58258
rect 379144 51258 379186 51494
rect 379422 51258 379464 51494
rect 379144 44494 379464 51258
rect 379144 44258 379186 44494
rect 379422 44258 379464 44494
rect 379144 37494 379464 44258
rect 379144 37258 379186 37494
rect 379422 37258 379464 37494
rect 379144 30494 379464 37258
rect 379144 30258 379186 30494
rect 379422 30258 379464 30494
rect 379144 23494 379464 30258
rect 379144 23258 379186 23494
rect 379422 23258 379464 23494
rect 379144 16494 379464 23258
rect 379144 16258 379186 16494
rect 379422 16258 379464 16494
rect 379144 9494 379464 16258
rect 379144 9258 379186 9494
rect 379422 9258 379464 9494
rect 379144 2494 379464 9258
rect 379144 2258 379186 2494
rect 379422 2258 379464 2494
rect 379144 -746 379464 2258
rect 379144 -982 379186 -746
rect 379422 -982 379464 -746
rect 379144 -1066 379464 -982
rect 379144 -1302 379186 -1066
rect 379422 -1302 379464 -1066
rect 379144 -2294 379464 -1302
rect 380876 706198 381196 706230
rect 380876 705962 380918 706198
rect 381154 705962 381196 706198
rect 380876 705878 381196 705962
rect 380876 705642 380918 705878
rect 381154 705642 381196 705878
rect 380876 696434 381196 705642
rect 380876 696198 380918 696434
rect 381154 696198 381196 696434
rect 380876 689434 381196 696198
rect 380876 689198 380918 689434
rect 381154 689198 381196 689434
rect 380876 682434 381196 689198
rect 380876 682198 380918 682434
rect 381154 682198 381196 682434
rect 380876 675434 381196 682198
rect 380876 675198 380918 675434
rect 381154 675198 381196 675434
rect 380876 668434 381196 675198
rect 380876 668198 380918 668434
rect 381154 668198 381196 668434
rect 380876 661434 381196 668198
rect 380876 661198 380918 661434
rect 381154 661198 381196 661434
rect 380876 654434 381196 661198
rect 380876 654198 380918 654434
rect 381154 654198 381196 654434
rect 380876 647434 381196 654198
rect 380876 647198 380918 647434
rect 381154 647198 381196 647434
rect 380876 640434 381196 647198
rect 380876 640198 380918 640434
rect 381154 640198 381196 640434
rect 380876 633434 381196 640198
rect 380876 633198 380918 633434
rect 381154 633198 381196 633434
rect 380876 626434 381196 633198
rect 380876 626198 380918 626434
rect 381154 626198 381196 626434
rect 380876 619434 381196 626198
rect 380876 619198 380918 619434
rect 381154 619198 381196 619434
rect 380876 612434 381196 619198
rect 380876 612198 380918 612434
rect 381154 612198 381196 612434
rect 380876 605434 381196 612198
rect 380876 605198 380918 605434
rect 381154 605198 381196 605434
rect 380876 598434 381196 605198
rect 380876 598198 380918 598434
rect 381154 598198 381196 598434
rect 380876 591434 381196 598198
rect 380876 591198 380918 591434
rect 381154 591198 381196 591434
rect 380876 584434 381196 591198
rect 380876 584198 380918 584434
rect 381154 584198 381196 584434
rect 380876 577434 381196 584198
rect 380876 577198 380918 577434
rect 381154 577198 381196 577434
rect 380876 570434 381196 577198
rect 380876 570198 380918 570434
rect 381154 570198 381196 570434
rect 380876 563434 381196 570198
rect 380876 563198 380918 563434
rect 381154 563198 381196 563434
rect 380876 556434 381196 563198
rect 380876 556198 380918 556434
rect 381154 556198 381196 556434
rect 380876 549434 381196 556198
rect 380876 549198 380918 549434
rect 381154 549198 381196 549434
rect 380876 542434 381196 549198
rect 380876 542198 380918 542434
rect 381154 542198 381196 542434
rect 380876 535434 381196 542198
rect 380876 535198 380918 535434
rect 381154 535198 381196 535434
rect 380876 528434 381196 535198
rect 380876 528198 380918 528434
rect 381154 528198 381196 528434
rect 380876 521434 381196 528198
rect 380876 521198 380918 521434
rect 381154 521198 381196 521434
rect 380876 514434 381196 521198
rect 380876 514198 380918 514434
rect 381154 514198 381196 514434
rect 380876 507434 381196 514198
rect 380876 507198 380918 507434
rect 381154 507198 381196 507434
rect 380876 500434 381196 507198
rect 380876 500198 380918 500434
rect 381154 500198 381196 500434
rect 380876 493434 381196 500198
rect 380876 493198 380918 493434
rect 381154 493198 381196 493434
rect 380876 486434 381196 493198
rect 380876 486198 380918 486434
rect 381154 486198 381196 486434
rect 380876 479434 381196 486198
rect 380876 479198 380918 479434
rect 381154 479198 381196 479434
rect 380876 472434 381196 479198
rect 380876 472198 380918 472434
rect 381154 472198 381196 472434
rect 380876 465434 381196 472198
rect 380876 465198 380918 465434
rect 381154 465198 381196 465434
rect 380876 458434 381196 465198
rect 380876 458198 380918 458434
rect 381154 458198 381196 458434
rect 380876 451434 381196 458198
rect 380876 451198 380918 451434
rect 381154 451198 381196 451434
rect 380876 444434 381196 451198
rect 380876 444198 380918 444434
rect 381154 444198 381196 444434
rect 380876 437434 381196 444198
rect 380876 437198 380918 437434
rect 381154 437198 381196 437434
rect 380876 430434 381196 437198
rect 380876 430198 380918 430434
rect 381154 430198 381196 430434
rect 380876 423434 381196 430198
rect 380876 423198 380918 423434
rect 381154 423198 381196 423434
rect 380876 416434 381196 423198
rect 380876 416198 380918 416434
rect 381154 416198 381196 416434
rect 380876 409434 381196 416198
rect 380876 409198 380918 409434
rect 381154 409198 381196 409434
rect 380876 402434 381196 409198
rect 380876 402198 380918 402434
rect 381154 402198 381196 402434
rect 380876 395434 381196 402198
rect 380876 395198 380918 395434
rect 381154 395198 381196 395434
rect 380876 388434 381196 395198
rect 380876 388198 380918 388434
rect 381154 388198 381196 388434
rect 380876 381434 381196 388198
rect 380876 381198 380918 381434
rect 381154 381198 381196 381434
rect 380876 374434 381196 381198
rect 380876 374198 380918 374434
rect 381154 374198 381196 374434
rect 380876 367434 381196 374198
rect 380876 367198 380918 367434
rect 381154 367198 381196 367434
rect 380876 360434 381196 367198
rect 380876 360198 380918 360434
rect 381154 360198 381196 360434
rect 380876 353434 381196 360198
rect 380876 353198 380918 353434
rect 381154 353198 381196 353434
rect 380876 346434 381196 353198
rect 380876 346198 380918 346434
rect 381154 346198 381196 346434
rect 380876 339434 381196 346198
rect 380876 339198 380918 339434
rect 381154 339198 381196 339434
rect 380876 332434 381196 339198
rect 380876 332198 380918 332434
rect 381154 332198 381196 332434
rect 380876 325434 381196 332198
rect 380876 325198 380918 325434
rect 381154 325198 381196 325434
rect 380876 318434 381196 325198
rect 380876 318198 380918 318434
rect 381154 318198 381196 318434
rect 380876 311434 381196 318198
rect 380876 311198 380918 311434
rect 381154 311198 381196 311434
rect 380876 304434 381196 311198
rect 380876 304198 380918 304434
rect 381154 304198 381196 304434
rect 380876 297434 381196 304198
rect 380876 297198 380918 297434
rect 381154 297198 381196 297434
rect 380876 290434 381196 297198
rect 380876 290198 380918 290434
rect 381154 290198 381196 290434
rect 380876 283434 381196 290198
rect 380876 283198 380918 283434
rect 381154 283198 381196 283434
rect 380876 276434 381196 283198
rect 380876 276198 380918 276434
rect 381154 276198 381196 276434
rect 380876 269434 381196 276198
rect 380876 269198 380918 269434
rect 381154 269198 381196 269434
rect 380876 262434 381196 269198
rect 380876 262198 380918 262434
rect 381154 262198 381196 262434
rect 380876 255434 381196 262198
rect 380876 255198 380918 255434
rect 381154 255198 381196 255434
rect 380876 248434 381196 255198
rect 380876 248198 380918 248434
rect 381154 248198 381196 248434
rect 380876 241434 381196 248198
rect 380876 241198 380918 241434
rect 381154 241198 381196 241434
rect 380876 234434 381196 241198
rect 380876 234198 380918 234434
rect 381154 234198 381196 234434
rect 380876 227434 381196 234198
rect 380876 227198 380918 227434
rect 381154 227198 381196 227434
rect 380876 220434 381196 227198
rect 380876 220198 380918 220434
rect 381154 220198 381196 220434
rect 380876 213434 381196 220198
rect 380876 213198 380918 213434
rect 381154 213198 381196 213434
rect 380876 206434 381196 213198
rect 380876 206198 380918 206434
rect 381154 206198 381196 206434
rect 380876 199434 381196 206198
rect 380876 199198 380918 199434
rect 381154 199198 381196 199434
rect 380876 192434 381196 199198
rect 380876 192198 380918 192434
rect 381154 192198 381196 192434
rect 380876 185434 381196 192198
rect 380876 185198 380918 185434
rect 381154 185198 381196 185434
rect 380876 178434 381196 185198
rect 380876 178198 380918 178434
rect 381154 178198 381196 178434
rect 380876 171434 381196 178198
rect 380876 171198 380918 171434
rect 381154 171198 381196 171434
rect 380876 164434 381196 171198
rect 380876 164198 380918 164434
rect 381154 164198 381196 164434
rect 380876 157434 381196 164198
rect 380876 157198 380918 157434
rect 381154 157198 381196 157434
rect 380876 150434 381196 157198
rect 380876 150198 380918 150434
rect 381154 150198 381196 150434
rect 380876 143434 381196 150198
rect 380876 143198 380918 143434
rect 381154 143198 381196 143434
rect 380876 136434 381196 143198
rect 380876 136198 380918 136434
rect 381154 136198 381196 136434
rect 380876 129434 381196 136198
rect 380876 129198 380918 129434
rect 381154 129198 381196 129434
rect 380876 122434 381196 129198
rect 380876 122198 380918 122434
rect 381154 122198 381196 122434
rect 380876 115434 381196 122198
rect 380876 115198 380918 115434
rect 381154 115198 381196 115434
rect 380876 108434 381196 115198
rect 380876 108198 380918 108434
rect 381154 108198 381196 108434
rect 380876 101434 381196 108198
rect 380876 101198 380918 101434
rect 381154 101198 381196 101434
rect 380876 94434 381196 101198
rect 380876 94198 380918 94434
rect 381154 94198 381196 94434
rect 380876 87434 381196 94198
rect 380876 87198 380918 87434
rect 381154 87198 381196 87434
rect 380876 80434 381196 87198
rect 380876 80198 380918 80434
rect 381154 80198 381196 80434
rect 380876 73434 381196 80198
rect 380876 73198 380918 73434
rect 381154 73198 381196 73434
rect 380876 66434 381196 73198
rect 380876 66198 380918 66434
rect 381154 66198 381196 66434
rect 380876 59434 381196 66198
rect 380876 59198 380918 59434
rect 381154 59198 381196 59434
rect 380876 52434 381196 59198
rect 380876 52198 380918 52434
rect 381154 52198 381196 52434
rect 380876 45434 381196 52198
rect 380876 45198 380918 45434
rect 381154 45198 381196 45434
rect 380876 38434 381196 45198
rect 380876 38198 380918 38434
rect 381154 38198 381196 38434
rect 380876 31434 381196 38198
rect 380876 31198 380918 31434
rect 381154 31198 381196 31434
rect 380876 24434 381196 31198
rect 380876 24198 380918 24434
rect 381154 24198 381196 24434
rect 380876 17434 381196 24198
rect 380876 17198 380918 17434
rect 381154 17198 381196 17434
rect 380876 10434 381196 17198
rect 380876 10198 380918 10434
rect 381154 10198 381196 10434
rect 380876 3434 381196 10198
rect 380876 3198 380918 3434
rect 381154 3198 381196 3434
rect 380876 -1706 381196 3198
rect 380876 -1942 380918 -1706
rect 381154 -1942 381196 -1706
rect 380876 -2026 381196 -1942
rect 380876 -2262 380918 -2026
rect 381154 -2262 381196 -2026
rect 380876 -2294 381196 -2262
rect 386144 705238 386464 706230
rect 386144 705002 386186 705238
rect 386422 705002 386464 705238
rect 386144 704918 386464 705002
rect 386144 704682 386186 704918
rect 386422 704682 386464 704918
rect 386144 695494 386464 704682
rect 386144 695258 386186 695494
rect 386422 695258 386464 695494
rect 386144 688494 386464 695258
rect 386144 688258 386186 688494
rect 386422 688258 386464 688494
rect 386144 681494 386464 688258
rect 386144 681258 386186 681494
rect 386422 681258 386464 681494
rect 386144 674494 386464 681258
rect 386144 674258 386186 674494
rect 386422 674258 386464 674494
rect 386144 667494 386464 674258
rect 386144 667258 386186 667494
rect 386422 667258 386464 667494
rect 386144 660494 386464 667258
rect 386144 660258 386186 660494
rect 386422 660258 386464 660494
rect 386144 653494 386464 660258
rect 386144 653258 386186 653494
rect 386422 653258 386464 653494
rect 386144 646494 386464 653258
rect 386144 646258 386186 646494
rect 386422 646258 386464 646494
rect 386144 639494 386464 646258
rect 386144 639258 386186 639494
rect 386422 639258 386464 639494
rect 386144 632494 386464 639258
rect 386144 632258 386186 632494
rect 386422 632258 386464 632494
rect 386144 625494 386464 632258
rect 386144 625258 386186 625494
rect 386422 625258 386464 625494
rect 386144 618494 386464 625258
rect 386144 618258 386186 618494
rect 386422 618258 386464 618494
rect 386144 611494 386464 618258
rect 386144 611258 386186 611494
rect 386422 611258 386464 611494
rect 386144 604494 386464 611258
rect 386144 604258 386186 604494
rect 386422 604258 386464 604494
rect 386144 597494 386464 604258
rect 386144 597258 386186 597494
rect 386422 597258 386464 597494
rect 386144 590494 386464 597258
rect 386144 590258 386186 590494
rect 386422 590258 386464 590494
rect 386144 583494 386464 590258
rect 386144 583258 386186 583494
rect 386422 583258 386464 583494
rect 386144 576494 386464 583258
rect 386144 576258 386186 576494
rect 386422 576258 386464 576494
rect 386144 569494 386464 576258
rect 386144 569258 386186 569494
rect 386422 569258 386464 569494
rect 386144 562494 386464 569258
rect 386144 562258 386186 562494
rect 386422 562258 386464 562494
rect 386144 555494 386464 562258
rect 386144 555258 386186 555494
rect 386422 555258 386464 555494
rect 386144 548494 386464 555258
rect 386144 548258 386186 548494
rect 386422 548258 386464 548494
rect 386144 541494 386464 548258
rect 386144 541258 386186 541494
rect 386422 541258 386464 541494
rect 386144 534494 386464 541258
rect 386144 534258 386186 534494
rect 386422 534258 386464 534494
rect 386144 527494 386464 534258
rect 386144 527258 386186 527494
rect 386422 527258 386464 527494
rect 386144 520494 386464 527258
rect 386144 520258 386186 520494
rect 386422 520258 386464 520494
rect 386144 513494 386464 520258
rect 386144 513258 386186 513494
rect 386422 513258 386464 513494
rect 386144 506494 386464 513258
rect 386144 506258 386186 506494
rect 386422 506258 386464 506494
rect 386144 499494 386464 506258
rect 386144 499258 386186 499494
rect 386422 499258 386464 499494
rect 386144 492494 386464 499258
rect 386144 492258 386186 492494
rect 386422 492258 386464 492494
rect 386144 485494 386464 492258
rect 386144 485258 386186 485494
rect 386422 485258 386464 485494
rect 386144 478494 386464 485258
rect 386144 478258 386186 478494
rect 386422 478258 386464 478494
rect 386144 471494 386464 478258
rect 386144 471258 386186 471494
rect 386422 471258 386464 471494
rect 386144 464494 386464 471258
rect 386144 464258 386186 464494
rect 386422 464258 386464 464494
rect 386144 457494 386464 464258
rect 386144 457258 386186 457494
rect 386422 457258 386464 457494
rect 386144 450494 386464 457258
rect 386144 450258 386186 450494
rect 386422 450258 386464 450494
rect 386144 443494 386464 450258
rect 386144 443258 386186 443494
rect 386422 443258 386464 443494
rect 386144 436494 386464 443258
rect 386144 436258 386186 436494
rect 386422 436258 386464 436494
rect 386144 429494 386464 436258
rect 386144 429258 386186 429494
rect 386422 429258 386464 429494
rect 386144 422494 386464 429258
rect 386144 422258 386186 422494
rect 386422 422258 386464 422494
rect 386144 415494 386464 422258
rect 386144 415258 386186 415494
rect 386422 415258 386464 415494
rect 386144 408494 386464 415258
rect 386144 408258 386186 408494
rect 386422 408258 386464 408494
rect 386144 401494 386464 408258
rect 386144 401258 386186 401494
rect 386422 401258 386464 401494
rect 386144 394494 386464 401258
rect 386144 394258 386186 394494
rect 386422 394258 386464 394494
rect 386144 387494 386464 394258
rect 386144 387258 386186 387494
rect 386422 387258 386464 387494
rect 386144 380494 386464 387258
rect 386144 380258 386186 380494
rect 386422 380258 386464 380494
rect 386144 373494 386464 380258
rect 386144 373258 386186 373494
rect 386422 373258 386464 373494
rect 386144 366494 386464 373258
rect 386144 366258 386186 366494
rect 386422 366258 386464 366494
rect 386144 359494 386464 366258
rect 386144 359258 386186 359494
rect 386422 359258 386464 359494
rect 386144 352494 386464 359258
rect 386144 352258 386186 352494
rect 386422 352258 386464 352494
rect 386144 345494 386464 352258
rect 386144 345258 386186 345494
rect 386422 345258 386464 345494
rect 386144 338494 386464 345258
rect 386144 338258 386186 338494
rect 386422 338258 386464 338494
rect 386144 331494 386464 338258
rect 386144 331258 386186 331494
rect 386422 331258 386464 331494
rect 386144 324494 386464 331258
rect 386144 324258 386186 324494
rect 386422 324258 386464 324494
rect 386144 317494 386464 324258
rect 386144 317258 386186 317494
rect 386422 317258 386464 317494
rect 386144 310494 386464 317258
rect 386144 310258 386186 310494
rect 386422 310258 386464 310494
rect 386144 303494 386464 310258
rect 386144 303258 386186 303494
rect 386422 303258 386464 303494
rect 386144 296494 386464 303258
rect 386144 296258 386186 296494
rect 386422 296258 386464 296494
rect 386144 289494 386464 296258
rect 386144 289258 386186 289494
rect 386422 289258 386464 289494
rect 386144 282494 386464 289258
rect 386144 282258 386186 282494
rect 386422 282258 386464 282494
rect 386144 275494 386464 282258
rect 386144 275258 386186 275494
rect 386422 275258 386464 275494
rect 386144 268494 386464 275258
rect 386144 268258 386186 268494
rect 386422 268258 386464 268494
rect 386144 261494 386464 268258
rect 386144 261258 386186 261494
rect 386422 261258 386464 261494
rect 386144 254494 386464 261258
rect 386144 254258 386186 254494
rect 386422 254258 386464 254494
rect 386144 247494 386464 254258
rect 386144 247258 386186 247494
rect 386422 247258 386464 247494
rect 386144 240494 386464 247258
rect 386144 240258 386186 240494
rect 386422 240258 386464 240494
rect 386144 233494 386464 240258
rect 386144 233258 386186 233494
rect 386422 233258 386464 233494
rect 386144 226494 386464 233258
rect 386144 226258 386186 226494
rect 386422 226258 386464 226494
rect 386144 219494 386464 226258
rect 386144 219258 386186 219494
rect 386422 219258 386464 219494
rect 386144 212494 386464 219258
rect 386144 212258 386186 212494
rect 386422 212258 386464 212494
rect 386144 205494 386464 212258
rect 386144 205258 386186 205494
rect 386422 205258 386464 205494
rect 386144 198494 386464 205258
rect 386144 198258 386186 198494
rect 386422 198258 386464 198494
rect 386144 191494 386464 198258
rect 386144 191258 386186 191494
rect 386422 191258 386464 191494
rect 386144 184494 386464 191258
rect 386144 184258 386186 184494
rect 386422 184258 386464 184494
rect 386144 177494 386464 184258
rect 386144 177258 386186 177494
rect 386422 177258 386464 177494
rect 386144 170494 386464 177258
rect 386144 170258 386186 170494
rect 386422 170258 386464 170494
rect 386144 163494 386464 170258
rect 386144 163258 386186 163494
rect 386422 163258 386464 163494
rect 386144 156494 386464 163258
rect 386144 156258 386186 156494
rect 386422 156258 386464 156494
rect 386144 149494 386464 156258
rect 386144 149258 386186 149494
rect 386422 149258 386464 149494
rect 386144 142494 386464 149258
rect 386144 142258 386186 142494
rect 386422 142258 386464 142494
rect 386144 135494 386464 142258
rect 386144 135258 386186 135494
rect 386422 135258 386464 135494
rect 386144 128494 386464 135258
rect 386144 128258 386186 128494
rect 386422 128258 386464 128494
rect 386144 121494 386464 128258
rect 386144 121258 386186 121494
rect 386422 121258 386464 121494
rect 386144 114494 386464 121258
rect 386144 114258 386186 114494
rect 386422 114258 386464 114494
rect 386144 107494 386464 114258
rect 386144 107258 386186 107494
rect 386422 107258 386464 107494
rect 386144 100494 386464 107258
rect 386144 100258 386186 100494
rect 386422 100258 386464 100494
rect 386144 93494 386464 100258
rect 386144 93258 386186 93494
rect 386422 93258 386464 93494
rect 386144 86494 386464 93258
rect 386144 86258 386186 86494
rect 386422 86258 386464 86494
rect 386144 79494 386464 86258
rect 386144 79258 386186 79494
rect 386422 79258 386464 79494
rect 386144 72494 386464 79258
rect 386144 72258 386186 72494
rect 386422 72258 386464 72494
rect 386144 65494 386464 72258
rect 386144 65258 386186 65494
rect 386422 65258 386464 65494
rect 386144 58494 386464 65258
rect 386144 58258 386186 58494
rect 386422 58258 386464 58494
rect 386144 51494 386464 58258
rect 386144 51258 386186 51494
rect 386422 51258 386464 51494
rect 386144 44494 386464 51258
rect 386144 44258 386186 44494
rect 386422 44258 386464 44494
rect 386144 37494 386464 44258
rect 386144 37258 386186 37494
rect 386422 37258 386464 37494
rect 386144 30494 386464 37258
rect 386144 30258 386186 30494
rect 386422 30258 386464 30494
rect 386144 23494 386464 30258
rect 386144 23258 386186 23494
rect 386422 23258 386464 23494
rect 386144 16494 386464 23258
rect 386144 16258 386186 16494
rect 386422 16258 386464 16494
rect 386144 9494 386464 16258
rect 386144 9258 386186 9494
rect 386422 9258 386464 9494
rect 386144 2494 386464 9258
rect 386144 2258 386186 2494
rect 386422 2258 386464 2494
rect 386144 -746 386464 2258
rect 386144 -982 386186 -746
rect 386422 -982 386464 -746
rect 386144 -1066 386464 -982
rect 386144 -1302 386186 -1066
rect 386422 -1302 386464 -1066
rect 386144 -2294 386464 -1302
rect 387876 706198 388196 706230
rect 387876 705962 387918 706198
rect 388154 705962 388196 706198
rect 387876 705878 388196 705962
rect 387876 705642 387918 705878
rect 388154 705642 388196 705878
rect 387876 696434 388196 705642
rect 387876 696198 387918 696434
rect 388154 696198 388196 696434
rect 387876 689434 388196 696198
rect 387876 689198 387918 689434
rect 388154 689198 388196 689434
rect 387876 682434 388196 689198
rect 387876 682198 387918 682434
rect 388154 682198 388196 682434
rect 387876 675434 388196 682198
rect 387876 675198 387918 675434
rect 388154 675198 388196 675434
rect 387876 668434 388196 675198
rect 387876 668198 387918 668434
rect 388154 668198 388196 668434
rect 387876 661434 388196 668198
rect 387876 661198 387918 661434
rect 388154 661198 388196 661434
rect 387876 654434 388196 661198
rect 387876 654198 387918 654434
rect 388154 654198 388196 654434
rect 387876 647434 388196 654198
rect 387876 647198 387918 647434
rect 388154 647198 388196 647434
rect 387876 640434 388196 647198
rect 387876 640198 387918 640434
rect 388154 640198 388196 640434
rect 387876 633434 388196 640198
rect 387876 633198 387918 633434
rect 388154 633198 388196 633434
rect 387876 626434 388196 633198
rect 387876 626198 387918 626434
rect 388154 626198 388196 626434
rect 387876 619434 388196 626198
rect 387876 619198 387918 619434
rect 388154 619198 388196 619434
rect 387876 612434 388196 619198
rect 387876 612198 387918 612434
rect 388154 612198 388196 612434
rect 387876 605434 388196 612198
rect 387876 605198 387918 605434
rect 388154 605198 388196 605434
rect 387876 598434 388196 605198
rect 387876 598198 387918 598434
rect 388154 598198 388196 598434
rect 387876 591434 388196 598198
rect 387876 591198 387918 591434
rect 388154 591198 388196 591434
rect 387876 584434 388196 591198
rect 387876 584198 387918 584434
rect 388154 584198 388196 584434
rect 387876 577434 388196 584198
rect 387876 577198 387918 577434
rect 388154 577198 388196 577434
rect 387876 570434 388196 577198
rect 387876 570198 387918 570434
rect 388154 570198 388196 570434
rect 387876 563434 388196 570198
rect 387876 563198 387918 563434
rect 388154 563198 388196 563434
rect 387876 556434 388196 563198
rect 387876 556198 387918 556434
rect 388154 556198 388196 556434
rect 387876 549434 388196 556198
rect 387876 549198 387918 549434
rect 388154 549198 388196 549434
rect 387876 542434 388196 549198
rect 387876 542198 387918 542434
rect 388154 542198 388196 542434
rect 387876 535434 388196 542198
rect 387876 535198 387918 535434
rect 388154 535198 388196 535434
rect 387876 528434 388196 535198
rect 387876 528198 387918 528434
rect 388154 528198 388196 528434
rect 387876 521434 388196 528198
rect 387876 521198 387918 521434
rect 388154 521198 388196 521434
rect 387876 514434 388196 521198
rect 387876 514198 387918 514434
rect 388154 514198 388196 514434
rect 387876 507434 388196 514198
rect 387876 507198 387918 507434
rect 388154 507198 388196 507434
rect 387876 500434 388196 507198
rect 387876 500198 387918 500434
rect 388154 500198 388196 500434
rect 387876 493434 388196 500198
rect 387876 493198 387918 493434
rect 388154 493198 388196 493434
rect 387876 486434 388196 493198
rect 387876 486198 387918 486434
rect 388154 486198 388196 486434
rect 387876 479434 388196 486198
rect 387876 479198 387918 479434
rect 388154 479198 388196 479434
rect 387876 472434 388196 479198
rect 387876 472198 387918 472434
rect 388154 472198 388196 472434
rect 387876 465434 388196 472198
rect 387876 465198 387918 465434
rect 388154 465198 388196 465434
rect 387876 458434 388196 465198
rect 387876 458198 387918 458434
rect 388154 458198 388196 458434
rect 387876 451434 388196 458198
rect 387876 451198 387918 451434
rect 388154 451198 388196 451434
rect 387876 444434 388196 451198
rect 387876 444198 387918 444434
rect 388154 444198 388196 444434
rect 387876 437434 388196 444198
rect 387876 437198 387918 437434
rect 388154 437198 388196 437434
rect 387876 430434 388196 437198
rect 387876 430198 387918 430434
rect 388154 430198 388196 430434
rect 387876 423434 388196 430198
rect 387876 423198 387918 423434
rect 388154 423198 388196 423434
rect 387876 416434 388196 423198
rect 387876 416198 387918 416434
rect 388154 416198 388196 416434
rect 387876 409434 388196 416198
rect 387876 409198 387918 409434
rect 388154 409198 388196 409434
rect 387876 402434 388196 409198
rect 387876 402198 387918 402434
rect 388154 402198 388196 402434
rect 387876 395434 388196 402198
rect 387876 395198 387918 395434
rect 388154 395198 388196 395434
rect 387876 388434 388196 395198
rect 387876 388198 387918 388434
rect 388154 388198 388196 388434
rect 387876 381434 388196 388198
rect 387876 381198 387918 381434
rect 388154 381198 388196 381434
rect 387876 374434 388196 381198
rect 387876 374198 387918 374434
rect 388154 374198 388196 374434
rect 387876 367434 388196 374198
rect 387876 367198 387918 367434
rect 388154 367198 388196 367434
rect 387876 360434 388196 367198
rect 387876 360198 387918 360434
rect 388154 360198 388196 360434
rect 387876 353434 388196 360198
rect 387876 353198 387918 353434
rect 388154 353198 388196 353434
rect 387876 346434 388196 353198
rect 387876 346198 387918 346434
rect 388154 346198 388196 346434
rect 387876 339434 388196 346198
rect 387876 339198 387918 339434
rect 388154 339198 388196 339434
rect 387876 332434 388196 339198
rect 387876 332198 387918 332434
rect 388154 332198 388196 332434
rect 387876 325434 388196 332198
rect 387876 325198 387918 325434
rect 388154 325198 388196 325434
rect 387876 318434 388196 325198
rect 387876 318198 387918 318434
rect 388154 318198 388196 318434
rect 387876 311434 388196 318198
rect 387876 311198 387918 311434
rect 388154 311198 388196 311434
rect 387876 304434 388196 311198
rect 387876 304198 387918 304434
rect 388154 304198 388196 304434
rect 387876 297434 388196 304198
rect 387876 297198 387918 297434
rect 388154 297198 388196 297434
rect 387876 290434 388196 297198
rect 387876 290198 387918 290434
rect 388154 290198 388196 290434
rect 387876 283434 388196 290198
rect 387876 283198 387918 283434
rect 388154 283198 388196 283434
rect 387876 276434 388196 283198
rect 387876 276198 387918 276434
rect 388154 276198 388196 276434
rect 387876 269434 388196 276198
rect 387876 269198 387918 269434
rect 388154 269198 388196 269434
rect 387876 262434 388196 269198
rect 387876 262198 387918 262434
rect 388154 262198 388196 262434
rect 387876 255434 388196 262198
rect 387876 255198 387918 255434
rect 388154 255198 388196 255434
rect 387876 248434 388196 255198
rect 387876 248198 387918 248434
rect 388154 248198 388196 248434
rect 387876 241434 388196 248198
rect 387876 241198 387918 241434
rect 388154 241198 388196 241434
rect 387876 234434 388196 241198
rect 387876 234198 387918 234434
rect 388154 234198 388196 234434
rect 387876 227434 388196 234198
rect 387876 227198 387918 227434
rect 388154 227198 388196 227434
rect 387876 220434 388196 227198
rect 387876 220198 387918 220434
rect 388154 220198 388196 220434
rect 387876 213434 388196 220198
rect 387876 213198 387918 213434
rect 388154 213198 388196 213434
rect 387876 206434 388196 213198
rect 387876 206198 387918 206434
rect 388154 206198 388196 206434
rect 387876 199434 388196 206198
rect 387876 199198 387918 199434
rect 388154 199198 388196 199434
rect 387876 192434 388196 199198
rect 387876 192198 387918 192434
rect 388154 192198 388196 192434
rect 387876 185434 388196 192198
rect 387876 185198 387918 185434
rect 388154 185198 388196 185434
rect 387876 178434 388196 185198
rect 387876 178198 387918 178434
rect 388154 178198 388196 178434
rect 387876 171434 388196 178198
rect 387876 171198 387918 171434
rect 388154 171198 388196 171434
rect 387876 164434 388196 171198
rect 387876 164198 387918 164434
rect 388154 164198 388196 164434
rect 387876 157434 388196 164198
rect 387876 157198 387918 157434
rect 388154 157198 388196 157434
rect 387876 150434 388196 157198
rect 387876 150198 387918 150434
rect 388154 150198 388196 150434
rect 387876 143434 388196 150198
rect 387876 143198 387918 143434
rect 388154 143198 388196 143434
rect 387876 136434 388196 143198
rect 387876 136198 387918 136434
rect 388154 136198 388196 136434
rect 387876 129434 388196 136198
rect 387876 129198 387918 129434
rect 388154 129198 388196 129434
rect 387876 122434 388196 129198
rect 387876 122198 387918 122434
rect 388154 122198 388196 122434
rect 387876 115434 388196 122198
rect 387876 115198 387918 115434
rect 388154 115198 388196 115434
rect 387876 108434 388196 115198
rect 387876 108198 387918 108434
rect 388154 108198 388196 108434
rect 387876 101434 388196 108198
rect 387876 101198 387918 101434
rect 388154 101198 388196 101434
rect 387876 94434 388196 101198
rect 387876 94198 387918 94434
rect 388154 94198 388196 94434
rect 387876 87434 388196 94198
rect 387876 87198 387918 87434
rect 388154 87198 388196 87434
rect 387876 80434 388196 87198
rect 387876 80198 387918 80434
rect 388154 80198 388196 80434
rect 387876 73434 388196 80198
rect 387876 73198 387918 73434
rect 388154 73198 388196 73434
rect 387876 66434 388196 73198
rect 387876 66198 387918 66434
rect 388154 66198 388196 66434
rect 387876 59434 388196 66198
rect 387876 59198 387918 59434
rect 388154 59198 388196 59434
rect 387876 52434 388196 59198
rect 387876 52198 387918 52434
rect 388154 52198 388196 52434
rect 387876 45434 388196 52198
rect 387876 45198 387918 45434
rect 388154 45198 388196 45434
rect 387876 38434 388196 45198
rect 387876 38198 387918 38434
rect 388154 38198 388196 38434
rect 387876 31434 388196 38198
rect 387876 31198 387918 31434
rect 388154 31198 388196 31434
rect 387876 24434 388196 31198
rect 387876 24198 387918 24434
rect 388154 24198 388196 24434
rect 387876 17434 388196 24198
rect 387876 17198 387918 17434
rect 388154 17198 388196 17434
rect 387876 10434 388196 17198
rect 387876 10198 387918 10434
rect 388154 10198 388196 10434
rect 387876 3434 388196 10198
rect 387876 3198 387918 3434
rect 388154 3198 388196 3434
rect 387876 -1706 388196 3198
rect 387876 -1942 387918 -1706
rect 388154 -1942 388196 -1706
rect 387876 -2026 388196 -1942
rect 387876 -2262 387918 -2026
rect 388154 -2262 388196 -2026
rect 387876 -2294 388196 -2262
rect 393144 705238 393464 706230
rect 393144 705002 393186 705238
rect 393422 705002 393464 705238
rect 393144 704918 393464 705002
rect 393144 704682 393186 704918
rect 393422 704682 393464 704918
rect 393144 695494 393464 704682
rect 393144 695258 393186 695494
rect 393422 695258 393464 695494
rect 393144 688494 393464 695258
rect 393144 688258 393186 688494
rect 393422 688258 393464 688494
rect 393144 681494 393464 688258
rect 393144 681258 393186 681494
rect 393422 681258 393464 681494
rect 393144 674494 393464 681258
rect 393144 674258 393186 674494
rect 393422 674258 393464 674494
rect 393144 667494 393464 674258
rect 393144 667258 393186 667494
rect 393422 667258 393464 667494
rect 393144 660494 393464 667258
rect 393144 660258 393186 660494
rect 393422 660258 393464 660494
rect 393144 653494 393464 660258
rect 393144 653258 393186 653494
rect 393422 653258 393464 653494
rect 393144 646494 393464 653258
rect 393144 646258 393186 646494
rect 393422 646258 393464 646494
rect 393144 639494 393464 646258
rect 393144 639258 393186 639494
rect 393422 639258 393464 639494
rect 393144 632494 393464 639258
rect 393144 632258 393186 632494
rect 393422 632258 393464 632494
rect 393144 625494 393464 632258
rect 393144 625258 393186 625494
rect 393422 625258 393464 625494
rect 393144 618494 393464 625258
rect 393144 618258 393186 618494
rect 393422 618258 393464 618494
rect 393144 611494 393464 618258
rect 393144 611258 393186 611494
rect 393422 611258 393464 611494
rect 393144 604494 393464 611258
rect 393144 604258 393186 604494
rect 393422 604258 393464 604494
rect 393144 597494 393464 604258
rect 393144 597258 393186 597494
rect 393422 597258 393464 597494
rect 393144 590494 393464 597258
rect 393144 590258 393186 590494
rect 393422 590258 393464 590494
rect 393144 583494 393464 590258
rect 393144 583258 393186 583494
rect 393422 583258 393464 583494
rect 393144 576494 393464 583258
rect 393144 576258 393186 576494
rect 393422 576258 393464 576494
rect 393144 569494 393464 576258
rect 393144 569258 393186 569494
rect 393422 569258 393464 569494
rect 393144 562494 393464 569258
rect 393144 562258 393186 562494
rect 393422 562258 393464 562494
rect 393144 555494 393464 562258
rect 393144 555258 393186 555494
rect 393422 555258 393464 555494
rect 393144 548494 393464 555258
rect 393144 548258 393186 548494
rect 393422 548258 393464 548494
rect 393144 541494 393464 548258
rect 393144 541258 393186 541494
rect 393422 541258 393464 541494
rect 393144 534494 393464 541258
rect 393144 534258 393186 534494
rect 393422 534258 393464 534494
rect 393144 527494 393464 534258
rect 393144 527258 393186 527494
rect 393422 527258 393464 527494
rect 393144 520494 393464 527258
rect 393144 520258 393186 520494
rect 393422 520258 393464 520494
rect 393144 513494 393464 520258
rect 393144 513258 393186 513494
rect 393422 513258 393464 513494
rect 393144 506494 393464 513258
rect 393144 506258 393186 506494
rect 393422 506258 393464 506494
rect 393144 499494 393464 506258
rect 393144 499258 393186 499494
rect 393422 499258 393464 499494
rect 393144 492494 393464 499258
rect 393144 492258 393186 492494
rect 393422 492258 393464 492494
rect 393144 485494 393464 492258
rect 393144 485258 393186 485494
rect 393422 485258 393464 485494
rect 393144 478494 393464 485258
rect 393144 478258 393186 478494
rect 393422 478258 393464 478494
rect 393144 471494 393464 478258
rect 393144 471258 393186 471494
rect 393422 471258 393464 471494
rect 393144 464494 393464 471258
rect 393144 464258 393186 464494
rect 393422 464258 393464 464494
rect 393144 457494 393464 464258
rect 393144 457258 393186 457494
rect 393422 457258 393464 457494
rect 393144 450494 393464 457258
rect 393144 450258 393186 450494
rect 393422 450258 393464 450494
rect 393144 443494 393464 450258
rect 393144 443258 393186 443494
rect 393422 443258 393464 443494
rect 393144 436494 393464 443258
rect 393144 436258 393186 436494
rect 393422 436258 393464 436494
rect 393144 429494 393464 436258
rect 393144 429258 393186 429494
rect 393422 429258 393464 429494
rect 393144 422494 393464 429258
rect 393144 422258 393186 422494
rect 393422 422258 393464 422494
rect 393144 415494 393464 422258
rect 393144 415258 393186 415494
rect 393422 415258 393464 415494
rect 393144 408494 393464 415258
rect 393144 408258 393186 408494
rect 393422 408258 393464 408494
rect 393144 401494 393464 408258
rect 393144 401258 393186 401494
rect 393422 401258 393464 401494
rect 393144 394494 393464 401258
rect 393144 394258 393186 394494
rect 393422 394258 393464 394494
rect 393144 387494 393464 394258
rect 393144 387258 393186 387494
rect 393422 387258 393464 387494
rect 393144 380494 393464 387258
rect 393144 380258 393186 380494
rect 393422 380258 393464 380494
rect 393144 373494 393464 380258
rect 393144 373258 393186 373494
rect 393422 373258 393464 373494
rect 393144 366494 393464 373258
rect 393144 366258 393186 366494
rect 393422 366258 393464 366494
rect 393144 359494 393464 366258
rect 393144 359258 393186 359494
rect 393422 359258 393464 359494
rect 393144 352494 393464 359258
rect 393144 352258 393186 352494
rect 393422 352258 393464 352494
rect 393144 345494 393464 352258
rect 393144 345258 393186 345494
rect 393422 345258 393464 345494
rect 393144 338494 393464 345258
rect 393144 338258 393186 338494
rect 393422 338258 393464 338494
rect 393144 331494 393464 338258
rect 393144 331258 393186 331494
rect 393422 331258 393464 331494
rect 393144 324494 393464 331258
rect 393144 324258 393186 324494
rect 393422 324258 393464 324494
rect 393144 317494 393464 324258
rect 393144 317258 393186 317494
rect 393422 317258 393464 317494
rect 393144 310494 393464 317258
rect 393144 310258 393186 310494
rect 393422 310258 393464 310494
rect 393144 303494 393464 310258
rect 393144 303258 393186 303494
rect 393422 303258 393464 303494
rect 393144 296494 393464 303258
rect 393144 296258 393186 296494
rect 393422 296258 393464 296494
rect 393144 289494 393464 296258
rect 393144 289258 393186 289494
rect 393422 289258 393464 289494
rect 393144 282494 393464 289258
rect 393144 282258 393186 282494
rect 393422 282258 393464 282494
rect 393144 275494 393464 282258
rect 393144 275258 393186 275494
rect 393422 275258 393464 275494
rect 393144 268494 393464 275258
rect 393144 268258 393186 268494
rect 393422 268258 393464 268494
rect 393144 261494 393464 268258
rect 393144 261258 393186 261494
rect 393422 261258 393464 261494
rect 393144 254494 393464 261258
rect 393144 254258 393186 254494
rect 393422 254258 393464 254494
rect 393144 247494 393464 254258
rect 393144 247258 393186 247494
rect 393422 247258 393464 247494
rect 393144 240494 393464 247258
rect 393144 240258 393186 240494
rect 393422 240258 393464 240494
rect 393144 233494 393464 240258
rect 393144 233258 393186 233494
rect 393422 233258 393464 233494
rect 393144 226494 393464 233258
rect 393144 226258 393186 226494
rect 393422 226258 393464 226494
rect 393144 219494 393464 226258
rect 393144 219258 393186 219494
rect 393422 219258 393464 219494
rect 393144 212494 393464 219258
rect 393144 212258 393186 212494
rect 393422 212258 393464 212494
rect 393144 205494 393464 212258
rect 393144 205258 393186 205494
rect 393422 205258 393464 205494
rect 393144 198494 393464 205258
rect 393144 198258 393186 198494
rect 393422 198258 393464 198494
rect 393144 191494 393464 198258
rect 393144 191258 393186 191494
rect 393422 191258 393464 191494
rect 393144 184494 393464 191258
rect 393144 184258 393186 184494
rect 393422 184258 393464 184494
rect 393144 177494 393464 184258
rect 393144 177258 393186 177494
rect 393422 177258 393464 177494
rect 393144 170494 393464 177258
rect 393144 170258 393186 170494
rect 393422 170258 393464 170494
rect 393144 163494 393464 170258
rect 393144 163258 393186 163494
rect 393422 163258 393464 163494
rect 393144 156494 393464 163258
rect 393144 156258 393186 156494
rect 393422 156258 393464 156494
rect 393144 149494 393464 156258
rect 393144 149258 393186 149494
rect 393422 149258 393464 149494
rect 393144 142494 393464 149258
rect 393144 142258 393186 142494
rect 393422 142258 393464 142494
rect 393144 135494 393464 142258
rect 393144 135258 393186 135494
rect 393422 135258 393464 135494
rect 393144 128494 393464 135258
rect 393144 128258 393186 128494
rect 393422 128258 393464 128494
rect 393144 121494 393464 128258
rect 393144 121258 393186 121494
rect 393422 121258 393464 121494
rect 393144 114494 393464 121258
rect 393144 114258 393186 114494
rect 393422 114258 393464 114494
rect 393144 107494 393464 114258
rect 393144 107258 393186 107494
rect 393422 107258 393464 107494
rect 393144 100494 393464 107258
rect 393144 100258 393186 100494
rect 393422 100258 393464 100494
rect 393144 93494 393464 100258
rect 393144 93258 393186 93494
rect 393422 93258 393464 93494
rect 393144 86494 393464 93258
rect 393144 86258 393186 86494
rect 393422 86258 393464 86494
rect 393144 79494 393464 86258
rect 393144 79258 393186 79494
rect 393422 79258 393464 79494
rect 393144 72494 393464 79258
rect 393144 72258 393186 72494
rect 393422 72258 393464 72494
rect 393144 65494 393464 72258
rect 393144 65258 393186 65494
rect 393422 65258 393464 65494
rect 393144 58494 393464 65258
rect 393144 58258 393186 58494
rect 393422 58258 393464 58494
rect 393144 51494 393464 58258
rect 393144 51258 393186 51494
rect 393422 51258 393464 51494
rect 393144 44494 393464 51258
rect 393144 44258 393186 44494
rect 393422 44258 393464 44494
rect 393144 37494 393464 44258
rect 393144 37258 393186 37494
rect 393422 37258 393464 37494
rect 393144 30494 393464 37258
rect 393144 30258 393186 30494
rect 393422 30258 393464 30494
rect 393144 23494 393464 30258
rect 393144 23258 393186 23494
rect 393422 23258 393464 23494
rect 393144 16494 393464 23258
rect 393144 16258 393186 16494
rect 393422 16258 393464 16494
rect 393144 9494 393464 16258
rect 393144 9258 393186 9494
rect 393422 9258 393464 9494
rect 393144 2494 393464 9258
rect 393144 2258 393186 2494
rect 393422 2258 393464 2494
rect 393144 -746 393464 2258
rect 393144 -982 393186 -746
rect 393422 -982 393464 -746
rect 393144 -1066 393464 -982
rect 393144 -1302 393186 -1066
rect 393422 -1302 393464 -1066
rect 393144 -2294 393464 -1302
rect 394876 706198 395196 706230
rect 394876 705962 394918 706198
rect 395154 705962 395196 706198
rect 394876 705878 395196 705962
rect 394876 705642 394918 705878
rect 395154 705642 395196 705878
rect 394876 696434 395196 705642
rect 394876 696198 394918 696434
rect 395154 696198 395196 696434
rect 394876 689434 395196 696198
rect 394876 689198 394918 689434
rect 395154 689198 395196 689434
rect 394876 682434 395196 689198
rect 394876 682198 394918 682434
rect 395154 682198 395196 682434
rect 394876 675434 395196 682198
rect 394876 675198 394918 675434
rect 395154 675198 395196 675434
rect 394876 668434 395196 675198
rect 394876 668198 394918 668434
rect 395154 668198 395196 668434
rect 394876 661434 395196 668198
rect 394876 661198 394918 661434
rect 395154 661198 395196 661434
rect 394876 654434 395196 661198
rect 394876 654198 394918 654434
rect 395154 654198 395196 654434
rect 394876 647434 395196 654198
rect 394876 647198 394918 647434
rect 395154 647198 395196 647434
rect 394876 640434 395196 647198
rect 394876 640198 394918 640434
rect 395154 640198 395196 640434
rect 394876 633434 395196 640198
rect 394876 633198 394918 633434
rect 395154 633198 395196 633434
rect 394876 626434 395196 633198
rect 394876 626198 394918 626434
rect 395154 626198 395196 626434
rect 394876 619434 395196 626198
rect 394876 619198 394918 619434
rect 395154 619198 395196 619434
rect 394876 612434 395196 619198
rect 394876 612198 394918 612434
rect 395154 612198 395196 612434
rect 394876 605434 395196 612198
rect 394876 605198 394918 605434
rect 395154 605198 395196 605434
rect 394876 598434 395196 605198
rect 394876 598198 394918 598434
rect 395154 598198 395196 598434
rect 394876 591434 395196 598198
rect 394876 591198 394918 591434
rect 395154 591198 395196 591434
rect 394876 584434 395196 591198
rect 394876 584198 394918 584434
rect 395154 584198 395196 584434
rect 394876 577434 395196 584198
rect 394876 577198 394918 577434
rect 395154 577198 395196 577434
rect 394876 570434 395196 577198
rect 394876 570198 394918 570434
rect 395154 570198 395196 570434
rect 394876 563434 395196 570198
rect 394876 563198 394918 563434
rect 395154 563198 395196 563434
rect 394876 556434 395196 563198
rect 394876 556198 394918 556434
rect 395154 556198 395196 556434
rect 394876 549434 395196 556198
rect 394876 549198 394918 549434
rect 395154 549198 395196 549434
rect 394876 542434 395196 549198
rect 394876 542198 394918 542434
rect 395154 542198 395196 542434
rect 394876 535434 395196 542198
rect 394876 535198 394918 535434
rect 395154 535198 395196 535434
rect 394876 528434 395196 535198
rect 394876 528198 394918 528434
rect 395154 528198 395196 528434
rect 394876 521434 395196 528198
rect 394876 521198 394918 521434
rect 395154 521198 395196 521434
rect 394876 514434 395196 521198
rect 394876 514198 394918 514434
rect 395154 514198 395196 514434
rect 394876 507434 395196 514198
rect 394876 507198 394918 507434
rect 395154 507198 395196 507434
rect 394876 500434 395196 507198
rect 394876 500198 394918 500434
rect 395154 500198 395196 500434
rect 394876 493434 395196 500198
rect 394876 493198 394918 493434
rect 395154 493198 395196 493434
rect 394876 486434 395196 493198
rect 394876 486198 394918 486434
rect 395154 486198 395196 486434
rect 394876 479434 395196 486198
rect 394876 479198 394918 479434
rect 395154 479198 395196 479434
rect 394876 472434 395196 479198
rect 394876 472198 394918 472434
rect 395154 472198 395196 472434
rect 394876 465434 395196 472198
rect 394876 465198 394918 465434
rect 395154 465198 395196 465434
rect 394876 458434 395196 465198
rect 394876 458198 394918 458434
rect 395154 458198 395196 458434
rect 394876 451434 395196 458198
rect 394876 451198 394918 451434
rect 395154 451198 395196 451434
rect 394876 444434 395196 451198
rect 394876 444198 394918 444434
rect 395154 444198 395196 444434
rect 394876 437434 395196 444198
rect 394876 437198 394918 437434
rect 395154 437198 395196 437434
rect 394876 430434 395196 437198
rect 394876 430198 394918 430434
rect 395154 430198 395196 430434
rect 394876 423434 395196 430198
rect 394876 423198 394918 423434
rect 395154 423198 395196 423434
rect 394876 416434 395196 423198
rect 394876 416198 394918 416434
rect 395154 416198 395196 416434
rect 394876 409434 395196 416198
rect 394876 409198 394918 409434
rect 395154 409198 395196 409434
rect 394876 402434 395196 409198
rect 394876 402198 394918 402434
rect 395154 402198 395196 402434
rect 394876 395434 395196 402198
rect 394876 395198 394918 395434
rect 395154 395198 395196 395434
rect 394876 388434 395196 395198
rect 394876 388198 394918 388434
rect 395154 388198 395196 388434
rect 394876 381434 395196 388198
rect 394876 381198 394918 381434
rect 395154 381198 395196 381434
rect 394876 374434 395196 381198
rect 394876 374198 394918 374434
rect 395154 374198 395196 374434
rect 394876 367434 395196 374198
rect 394876 367198 394918 367434
rect 395154 367198 395196 367434
rect 394876 360434 395196 367198
rect 394876 360198 394918 360434
rect 395154 360198 395196 360434
rect 394876 353434 395196 360198
rect 394876 353198 394918 353434
rect 395154 353198 395196 353434
rect 394876 346434 395196 353198
rect 394876 346198 394918 346434
rect 395154 346198 395196 346434
rect 394876 339434 395196 346198
rect 394876 339198 394918 339434
rect 395154 339198 395196 339434
rect 394876 332434 395196 339198
rect 394876 332198 394918 332434
rect 395154 332198 395196 332434
rect 394876 325434 395196 332198
rect 394876 325198 394918 325434
rect 395154 325198 395196 325434
rect 394876 318434 395196 325198
rect 394876 318198 394918 318434
rect 395154 318198 395196 318434
rect 394876 311434 395196 318198
rect 394876 311198 394918 311434
rect 395154 311198 395196 311434
rect 394876 304434 395196 311198
rect 394876 304198 394918 304434
rect 395154 304198 395196 304434
rect 394876 297434 395196 304198
rect 394876 297198 394918 297434
rect 395154 297198 395196 297434
rect 394876 290434 395196 297198
rect 394876 290198 394918 290434
rect 395154 290198 395196 290434
rect 394876 283434 395196 290198
rect 394876 283198 394918 283434
rect 395154 283198 395196 283434
rect 394876 276434 395196 283198
rect 394876 276198 394918 276434
rect 395154 276198 395196 276434
rect 394876 269434 395196 276198
rect 394876 269198 394918 269434
rect 395154 269198 395196 269434
rect 394876 262434 395196 269198
rect 394876 262198 394918 262434
rect 395154 262198 395196 262434
rect 394876 255434 395196 262198
rect 394876 255198 394918 255434
rect 395154 255198 395196 255434
rect 394876 248434 395196 255198
rect 394876 248198 394918 248434
rect 395154 248198 395196 248434
rect 394876 241434 395196 248198
rect 394876 241198 394918 241434
rect 395154 241198 395196 241434
rect 394876 234434 395196 241198
rect 394876 234198 394918 234434
rect 395154 234198 395196 234434
rect 394876 227434 395196 234198
rect 394876 227198 394918 227434
rect 395154 227198 395196 227434
rect 394876 220434 395196 227198
rect 394876 220198 394918 220434
rect 395154 220198 395196 220434
rect 394876 213434 395196 220198
rect 394876 213198 394918 213434
rect 395154 213198 395196 213434
rect 394876 206434 395196 213198
rect 394876 206198 394918 206434
rect 395154 206198 395196 206434
rect 394876 199434 395196 206198
rect 394876 199198 394918 199434
rect 395154 199198 395196 199434
rect 394876 192434 395196 199198
rect 394876 192198 394918 192434
rect 395154 192198 395196 192434
rect 394876 185434 395196 192198
rect 394876 185198 394918 185434
rect 395154 185198 395196 185434
rect 394876 178434 395196 185198
rect 394876 178198 394918 178434
rect 395154 178198 395196 178434
rect 394876 171434 395196 178198
rect 394876 171198 394918 171434
rect 395154 171198 395196 171434
rect 394876 164434 395196 171198
rect 394876 164198 394918 164434
rect 395154 164198 395196 164434
rect 394876 157434 395196 164198
rect 394876 157198 394918 157434
rect 395154 157198 395196 157434
rect 394876 150434 395196 157198
rect 394876 150198 394918 150434
rect 395154 150198 395196 150434
rect 394876 143434 395196 150198
rect 394876 143198 394918 143434
rect 395154 143198 395196 143434
rect 394876 136434 395196 143198
rect 394876 136198 394918 136434
rect 395154 136198 395196 136434
rect 394876 129434 395196 136198
rect 394876 129198 394918 129434
rect 395154 129198 395196 129434
rect 394876 122434 395196 129198
rect 394876 122198 394918 122434
rect 395154 122198 395196 122434
rect 394876 115434 395196 122198
rect 394876 115198 394918 115434
rect 395154 115198 395196 115434
rect 394876 108434 395196 115198
rect 394876 108198 394918 108434
rect 395154 108198 395196 108434
rect 394876 101434 395196 108198
rect 394876 101198 394918 101434
rect 395154 101198 395196 101434
rect 394876 94434 395196 101198
rect 394876 94198 394918 94434
rect 395154 94198 395196 94434
rect 394876 87434 395196 94198
rect 394876 87198 394918 87434
rect 395154 87198 395196 87434
rect 394876 80434 395196 87198
rect 394876 80198 394918 80434
rect 395154 80198 395196 80434
rect 394876 73434 395196 80198
rect 394876 73198 394918 73434
rect 395154 73198 395196 73434
rect 394876 66434 395196 73198
rect 394876 66198 394918 66434
rect 395154 66198 395196 66434
rect 394876 59434 395196 66198
rect 394876 59198 394918 59434
rect 395154 59198 395196 59434
rect 394876 52434 395196 59198
rect 394876 52198 394918 52434
rect 395154 52198 395196 52434
rect 394876 45434 395196 52198
rect 394876 45198 394918 45434
rect 395154 45198 395196 45434
rect 394876 38434 395196 45198
rect 394876 38198 394918 38434
rect 395154 38198 395196 38434
rect 394876 31434 395196 38198
rect 394876 31198 394918 31434
rect 395154 31198 395196 31434
rect 394876 24434 395196 31198
rect 394876 24198 394918 24434
rect 395154 24198 395196 24434
rect 394876 17434 395196 24198
rect 394876 17198 394918 17434
rect 395154 17198 395196 17434
rect 394876 10434 395196 17198
rect 394876 10198 394918 10434
rect 395154 10198 395196 10434
rect 394876 3434 395196 10198
rect 394876 3198 394918 3434
rect 395154 3198 395196 3434
rect 394876 -1706 395196 3198
rect 394876 -1942 394918 -1706
rect 395154 -1942 395196 -1706
rect 394876 -2026 395196 -1942
rect 394876 -2262 394918 -2026
rect 395154 -2262 395196 -2026
rect 394876 -2294 395196 -2262
rect 400144 705238 400464 706230
rect 400144 705002 400186 705238
rect 400422 705002 400464 705238
rect 400144 704918 400464 705002
rect 400144 704682 400186 704918
rect 400422 704682 400464 704918
rect 400144 695494 400464 704682
rect 400144 695258 400186 695494
rect 400422 695258 400464 695494
rect 400144 688494 400464 695258
rect 400144 688258 400186 688494
rect 400422 688258 400464 688494
rect 400144 681494 400464 688258
rect 400144 681258 400186 681494
rect 400422 681258 400464 681494
rect 400144 674494 400464 681258
rect 400144 674258 400186 674494
rect 400422 674258 400464 674494
rect 400144 667494 400464 674258
rect 400144 667258 400186 667494
rect 400422 667258 400464 667494
rect 400144 660494 400464 667258
rect 400144 660258 400186 660494
rect 400422 660258 400464 660494
rect 400144 653494 400464 660258
rect 400144 653258 400186 653494
rect 400422 653258 400464 653494
rect 400144 646494 400464 653258
rect 400144 646258 400186 646494
rect 400422 646258 400464 646494
rect 400144 639494 400464 646258
rect 400144 639258 400186 639494
rect 400422 639258 400464 639494
rect 400144 632494 400464 639258
rect 400144 632258 400186 632494
rect 400422 632258 400464 632494
rect 400144 625494 400464 632258
rect 400144 625258 400186 625494
rect 400422 625258 400464 625494
rect 400144 618494 400464 625258
rect 400144 618258 400186 618494
rect 400422 618258 400464 618494
rect 400144 611494 400464 618258
rect 400144 611258 400186 611494
rect 400422 611258 400464 611494
rect 400144 604494 400464 611258
rect 400144 604258 400186 604494
rect 400422 604258 400464 604494
rect 400144 597494 400464 604258
rect 400144 597258 400186 597494
rect 400422 597258 400464 597494
rect 400144 590494 400464 597258
rect 400144 590258 400186 590494
rect 400422 590258 400464 590494
rect 400144 583494 400464 590258
rect 400144 583258 400186 583494
rect 400422 583258 400464 583494
rect 400144 576494 400464 583258
rect 400144 576258 400186 576494
rect 400422 576258 400464 576494
rect 400144 569494 400464 576258
rect 400144 569258 400186 569494
rect 400422 569258 400464 569494
rect 400144 562494 400464 569258
rect 400144 562258 400186 562494
rect 400422 562258 400464 562494
rect 400144 555494 400464 562258
rect 400144 555258 400186 555494
rect 400422 555258 400464 555494
rect 400144 548494 400464 555258
rect 400144 548258 400186 548494
rect 400422 548258 400464 548494
rect 400144 541494 400464 548258
rect 400144 541258 400186 541494
rect 400422 541258 400464 541494
rect 400144 534494 400464 541258
rect 400144 534258 400186 534494
rect 400422 534258 400464 534494
rect 400144 527494 400464 534258
rect 400144 527258 400186 527494
rect 400422 527258 400464 527494
rect 400144 520494 400464 527258
rect 400144 520258 400186 520494
rect 400422 520258 400464 520494
rect 400144 513494 400464 520258
rect 400144 513258 400186 513494
rect 400422 513258 400464 513494
rect 400144 506494 400464 513258
rect 400144 506258 400186 506494
rect 400422 506258 400464 506494
rect 400144 499494 400464 506258
rect 400144 499258 400186 499494
rect 400422 499258 400464 499494
rect 400144 492494 400464 499258
rect 400144 492258 400186 492494
rect 400422 492258 400464 492494
rect 400144 485494 400464 492258
rect 400144 485258 400186 485494
rect 400422 485258 400464 485494
rect 400144 478494 400464 485258
rect 400144 478258 400186 478494
rect 400422 478258 400464 478494
rect 400144 471494 400464 478258
rect 400144 471258 400186 471494
rect 400422 471258 400464 471494
rect 400144 464494 400464 471258
rect 400144 464258 400186 464494
rect 400422 464258 400464 464494
rect 400144 457494 400464 464258
rect 400144 457258 400186 457494
rect 400422 457258 400464 457494
rect 400144 450494 400464 457258
rect 400144 450258 400186 450494
rect 400422 450258 400464 450494
rect 400144 443494 400464 450258
rect 400144 443258 400186 443494
rect 400422 443258 400464 443494
rect 400144 436494 400464 443258
rect 400144 436258 400186 436494
rect 400422 436258 400464 436494
rect 400144 429494 400464 436258
rect 400144 429258 400186 429494
rect 400422 429258 400464 429494
rect 400144 422494 400464 429258
rect 400144 422258 400186 422494
rect 400422 422258 400464 422494
rect 400144 415494 400464 422258
rect 400144 415258 400186 415494
rect 400422 415258 400464 415494
rect 400144 408494 400464 415258
rect 400144 408258 400186 408494
rect 400422 408258 400464 408494
rect 400144 401494 400464 408258
rect 400144 401258 400186 401494
rect 400422 401258 400464 401494
rect 400144 394494 400464 401258
rect 400144 394258 400186 394494
rect 400422 394258 400464 394494
rect 400144 387494 400464 394258
rect 400144 387258 400186 387494
rect 400422 387258 400464 387494
rect 400144 380494 400464 387258
rect 400144 380258 400186 380494
rect 400422 380258 400464 380494
rect 400144 373494 400464 380258
rect 400144 373258 400186 373494
rect 400422 373258 400464 373494
rect 400144 366494 400464 373258
rect 400144 366258 400186 366494
rect 400422 366258 400464 366494
rect 400144 359494 400464 366258
rect 400144 359258 400186 359494
rect 400422 359258 400464 359494
rect 400144 352494 400464 359258
rect 400144 352258 400186 352494
rect 400422 352258 400464 352494
rect 400144 345494 400464 352258
rect 400144 345258 400186 345494
rect 400422 345258 400464 345494
rect 400144 338494 400464 345258
rect 400144 338258 400186 338494
rect 400422 338258 400464 338494
rect 400144 331494 400464 338258
rect 400144 331258 400186 331494
rect 400422 331258 400464 331494
rect 400144 324494 400464 331258
rect 400144 324258 400186 324494
rect 400422 324258 400464 324494
rect 400144 317494 400464 324258
rect 400144 317258 400186 317494
rect 400422 317258 400464 317494
rect 400144 310494 400464 317258
rect 400144 310258 400186 310494
rect 400422 310258 400464 310494
rect 400144 303494 400464 310258
rect 400144 303258 400186 303494
rect 400422 303258 400464 303494
rect 400144 296494 400464 303258
rect 400144 296258 400186 296494
rect 400422 296258 400464 296494
rect 400144 289494 400464 296258
rect 400144 289258 400186 289494
rect 400422 289258 400464 289494
rect 400144 282494 400464 289258
rect 400144 282258 400186 282494
rect 400422 282258 400464 282494
rect 400144 275494 400464 282258
rect 400144 275258 400186 275494
rect 400422 275258 400464 275494
rect 400144 268494 400464 275258
rect 400144 268258 400186 268494
rect 400422 268258 400464 268494
rect 400144 261494 400464 268258
rect 400144 261258 400186 261494
rect 400422 261258 400464 261494
rect 400144 254494 400464 261258
rect 400144 254258 400186 254494
rect 400422 254258 400464 254494
rect 400144 247494 400464 254258
rect 400144 247258 400186 247494
rect 400422 247258 400464 247494
rect 400144 240494 400464 247258
rect 400144 240258 400186 240494
rect 400422 240258 400464 240494
rect 400144 233494 400464 240258
rect 400144 233258 400186 233494
rect 400422 233258 400464 233494
rect 400144 226494 400464 233258
rect 400144 226258 400186 226494
rect 400422 226258 400464 226494
rect 400144 219494 400464 226258
rect 400144 219258 400186 219494
rect 400422 219258 400464 219494
rect 400144 212494 400464 219258
rect 400144 212258 400186 212494
rect 400422 212258 400464 212494
rect 400144 205494 400464 212258
rect 400144 205258 400186 205494
rect 400422 205258 400464 205494
rect 400144 198494 400464 205258
rect 400144 198258 400186 198494
rect 400422 198258 400464 198494
rect 400144 191494 400464 198258
rect 400144 191258 400186 191494
rect 400422 191258 400464 191494
rect 400144 184494 400464 191258
rect 400144 184258 400186 184494
rect 400422 184258 400464 184494
rect 400144 177494 400464 184258
rect 400144 177258 400186 177494
rect 400422 177258 400464 177494
rect 400144 170494 400464 177258
rect 400144 170258 400186 170494
rect 400422 170258 400464 170494
rect 400144 163494 400464 170258
rect 400144 163258 400186 163494
rect 400422 163258 400464 163494
rect 400144 156494 400464 163258
rect 400144 156258 400186 156494
rect 400422 156258 400464 156494
rect 400144 149494 400464 156258
rect 400144 149258 400186 149494
rect 400422 149258 400464 149494
rect 400144 142494 400464 149258
rect 400144 142258 400186 142494
rect 400422 142258 400464 142494
rect 400144 135494 400464 142258
rect 400144 135258 400186 135494
rect 400422 135258 400464 135494
rect 400144 128494 400464 135258
rect 400144 128258 400186 128494
rect 400422 128258 400464 128494
rect 400144 121494 400464 128258
rect 400144 121258 400186 121494
rect 400422 121258 400464 121494
rect 400144 114494 400464 121258
rect 400144 114258 400186 114494
rect 400422 114258 400464 114494
rect 400144 107494 400464 114258
rect 400144 107258 400186 107494
rect 400422 107258 400464 107494
rect 400144 100494 400464 107258
rect 400144 100258 400186 100494
rect 400422 100258 400464 100494
rect 400144 93494 400464 100258
rect 400144 93258 400186 93494
rect 400422 93258 400464 93494
rect 400144 86494 400464 93258
rect 400144 86258 400186 86494
rect 400422 86258 400464 86494
rect 400144 79494 400464 86258
rect 400144 79258 400186 79494
rect 400422 79258 400464 79494
rect 400144 72494 400464 79258
rect 400144 72258 400186 72494
rect 400422 72258 400464 72494
rect 400144 65494 400464 72258
rect 400144 65258 400186 65494
rect 400422 65258 400464 65494
rect 400144 58494 400464 65258
rect 400144 58258 400186 58494
rect 400422 58258 400464 58494
rect 400144 51494 400464 58258
rect 400144 51258 400186 51494
rect 400422 51258 400464 51494
rect 400144 44494 400464 51258
rect 400144 44258 400186 44494
rect 400422 44258 400464 44494
rect 400144 37494 400464 44258
rect 400144 37258 400186 37494
rect 400422 37258 400464 37494
rect 400144 30494 400464 37258
rect 400144 30258 400186 30494
rect 400422 30258 400464 30494
rect 400144 23494 400464 30258
rect 400144 23258 400186 23494
rect 400422 23258 400464 23494
rect 400144 16494 400464 23258
rect 400144 16258 400186 16494
rect 400422 16258 400464 16494
rect 400144 9494 400464 16258
rect 400144 9258 400186 9494
rect 400422 9258 400464 9494
rect 400144 2494 400464 9258
rect 400144 2258 400186 2494
rect 400422 2258 400464 2494
rect 400144 -746 400464 2258
rect 400144 -982 400186 -746
rect 400422 -982 400464 -746
rect 400144 -1066 400464 -982
rect 400144 -1302 400186 -1066
rect 400422 -1302 400464 -1066
rect 400144 -2294 400464 -1302
rect 401876 706198 402196 706230
rect 401876 705962 401918 706198
rect 402154 705962 402196 706198
rect 401876 705878 402196 705962
rect 401876 705642 401918 705878
rect 402154 705642 402196 705878
rect 401876 696434 402196 705642
rect 401876 696198 401918 696434
rect 402154 696198 402196 696434
rect 401876 689434 402196 696198
rect 401876 689198 401918 689434
rect 402154 689198 402196 689434
rect 401876 682434 402196 689198
rect 401876 682198 401918 682434
rect 402154 682198 402196 682434
rect 401876 675434 402196 682198
rect 401876 675198 401918 675434
rect 402154 675198 402196 675434
rect 401876 668434 402196 675198
rect 401876 668198 401918 668434
rect 402154 668198 402196 668434
rect 401876 661434 402196 668198
rect 401876 661198 401918 661434
rect 402154 661198 402196 661434
rect 401876 654434 402196 661198
rect 401876 654198 401918 654434
rect 402154 654198 402196 654434
rect 401876 647434 402196 654198
rect 401876 647198 401918 647434
rect 402154 647198 402196 647434
rect 401876 640434 402196 647198
rect 401876 640198 401918 640434
rect 402154 640198 402196 640434
rect 401876 633434 402196 640198
rect 401876 633198 401918 633434
rect 402154 633198 402196 633434
rect 401876 626434 402196 633198
rect 401876 626198 401918 626434
rect 402154 626198 402196 626434
rect 401876 619434 402196 626198
rect 401876 619198 401918 619434
rect 402154 619198 402196 619434
rect 401876 612434 402196 619198
rect 401876 612198 401918 612434
rect 402154 612198 402196 612434
rect 401876 605434 402196 612198
rect 401876 605198 401918 605434
rect 402154 605198 402196 605434
rect 401876 598434 402196 605198
rect 401876 598198 401918 598434
rect 402154 598198 402196 598434
rect 401876 591434 402196 598198
rect 401876 591198 401918 591434
rect 402154 591198 402196 591434
rect 401876 584434 402196 591198
rect 401876 584198 401918 584434
rect 402154 584198 402196 584434
rect 401876 577434 402196 584198
rect 401876 577198 401918 577434
rect 402154 577198 402196 577434
rect 401876 570434 402196 577198
rect 401876 570198 401918 570434
rect 402154 570198 402196 570434
rect 401876 563434 402196 570198
rect 401876 563198 401918 563434
rect 402154 563198 402196 563434
rect 401876 556434 402196 563198
rect 401876 556198 401918 556434
rect 402154 556198 402196 556434
rect 401876 549434 402196 556198
rect 401876 549198 401918 549434
rect 402154 549198 402196 549434
rect 401876 542434 402196 549198
rect 401876 542198 401918 542434
rect 402154 542198 402196 542434
rect 401876 535434 402196 542198
rect 401876 535198 401918 535434
rect 402154 535198 402196 535434
rect 401876 528434 402196 535198
rect 401876 528198 401918 528434
rect 402154 528198 402196 528434
rect 401876 521434 402196 528198
rect 401876 521198 401918 521434
rect 402154 521198 402196 521434
rect 401876 514434 402196 521198
rect 401876 514198 401918 514434
rect 402154 514198 402196 514434
rect 401876 507434 402196 514198
rect 401876 507198 401918 507434
rect 402154 507198 402196 507434
rect 401876 500434 402196 507198
rect 401876 500198 401918 500434
rect 402154 500198 402196 500434
rect 401876 493434 402196 500198
rect 401876 493198 401918 493434
rect 402154 493198 402196 493434
rect 401876 486434 402196 493198
rect 401876 486198 401918 486434
rect 402154 486198 402196 486434
rect 401876 479434 402196 486198
rect 401876 479198 401918 479434
rect 402154 479198 402196 479434
rect 401876 472434 402196 479198
rect 401876 472198 401918 472434
rect 402154 472198 402196 472434
rect 401876 465434 402196 472198
rect 401876 465198 401918 465434
rect 402154 465198 402196 465434
rect 401876 458434 402196 465198
rect 401876 458198 401918 458434
rect 402154 458198 402196 458434
rect 401876 451434 402196 458198
rect 401876 451198 401918 451434
rect 402154 451198 402196 451434
rect 401876 444434 402196 451198
rect 401876 444198 401918 444434
rect 402154 444198 402196 444434
rect 401876 437434 402196 444198
rect 401876 437198 401918 437434
rect 402154 437198 402196 437434
rect 401876 430434 402196 437198
rect 401876 430198 401918 430434
rect 402154 430198 402196 430434
rect 401876 423434 402196 430198
rect 401876 423198 401918 423434
rect 402154 423198 402196 423434
rect 401876 416434 402196 423198
rect 401876 416198 401918 416434
rect 402154 416198 402196 416434
rect 401876 409434 402196 416198
rect 401876 409198 401918 409434
rect 402154 409198 402196 409434
rect 401876 402434 402196 409198
rect 401876 402198 401918 402434
rect 402154 402198 402196 402434
rect 401876 395434 402196 402198
rect 401876 395198 401918 395434
rect 402154 395198 402196 395434
rect 401876 388434 402196 395198
rect 401876 388198 401918 388434
rect 402154 388198 402196 388434
rect 401876 381434 402196 388198
rect 401876 381198 401918 381434
rect 402154 381198 402196 381434
rect 401876 374434 402196 381198
rect 401876 374198 401918 374434
rect 402154 374198 402196 374434
rect 401876 367434 402196 374198
rect 401876 367198 401918 367434
rect 402154 367198 402196 367434
rect 401876 360434 402196 367198
rect 401876 360198 401918 360434
rect 402154 360198 402196 360434
rect 401876 353434 402196 360198
rect 401876 353198 401918 353434
rect 402154 353198 402196 353434
rect 401876 346434 402196 353198
rect 401876 346198 401918 346434
rect 402154 346198 402196 346434
rect 401876 339434 402196 346198
rect 401876 339198 401918 339434
rect 402154 339198 402196 339434
rect 401876 332434 402196 339198
rect 401876 332198 401918 332434
rect 402154 332198 402196 332434
rect 401876 325434 402196 332198
rect 401876 325198 401918 325434
rect 402154 325198 402196 325434
rect 401876 318434 402196 325198
rect 401876 318198 401918 318434
rect 402154 318198 402196 318434
rect 401876 311434 402196 318198
rect 401876 311198 401918 311434
rect 402154 311198 402196 311434
rect 401876 304434 402196 311198
rect 401876 304198 401918 304434
rect 402154 304198 402196 304434
rect 401876 297434 402196 304198
rect 401876 297198 401918 297434
rect 402154 297198 402196 297434
rect 401876 290434 402196 297198
rect 401876 290198 401918 290434
rect 402154 290198 402196 290434
rect 401876 283434 402196 290198
rect 401876 283198 401918 283434
rect 402154 283198 402196 283434
rect 401876 276434 402196 283198
rect 401876 276198 401918 276434
rect 402154 276198 402196 276434
rect 401876 269434 402196 276198
rect 401876 269198 401918 269434
rect 402154 269198 402196 269434
rect 401876 262434 402196 269198
rect 401876 262198 401918 262434
rect 402154 262198 402196 262434
rect 401876 255434 402196 262198
rect 401876 255198 401918 255434
rect 402154 255198 402196 255434
rect 401876 248434 402196 255198
rect 401876 248198 401918 248434
rect 402154 248198 402196 248434
rect 401876 241434 402196 248198
rect 401876 241198 401918 241434
rect 402154 241198 402196 241434
rect 401876 234434 402196 241198
rect 401876 234198 401918 234434
rect 402154 234198 402196 234434
rect 401876 227434 402196 234198
rect 401876 227198 401918 227434
rect 402154 227198 402196 227434
rect 401876 220434 402196 227198
rect 401876 220198 401918 220434
rect 402154 220198 402196 220434
rect 401876 213434 402196 220198
rect 401876 213198 401918 213434
rect 402154 213198 402196 213434
rect 401876 206434 402196 213198
rect 401876 206198 401918 206434
rect 402154 206198 402196 206434
rect 401876 199434 402196 206198
rect 401876 199198 401918 199434
rect 402154 199198 402196 199434
rect 401876 192434 402196 199198
rect 401876 192198 401918 192434
rect 402154 192198 402196 192434
rect 401876 185434 402196 192198
rect 401876 185198 401918 185434
rect 402154 185198 402196 185434
rect 401876 178434 402196 185198
rect 401876 178198 401918 178434
rect 402154 178198 402196 178434
rect 401876 171434 402196 178198
rect 401876 171198 401918 171434
rect 402154 171198 402196 171434
rect 401876 164434 402196 171198
rect 401876 164198 401918 164434
rect 402154 164198 402196 164434
rect 401876 157434 402196 164198
rect 401876 157198 401918 157434
rect 402154 157198 402196 157434
rect 401876 150434 402196 157198
rect 401876 150198 401918 150434
rect 402154 150198 402196 150434
rect 401876 143434 402196 150198
rect 401876 143198 401918 143434
rect 402154 143198 402196 143434
rect 401876 136434 402196 143198
rect 401876 136198 401918 136434
rect 402154 136198 402196 136434
rect 401876 129434 402196 136198
rect 401876 129198 401918 129434
rect 402154 129198 402196 129434
rect 401876 122434 402196 129198
rect 401876 122198 401918 122434
rect 402154 122198 402196 122434
rect 401876 115434 402196 122198
rect 401876 115198 401918 115434
rect 402154 115198 402196 115434
rect 401876 108434 402196 115198
rect 401876 108198 401918 108434
rect 402154 108198 402196 108434
rect 401876 101434 402196 108198
rect 401876 101198 401918 101434
rect 402154 101198 402196 101434
rect 401876 94434 402196 101198
rect 401876 94198 401918 94434
rect 402154 94198 402196 94434
rect 401876 87434 402196 94198
rect 401876 87198 401918 87434
rect 402154 87198 402196 87434
rect 401876 80434 402196 87198
rect 401876 80198 401918 80434
rect 402154 80198 402196 80434
rect 401876 73434 402196 80198
rect 401876 73198 401918 73434
rect 402154 73198 402196 73434
rect 401876 66434 402196 73198
rect 401876 66198 401918 66434
rect 402154 66198 402196 66434
rect 401876 59434 402196 66198
rect 401876 59198 401918 59434
rect 402154 59198 402196 59434
rect 401876 52434 402196 59198
rect 401876 52198 401918 52434
rect 402154 52198 402196 52434
rect 401876 45434 402196 52198
rect 401876 45198 401918 45434
rect 402154 45198 402196 45434
rect 401876 38434 402196 45198
rect 401876 38198 401918 38434
rect 402154 38198 402196 38434
rect 401876 31434 402196 38198
rect 401876 31198 401918 31434
rect 402154 31198 402196 31434
rect 401876 24434 402196 31198
rect 401876 24198 401918 24434
rect 402154 24198 402196 24434
rect 401876 17434 402196 24198
rect 401876 17198 401918 17434
rect 402154 17198 402196 17434
rect 401876 10434 402196 17198
rect 401876 10198 401918 10434
rect 402154 10198 402196 10434
rect 401876 3434 402196 10198
rect 401876 3198 401918 3434
rect 402154 3198 402196 3434
rect 401876 -1706 402196 3198
rect 401876 -1942 401918 -1706
rect 402154 -1942 402196 -1706
rect 401876 -2026 402196 -1942
rect 401876 -2262 401918 -2026
rect 402154 -2262 402196 -2026
rect 401876 -2294 402196 -2262
rect 407144 705238 407464 706230
rect 407144 705002 407186 705238
rect 407422 705002 407464 705238
rect 407144 704918 407464 705002
rect 407144 704682 407186 704918
rect 407422 704682 407464 704918
rect 407144 695494 407464 704682
rect 407144 695258 407186 695494
rect 407422 695258 407464 695494
rect 407144 688494 407464 695258
rect 407144 688258 407186 688494
rect 407422 688258 407464 688494
rect 407144 681494 407464 688258
rect 407144 681258 407186 681494
rect 407422 681258 407464 681494
rect 407144 674494 407464 681258
rect 407144 674258 407186 674494
rect 407422 674258 407464 674494
rect 407144 667494 407464 674258
rect 407144 667258 407186 667494
rect 407422 667258 407464 667494
rect 407144 660494 407464 667258
rect 407144 660258 407186 660494
rect 407422 660258 407464 660494
rect 407144 653494 407464 660258
rect 407144 653258 407186 653494
rect 407422 653258 407464 653494
rect 407144 646494 407464 653258
rect 407144 646258 407186 646494
rect 407422 646258 407464 646494
rect 407144 639494 407464 646258
rect 407144 639258 407186 639494
rect 407422 639258 407464 639494
rect 407144 632494 407464 639258
rect 407144 632258 407186 632494
rect 407422 632258 407464 632494
rect 407144 625494 407464 632258
rect 407144 625258 407186 625494
rect 407422 625258 407464 625494
rect 407144 618494 407464 625258
rect 407144 618258 407186 618494
rect 407422 618258 407464 618494
rect 407144 611494 407464 618258
rect 407144 611258 407186 611494
rect 407422 611258 407464 611494
rect 407144 604494 407464 611258
rect 407144 604258 407186 604494
rect 407422 604258 407464 604494
rect 407144 597494 407464 604258
rect 407144 597258 407186 597494
rect 407422 597258 407464 597494
rect 407144 590494 407464 597258
rect 407144 590258 407186 590494
rect 407422 590258 407464 590494
rect 407144 583494 407464 590258
rect 407144 583258 407186 583494
rect 407422 583258 407464 583494
rect 407144 576494 407464 583258
rect 407144 576258 407186 576494
rect 407422 576258 407464 576494
rect 407144 569494 407464 576258
rect 407144 569258 407186 569494
rect 407422 569258 407464 569494
rect 407144 562494 407464 569258
rect 407144 562258 407186 562494
rect 407422 562258 407464 562494
rect 407144 555494 407464 562258
rect 407144 555258 407186 555494
rect 407422 555258 407464 555494
rect 407144 548494 407464 555258
rect 407144 548258 407186 548494
rect 407422 548258 407464 548494
rect 407144 541494 407464 548258
rect 407144 541258 407186 541494
rect 407422 541258 407464 541494
rect 407144 534494 407464 541258
rect 407144 534258 407186 534494
rect 407422 534258 407464 534494
rect 407144 527494 407464 534258
rect 407144 527258 407186 527494
rect 407422 527258 407464 527494
rect 407144 520494 407464 527258
rect 407144 520258 407186 520494
rect 407422 520258 407464 520494
rect 407144 513494 407464 520258
rect 407144 513258 407186 513494
rect 407422 513258 407464 513494
rect 407144 506494 407464 513258
rect 407144 506258 407186 506494
rect 407422 506258 407464 506494
rect 407144 499494 407464 506258
rect 407144 499258 407186 499494
rect 407422 499258 407464 499494
rect 407144 492494 407464 499258
rect 407144 492258 407186 492494
rect 407422 492258 407464 492494
rect 407144 485494 407464 492258
rect 407144 485258 407186 485494
rect 407422 485258 407464 485494
rect 407144 478494 407464 485258
rect 407144 478258 407186 478494
rect 407422 478258 407464 478494
rect 407144 471494 407464 478258
rect 407144 471258 407186 471494
rect 407422 471258 407464 471494
rect 407144 464494 407464 471258
rect 407144 464258 407186 464494
rect 407422 464258 407464 464494
rect 407144 457494 407464 464258
rect 407144 457258 407186 457494
rect 407422 457258 407464 457494
rect 407144 450494 407464 457258
rect 407144 450258 407186 450494
rect 407422 450258 407464 450494
rect 407144 443494 407464 450258
rect 407144 443258 407186 443494
rect 407422 443258 407464 443494
rect 407144 436494 407464 443258
rect 407144 436258 407186 436494
rect 407422 436258 407464 436494
rect 407144 429494 407464 436258
rect 407144 429258 407186 429494
rect 407422 429258 407464 429494
rect 407144 422494 407464 429258
rect 407144 422258 407186 422494
rect 407422 422258 407464 422494
rect 407144 415494 407464 422258
rect 407144 415258 407186 415494
rect 407422 415258 407464 415494
rect 407144 408494 407464 415258
rect 407144 408258 407186 408494
rect 407422 408258 407464 408494
rect 407144 401494 407464 408258
rect 407144 401258 407186 401494
rect 407422 401258 407464 401494
rect 407144 394494 407464 401258
rect 407144 394258 407186 394494
rect 407422 394258 407464 394494
rect 407144 387494 407464 394258
rect 407144 387258 407186 387494
rect 407422 387258 407464 387494
rect 407144 380494 407464 387258
rect 407144 380258 407186 380494
rect 407422 380258 407464 380494
rect 407144 373494 407464 380258
rect 407144 373258 407186 373494
rect 407422 373258 407464 373494
rect 407144 366494 407464 373258
rect 407144 366258 407186 366494
rect 407422 366258 407464 366494
rect 407144 359494 407464 366258
rect 407144 359258 407186 359494
rect 407422 359258 407464 359494
rect 407144 352494 407464 359258
rect 407144 352258 407186 352494
rect 407422 352258 407464 352494
rect 407144 345494 407464 352258
rect 407144 345258 407186 345494
rect 407422 345258 407464 345494
rect 407144 338494 407464 345258
rect 407144 338258 407186 338494
rect 407422 338258 407464 338494
rect 407144 331494 407464 338258
rect 407144 331258 407186 331494
rect 407422 331258 407464 331494
rect 407144 324494 407464 331258
rect 407144 324258 407186 324494
rect 407422 324258 407464 324494
rect 407144 317494 407464 324258
rect 407144 317258 407186 317494
rect 407422 317258 407464 317494
rect 407144 310494 407464 317258
rect 407144 310258 407186 310494
rect 407422 310258 407464 310494
rect 407144 303494 407464 310258
rect 407144 303258 407186 303494
rect 407422 303258 407464 303494
rect 407144 296494 407464 303258
rect 407144 296258 407186 296494
rect 407422 296258 407464 296494
rect 407144 289494 407464 296258
rect 407144 289258 407186 289494
rect 407422 289258 407464 289494
rect 407144 282494 407464 289258
rect 407144 282258 407186 282494
rect 407422 282258 407464 282494
rect 407144 275494 407464 282258
rect 407144 275258 407186 275494
rect 407422 275258 407464 275494
rect 407144 268494 407464 275258
rect 407144 268258 407186 268494
rect 407422 268258 407464 268494
rect 407144 261494 407464 268258
rect 407144 261258 407186 261494
rect 407422 261258 407464 261494
rect 407144 254494 407464 261258
rect 407144 254258 407186 254494
rect 407422 254258 407464 254494
rect 407144 247494 407464 254258
rect 407144 247258 407186 247494
rect 407422 247258 407464 247494
rect 407144 240494 407464 247258
rect 407144 240258 407186 240494
rect 407422 240258 407464 240494
rect 407144 233494 407464 240258
rect 407144 233258 407186 233494
rect 407422 233258 407464 233494
rect 407144 226494 407464 233258
rect 407144 226258 407186 226494
rect 407422 226258 407464 226494
rect 407144 219494 407464 226258
rect 407144 219258 407186 219494
rect 407422 219258 407464 219494
rect 407144 212494 407464 219258
rect 407144 212258 407186 212494
rect 407422 212258 407464 212494
rect 407144 205494 407464 212258
rect 407144 205258 407186 205494
rect 407422 205258 407464 205494
rect 407144 198494 407464 205258
rect 407144 198258 407186 198494
rect 407422 198258 407464 198494
rect 407144 191494 407464 198258
rect 407144 191258 407186 191494
rect 407422 191258 407464 191494
rect 407144 184494 407464 191258
rect 407144 184258 407186 184494
rect 407422 184258 407464 184494
rect 407144 177494 407464 184258
rect 407144 177258 407186 177494
rect 407422 177258 407464 177494
rect 407144 170494 407464 177258
rect 407144 170258 407186 170494
rect 407422 170258 407464 170494
rect 407144 163494 407464 170258
rect 407144 163258 407186 163494
rect 407422 163258 407464 163494
rect 407144 156494 407464 163258
rect 407144 156258 407186 156494
rect 407422 156258 407464 156494
rect 407144 149494 407464 156258
rect 407144 149258 407186 149494
rect 407422 149258 407464 149494
rect 407144 142494 407464 149258
rect 407144 142258 407186 142494
rect 407422 142258 407464 142494
rect 407144 135494 407464 142258
rect 407144 135258 407186 135494
rect 407422 135258 407464 135494
rect 407144 128494 407464 135258
rect 407144 128258 407186 128494
rect 407422 128258 407464 128494
rect 407144 121494 407464 128258
rect 407144 121258 407186 121494
rect 407422 121258 407464 121494
rect 407144 114494 407464 121258
rect 407144 114258 407186 114494
rect 407422 114258 407464 114494
rect 407144 107494 407464 114258
rect 407144 107258 407186 107494
rect 407422 107258 407464 107494
rect 407144 100494 407464 107258
rect 407144 100258 407186 100494
rect 407422 100258 407464 100494
rect 407144 93494 407464 100258
rect 407144 93258 407186 93494
rect 407422 93258 407464 93494
rect 407144 86494 407464 93258
rect 407144 86258 407186 86494
rect 407422 86258 407464 86494
rect 407144 79494 407464 86258
rect 407144 79258 407186 79494
rect 407422 79258 407464 79494
rect 407144 72494 407464 79258
rect 407144 72258 407186 72494
rect 407422 72258 407464 72494
rect 407144 65494 407464 72258
rect 407144 65258 407186 65494
rect 407422 65258 407464 65494
rect 407144 58494 407464 65258
rect 407144 58258 407186 58494
rect 407422 58258 407464 58494
rect 407144 51494 407464 58258
rect 407144 51258 407186 51494
rect 407422 51258 407464 51494
rect 407144 44494 407464 51258
rect 407144 44258 407186 44494
rect 407422 44258 407464 44494
rect 407144 37494 407464 44258
rect 407144 37258 407186 37494
rect 407422 37258 407464 37494
rect 407144 30494 407464 37258
rect 407144 30258 407186 30494
rect 407422 30258 407464 30494
rect 407144 23494 407464 30258
rect 407144 23258 407186 23494
rect 407422 23258 407464 23494
rect 407144 16494 407464 23258
rect 407144 16258 407186 16494
rect 407422 16258 407464 16494
rect 407144 9494 407464 16258
rect 407144 9258 407186 9494
rect 407422 9258 407464 9494
rect 407144 2494 407464 9258
rect 407144 2258 407186 2494
rect 407422 2258 407464 2494
rect 407144 -746 407464 2258
rect 407144 -982 407186 -746
rect 407422 -982 407464 -746
rect 407144 -1066 407464 -982
rect 407144 -1302 407186 -1066
rect 407422 -1302 407464 -1066
rect 407144 -2294 407464 -1302
rect 408876 706198 409196 706230
rect 408876 705962 408918 706198
rect 409154 705962 409196 706198
rect 408876 705878 409196 705962
rect 408876 705642 408918 705878
rect 409154 705642 409196 705878
rect 408876 696434 409196 705642
rect 408876 696198 408918 696434
rect 409154 696198 409196 696434
rect 408876 689434 409196 696198
rect 408876 689198 408918 689434
rect 409154 689198 409196 689434
rect 408876 682434 409196 689198
rect 408876 682198 408918 682434
rect 409154 682198 409196 682434
rect 408876 675434 409196 682198
rect 408876 675198 408918 675434
rect 409154 675198 409196 675434
rect 408876 668434 409196 675198
rect 408876 668198 408918 668434
rect 409154 668198 409196 668434
rect 408876 661434 409196 668198
rect 408876 661198 408918 661434
rect 409154 661198 409196 661434
rect 408876 654434 409196 661198
rect 408876 654198 408918 654434
rect 409154 654198 409196 654434
rect 408876 647434 409196 654198
rect 408876 647198 408918 647434
rect 409154 647198 409196 647434
rect 408876 640434 409196 647198
rect 408876 640198 408918 640434
rect 409154 640198 409196 640434
rect 408876 633434 409196 640198
rect 408876 633198 408918 633434
rect 409154 633198 409196 633434
rect 408876 626434 409196 633198
rect 408876 626198 408918 626434
rect 409154 626198 409196 626434
rect 408876 619434 409196 626198
rect 408876 619198 408918 619434
rect 409154 619198 409196 619434
rect 408876 612434 409196 619198
rect 408876 612198 408918 612434
rect 409154 612198 409196 612434
rect 408876 605434 409196 612198
rect 408876 605198 408918 605434
rect 409154 605198 409196 605434
rect 408876 598434 409196 605198
rect 408876 598198 408918 598434
rect 409154 598198 409196 598434
rect 408876 591434 409196 598198
rect 408876 591198 408918 591434
rect 409154 591198 409196 591434
rect 408876 584434 409196 591198
rect 408876 584198 408918 584434
rect 409154 584198 409196 584434
rect 408876 577434 409196 584198
rect 408876 577198 408918 577434
rect 409154 577198 409196 577434
rect 408876 570434 409196 577198
rect 408876 570198 408918 570434
rect 409154 570198 409196 570434
rect 408876 563434 409196 570198
rect 408876 563198 408918 563434
rect 409154 563198 409196 563434
rect 408876 556434 409196 563198
rect 408876 556198 408918 556434
rect 409154 556198 409196 556434
rect 408876 549434 409196 556198
rect 408876 549198 408918 549434
rect 409154 549198 409196 549434
rect 408876 542434 409196 549198
rect 408876 542198 408918 542434
rect 409154 542198 409196 542434
rect 408876 535434 409196 542198
rect 408876 535198 408918 535434
rect 409154 535198 409196 535434
rect 408876 528434 409196 535198
rect 408876 528198 408918 528434
rect 409154 528198 409196 528434
rect 408876 521434 409196 528198
rect 408876 521198 408918 521434
rect 409154 521198 409196 521434
rect 408876 514434 409196 521198
rect 408876 514198 408918 514434
rect 409154 514198 409196 514434
rect 408876 507434 409196 514198
rect 408876 507198 408918 507434
rect 409154 507198 409196 507434
rect 408876 500434 409196 507198
rect 408876 500198 408918 500434
rect 409154 500198 409196 500434
rect 408876 493434 409196 500198
rect 408876 493198 408918 493434
rect 409154 493198 409196 493434
rect 408876 486434 409196 493198
rect 408876 486198 408918 486434
rect 409154 486198 409196 486434
rect 408876 479434 409196 486198
rect 408876 479198 408918 479434
rect 409154 479198 409196 479434
rect 408876 472434 409196 479198
rect 408876 472198 408918 472434
rect 409154 472198 409196 472434
rect 408876 465434 409196 472198
rect 408876 465198 408918 465434
rect 409154 465198 409196 465434
rect 408876 458434 409196 465198
rect 408876 458198 408918 458434
rect 409154 458198 409196 458434
rect 408876 451434 409196 458198
rect 408876 451198 408918 451434
rect 409154 451198 409196 451434
rect 408876 444434 409196 451198
rect 408876 444198 408918 444434
rect 409154 444198 409196 444434
rect 408876 437434 409196 444198
rect 408876 437198 408918 437434
rect 409154 437198 409196 437434
rect 408876 430434 409196 437198
rect 408876 430198 408918 430434
rect 409154 430198 409196 430434
rect 408876 423434 409196 430198
rect 408876 423198 408918 423434
rect 409154 423198 409196 423434
rect 408876 416434 409196 423198
rect 408876 416198 408918 416434
rect 409154 416198 409196 416434
rect 408876 409434 409196 416198
rect 408876 409198 408918 409434
rect 409154 409198 409196 409434
rect 408876 402434 409196 409198
rect 408876 402198 408918 402434
rect 409154 402198 409196 402434
rect 408876 395434 409196 402198
rect 408876 395198 408918 395434
rect 409154 395198 409196 395434
rect 408876 388434 409196 395198
rect 408876 388198 408918 388434
rect 409154 388198 409196 388434
rect 408876 381434 409196 388198
rect 408876 381198 408918 381434
rect 409154 381198 409196 381434
rect 408876 374434 409196 381198
rect 408876 374198 408918 374434
rect 409154 374198 409196 374434
rect 408876 367434 409196 374198
rect 408876 367198 408918 367434
rect 409154 367198 409196 367434
rect 408876 360434 409196 367198
rect 408876 360198 408918 360434
rect 409154 360198 409196 360434
rect 408876 353434 409196 360198
rect 408876 353198 408918 353434
rect 409154 353198 409196 353434
rect 408876 346434 409196 353198
rect 408876 346198 408918 346434
rect 409154 346198 409196 346434
rect 408876 339434 409196 346198
rect 408876 339198 408918 339434
rect 409154 339198 409196 339434
rect 408876 332434 409196 339198
rect 408876 332198 408918 332434
rect 409154 332198 409196 332434
rect 408876 325434 409196 332198
rect 408876 325198 408918 325434
rect 409154 325198 409196 325434
rect 408876 318434 409196 325198
rect 408876 318198 408918 318434
rect 409154 318198 409196 318434
rect 408876 311434 409196 318198
rect 408876 311198 408918 311434
rect 409154 311198 409196 311434
rect 408876 304434 409196 311198
rect 408876 304198 408918 304434
rect 409154 304198 409196 304434
rect 408876 297434 409196 304198
rect 408876 297198 408918 297434
rect 409154 297198 409196 297434
rect 408876 290434 409196 297198
rect 408876 290198 408918 290434
rect 409154 290198 409196 290434
rect 408876 283434 409196 290198
rect 408876 283198 408918 283434
rect 409154 283198 409196 283434
rect 408876 276434 409196 283198
rect 408876 276198 408918 276434
rect 409154 276198 409196 276434
rect 408876 269434 409196 276198
rect 408876 269198 408918 269434
rect 409154 269198 409196 269434
rect 408876 262434 409196 269198
rect 408876 262198 408918 262434
rect 409154 262198 409196 262434
rect 408876 255434 409196 262198
rect 408876 255198 408918 255434
rect 409154 255198 409196 255434
rect 408876 248434 409196 255198
rect 408876 248198 408918 248434
rect 409154 248198 409196 248434
rect 408876 241434 409196 248198
rect 408876 241198 408918 241434
rect 409154 241198 409196 241434
rect 408876 234434 409196 241198
rect 408876 234198 408918 234434
rect 409154 234198 409196 234434
rect 408876 227434 409196 234198
rect 408876 227198 408918 227434
rect 409154 227198 409196 227434
rect 408876 220434 409196 227198
rect 408876 220198 408918 220434
rect 409154 220198 409196 220434
rect 408876 213434 409196 220198
rect 408876 213198 408918 213434
rect 409154 213198 409196 213434
rect 408876 206434 409196 213198
rect 408876 206198 408918 206434
rect 409154 206198 409196 206434
rect 408876 199434 409196 206198
rect 408876 199198 408918 199434
rect 409154 199198 409196 199434
rect 408876 192434 409196 199198
rect 408876 192198 408918 192434
rect 409154 192198 409196 192434
rect 408876 185434 409196 192198
rect 408876 185198 408918 185434
rect 409154 185198 409196 185434
rect 408876 178434 409196 185198
rect 408876 178198 408918 178434
rect 409154 178198 409196 178434
rect 408876 171434 409196 178198
rect 408876 171198 408918 171434
rect 409154 171198 409196 171434
rect 408876 164434 409196 171198
rect 408876 164198 408918 164434
rect 409154 164198 409196 164434
rect 408876 157434 409196 164198
rect 408876 157198 408918 157434
rect 409154 157198 409196 157434
rect 408876 150434 409196 157198
rect 408876 150198 408918 150434
rect 409154 150198 409196 150434
rect 408876 143434 409196 150198
rect 408876 143198 408918 143434
rect 409154 143198 409196 143434
rect 408876 136434 409196 143198
rect 408876 136198 408918 136434
rect 409154 136198 409196 136434
rect 408876 129434 409196 136198
rect 408876 129198 408918 129434
rect 409154 129198 409196 129434
rect 408876 122434 409196 129198
rect 408876 122198 408918 122434
rect 409154 122198 409196 122434
rect 408876 115434 409196 122198
rect 408876 115198 408918 115434
rect 409154 115198 409196 115434
rect 408876 108434 409196 115198
rect 408876 108198 408918 108434
rect 409154 108198 409196 108434
rect 408876 101434 409196 108198
rect 408876 101198 408918 101434
rect 409154 101198 409196 101434
rect 408876 94434 409196 101198
rect 408876 94198 408918 94434
rect 409154 94198 409196 94434
rect 408876 87434 409196 94198
rect 408876 87198 408918 87434
rect 409154 87198 409196 87434
rect 408876 80434 409196 87198
rect 408876 80198 408918 80434
rect 409154 80198 409196 80434
rect 408876 73434 409196 80198
rect 408876 73198 408918 73434
rect 409154 73198 409196 73434
rect 408876 66434 409196 73198
rect 408876 66198 408918 66434
rect 409154 66198 409196 66434
rect 408876 59434 409196 66198
rect 408876 59198 408918 59434
rect 409154 59198 409196 59434
rect 408876 52434 409196 59198
rect 408876 52198 408918 52434
rect 409154 52198 409196 52434
rect 408876 45434 409196 52198
rect 408876 45198 408918 45434
rect 409154 45198 409196 45434
rect 408876 38434 409196 45198
rect 408876 38198 408918 38434
rect 409154 38198 409196 38434
rect 408876 31434 409196 38198
rect 408876 31198 408918 31434
rect 409154 31198 409196 31434
rect 408876 24434 409196 31198
rect 408876 24198 408918 24434
rect 409154 24198 409196 24434
rect 408876 17434 409196 24198
rect 408876 17198 408918 17434
rect 409154 17198 409196 17434
rect 408876 10434 409196 17198
rect 408876 10198 408918 10434
rect 409154 10198 409196 10434
rect 408876 3434 409196 10198
rect 408876 3198 408918 3434
rect 409154 3198 409196 3434
rect 408876 -1706 409196 3198
rect 408876 -1942 408918 -1706
rect 409154 -1942 409196 -1706
rect 408876 -2026 409196 -1942
rect 408876 -2262 408918 -2026
rect 409154 -2262 409196 -2026
rect 408876 -2294 409196 -2262
rect 414144 705238 414464 706230
rect 414144 705002 414186 705238
rect 414422 705002 414464 705238
rect 414144 704918 414464 705002
rect 414144 704682 414186 704918
rect 414422 704682 414464 704918
rect 414144 695494 414464 704682
rect 414144 695258 414186 695494
rect 414422 695258 414464 695494
rect 414144 688494 414464 695258
rect 414144 688258 414186 688494
rect 414422 688258 414464 688494
rect 414144 681494 414464 688258
rect 414144 681258 414186 681494
rect 414422 681258 414464 681494
rect 414144 674494 414464 681258
rect 414144 674258 414186 674494
rect 414422 674258 414464 674494
rect 414144 667494 414464 674258
rect 414144 667258 414186 667494
rect 414422 667258 414464 667494
rect 414144 660494 414464 667258
rect 414144 660258 414186 660494
rect 414422 660258 414464 660494
rect 414144 653494 414464 660258
rect 414144 653258 414186 653494
rect 414422 653258 414464 653494
rect 414144 646494 414464 653258
rect 414144 646258 414186 646494
rect 414422 646258 414464 646494
rect 414144 639494 414464 646258
rect 414144 639258 414186 639494
rect 414422 639258 414464 639494
rect 414144 632494 414464 639258
rect 414144 632258 414186 632494
rect 414422 632258 414464 632494
rect 414144 625494 414464 632258
rect 414144 625258 414186 625494
rect 414422 625258 414464 625494
rect 414144 618494 414464 625258
rect 414144 618258 414186 618494
rect 414422 618258 414464 618494
rect 414144 611494 414464 618258
rect 414144 611258 414186 611494
rect 414422 611258 414464 611494
rect 414144 604494 414464 611258
rect 414144 604258 414186 604494
rect 414422 604258 414464 604494
rect 414144 597494 414464 604258
rect 414144 597258 414186 597494
rect 414422 597258 414464 597494
rect 414144 590494 414464 597258
rect 414144 590258 414186 590494
rect 414422 590258 414464 590494
rect 414144 583494 414464 590258
rect 414144 583258 414186 583494
rect 414422 583258 414464 583494
rect 414144 576494 414464 583258
rect 414144 576258 414186 576494
rect 414422 576258 414464 576494
rect 414144 569494 414464 576258
rect 414144 569258 414186 569494
rect 414422 569258 414464 569494
rect 414144 562494 414464 569258
rect 414144 562258 414186 562494
rect 414422 562258 414464 562494
rect 414144 555494 414464 562258
rect 414144 555258 414186 555494
rect 414422 555258 414464 555494
rect 414144 548494 414464 555258
rect 414144 548258 414186 548494
rect 414422 548258 414464 548494
rect 414144 541494 414464 548258
rect 414144 541258 414186 541494
rect 414422 541258 414464 541494
rect 414144 534494 414464 541258
rect 414144 534258 414186 534494
rect 414422 534258 414464 534494
rect 414144 527494 414464 534258
rect 414144 527258 414186 527494
rect 414422 527258 414464 527494
rect 414144 520494 414464 527258
rect 414144 520258 414186 520494
rect 414422 520258 414464 520494
rect 414144 513494 414464 520258
rect 414144 513258 414186 513494
rect 414422 513258 414464 513494
rect 414144 506494 414464 513258
rect 414144 506258 414186 506494
rect 414422 506258 414464 506494
rect 414144 499494 414464 506258
rect 414144 499258 414186 499494
rect 414422 499258 414464 499494
rect 414144 492494 414464 499258
rect 414144 492258 414186 492494
rect 414422 492258 414464 492494
rect 414144 485494 414464 492258
rect 414144 485258 414186 485494
rect 414422 485258 414464 485494
rect 414144 478494 414464 485258
rect 414144 478258 414186 478494
rect 414422 478258 414464 478494
rect 414144 471494 414464 478258
rect 414144 471258 414186 471494
rect 414422 471258 414464 471494
rect 414144 464494 414464 471258
rect 414144 464258 414186 464494
rect 414422 464258 414464 464494
rect 414144 457494 414464 464258
rect 414144 457258 414186 457494
rect 414422 457258 414464 457494
rect 414144 450494 414464 457258
rect 414144 450258 414186 450494
rect 414422 450258 414464 450494
rect 414144 443494 414464 450258
rect 414144 443258 414186 443494
rect 414422 443258 414464 443494
rect 414144 436494 414464 443258
rect 414144 436258 414186 436494
rect 414422 436258 414464 436494
rect 414144 429494 414464 436258
rect 414144 429258 414186 429494
rect 414422 429258 414464 429494
rect 414144 422494 414464 429258
rect 414144 422258 414186 422494
rect 414422 422258 414464 422494
rect 414144 415494 414464 422258
rect 414144 415258 414186 415494
rect 414422 415258 414464 415494
rect 414144 408494 414464 415258
rect 414144 408258 414186 408494
rect 414422 408258 414464 408494
rect 414144 401494 414464 408258
rect 414144 401258 414186 401494
rect 414422 401258 414464 401494
rect 414144 394494 414464 401258
rect 414144 394258 414186 394494
rect 414422 394258 414464 394494
rect 414144 387494 414464 394258
rect 414144 387258 414186 387494
rect 414422 387258 414464 387494
rect 414144 380494 414464 387258
rect 414144 380258 414186 380494
rect 414422 380258 414464 380494
rect 414144 373494 414464 380258
rect 414144 373258 414186 373494
rect 414422 373258 414464 373494
rect 414144 366494 414464 373258
rect 414144 366258 414186 366494
rect 414422 366258 414464 366494
rect 414144 359494 414464 366258
rect 414144 359258 414186 359494
rect 414422 359258 414464 359494
rect 414144 352494 414464 359258
rect 414144 352258 414186 352494
rect 414422 352258 414464 352494
rect 414144 345494 414464 352258
rect 414144 345258 414186 345494
rect 414422 345258 414464 345494
rect 414144 338494 414464 345258
rect 414144 338258 414186 338494
rect 414422 338258 414464 338494
rect 414144 331494 414464 338258
rect 414144 331258 414186 331494
rect 414422 331258 414464 331494
rect 414144 324494 414464 331258
rect 414144 324258 414186 324494
rect 414422 324258 414464 324494
rect 414144 317494 414464 324258
rect 414144 317258 414186 317494
rect 414422 317258 414464 317494
rect 414144 310494 414464 317258
rect 414144 310258 414186 310494
rect 414422 310258 414464 310494
rect 414144 303494 414464 310258
rect 414144 303258 414186 303494
rect 414422 303258 414464 303494
rect 414144 296494 414464 303258
rect 414144 296258 414186 296494
rect 414422 296258 414464 296494
rect 414144 289494 414464 296258
rect 414144 289258 414186 289494
rect 414422 289258 414464 289494
rect 414144 282494 414464 289258
rect 414144 282258 414186 282494
rect 414422 282258 414464 282494
rect 414144 275494 414464 282258
rect 414144 275258 414186 275494
rect 414422 275258 414464 275494
rect 414144 268494 414464 275258
rect 414144 268258 414186 268494
rect 414422 268258 414464 268494
rect 414144 261494 414464 268258
rect 414144 261258 414186 261494
rect 414422 261258 414464 261494
rect 414144 254494 414464 261258
rect 414144 254258 414186 254494
rect 414422 254258 414464 254494
rect 414144 247494 414464 254258
rect 414144 247258 414186 247494
rect 414422 247258 414464 247494
rect 414144 240494 414464 247258
rect 414144 240258 414186 240494
rect 414422 240258 414464 240494
rect 414144 233494 414464 240258
rect 414144 233258 414186 233494
rect 414422 233258 414464 233494
rect 414144 226494 414464 233258
rect 414144 226258 414186 226494
rect 414422 226258 414464 226494
rect 414144 219494 414464 226258
rect 414144 219258 414186 219494
rect 414422 219258 414464 219494
rect 414144 212494 414464 219258
rect 414144 212258 414186 212494
rect 414422 212258 414464 212494
rect 414144 205494 414464 212258
rect 414144 205258 414186 205494
rect 414422 205258 414464 205494
rect 414144 198494 414464 205258
rect 414144 198258 414186 198494
rect 414422 198258 414464 198494
rect 414144 191494 414464 198258
rect 414144 191258 414186 191494
rect 414422 191258 414464 191494
rect 414144 184494 414464 191258
rect 414144 184258 414186 184494
rect 414422 184258 414464 184494
rect 414144 177494 414464 184258
rect 414144 177258 414186 177494
rect 414422 177258 414464 177494
rect 414144 170494 414464 177258
rect 414144 170258 414186 170494
rect 414422 170258 414464 170494
rect 414144 163494 414464 170258
rect 414144 163258 414186 163494
rect 414422 163258 414464 163494
rect 414144 156494 414464 163258
rect 414144 156258 414186 156494
rect 414422 156258 414464 156494
rect 414144 149494 414464 156258
rect 414144 149258 414186 149494
rect 414422 149258 414464 149494
rect 414144 142494 414464 149258
rect 414144 142258 414186 142494
rect 414422 142258 414464 142494
rect 414144 135494 414464 142258
rect 414144 135258 414186 135494
rect 414422 135258 414464 135494
rect 414144 128494 414464 135258
rect 414144 128258 414186 128494
rect 414422 128258 414464 128494
rect 414144 121494 414464 128258
rect 414144 121258 414186 121494
rect 414422 121258 414464 121494
rect 414144 114494 414464 121258
rect 414144 114258 414186 114494
rect 414422 114258 414464 114494
rect 414144 107494 414464 114258
rect 414144 107258 414186 107494
rect 414422 107258 414464 107494
rect 414144 100494 414464 107258
rect 414144 100258 414186 100494
rect 414422 100258 414464 100494
rect 414144 93494 414464 100258
rect 414144 93258 414186 93494
rect 414422 93258 414464 93494
rect 414144 86494 414464 93258
rect 414144 86258 414186 86494
rect 414422 86258 414464 86494
rect 414144 79494 414464 86258
rect 414144 79258 414186 79494
rect 414422 79258 414464 79494
rect 414144 72494 414464 79258
rect 414144 72258 414186 72494
rect 414422 72258 414464 72494
rect 414144 65494 414464 72258
rect 414144 65258 414186 65494
rect 414422 65258 414464 65494
rect 414144 58494 414464 65258
rect 414144 58258 414186 58494
rect 414422 58258 414464 58494
rect 414144 51494 414464 58258
rect 414144 51258 414186 51494
rect 414422 51258 414464 51494
rect 414144 44494 414464 51258
rect 414144 44258 414186 44494
rect 414422 44258 414464 44494
rect 414144 37494 414464 44258
rect 414144 37258 414186 37494
rect 414422 37258 414464 37494
rect 414144 30494 414464 37258
rect 414144 30258 414186 30494
rect 414422 30258 414464 30494
rect 414144 23494 414464 30258
rect 414144 23258 414186 23494
rect 414422 23258 414464 23494
rect 414144 16494 414464 23258
rect 414144 16258 414186 16494
rect 414422 16258 414464 16494
rect 414144 9494 414464 16258
rect 414144 9258 414186 9494
rect 414422 9258 414464 9494
rect 414144 2494 414464 9258
rect 414144 2258 414186 2494
rect 414422 2258 414464 2494
rect 414144 -746 414464 2258
rect 414144 -982 414186 -746
rect 414422 -982 414464 -746
rect 414144 -1066 414464 -982
rect 414144 -1302 414186 -1066
rect 414422 -1302 414464 -1066
rect 414144 -2294 414464 -1302
rect 415876 706198 416196 706230
rect 415876 705962 415918 706198
rect 416154 705962 416196 706198
rect 415876 705878 416196 705962
rect 415876 705642 415918 705878
rect 416154 705642 416196 705878
rect 415876 696434 416196 705642
rect 415876 696198 415918 696434
rect 416154 696198 416196 696434
rect 415876 689434 416196 696198
rect 415876 689198 415918 689434
rect 416154 689198 416196 689434
rect 415876 682434 416196 689198
rect 415876 682198 415918 682434
rect 416154 682198 416196 682434
rect 415876 675434 416196 682198
rect 415876 675198 415918 675434
rect 416154 675198 416196 675434
rect 415876 668434 416196 675198
rect 415876 668198 415918 668434
rect 416154 668198 416196 668434
rect 415876 661434 416196 668198
rect 415876 661198 415918 661434
rect 416154 661198 416196 661434
rect 415876 654434 416196 661198
rect 415876 654198 415918 654434
rect 416154 654198 416196 654434
rect 415876 647434 416196 654198
rect 415876 647198 415918 647434
rect 416154 647198 416196 647434
rect 415876 640434 416196 647198
rect 415876 640198 415918 640434
rect 416154 640198 416196 640434
rect 415876 633434 416196 640198
rect 415876 633198 415918 633434
rect 416154 633198 416196 633434
rect 415876 626434 416196 633198
rect 415876 626198 415918 626434
rect 416154 626198 416196 626434
rect 415876 619434 416196 626198
rect 415876 619198 415918 619434
rect 416154 619198 416196 619434
rect 415876 612434 416196 619198
rect 415876 612198 415918 612434
rect 416154 612198 416196 612434
rect 415876 605434 416196 612198
rect 415876 605198 415918 605434
rect 416154 605198 416196 605434
rect 415876 598434 416196 605198
rect 415876 598198 415918 598434
rect 416154 598198 416196 598434
rect 415876 591434 416196 598198
rect 415876 591198 415918 591434
rect 416154 591198 416196 591434
rect 415876 584434 416196 591198
rect 415876 584198 415918 584434
rect 416154 584198 416196 584434
rect 415876 577434 416196 584198
rect 415876 577198 415918 577434
rect 416154 577198 416196 577434
rect 415876 570434 416196 577198
rect 415876 570198 415918 570434
rect 416154 570198 416196 570434
rect 415876 563434 416196 570198
rect 415876 563198 415918 563434
rect 416154 563198 416196 563434
rect 415876 556434 416196 563198
rect 415876 556198 415918 556434
rect 416154 556198 416196 556434
rect 415876 549434 416196 556198
rect 415876 549198 415918 549434
rect 416154 549198 416196 549434
rect 415876 542434 416196 549198
rect 415876 542198 415918 542434
rect 416154 542198 416196 542434
rect 415876 535434 416196 542198
rect 415876 535198 415918 535434
rect 416154 535198 416196 535434
rect 415876 528434 416196 535198
rect 415876 528198 415918 528434
rect 416154 528198 416196 528434
rect 415876 521434 416196 528198
rect 415876 521198 415918 521434
rect 416154 521198 416196 521434
rect 415876 514434 416196 521198
rect 415876 514198 415918 514434
rect 416154 514198 416196 514434
rect 415876 507434 416196 514198
rect 415876 507198 415918 507434
rect 416154 507198 416196 507434
rect 415876 500434 416196 507198
rect 415876 500198 415918 500434
rect 416154 500198 416196 500434
rect 415876 493434 416196 500198
rect 415876 493198 415918 493434
rect 416154 493198 416196 493434
rect 415876 486434 416196 493198
rect 415876 486198 415918 486434
rect 416154 486198 416196 486434
rect 415876 479434 416196 486198
rect 415876 479198 415918 479434
rect 416154 479198 416196 479434
rect 415876 472434 416196 479198
rect 415876 472198 415918 472434
rect 416154 472198 416196 472434
rect 415876 465434 416196 472198
rect 415876 465198 415918 465434
rect 416154 465198 416196 465434
rect 415876 458434 416196 465198
rect 415876 458198 415918 458434
rect 416154 458198 416196 458434
rect 415876 451434 416196 458198
rect 415876 451198 415918 451434
rect 416154 451198 416196 451434
rect 415876 444434 416196 451198
rect 415876 444198 415918 444434
rect 416154 444198 416196 444434
rect 415876 437434 416196 444198
rect 415876 437198 415918 437434
rect 416154 437198 416196 437434
rect 415876 430434 416196 437198
rect 415876 430198 415918 430434
rect 416154 430198 416196 430434
rect 415876 423434 416196 430198
rect 415876 423198 415918 423434
rect 416154 423198 416196 423434
rect 415876 416434 416196 423198
rect 415876 416198 415918 416434
rect 416154 416198 416196 416434
rect 415876 409434 416196 416198
rect 415876 409198 415918 409434
rect 416154 409198 416196 409434
rect 415876 402434 416196 409198
rect 415876 402198 415918 402434
rect 416154 402198 416196 402434
rect 415876 395434 416196 402198
rect 415876 395198 415918 395434
rect 416154 395198 416196 395434
rect 415876 388434 416196 395198
rect 415876 388198 415918 388434
rect 416154 388198 416196 388434
rect 415876 381434 416196 388198
rect 415876 381198 415918 381434
rect 416154 381198 416196 381434
rect 415876 374434 416196 381198
rect 415876 374198 415918 374434
rect 416154 374198 416196 374434
rect 415876 367434 416196 374198
rect 415876 367198 415918 367434
rect 416154 367198 416196 367434
rect 415876 360434 416196 367198
rect 415876 360198 415918 360434
rect 416154 360198 416196 360434
rect 415876 353434 416196 360198
rect 415876 353198 415918 353434
rect 416154 353198 416196 353434
rect 415876 346434 416196 353198
rect 415876 346198 415918 346434
rect 416154 346198 416196 346434
rect 415876 339434 416196 346198
rect 415876 339198 415918 339434
rect 416154 339198 416196 339434
rect 415876 332434 416196 339198
rect 415876 332198 415918 332434
rect 416154 332198 416196 332434
rect 415876 325434 416196 332198
rect 415876 325198 415918 325434
rect 416154 325198 416196 325434
rect 415876 318434 416196 325198
rect 415876 318198 415918 318434
rect 416154 318198 416196 318434
rect 415876 311434 416196 318198
rect 415876 311198 415918 311434
rect 416154 311198 416196 311434
rect 415876 304434 416196 311198
rect 415876 304198 415918 304434
rect 416154 304198 416196 304434
rect 415876 297434 416196 304198
rect 415876 297198 415918 297434
rect 416154 297198 416196 297434
rect 415876 290434 416196 297198
rect 415876 290198 415918 290434
rect 416154 290198 416196 290434
rect 415876 283434 416196 290198
rect 415876 283198 415918 283434
rect 416154 283198 416196 283434
rect 415876 276434 416196 283198
rect 415876 276198 415918 276434
rect 416154 276198 416196 276434
rect 415876 269434 416196 276198
rect 415876 269198 415918 269434
rect 416154 269198 416196 269434
rect 415876 262434 416196 269198
rect 415876 262198 415918 262434
rect 416154 262198 416196 262434
rect 415876 255434 416196 262198
rect 415876 255198 415918 255434
rect 416154 255198 416196 255434
rect 415876 248434 416196 255198
rect 415876 248198 415918 248434
rect 416154 248198 416196 248434
rect 415876 241434 416196 248198
rect 415876 241198 415918 241434
rect 416154 241198 416196 241434
rect 415876 234434 416196 241198
rect 415876 234198 415918 234434
rect 416154 234198 416196 234434
rect 415876 227434 416196 234198
rect 415876 227198 415918 227434
rect 416154 227198 416196 227434
rect 415876 220434 416196 227198
rect 415876 220198 415918 220434
rect 416154 220198 416196 220434
rect 415876 213434 416196 220198
rect 415876 213198 415918 213434
rect 416154 213198 416196 213434
rect 415876 206434 416196 213198
rect 415876 206198 415918 206434
rect 416154 206198 416196 206434
rect 415876 199434 416196 206198
rect 415876 199198 415918 199434
rect 416154 199198 416196 199434
rect 415876 192434 416196 199198
rect 415876 192198 415918 192434
rect 416154 192198 416196 192434
rect 415876 185434 416196 192198
rect 415876 185198 415918 185434
rect 416154 185198 416196 185434
rect 415876 178434 416196 185198
rect 415876 178198 415918 178434
rect 416154 178198 416196 178434
rect 415876 171434 416196 178198
rect 415876 171198 415918 171434
rect 416154 171198 416196 171434
rect 415876 164434 416196 171198
rect 415876 164198 415918 164434
rect 416154 164198 416196 164434
rect 415876 157434 416196 164198
rect 415876 157198 415918 157434
rect 416154 157198 416196 157434
rect 415876 150434 416196 157198
rect 415876 150198 415918 150434
rect 416154 150198 416196 150434
rect 415876 143434 416196 150198
rect 415876 143198 415918 143434
rect 416154 143198 416196 143434
rect 415876 136434 416196 143198
rect 415876 136198 415918 136434
rect 416154 136198 416196 136434
rect 415876 129434 416196 136198
rect 415876 129198 415918 129434
rect 416154 129198 416196 129434
rect 415876 122434 416196 129198
rect 415876 122198 415918 122434
rect 416154 122198 416196 122434
rect 415876 115434 416196 122198
rect 415876 115198 415918 115434
rect 416154 115198 416196 115434
rect 415876 108434 416196 115198
rect 415876 108198 415918 108434
rect 416154 108198 416196 108434
rect 415876 101434 416196 108198
rect 415876 101198 415918 101434
rect 416154 101198 416196 101434
rect 415876 94434 416196 101198
rect 415876 94198 415918 94434
rect 416154 94198 416196 94434
rect 415876 87434 416196 94198
rect 415876 87198 415918 87434
rect 416154 87198 416196 87434
rect 415876 80434 416196 87198
rect 415876 80198 415918 80434
rect 416154 80198 416196 80434
rect 415876 73434 416196 80198
rect 415876 73198 415918 73434
rect 416154 73198 416196 73434
rect 415876 66434 416196 73198
rect 415876 66198 415918 66434
rect 416154 66198 416196 66434
rect 415876 59434 416196 66198
rect 415876 59198 415918 59434
rect 416154 59198 416196 59434
rect 415876 52434 416196 59198
rect 415876 52198 415918 52434
rect 416154 52198 416196 52434
rect 415876 45434 416196 52198
rect 415876 45198 415918 45434
rect 416154 45198 416196 45434
rect 415876 38434 416196 45198
rect 415876 38198 415918 38434
rect 416154 38198 416196 38434
rect 415876 31434 416196 38198
rect 415876 31198 415918 31434
rect 416154 31198 416196 31434
rect 415876 24434 416196 31198
rect 415876 24198 415918 24434
rect 416154 24198 416196 24434
rect 415876 17434 416196 24198
rect 415876 17198 415918 17434
rect 416154 17198 416196 17434
rect 415876 10434 416196 17198
rect 415876 10198 415918 10434
rect 416154 10198 416196 10434
rect 415876 3434 416196 10198
rect 415876 3198 415918 3434
rect 416154 3198 416196 3434
rect 415876 -1706 416196 3198
rect 415876 -1942 415918 -1706
rect 416154 -1942 416196 -1706
rect 415876 -2026 416196 -1942
rect 415876 -2262 415918 -2026
rect 416154 -2262 416196 -2026
rect 415876 -2294 416196 -2262
rect 421144 705238 421464 706230
rect 421144 705002 421186 705238
rect 421422 705002 421464 705238
rect 421144 704918 421464 705002
rect 421144 704682 421186 704918
rect 421422 704682 421464 704918
rect 421144 695494 421464 704682
rect 421144 695258 421186 695494
rect 421422 695258 421464 695494
rect 421144 688494 421464 695258
rect 421144 688258 421186 688494
rect 421422 688258 421464 688494
rect 421144 681494 421464 688258
rect 421144 681258 421186 681494
rect 421422 681258 421464 681494
rect 421144 674494 421464 681258
rect 421144 674258 421186 674494
rect 421422 674258 421464 674494
rect 421144 667494 421464 674258
rect 421144 667258 421186 667494
rect 421422 667258 421464 667494
rect 421144 660494 421464 667258
rect 421144 660258 421186 660494
rect 421422 660258 421464 660494
rect 421144 653494 421464 660258
rect 421144 653258 421186 653494
rect 421422 653258 421464 653494
rect 421144 646494 421464 653258
rect 421144 646258 421186 646494
rect 421422 646258 421464 646494
rect 421144 639494 421464 646258
rect 421144 639258 421186 639494
rect 421422 639258 421464 639494
rect 421144 632494 421464 639258
rect 421144 632258 421186 632494
rect 421422 632258 421464 632494
rect 421144 625494 421464 632258
rect 421144 625258 421186 625494
rect 421422 625258 421464 625494
rect 421144 618494 421464 625258
rect 421144 618258 421186 618494
rect 421422 618258 421464 618494
rect 421144 611494 421464 618258
rect 421144 611258 421186 611494
rect 421422 611258 421464 611494
rect 421144 604494 421464 611258
rect 421144 604258 421186 604494
rect 421422 604258 421464 604494
rect 421144 597494 421464 604258
rect 421144 597258 421186 597494
rect 421422 597258 421464 597494
rect 421144 590494 421464 597258
rect 421144 590258 421186 590494
rect 421422 590258 421464 590494
rect 421144 583494 421464 590258
rect 421144 583258 421186 583494
rect 421422 583258 421464 583494
rect 421144 576494 421464 583258
rect 421144 576258 421186 576494
rect 421422 576258 421464 576494
rect 421144 569494 421464 576258
rect 421144 569258 421186 569494
rect 421422 569258 421464 569494
rect 421144 562494 421464 569258
rect 421144 562258 421186 562494
rect 421422 562258 421464 562494
rect 421144 555494 421464 562258
rect 421144 555258 421186 555494
rect 421422 555258 421464 555494
rect 421144 548494 421464 555258
rect 421144 548258 421186 548494
rect 421422 548258 421464 548494
rect 421144 541494 421464 548258
rect 421144 541258 421186 541494
rect 421422 541258 421464 541494
rect 421144 534494 421464 541258
rect 421144 534258 421186 534494
rect 421422 534258 421464 534494
rect 421144 527494 421464 534258
rect 421144 527258 421186 527494
rect 421422 527258 421464 527494
rect 421144 520494 421464 527258
rect 421144 520258 421186 520494
rect 421422 520258 421464 520494
rect 421144 513494 421464 520258
rect 421144 513258 421186 513494
rect 421422 513258 421464 513494
rect 421144 506494 421464 513258
rect 421144 506258 421186 506494
rect 421422 506258 421464 506494
rect 421144 499494 421464 506258
rect 421144 499258 421186 499494
rect 421422 499258 421464 499494
rect 421144 492494 421464 499258
rect 421144 492258 421186 492494
rect 421422 492258 421464 492494
rect 421144 485494 421464 492258
rect 421144 485258 421186 485494
rect 421422 485258 421464 485494
rect 421144 478494 421464 485258
rect 421144 478258 421186 478494
rect 421422 478258 421464 478494
rect 421144 471494 421464 478258
rect 421144 471258 421186 471494
rect 421422 471258 421464 471494
rect 421144 464494 421464 471258
rect 421144 464258 421186 464494
rect 421422 464258 421464 464494
rect 421144 457494 421464 464258
rect 421144 457258 421186 457494
rect 421422 457258 421464 457494
rect 421144 450494 421464 457258
rect 421144 450258 421186 450494
rect 421422 450258 421464 450494
rect 421144 443494 421464 450258
rect 421144 443258 421186 443494
rect 421422 443258 421464 443494
rect 421144 436494 421464 443258
rect 421144 436258 421186 436494
rect 421422 436258 421464 436494
rect 421144 429494 421464 436258
rect 421144 429258 421186 429494
rect 421422 429258 421464 429494
rect 421144 422494 421464 429258
rect 421144 422258 421186 422494
rect 421422 422258 421464 422494
rect 421144 415494 421464 422258
rect 421144 415258 421186 415494
rect 421422 415258 421464 415494
rect 421144 408494 421464 415258
rect 421144 408258 421186 408494
rect 421422 408258 421464 408494
rect 421144 401494 421464 408258
rect 421144 401258 421186 401494
rect 421422 401258 421464 401494
rect 421144 394494 421464 401258
rect 421144 394258 421186 394494
rect 421422 394258 421464 394494
rect 421144 387494 421464 394258
rect 421144 387258 421186 387494
rect 421422 387258 421464 387494
rect 421144 380494 421464 387258
rect 421144 380258 421186 380494
rect 421422 380258 421464 380494
rect 421144 373494 421464 380258
rect 421144 373258 421186 373494
rect 421422 373258 421464 373494
rect 421144 366494 421464 373258
rect 421144 366258 421186 366494
rect 421422 366258 421464 366494
rect 421144 359494 421464 366258
rect 421144 359258 421186 359494
rect 421422 359258 421464 359494
rect 421144 352494 421464 359258
rect 421144 352258 421186 352494
rect 421422 352258 421464 352494
rect 421144 345494 421464 352258
rect 421144 345258 421186 345494
rect 421422 345258 421464 345494
rect 421144 338494 421464 345258
rect 421144 338258 421186 338494
rect 421422 338258 421464 338494
rect 421144 331494 421464 338258
rect 421144 331258 421186 331494
rect 421422 331258 421464 331494
rect 421144 324494 421464 331258
rect 421144 324258 421186 324494
rect 421422 324258 421464 324494
rect 421144 317494 421464 324258
rect 421144 317258 421186 317494
rect 421422 317258 421464 317494
rect 421144 310494 421464 317258
rect 421144 310258 421186 310494
rect 421422 310258 421464 310494
rect 421144 303494 421464 310258
rect 421144 303258 421186 303494
rect 421422 303258 421464 303494
rect 421144 296494 421464 303258
rect 421144 296258 421186 296494
rect 421422 296258 421464 296494
rect 421144 289494 421464 296258
rect 421144 289258 421186 289494
rect 421422 289258 421464 289494
rect 421144 282494 421464 289258
rect 421144 282258 421186 282494
rect 421422 282258 421464 282494
rect 421144 275494 421464 282258
rect 421144 275258 421186 275494
rect 421422 275258 421464 275494
rect 421144 268494 421464 275258
rect 421144 268258 421186 268494
rect 421422 268258 421464 268494
rect 421144 261494 421464 268258
rect 421144 261258 421186 261494
rect 421422 261258 421464 261494
rect 421144 254494 421464 261258
rect 421144 254258 421186 254494
rect 421422 254258 421464 254494
rect 421144 247494 421464 254258
rect 421144 247258 421186 247494
rect 421422 247258 421464 247494
rect 421144 240494 421464 247258
rect 421144 240258 421186 240494
rect 421422 240258 421464 240494
rect 421144 233494 421464 240258
rect 421144 233258 421186 233494
rect 421422 233258 421464 233494
rect 421144 226494 421464 233258
rect 421144 226258 421186 226494
rect 421422 226258 421464 226494
rect 421144 219494 421464 226258
rect 421144 219258 421186 219494
rect 421422 219258 421464 219494
rect 421144 212494 421464 219258
rect 421144 212258 421186 212494
rect 421422 212258 421464 212494
rect 421144 205494 421464 212258
rect 421144 205258 421186 205494
rect 421422 205258 421464 205494
rect 421144 198494 421464 205258
rect 421144 198258 421186 198494
rect 421422 198258 421464 198494
rect 421144 191494 421464 198258
rect 421144 191258 421186 191494
rect 421422 191258 421464 191494
rect 421144 184494 421464 191258
rect 421144 184258 421186 184494
rect 421422 184258 421464 184494
rect 421144 177494 421464 184258
rect 421144 177258 421186 177494
rect 421422 177258 421464 177494
rect 421144 170494 421464 177258
rect 421144 170258 421186 170494
rect 421422 170258 421464 170494
rect 421144 163494 421464 170258
rect 421144 163258 421186 163494
rect 421422 163258 421464 163494
rect 421144 156494 421464 163258
rect 421144 156258 421186 156494
rect 421422 156258 421464 156494
rect 421144 149494 421464 156258
rect 421144 149258 421186 149494
rect 421422 149258 421464 149494
rect 421144 142494 421464 149258
rect 421144 142258 421186 142494
rect 421422 142258 421464 142494
rect 421144 135494 421464 142258
rect 421144 135258 421186 135494
rect 421422 135258 421464 135494
rect 421144 128494 421464 135258
rect 421144 128258 421186 128494
rect 421422 128258 421464 128494
rect 421144 121494 421464 128258
rect 421144 121258 421186 121494
rect 421422 121258 421464 121494
rect 421144 114494 421464 121258
rect 421144 114258 421186 114494
rect 421422 114258 421464 114494
rect 421144 107494 421464 114258
rect 421144 107258 421186 107494
rect 421422 107258 421464 107494
rect 421144 100494 421464 107258
rect 421144 100258 421186 100494
rect 421422 100258 421464 100494
rect 421144 93494 421464 100258
rect 421144 93258 421186 93494
rect 421422 93258 421464 93494
rect 421144 86494 421464 93258
rect 421144 86258 421186 86494
rect 421422 86258 421464 86494
rect 421144 79494 421464 86258
rect 421144 79258 421186 79494
rect 421422 79258 421464 79494
rect 421144 72494 421464 79258
rect 421144 72258 421186 72494
rect 421422 72258 421464 72494
rect 421144 65494 421464 72258
rect 421144 65258 421186 65494
rect 421422 65258 421464 65494
rect 421144 58494 421464 65258
rect 421144 58258 421186 58494
rect 421422 58258 421464 58494
rect 421144 51494 421464 58258
rect 421144 51258 421186 51494
rect 421422 51258 421464 51494
rect 421144 44494 421464 51258
rect 421144 44258 421186 44494
rect 421422 44258 421464 44494
rect 421144 37494 421464 44258
rect 421144 37258 421186 37494
rect 421422 37258 421464 37494
rect 421144 30494 421464 37258
rect 421144 30258 421186 30494
rect 421422 30258 421464 30494
rect 421144 23494 421464 30258
rect 421144 23258 421186 23494
rect 421422 23258 421464 23494
rect 421144 16494 421464 23258
rect 421144 16258 421186 16494
rect 421422 16258 421464 16494
rect 421144 9494 421464 16258
rect 421144 9258 421186 9494
rect 421422 9258 421464 9494
rect 421144 2494 421464 9258
rect 421144 2258 421186 2494
rect 421422 2258 421464 2494
rect 421144 -746 421464 2258
rect 421144 -982 421186 -746
rect 421422 -982 421464 -746
rect 421144 -1066 421464 -982
rect 421144 -1302 421186 -1066
rect 421422 -1302 421464 -1066
rect 421144 -2294 421464 -1302
rect 422876 706198 423196 706230
rect 422876 705962 422918 706198
rect 423154 705962 423196 706198
rect 422876 705878 423196 705962
rect 422876 705642 422918 705878
rect 423154 705642 423196 705878
rect 422876 696434 423196 705642
rect 422876 696198 422918 696434
rect 423154 696198 423196 696434
rect 422876 689434 423196 696198
rect 422876 689198 422918 689434
rect 423154 689198 423196 689434
rect 422876 682434 423196 689198
rect 422876 682198 422918 682434
rect 423154 682198 423196 682434
rect 422876 675434 423196 682198
rect 422876 675198 422918 675434
rect 423154 675198 423196 675434
rect 422876 668434 423196 675198
rect 422876 668198 422918 668434
rect 423154 668198 423196 668434
rect 422876 661434 423196 668198
rect 422876 661198 422918 661434
rect 423154 661198 423196 661434
rect 422876 654434 423196 661198
rect 422876 654198 422918 654434
rect 423154 654198 423196 654434
rect 422876 647434 423196 654198
rect 422876 647198 422918 647434
rect 423154 647198 423196 647434
rect 422876 640434 423196 647198
rect 422876 640198 422918 640434
rect 423154 640198 423196 640434
rect 422876 633434 423196 640198
rect 422876 633198 422918 633434
rect 423154 633198 423196 633434
rect 422876 626434 423196 633198
rect 422876 626198 422918 626434
rect 423154 626198 423196 626434
rect 422876 619434 423196 626198
rect 422876 619198 422918 619434
rect 423154 619198 423196 619434
rect 422876 612434 423196 619198
rect 422876 612198 422918 612434
rect 423154 612198 423196 612434
rect 422876 605434 423196 612198
rect 422876 605198 422918 605434
rect 423154 605198 423196 605434
rect 422876 598434 423196 605198
rect 422876 598198 422918 598434
rect 423154 598198 423196 598434
rect 422876 591434 423196 598198
rect 422876 591198 422918 591434
rect 423154 591198 423196 591434
rect 422876 584434 423196 591198
rect 422876 584198 422918 584434
rect 423154 584198 423196 584434
rect 422876 577434 423196 584198
rect 422876 577198 422918 577434
rect 423154 577198 423196 577434
rect 422876 570434 423196 577198
rect 422876 570198 422918 570434
rect 423154 570198 423196 570434
rect 422876 563434 423196 570198
rect 422876 563198 422918 563434
rect 423154 563198 423196 563434
rect 422876 556434 423196 563198
rect 422876 556198 422918 556434
rect 423154 556198 423196 556434
rect 422876 549434 423196 556198
rect 422876 549198 422918 549434
rect 423154 549198 423196 549434
rect 422876 542434 423196 549198
rect 422876 542198 422918 542434
rect 423154 542198 423196 542434
rect 422876 535434 423196 542198
rect 422876 535198 422918 535434
rect 423154 535198 423196 535434
rect 422876 528434 423196 535198
rect 422876 528198 422918 528434
rect 423154 528198 423196 528434
rect 422876 521434 423196 528198
rect 422876 521198 422918 521434
rect 423154 521198 423196 521434
rect 422876 514434 423196 521198
rect 422876 514198 422918 514434
rect 423154 514198 423196 514434
rect 422876 507434 423196 514198
rect 422876 507198 422918 507434
rect 423154 507198 423196 507434
rect 422876 500434 423196 507198
rect 422876 500198 422918 500434
rect 423154 500198 423196 500434
rect 422876 493434 423196 500198
rect 422876 493198 422918 493434
rect 423154 493198 423196 493434
rect 422876 486434 423196 493198
rect 422876 486198 422918 486434
rect 423154 486198 423196 486434
rect 422876 479434 423196 486198
rect 422876 479198 422918 479434
rect 423154 479198 423196 479434
rect 422876 472434 423196 479198
rect 422876 472198 422918 472434
rect 423154 472198 423196 472434
rect 422876 465434 423196 472198
rect 422876 465198 422918 465434
rect 423154 465198 423196 465434
rect 422876 458434 423196 465198
rect 422876 458198 422918 458434
rect 423154 458198 423196 458434
rect 422876 451434 423196 458198
rect 422876 451198 422918 451434
rect 423154 451198 423196 451434
rect 422876 444434 423196 451198
rect 422876 444198 422918 444434
rect 423154 444198 423196 444434
rect 422876 437434 423196 444198
rect 422876 437198 422918 437434
rect 423154 437198 423196 437434
rect 422876 430434 423196 437198
rect 422876 430198 422918 430434
rect 423154 430198 423196 430434
rect 422876 423434 423196 430198
rect 422876 423198 422918 423434
rect 423154 423198 423196 423434
rect 422876 416434 423196 423198
rect 422876 416198 422918 416434
rect 423154 416198 423196 416434
rect 422876 409434 423196 416198
rect 422876 409198 422918 409434
rect 423154 409198 423196 409434
rect 422876 402434 423196 409198
rect 422876 402198 422918 402434
rect 423154 402198 423196 402434
rect 422876 395434 423196 402198
rect 422876 395198 422918 395434
rect 423154 395198 423196 395434
rect 422876 388434 423196 395198
rect 422876 388198 422918 388434
rect 423154 388198 423196 388434
rect 422876 381434 423196 388198
rect 422876 381198 422918 381434
rect 423154 381198 423196 381434
rect 422876 374434 423196 381198
rect 422876 374198 422918 374434
rect 423154 374198 423196 374434
rect 422876 367434 423196 374198
rect 422876 367198 422918 367434
rect 423154 367198 423196 367434
rect 422876 360434 423196 367198
rect 422876 360198 422918 360434
rect 423154 360198 423196 360434
rect 422876 353434 423196 360198
rect 422876 353198 422918 353434
rect 423154 353198 423196 353434
rect 422876 346434 423196 353198
rect 422876 346198 422918 346434
rect 423154 346198 423196 346434
rect 422876 339434 423196 346198
rect 422876 339198 422918 339434
rect 423154 339198 423196 339434
rect 422876 332434 423196 339198
rect 422876 332198 422918 332434
rect 423154 332198 423196 332434
rect 422876 325434 423196 332198
rect 422876 325198 422918 325434
rect 423154 325198 423196 325434
rect 422876 318434 423196 325198
rect 422876 318198 422918 318434
rect 423154 318198 423196 318434
rect 422876 311434 423196 318198
rect 422876 311198 422918 311434
rect 423154 311198 423196 311434
rect 422876 304434 423196 311198
rect 422876 304198 422918 304434
rect 423154 304198 423196 304434
rect 422876 297434 423196 304198
rect 422876 297198 422918 297434
rect 423154 297198 423196 297434
rect 422876 290434 423196 297198
rect 422876 290198 422918 290434
rect 423154 290198 423196 290434
rect 422876 283434 423196 290198
rect 422876 283198 422918 283434
rect 423154 283198 423196 283434
rect 422876 276434 423196 283198
rect 422876 276198 422918 276434
rect 423154 276198 423196 276434
rect 422876 269434 423196 276198
rect 422876 269198 422918 269434
rect 423154 269198 423196 269434
rect 422876 262434 423196 269198
rect 422876 262198 422918 262434
rect 423154 262198 423196 262434
rect 422876 255434 423196 262198
rect 422876 255198 422918 255434
rect 423154 255198 423196 255434
rect 422876 248434 423196 255198
rect 422876 248198 422918 248434
rect 423154 248198 423196 248434
rect 422876 241434 423196 248198
rect 422876 241198 422918 241434
rect 423154 241198 423196 241434
rect 422876 234434 423196 241198
rect 422876 234198 422918 234434
rect 423154 234198 423196 234434
rect 422876 227434 423196 234198
rect 422876 227198 422918 227434
rect 423154 227198 423196 227434
rect 422876 220434 423196 227198
rect 422876 220198 422918 220434
rect 423154 220198 423196 220434
rect 422876 213434 423196 220198
rect 422876 213198 422918 213434
rect 423154 213198 423196 213434
rect 422876 206434 423196 213198
rect 422876 206198 422918 206434
rect 423154 206198 423196 206434
rect 422876 199434 423196 206198
rect 422876 199198 422918 199434
rect 423154 199198 423196 199434
rect 422876 192434 423196 199198
rect 422876 192198 422918 192434
rect 423154 192198 423196 192434
rect 422876 185434 423196 192198
rect 422876 185198 422918 185434
rect 423154 185198 423196 185434
rect 422876 178434 423196 185198
rect 422876 178198 422918 178434
rect 423154 178198 423196 178434
rect 422876 171434 423196 178198
rect 422876 171198 422918 171434
rect 423154 171198 423196 171434
rect 422876 164434 423196 171198
rect 422876 164198 422918 164434
rect 423154 164198 423196 164434
rect 422876 157434 423196 164198
rect 422876 157198 422918 157434
rect 423154 157198 423196 157434
rect 422876 150434 423196 157198
rect 422876 150198 422918 150434
rect 423154 150198 423196 150434
rect 422876 143434 423196 150198
rect 422876 143198 422918 143434
rect 423154 143198 423196 143434
rect 422876 136434 423196 143198
rect 422876 136198 422918 136434
rect 423154 136198 423196 136434
rect 422876 129434 423196 136198
rect 422876 129198 422918 129434
rect 423154 129198 423196 129434
rect 422876 122434 423196 129198
rect 422876 122198 422918 122434
rect 423154 122198 423196 122434
rect 422876 115434 423196 122198
rect 422876 115198 422918 115434
rect 423154 115198 423196 115434
rect 422876 108434 423196 115198
rect 422876 108198 422918 108434
rect 423154 108198 423196 108434
rect 422876 101434 423196 108198
rect 422876 101198 422918 101434
rect 423154 101198 423196 101434
rect 422876 94434 423196 101198
rect 422876 94198 422918 94434
rect 423154 94198 423196 94434
rect 422876 87434 423196 94198
rect 422876 87198 422918 87434
rect 423154 87198 423196 87434
rect 422876 80434 423196 87198
rect 422876 80198 422918 80434
rect 423154 80198 423196 80434
rect 422876 73434 423196 80198
rect 422876 73198 422918 73434
rect 423154 73198 423196 73434
rect 422876 66434 423196 73198
rect 422876 66198 422918 66434
rect 423154 66198 423196 66434
rect 422876 59434 423196 66198
rect 422876 59198 422918 59434
rect 423154 59198 423196 59434
rect 422876 52434 423196 59198
rect 422876 52198 422918 52434
rect 423154 52198 423196 52434
rect 422876 45434 423196 52198
rect 422876 45198 422918 45434
rect 423154 45198 423196 45434
rect 422876 38434 423196 45198
rect 422876 38198 422918 38434
rect 423154 38198 423196 38434
rect 422876 31434 423196 38198
rect 422876 31198 422918 31434
rect 423154 31198 423196 31434
rect 422876 24434 423196 31198
rect 422876 24198 422918 24434
rect 423154 24198 423196 24434
rect 422876 17434 423196 24198
rect 422876 17198 422918 17434
rect 423154 17198 423196 17434
rect 422876 10434 423196 17198
rect 422876 10198 422918 10434
rect 423154 10198 423196 10434
rect 422876 3434 423196 10198
rect 422876 3198 422918 3434
rect 423154 3198 423196 3434
rect 422876 -1706 423196 3198
rect 422876 -1942 422918 -1706
rect 423154 -1942 423196 -1706
rect 422876 -2026 423196 -1942
rect 422876 -2262 422918 -2026
rect 423154 -2262 423196 -2026
rect 422876 -2294 423196 -2262
rect 428144 705238 428464 706230
rect 428144 705002 428186 705238
rect 428422 705002 428464 705238
rect 428144 704918 428464 705002
rect 428144 704682 428186 704918
rect 428422 704682 428464 704918
rect 428144 695494 428464 704682
rect 428144 695258 428186 695494
rect 428422 695258 428464 695494
rect 428144 688494 428464 695258
rect 428144 688258 428186 688494
rect 428422 688258 428464 688494
rect 428144 681494 428464 688258
rect 428144 681258 428186 681494
rect 428422 681258 428464 681494
rect 428144 674494 428464 681258
rect 428144 674258 428186 674494
rect 428422 674258 428464 674494
rect 428144 667494 428464 674258
rect 428144 667258 428186 667494
rect 428422 667258 428464 667494
rect 428144 660494 428464 667258
rect 428144 660258 428186 660494
rect 428422 660258 428464 660494
rect 428144 653494 428464 660258
rect 428144 653258 428186 653494
rect 428422 653258 428464 653494
rect 428144 646494 428464 653258
rect 428144 646258 428186 646494
rect 428422 646258 428464 646494
rect 428144 639494 428464 646258
rect 428144 639258 428186 639494
rect 428422 639258 428464 639494
rect 428144 632494 428464 639258
rect 428144 632258 428186 632494
rect 428422 632258 428464 632494
rect 428144 625494 428464 632258
rect 428144 625258 428186 625494
rect 428422 625258 428464 625494
rect 428144 618494 428464 625258
rect 428144 618258 428186 618494
rect 428422 618258 428464 618494
rect 428144 611494 428464 618258
rect 428144 611258 428186 611494
rect 428422 611258 428464 611494
rect 428144 604494 428464 611258
rect 428144 604258 428186 604494
rect 428422 604258 428464 604494
rect 428144 597494 428464 604258
rect 428144 597258 428186 597494
rect 428422 597258 428464 597494
rect 428144 590494 428464 597258
rect 428144 590258 428186 590494
rect 428422 590258 428464 590494
rect 428144 583494 428464 590258
rect 428144 583258 428186 583494
rect 428422 583258 428464 583494
rect 428144 576494 428464 583258
rect 428144 576258 428186 576494
rect 428422 576258 428464 576494
rect 428144 569494 428464 576258
rect 428144 569258 428186 569494
rect 428422 569258 428464 569494
rect 428144 562494 428464 569258
rect 428144 562258 428186 562494
rect 428422 562258 428464 562494
rect 428144 555494 428464 562258
rect 428144 555258 428186 555494
rect 428422 555258 428464 555494
rect 428144 548494 428464 555258
rect 428144 548258 428186 548494
rect 428422 548258 428464 548494
rect 428144 541494 428464 548258
rect 428144 541258 428186 541494
rect 428422 541258 428464 541494
rect 428144 534494 428464 541258
rect 428144 534258 428186 534494
rect 428422 534258 428464 534494
rect 428144 527494 428464 534258
rect 428144 527258 428186 527494
rect 428422 527258 428464 527494
rect 428144 520494 428464 527258
rect 428144 520258 428186 520494
rect 428422 520258 428464 520494
rect 428144 513494 428464 520258
rect 428144 513258 428186 513494
rect 428422 513258 428464 513494
rect 428144 506494 428464 513258
rect 428144 506258 428186 506494
rect 428422 506258 428464 506494
rect 428144 499494 428464 506258
rect 428144 499258 428186 499494
rect 428422 499258 428464 499494
rect 428144 492494 428464 499258
rect 428144 492258 428186 492494
rect 428422 492258 428464 492494
rect 428144 485494 428464 492258
rect 428144 485258 428186 485494
rect 428422 485258 428464 485494
rect 428144 478494 428464 485258
rect 428144 478258 428186 478494
rect 428422 478258 428464 478494
rect 428144 471494 428464 478258
rect 428144 471258 428186 471494
rect 428422 471258 428464 471494
rect 428144 464494 428464 471258
rect 428144 464258 428186 464494
rect 428422 464258 428464 464494
rect 428144 457494 428464 464258
rect 428144 457258 428186 457494
rect 428422 457258 428464 457494
rect 428144 450494 428464 457258
rect 428144 450258 428186 450494
rect 428422 450258 428464 450494
rect 428144 443494 428464 450258
rect 428144 443258 428186 443494
rect 428422 443258 428464 443494
rect 428144 436494 428464 443258
rect 428144 436258 428186 436494
rect 428422 436258 428464 436494
rect 428144 429494 428464 436258
rect 428144 429258 428186 429494
rect 428422 429258 428464 429494
rect 428144 422494 428464 429258
rect 428144 422258 428186 422494
rect 428422 422258 428464 422494
rect 428144 415494 428464 422258
rect 428144 415258 428186 415494
rect 428422 415258 428464 415494
rect 428144 408494 428464 415258
rect 428144 408258 428186 408494
rect 428422 408258 428464 408494
rect 428144 401494 428464 408258
rect 428144 401258 428186 401494
rect 428422 401258 428464 401494
rect 428144 394494 428464 401258
rect 428144 394258 428186 394494
rect 428422 394258 428464 394494
rect 428144 387494 428464 394258
rect 428144 387258 428186 387494
rect 428422 387258 428464 387494
rect 428144 380494 428464 387258
rect 428144 380258 428186 380494
rect 428422 380258 428464 380494
rect 428144 373494 428464 380258
rect 428144 373258 428186 373494
rect 428422 373258 428464 373494
rect 428144 366494 428464 373258
rect 428144 366258 428186 366494
rect 428422 366258 428464 366494
rect 428144 359494 428464 366258
rect 428144 359258 428186 359494
rect 428422 359258 428464 359494
rect 428144 352494 428464 359258
rect 428144 352258 428186 352494
rect 428422 352258 428464 352494
rect 428144 345494 428464 352258
rect 428144 345258 428186 345494
rect 428422 345258 428464 345494
rect 428144 338494 428464 345258
rect 428144 338258 428186 338494
rect 428422 338258 428464 338494
rect 428144 331494 428464 338258
rect 428144 331258 428186 331494
rect 428422 331258 428464 331494
rect 428144 324494 428464 331258
rect 428144 324258 428186 324494
rect 428422 324258 428464 324494
rect 428144 317494 428464 324258
rect 428144 317258 428186 317494
rect 428422 317258 428464 317494
rect 428144 310494 428464 317258
rect 428144 310258 428186 310494
rect 428422 310258 428464 310494
rect 428144 303494 428464 310258
rect 428144 303258 428186 303494
rect 428422 303258 428464 303494
rect 428144 296494 428464 303258
rect 428144 296258 428186 296494
rect 428422 296258 428464 296494
rect 428144 289494 428464 296258
rect 428144 289258 428186 289494
rect 428422 289258 428464 289494
rect 428144 282494 428464 289258
rect 428144 282258 428186 282494
rect 428422 282258 428464 282494
rect 428144 275494 428464 282258
rect 428144 275258 428186 275494
rect 428422 275258 428464 275494
rect 428144 268494 428464 275258
rect 428144 268258 428186 268494
rect 428422 268258 428464 268494
rect 428144 261494 428464 268258
rect 428144 261258 428186 261494
rect 428422 261258 428464 261494
rect 428144 254494 428464 261258
rect 428144 254258 428186 254494
rect 428422 254258 428464 254494
rect 428144 247494 428464 254258
rect 428144 247258 428186 247494
rect 428422 247258 428464 247494
rect 428144 240494 428464 247258
rect 428144 240258 428186 240494
rect 428422 240258 428464 240494
rect 428144 233494 428464 240258
rect 428144 233258 428186 233494
rect 428422 233258 428464 233494
rect 428144 226494 428464 233258
rect 428144 226258 428186 226494
rect 428422 226258 428464 226494
rect 428144 219494 428464 226258
rect 428144 219258 428186 219494
rect 428422 219258 428464 219494
rect 428144 212494 428464 219258
rect 428144 212258 428186 212494
rect 428422 212258 428464 212494
rect 428144 205494 428464 212258
rect 428144 205258 428186 205494
rect 428422 205258 428464 205494
rect 428144 198494 428464 205258
rect 428144 198258 428186 198494
rect 428422 198258 428464 198494
rect 428144 191494 428464 198258
rect 428144 191258 428186 191494
rect 428422 191258 428464 191494
rect 428144 184494 428464 191258
rect 428144 184258 428186 184494
rect 428422 184258 428464 184494
rect 428144 177494 428464 184258
rect 428144 177258 428186 177494
rect 428422 177258 428464 177494
rect 428144 170494 428464 177258
rect 428144 170258 428186 170494
rect 428422 170258 428464 170494
rect 428144 163494 428464 170258
rect 428144 163258 428186 163494
rect 428422 163258 428464 163494
rect 428144 156494 428464 163258
rect 428144 156258 428186 156494
rect 428422 156258 428464 156494
rect 428144 149494 428464 156258
rect 428144 149258 428186 149494
rect 428422 149258 428464 149494
rect 428144 142494 428464 149258
rect 428144 142258 428186 142494
rect 428422 142258 428464 142494
rect 428144 135494 428464 142258
rect 428144 135258 428186 135494
rect 428422 135258 428464 135494
rect 428144 128494 428464 135258
rect 428144 128258 428186 128494
rect 428422 128258 428464 128494
rect 428144 121494 428464 128258
rect 428144 121258 428186 121494
rect 428422 121258 428464 121494
rect 428144 114494 428464 121258
rect 428144 114258 428186 114494
rect 428422 114258 428464 114494
rect 428144 107494 428464 114258
rect 428144 107258 428186 107494
rect 428422 107258 428464 107494
rect 428144 100494 428464 107258
rect 428144 100258 428186 100494
rect 428422 100258 428464 100494
rect 428144 93494 428464 100258
rect 428144 93258 428186 93494
rect 428422 93258 428464 93494
rect 428144 86494 428464 93258
rect 428144 86258 428186 86494
rect 428422 86258 428464 86494
rect 428144 79494 428464 86258
rect 428144 79258 428186 79494
rect 428422 79258 428464 79494
rect 428144 72494 428464 79258
rect 428144 72258 428186 72494
rect 428422 72258 428464 72494
rect 428144 65494 428464 72258
rect 428144 65258 428186 65494
rect 428422 65258 428464 65494
rect 428144 58494 428464 65258
rect 428144 58258 428186 58494
rect 428422 58258 428464 58494
rect 428144 51494 428464 58258
rect 428144 51258 428186 51494
rect 428422 51258 428464 51494
rect 428144 44494 428464 51258
rect 428144 44258 428186 44494
rect 428422 44258 428464 44494
rect 428144 37494 428464 44258
rect 428144 37258 428186 37494
rect 428422 37258 428464 37494
rect 428144 30494 428464 37258
rect 428144 30258 428186 30494
rect 428422 30258 428464 30494
rect 428144 23494 428464 30258
rect 428144 23258 428186 23494
rect 428422 23258 428464 23494
rect 428144 16494 428464 23258
rect 428144 16258 428186 16494
rect 428422 16258 428464 16494
rect 428144 9494 428464 16258
rect 428144 9258 428186 9494
rect 428422 9258 428464 9494
rect 428144 2494 428464 9258
rect 428144 2258 428186 2494
rect 428422 2258 428464 2494
rect 428144 -746 428464 2258
rect 428144 -982 428186 -746
rect 428422 -982 428464 -746
rect 428144 -1066 428464 -982
rect 428144 -1302 428186 -1066
rect 428422 -1302 428464 -1066
rect 428144 -2294 428464 -1302
rect 429876 706198 430196 706230
rect 429876 705962 429918 706198
rect 430154 705962 430196 706198
rect 429876 705878 430196 705962
rect 429876 705642 429918 705878
rect 430154 705642 430196 705878
rect 429876 696434 430196 705642
rect 429876 696198 429918 696434
rect 430154 696198 430196 696434
rect 429876 689434 430196 696198
rect 429876 689198 429918 689434
rect 430154 689198 430196 689434
rect 429876 682434 430196 689198
rect 429876 682198 429918 682434
rect 430154 682198 430196 682434
rect 429876 675434 430196 682198
rect 429876 675198 429918 675434
rect 430154 675198 430196 675434
rect 429876 668434 430196 675198
rect 429876 668198 429918 668434
rect 430154 668198 430196 668434
rect 429876 661434 430196 668198
rect 429876 661198 429918 661434
rect 430154 661198 430196 661434
rect 429876 654434 430196 661198
rect 429876 654198 429918 654434
rect 430154 654198 430196 654434
rect 429876 647434 430196 654198
rect 429876 647198 429918 647434
rect 430154 647198 430196 647434
rect 429876 640434 430196 647198
rect 429876 640198 429918 640434
rect 430154 640198 430196 640434
rect 429876 633434 430196 640198
rect 429876 633198 429918 633434
rect 430154 633198 430196 633434
rect 429876 626434 430196 633198
rect 429876 626198 429918 626434
rect 430154 626198 430196 626434
rect 429876 619434 430196 626198
rect 429876 619198 429918 619434
rect 430154 619198 430196 619434
rect 429876 612434 430196 619198
rect 429876 612198 429918 612434
rect 430154 612198 430196 612434
rect 429876 605434 430196 612198
rect 429876 605198 429918 605434
rect 430154 605198 430196 605434
rect 429876 598434 430196 605198
rect 429876 598198 429918 598434
rect 430154 598198 430196 598434
rect 429876 591434 430196 598198
rect 429876 591198 429918 591434
rect 430154 591198 430196 591434
rect 429876 584434 430196 591198
rect 429876 584198 429918 584434
rect 430154 584198 430196 584434
rect 429876 577434 430196 584198
rect 429876 577198 429918 577434
rect 430154 577198 430196 577434
rect 429876 570434 430196 577198
rect 429876 570198 429918 570434
rect 430154 570198 430196 570434
rect 429876 563434 430196 570198
rect 429876 563198 429918 563434
rect 430154 563198 430196 563434
rect 429876 556434 430196 563198
rect 429876 556198 429918 556434
rect 430154 556198 430196 556434
rect 429876 549434 430196 556198
rect 429876 549198 429918 549434
rect 430154 549198 430196 549434
rect 429876 542434 430196 549198
rect 429876 542198 429918 542434
rect 430154 542198 430196 542434
rect 429876 535434 430196 542198
rect 429876 535198 429918 535434
rect 430154 535198 430196 535434
rect 429876 528434 430196 535198
rect 429876 528198 429918 528434
rect 430154 528198 430196 528434
rect 429876 521434 430196 528198
rect 429876 521198 429918 521434
rect 430154 521198 430196 521434
rect 429876 514434 430196 521198
rect 429876 514198 429918 514434
rect 430154 514198 430196 514434
rect 429876 507434 430196 514198
rect 429876 507198 429918 507434
rect 430154 507198 430196 507434
rect 429876 500434 430196 507198
rect 429876 500198 429918 500434
rect 430154 500198 430196 500434
rect 429876 493434 430196 500198
rect 429876 493198 429918 493434
rect 430154 493198 430196 493434
rect 429876 486434 430196 493198
rect 429876 486198 429918 486434
rect 430154 486198 430196 486434
rect 429876 479434 430196 486198
rect 429876 479198 429918 479434
rect 430154 479198 430196 479434
rect 429876 472434 430196 479198
rect 429876 472198 429918 472434
rect 430154 472198 430196 472434
rect 429876 465434 430196 472198
rect 429876 465198 429918 465434
rect 430154 465198 430196 465434
rect 429876 458434 430196 465198
rect 429876 458198 429918 458434
rect 430154 458198 430196 458434
rect 429876 451434 430196 458198
rect 429876 451198 429918 451434
rect 430154 451198 430196 451434
rect 429876 444434 430196 451198
rect 429876 444198 429918 444434
rect 430154 444198 430196 444434
rect 429876 437434 430196 444198
rect 429876 437198 429918 437434
rect 430154 437198 430196 437434
rect 429876 430434 430196 437198
rect 429876 430198 429918 430434
rect 430154 430198 430196 430434
rect 429876 423434 430196 430198
rect 429876 423198 429918 423434
rect 430154 423198 430196 423434
rect 429876 416434 430196 423198
rect 429876 416198 429918 416434
rect 430154 416198 430196 416434
rect 429876 409434 430196 416198
rect 429876 409198 429918 409434
rect 430154 409198 430196 409434
rect 429876 402434 430196 409198
rect 429876 402198 429918 402434
rect 430154 402198 430196 402434
rect 429876 395434 430196 402198
rect 429876 395198 429918 395434
rect 430154 395198 430196 395434
rect 429876 388434 430196 395198
rect 429876 388198 429918 388434
rect 430154 388198 430196 388434
rect 429876 381434 430196 388198
rect 429876 381198 429918 381434
rect 430154 381198 430196 381434
rect 429876 374434 430196 381198
rect 429876 374198 429918 374434
rect 430154 374198 430196 374434
rect 429876 367434 430196 374198
rect 429876 367198 429918 367434
rect 430154 367198 430196 367434
rect 429876 360434 430196 367198
rect 429876 360198 429918 360434
rect 430154 360198 430196 360434
rect 429876 353434 430196 360198
rect 429876 353198 429918 353434
rect 430154 353198 430196 353434
rect 429876 346434 430196 353198
rect 429876 346198 429918 346434
rect 430154 346198 430196 346434
rect 429876 339434 430196 346198
rect 429876 339198 429918 339434
rect 430154 339198 430196 339434
rect 429876 332434 430196 339198
rect 429876 332198 429918 332434
rect 430154 332198 430196 332434
rect 429876 325434 430196 332198
rect 429876 325198 429918 325434
rect 430154 325198 430196 325434
rect 429876 318434 430196 325198
rect 429876 318198 429918 318434
rect 430154 318198 430196 318434
rect 429876 311434 430196 318198
rect 429876 311198 429918 311434
rect 430154 311198 430196 311434
rect 429876 304434 430196 311198
rect 429876 304198 429918 304434
rect 430154 304198 430196 304434
rect 429876 297434 430196 304198
rect 429876 297198 429918 297434
rect 430154 297198 430196 297434
rect 429876 290434 430196 297198
rect 429876 290198 429918 290434
rect 430154 290198 430196 290434
rect 429876 283434 430196 290198
rect 429876 283198 429918 283434
rect 430154 283198 430196 283434
rect 429876 276434 430196 283198
rect 429876 276198 429918 276434
rect 430154 276198 430196 276434
rect 429876 269434 430196 276198
rect 429876 269198 429918 269434
rect 430154 269198 430196 269434
rect 429876 262434 430196 269198
rect 429876 262198 429918 262434
rect 430154 262198 430196 262434
rect 429876 255434 430196 262198
rect 429876 255198 429918 255434
rect 430154 255198 430196 255434
rect 429876 248434 430196 255198
rect 429876 248198 429918 248434
rect 430154 248198 430196 248434
rect 429876 241434 430196 248198
rect 429876 241198 429918 241434
rect 430154 241198 430196 241434
rect 429876 234434 430196 241198
rect 429876 234198 429918 234434
rect 430154 234198 430196 234434
rect 429876 227434 430196 234198
rect 429876 227198 429918 227434
rect 430154 227198 430196 227434
rect 429876 220434 430196 227198
rect 429876 220198 429918 220434
rect 430154 220198 430196 220434
rect 429876 213434 430196 220198
rect 429876 213198 429918 213434
rect 430154 213198 430196 213434
rect 429876 206434 430196 213198
rect 429876 206198 429918 206434
rect 430154 206198 430196 206434
rect 429876 199434 430196 206198
rect 429876 199198 429918 199434
rect 430154 199198 430196 199434
rect 429876 192434 430196 199198
rect 429876 192198 429918 192434
rect 430154 192198 430196 192434
rect 429876 185434 430196 192198
rect 429876 185198 429918 185434
rect 430154 185198 430196 185434
rect 429876 178434 430196 185198
rect 429876 178198 429918 178434
rect 430154 178198 430196 178434
rect 429876 171434 430196 178198
rect 429876 171198 429918 171434
rect 430154 171198 430196 171434
rect 429876 164434 430196 171198
rect 429876 164198 429918 164434
rect 430154 164198 430196 164434
rect 429876 157434 430196 164198
rect 429876 157198 429918 157434
rect 430154 157198 430196 157434
rect 429876 150434 430196 157198
rect 429876 150198 429918 150434
rect 430154 150198 430196 150434
rect 429876 143434 430196 150198
rect 429876 143198 429918 143434
rect 430154 143198 430196 143434
rect 429876 136434 430196 143198
rect 429876 136198 429918 136434
rect 430154 136198 430196 136434
rect 429876 129434 430196 136198
rect 429876 129198 429918 129434
rect 430154 129198 430196 129434
rect 429876 122434 430196 129198
rect 429876 122198 429918 122434
rect 430154 122198 430196 122434
rect 429876 115434 430196 122198
rect 429876 115198 429918 115434
rect 430154 115198 430196 115434
rect 429876 108434 430196 115198
rect 429876 108198 429918 108434
rect 430154 108198 430196 108434
rect 429876 101434 430196 108198
rect 429876 101198 429918 101434
rect 430154 101198 430196 101434
rect 429876 94434 430196 101198
rect 429876 94198 429918 94434
rect 430154 94198 430196 94434
rect 429876 87434 430196 94198
rect 429876 87198 429918 87434
rect 430154 87198 430196 87434
rect 429876 80434 430196 87198
rect 429876 80198 429918 80434
rect 430154 80198 430196 80434
rect 429876 73434 430196 80198
rect 429876 73198 429918 73434
rect 430154 73198 430196 73434
rect 429876 66434 430196 73198
rect 429876 66198 429918 66434
rect 430154 66198 430196 66434
rect 429876 59434 430196 66198
rect 429876 59198 429918 59434
rect 430154 59198 430196 59434
rect 429876 52434 430196 59198
rect 429876 52198 429918 52434
rect 430154 52198 430196 52434
rect 429876 45434 430196 52198
rect 429876 45198 429918 45434
rect 430154 45198 430196 45434
rect 429876 38434 430196 45198
rect 429876 38198 429918 38434
rect 430154 38198 430196 38434
rect 429876 31434 430196 38198
rect 429876 31198 429918 31434
rect 430154 31198 430196 31434
rect 429876 24434 430196 31198
rect 429876 24198 429918 24434
rect 430154 24198 430196 24434
rect 429876 17434 430196 24198
rect 429876 17198 429918 17434
rect 430154 17198 430196 17434
rect 429876 10434 430196 17198
rect 429876 10198 429918 10434
rect 430154 10198 430196 10434
rect 429876 3434 430196 10198
rect 429876 3198 429918 3434
rect 430154 3198 430196 3434
rect 429876 -1706 430196 3198
rect 429876 -1942 429918 -1706
rect 430154 -1942 430196 -1706
rect 429876 -2026 430196 -1942
rect 429876 -2262 429918 -2026
rect 430154 -2262 430196 -2026
rect 429876 -2294 430196 -2262
rect 435144 705238 435464 706230
rect 435144 705002 435186 705238
rect 435422 705002 435464 705238
rect 435144 704918 435464 705002
rect 435144 704682 435186 704918
rect 435422 704682 435464 704918
rect 435144 695494 435464 704682
rect 435144 695258 435186 695494
rect 435422 695258 435464 695494
rect 435144 688494 435464 695258
rect 435144 688258 435186 688494
rect 435422 688258 435464 688494
rect 435144 681494 435464 688258
rect 435144 681258 435186 681494
rect 435422 681258 435464 681494
rect 435144 674494 435464 681258
rect 435144 674258 435186 674494
rect 435422 674258 435464 674494
rect 435144 667494 435464 674258
rect 435144 667258 435186 667494
rect 435422 667258 435464 667494
rect 435144 660494 435464 667258
rect 435144 660258 435186 660494
rect 435422 660258 435464 660494
rect 435144 653494 435464 660258
rect 435144 653258 435186 653494
rect 435422 653258 435464 653494
rect 435144 646494 435464 653258
rect 435144 646258 435186 646494
rect 435422 646258 435464 646494
rect 435144 639494 435464 646258
rect 435144 639258 435186 639494
rect 435422 639258 435464 639494
rect 435144 632494 435464 639258
rect 435144 632258 435186 632494
rect 435422 632258 435464 632494
rect 435144 625494 435464 632258
rect 435144 625258 435186 625494
rect 435422 625258 435464 625494
rect 435144 618494 435464 625258
rect 435144 618258 435186 618494
rect 435422 618258 435464 618494
rect 435144 611494 435464 618258
rect 435144 611258 435186 611494
rect 435422 611258 435464 611494
rect 435144 604494 435464 611258
rect 435144 604258 435186 604494
rect 435422 604258 435464 604494
rect 435144 597494 435464 604258
rect 435144 597258 435186 597494
rect 435422 597258 435464 597494
rect 435144 590494 435464 597258
rect 435144 590258 435186 590494
rect 435422 590258 435464 590494
rect 435144 583494 435464 590258
rect 435144 583258 435186 583494
rect 435422 583258 435464 583494
rect 435144 576494 435464 583258
rect 435144 576258 435186 576494
rect 435422 576258 435464 576494
rect 435144 569494 435464 576258
rect 435144 569258 435186 569494
rect 435422 569258 435464 569494
rect 435144 562494 435464 569258
rect 435144 562258 435186 562494
rect 435422 562258 435464 562494
rect 435144 555494 435464 562258
rect 435144 555258 435186 555494
rect 435422 555258 435464 555494
rect 435144 548494 435464 555258
rect 435144 548258 435186 548494
rect 435422 548258 435464 548494
rect 435144 541494 435464 548258
rect 435144 541258 435186 541494
rect 435422 541258 435464 541494
rect 435144 534494 435464 541258
rect 435144 534258 435186 534494
rect 435422 534258 435464 534494
rect 435144 527494 435464 534258
rect 435144 527258 435186 527494
rect 435422 527258 435464 527494
rect 435144 520494 435464 527258
rect 435144 520258 435186 520494
rect 435422 520258 435464 520494
rect 435144 513494 435464 520258
rect 435144 513258 435186 513494
rect 435422 513258 435464 513494
rect 435144 506494 435464 513258
rect 435144 506258 435186 506494
rect 435422 506258 435464 506494
rect 435144 499494 435464 506258
rect 435144 499258 435186 499494
rect 435422 499258 435464 499494
rect 435144 492494 435464 499258
rect 435144 492258 435186 492494
rect 435422 492258 435464 492494
rect 435144 485494 435464 492258
rect 435144 485258 435186 485494
rect 435422 485258 435464 485494
rect 435144 478494 435464 485258
rect 435144 478258 435186 478494
rect 435422 478258 435464 478494
rect 435144 471494 435464 478258
rect 435144 471258 435186 471494
rect 435422 471258 435464 471494
rect 435144 464494 435464 471258
rect 435144 464258 435186 464494
rect 435422 464258 435464 464494
rect 435144 457494 435464 464258
rect 435144 457258 435186 457494
rect 435422 457258 435464 457494
rect 435144 450494 435464 457258
rect 435144 450258 435186 450494
rect 435422 450258 435464 450494
rect 435144 443494 435464 450258
rect 435144 443258 435186 443494
rect 435422 443258 435464 443494
rect 435144 436494 435464 443258
rect 435144 436258 435186 436494
rect 435422 436258 435464 436494
rect 435144 429494 435464 436258
rect 435144 429258 435186 429494
rect 435422 429258 435464 429494
rect 435144 422494 435464 429258
rect 435144 422258 435186 422494
rect 435422 422258 435464 422494
rect 435144 415494 435464 422258
rect 435144 415258 435186 415494
rect 435422 415258 435464 415494
rect 435144 408494 435464 415258
rect 435144 408258 435186 408494
rect 435422 408258 435464 408494
rect 435144 401494 435464 408258
rect 435144 401258 435186 401494
rect 435422 401258 435464 401494
rect 435144 394494 435464 401258
rect 435144 394258 435186 394494
rect 435422 394258 435464 394494
rect 435144 387494 435464 394258
rect 435144 387258 435186 387494
rect 435422 387258 435464 387494
rect 435144 380494 435464 387258
rect 435144 380258 435186 380494
rect 435422 380258 435464 380494
rect 435144 373494 435464 380258
rect 435144 373258 435186 373494
rect 435422 373258 435464 373494
rect 435144 366494 435464 373258
rect 435144 366258 435186 366494
rect 435422 366258 435464 366494
rect 435144 359494 435464 366258
rect 435144 359258 435186 359494
rect 435422 359258 435464 359494
rect 435144 352494 435464 359258
rect 435144 352258 435186 352494
rect 435422 352258 435464 352494
rect 435144 345494 435464 352258
rect 435144 345258 435186 345494
rect 435422 345258 435464 345494
rect 435144 338494 435464 345258
rect 435144 338258 435186 338494
rect 435422 338258 435464 338494
rect 435144 331494 435464 338258
rect 435144 331258 435186 331494
rect 435422 331258 435464 331494
rect 435144 324494 435464 331258
rect 435144 324258 435186 324494
rect 435422 324258 435464 324494
rect 435144 317494 435464 324258
rect 435144 317258 435186 317494
rect 435422 317258 435464 317494
rect 435144 310494 435464 317258
rect 435144 310258 435186 310494
rect 435422 310258 435464 310494
rect 435144 303494 435464 310258
rect 435144 303258 435186 303494
rect 435422 303258 435464 303494
rect 435144 296494 435464 303258
rect 435144 296258 435186 296494
rect 435422 296258 435464 296494
rect 435144 289494 435464 296258
rect 435144 289258 435186 289494
rect 435422 289258 435464 289494
rect 435144 282494 435464 289258
rect 435144 282258 435186 282494
rect 435422 282258 435464 282494
rect 435144 275494 435464 282258
rect 435144 275258 435186 275494
rect 435422 275258 435464 275494
rect 435144 268494 435464 275258
rect 435144 268258 435186 268494
rect 435422 268258 435464 268494
rect 435144 261494 435464 268258
rect 435144 261258 435186 261494
rect 435422 261258 435464 261494
rect 435144 254494 435464 261258
rect 435144 254258 435186 254494
rect 435422 254258 435464 254494
rect 435144 247494 435464 254258
rect 435144 247258 435186 247494
rect 435422 247258 435464 247494
rect 435144 240494 435464 247258
rect 435144 240258 435186 240494
rect 435422 240258 435464 240494
rect 435144 233494 435464 240258
rect 435144 233258 435186 233494
rect 435422 233258 435464 233494
rect 435144 226494 435464 233258
rect 435144 226258 435186 226494
rect 435422 226258 435464 226494
rect 435144 219494 435464 226258
rect 435144 219258 435186 219494
rect 435422 219258 435464 219494
rect 435144 212494 435464 219258
rect 435144 212258 435186 212494
rect 435422 212258 435464 212494
rect 435144 205494 435464 212258
rect 435144 205258 435186 205494
rect 435422 205258 435464 205494
rect 435144 198494 435464 205258
rect 435144 198258 435186 198494
rect 435422 198258 435464 198494
rect 435144 191494 435464 198258
rect 435144 191258 435186 191494
rect 435422 191258 435464 191494
rect 435144 184494 435464 191258
rect 435144 184258 435186 184494
rect 435422 184258 435464 184494
rect 435144 177494 435464 184258
rect 435144 177258 435186 177494
rect 435422 177258 435464 177494
rect 435144 170494 435464 177258
rect 435144 170258 435186 170494
rect 435422 170258 435464 170494
rect 435144 163494 435464 170258
rect 435144 163258 435186 163494
rect 435422 163258 435464 163494
rect 435144 156494 435464 163258
rect 435144 156258 435186 156494
rect 435422 156258 435464 156494
rect 435144 149494 435464 156258
rect 435144 149258 435186 149494
rect 435422 149258 435464 149494
rect 435144 142494 435464 149258
rect 435144 142258 435186 142494
rect 435422 142258 435464 142494
rect 435144 135494 435464 142258
rect 435144 135258 435186 135494
rect 435422 135258 435464 135494
rect 435144 128494 435464 135258
rect 435144 128258 435186 128494
rect 435422 128258 435464 128494
rect 435144 121494 435464 128258
rect 435144 121258 435186 121494
rect 435422 121258 435464 121494
rect 435144 114494 435464 121258
rect 435144 114258 435186 114494
rect 435422 114258 435464 114494
rect 435144 107494 435464 114258
rect 435144 107258 435186 107494
rect 435422 107258 435464 107494
rect 435144 100494 435464 107258
rect 435144 100258 435186 100494
rect 435422 100258 435464 100494
rect 435144 93494 435464 100258
rect 435144 93258 435186 93494
rect 435422 93258 435464 93494
rect 435144 86494 435464 93258
rect 435144 86258 435186 86494
rect 435422 86258 435464 86494
rect 435144 79494 435464 86258
rect 435144 79258 435186 79494
rect 435422 79258 435464 79494
rect 435144 72494 435464 79258
rect 435144 72258 435186 72494
rect 435422 72258 435464 72494
rect 435144 65494 435464 72258
rect 435144 65258 435186 65494
rect 435422 65258 435464 65494
rect 435144 58494 435464 65258
rect 435144 58258 435186 58494
rect 435422 58258 435464 58494
rect 435144 51494 435464 58258
rect 435144 51258 435186 51494
rect 435422 51258 435464 51494
rect 435144 44494 435464 51258
rect 435144 44258 435186 44494
rect 435422 44258 435464 44494
rect 435144 37494 435464 44258
rect 435144 37258 435186 37494
rect 435422 37258 435464 37494
rect 435144 30494 435464 37258
rect 435144 30258 435186 30494
rect 435422 30258 435464 30494
rect 435144 23494 435464 30258
rect 435144 23258 435186 23494
rect 435422 23258 435464 23494
rect 435144 16494 435464 23258
rect 435144 16258 435186 16494
rect 435422 16258 435464 16494
rect 435144 9494 435464 16258
rect 435144 9258 435186 9494
rect 435422 9258 435464 9494
rect 435144 2494 435464 9258
rect 435144 2258 435186 2494
rect 435422 2258 435464 2494
rect 435144 -746 435464 2258
rect 435144 -982 435186 -746
rect 435422 -982 435464 -746
rect 435144 -1066 435464 -982
rect 435144 -1302 435186 -1066
rect 435422 -1302 435464 -1066
rect 435144 -2294 435464 -1302
rect 436876 706198 437196 706230
rect 436876 705962 436918 706198
rect 437154 705962 437196 706198
rect 436876 705878 437196 705962
rect 436876 705642 436918 705878
rect 437154 705642 437196 705878
rect 436876 696434 437196 705642
rect 436876 696198 436918 696434
rect 437154 696198 437196 696434
rect 436876 689434 437196 696198
rect 436876 689198 436918 689434
rect 437154 689198 437196 689434
rect 436876 682434 437196 689198
rect 436876 682198 436918 682434
rect 437154 682198 437196 682434
rect 436876 675434 437196 682198
rect 436876 675198 436918 675434
rect 437154 675198 437196 675434
rect 436876 668434 437196 675198
rect 436876 668198 436918 668434
rect 437154 668198 437196 668434
rect 436876 661434 437196 668198
rect 436876 661198 436918 661434
rect 437154 661198 437196 661434
rect 436876 654434 437196 661198
rect 436876 654198 436918 654434
rect 437154 654198 437196 654434
rect 436876 647434 437196 654198
rect 436876 647198 436918 647434
rect 437154 647198 437196 647434
rect 436876 640434 437196 647198
rect 436876 640198 436918 640434
rect 437154 640198 437196 640434
rect 436876 633434 437196 640198
rect 436876 633198 436918 633434
rect 437154 633198 437196 633434
rect 436876 626434 437196 633198
rect 436876 626198 436918 626434
rect 437154 626198 437196 626434
rect 436876 619434 437196 626198
rect 436876 619198 436918 619434
rect 437154 619198 437196 619434
rect 436876 612434 437196 619198
rect 436876 612198 436918 612434
rect 437154 612198 437196 612434
rect 436876 605434 437196 612198
rect 436876 605198 436918 605434
rect 437154 605198 437196 605434
rect 436876 598434 437196 605198
rect 436876 598198 436918 598434
rect 437154 598198 437196 598434
rect 436876 591434 437196 598198
rect 436876 591198 436918 591434
rect 437154 591198 437196 591434
rect 436876 584434 437196 591198
rect 436876 584198 436918 584434
rect 437154 584198 437196 584434
rect 436876 577434 437196 584198
rect 436876 577198 436918 577434
rect 437154 577198 437196 577434
rect 436876 570434 437196 577198
rect 436876 570198 436918 570434
rect 437154 570198 437196 570434
rect 436876 563434 437196 570198
rect 436876 563198 436918 563434
rect 437154 563198 437196 563434
rect 436876 556434 437196 563198
rect 436876 556198 436918 556434
rect 437154 556198 437196 556434
rect 436876 549434 437196 556198
rect 436876 549198 436918 549434
rect 437154 549198 437196 549434
rect 436876 542434 437196 549198
rect 436876 542198 436918 542434
rect 437154 542198 437196 542434
rect 436876 535434 437196 542198
rect 436876 535198 436918 535434
rect 437154 535198 437196 535434
rect 436876 528434 437196 535198
rect 436876 528198 436918 528434
rect 437154 528198 437196 528434
rect 436876 521434 437196 528198
rect 436876 521198 436918 521434
rect 437154 521198 437196 521434
rect 436876 514434 437196 521198
rect 436876 514198 436918 514434
rect 437154 514198 437196 514434
rect 436876 507434 437196 514198
rect 436876 507198 436918 507434
rect 437154 507198 437196 507434
rect 436876 500434 437196 507198
rect 436876 500198 436918 500434
rect 437154 500198 437196 500434
rect 436876 493434 437196 500198
rect 436876 493198 436918 493434
rect 437154 493198 437196 493434
rect 436876 486434 437196 493198
rect 436876 486198 436918 486434
rect 437154 486198 437196 486434
rect 436876 479434 437196 486198
rect 436876 479198 436918 479434
rect 437154 479198 437196 479434
rect 436876 472434 437196 479198
rect 436876 472198 436918 472434
rect 437154 472198 437196 472434
rect 436876 465434 437196 472198
rect 436876 465198 436918 465434
rect 437154 465198 437196 465434
rect 436876 458434 437196 465198
rect 436876 458198 436918 458434
rect 437154 458198 437196 458434
rect 436876 451434 437196 458198
rect 436876 451198 436918 451434
rect 437154 451198 437196 451434
rect 436876 444434 437196 451198
rect 436876 444198 436918 444434
rect 437154 444198 437196 444434
rect 436876 437434 437196 444198
rect 436876 437198 436918 437434
rect 437154 437198 437196 437434
rect 436876 430434 437196 437198
rect 436876 430198 436918 430434
rect 437154 430198 437196 430434
rect 436876 423434 437196 430198
rect 436876 423198 436918 423434
rect 437154 423198 437196 423434
rect 436876 416434 437196 423198
rect 436876 416198 436918 416434
rect 437154 416198 437196 416434
rect 436876 409434 437196 416198
rect 436876 409198 436918 409434
rect 437154 409198 437196 409434
rect 436876 402434 437196 409198
rect 436876 402198 436918 402434
rect 437154 402198 437196 402434
rect 436876 395434 437196 402198
rect 436876 395198 436918 395434
rect 437154 395198 437196 395434
rect 436876 388434 437196 395198
rect 436876 388198 436918 388434
rect 437154 388198 437196 388434
rect 436876 381434 437196 388198
rect 436876 381198 436918 381434
rect 437154 381198 437196 381434
rect 436876 374434 437196 381198
rect 436876 374198 436918 374434
rect 437154 374198 437196 374434
rect 436876 367434 437196 374198
rect 436876 367198 436918 367434
rect 437154 367198 437196 367434
rect 436876 360434 437196 367198
rect 436876 360198 436918 360434
rect 437154 360198 437196 360434
rect 436876 353434 437196 360198
rect 436876 353198 436918 353434
rect 437154 353198 437196 353434
rect 436876 346434 437196 353198
rect 436876 346198 436918 346434
rect 437154 346198 437196 346434
rect 436876 339434 437196 346198
rect 436876 339198 436918 339434
rect 437154 339198 437196 339434
rect 436876 332434 437196 339198
rect 436876 332198 436918 332434
rect 437154 332198 437196 332434
rect 436876 325434 437196 332198
rect 436876 325198 436918 325434
rect 437154 325198 437196 325434
rect 436876 318434 437196 325198
rect 436876 318198 436918 318434
rect 437154 318198 437196 318434
rect 436876 311434 437196 318198
rect 436876 311198 436918 311434
rect 437154 311198 437196 311434
rect 436876 304434 437196 311198
rect 436876 304198 436918 304434
rect 437154 304198 437196 304434
rect 436876 297434 437196 304198
rect 436876 297198 436918 297434
rect 437154 297198 437196 297434
rect 436876 290434 437196 297198
rect 436876 290198 436918 290434
rect 437154 290198 437196 290434
rect 436876 283434 437196 290198
rect 436876 283198 436918 283434
rect 437154 283198 437196 283434
rect 436876 276434 437196 283198
rect 436876 276198 436918 276434
rect 437154 276198 437196 276434
rect 436876 269434 437196 276198
rect 436876 269198 436918 269434
rect 437154 269198 437196 269434
rect 436876 262434 437196 269198
rect 436876 262198 436918 262434
rect 437154 262198 437196 262434
rect 436876 255434 437196 262198
rect 436876 255198 436918 255434
rect 437154 255198 437196 255434
rect 436876 248434 437196 255198
rect 436876 248198 436918 248434
rect 437154 248198 437196 248434
rect 436876 241434 437196 248198
rect 436876 241198 436918 241434
rect 437154 241198 437196 241434
rect 436876 234434 437196 241198
rect 436876 234198 436918 234434
rect 437154 234198 437196 234434
rect 436876 227434 437196 234198
rect 436876 227198 436918 227434
rect 437154 227198 437196 227434
rect 436876 220434 437196 227198
rect 436876 220198 436918 220434
rect 437154 220198 437196 220434
rect 436876 213434 437196 220198
rect 436876 213198 436918 213434
rect 437154 213198 437196 213434
rect 436876 206434 437196 213198
rect 436876 206198 436918 206434
rect 437154 206198 437196 206434
rect 436876 199434 437196 206198
rect 436876 199198 436918 199434
rect 437154 199198 437196 199434
rect 436876 192434 437196 199198
rect 436876 192198 436918 192434
rect 437154 192198 437196 192434
rect 436876 185434 437196 192198
rect 436876 185198 436918 185434
rect 437154 185198 437196 185434
rect 436876 178434 437196 185198
rect 436876 178198 436918 178434
rect 437154 178198 437196 178434
rect 436876 171434 437196 178198
rect 436876 171198 436918 171434
rect 437154 171198 437196 171434
rect 436876 164434 437196 171198
rect 436876 164198 436918 164434
rect 437154 164198 437196 164434
rect 436876 157434 437196 164198
rect 436876 157198 436918 157434
rect 437154 157198 437196 157434
rect 436876 150434 437196 157198
rect 436876 150198 436918 150434
rect 437154 150198 437196 150434
rect 436876 143434 437196 150198
rect 436876 143198 436918 143434
rect 437154 143198 437196 143434
rect 436876 136434 437196 143198
rect 436876 136198 436918 136434
rect 437154 136198 437196 136434
rect 436876 129434 437196 136198
rect 436876 129198 436918 129434
rect 437154 129198 437196 129434
rect 436876 122434 437196 129198
rect 436876 122198 436918 122434
rect 437154 122198 437196 122434
rect 436876 115434 437196 122198
rect 436876 115198 436918 115434
rect 437154 115198 437196 115434
rect 436876 108434 437196 115198
rect 436876 108198 436918 108434
rect 437154 108198 437196 108434
rect 436876 101434 437196 108198
rect 436876 101198 436918 101434
rect 437154 101198 437196 101434
rect 436876 94434 437196 101198
rect 436876 94198 436918 94434
rect 437154 94198 437196 94434
rect 436876 87434 437196 94198
rect 436876 87198 436918 87434
rect 437154 87198 437196 87434
rect 436876 80434 437196 87198
rect 436876 80198 436918 80434
rect 437154 80198 437196 80434
rect 436876 73434 437196 80198
rect 436876 73198 436918 73434
rect 437154 73198 437196 73434
rect 436876 66434 437196 73198
rect 436876 66198 436918 66434
rect 437154 66198 437196 66434
rect 436876 59434 437196 66198
rect 436876 59198 436918 59434
rect 437154 59198 437196 59434
rect 436876 52434 437196 59198
rect 436876 52198 436918 52434
rect 437154 52198 437196 52434
rect 436876 45434 437196 52198
rect 436876 45198 436918 45434
rect 437154 45198 437196 45434
rect 436876 38434 437196 45198
rect 436876 38198 436918 38434
rect 437154 38198 437196 38434
rect 436876 31434 437196 38198
rect 436876 31198 436918 31434
rect 437154 31198 437196 31434
rect 436876 24434 437196 31198
rect 436876 24198 436918 24434
rect 437154 24198 437196 24434
rect 436876 17434 437196 24198
rect 436876 17198 436918 17434
rect 437154 17198 437196 17434
rect 436876 10434 437196 17198
rect 436876 10198 436918 10434
rect 437154 10198 437196 10434
rect 436876 3434 437196 10198
rect 436876 3198 436918 3434
rect 437154 3198 437196 3434
rect 436876 -1706 437196 3198
rect 436876 -1942 436918 -1706
rect 437154 -1942 437196 -1706
rect 436876 -2026 437196 -1942
rect 436876 -2262 436918 -2026
rect 437154 -2262 437196 -2026
rect 436876 -2294 437196 -2262
rect 442144 705238 442464 706230
rect 442144 705002 442186 705238
rect 442422 705002 442464 705238
rect 442144 704918 442464 705002
rect 442144 704682 442186 704918
rect 442422 704682 442464 704918
rect 442144 695494 442464 704682
rect 442144 695258 442186 695494
rect 442422 695258 442464 695494
rect 442144 688494 442464 695258
rect 442144 688258 442186 688494
rect 442422 688258 442464 688494
rect 442144 681494 442464 688258
rect 442144 681258 442186 681494
rect 442422 681258 442464 681494
rect 442144 674494 442464 681258
rect 442144 674258 442186 674494
rect 442422 674258 442464 674494
rect 442144 667494 442464 674258
rect 442144 667258 442186 667494
rect 442422 667258 442464 667494
rect 442144 660494 442464 667258
rect 442144 660258 442186 660494
rect 442422 660258 442464 660494
rect 442144 653494 442464 660258
rect 442144 653258 442186 653494
rect 442422 653258 442464 653494
rect 442144 646494 442464 653258
rect 442144 646258 442186 646494
rect 442422 646258 442464 646494
rect 442144 639494 442464 646258
rect 442144 639258 442186 639494
rect 442422 639258 442464 639494
rect 442144 632494 442464 639258
rect 442144 632258 442186 632494
rect 442422 632258 442464 632494
rect 442144 625494 442464 632258
rect 442144 625258 442186 625494
rect 442422 625258 442464 625494
rect 442144 618494 442464 625258
rect 442144 618258 442186 618494
rect 442422 618258 442464 618494
rect 442144 611494 442464 618258
rect 442144 611258 442186 611494
rect 442422 611258 442464 611494
rect 442144 604494 442464 611258
rect 442144 604258 442186 604494
rect 442422 604258 442464 604494
rect 442144 597494 442464 604258
rect 442144 597258 442186 597494
rect 442422 597258 442464 597494
rect 442144 590494 442464 597258
rect 442144 590258 442186 590494
rect 442422 590258 442464 590494
rect 442144 583494 442464 590258
rect 442144 583258 442186 583494
rect 442422 583258 442464 583494
rect 442144 576494 442464 583258
rect 442144 576258 442186 576494
rect 442422 576258 442464 576494
rect 442144 569494 442464 576258
rect 442144 569258 442186 569494
rect 442422 569258 442464 569494
rect 442144 562494 442464 569258
rect 442144 562258 442186 562494
rect 442422 562258 442464 562494
rect 442144 555494 442464 562258
rect 442144 555258 442186 555494
rect 442422 555258 442464 555494
rect 442144 548494 442464 555258
rect 442144 548258 442186 548494
rect 442422 548258 442464 548494
rect 442144 541494 442464 548258
rect 442144 541258 442186 541494
rect 442422 541258 442464 541494
rect 442144 534494 442464 541258
rect 442144 534258 442186 534494
rect 442422 534258 442464 534494
rect 442144 527494 442464 534258
rect 442144 527258 442186 527494
rect 442422 527258 442464 527494
rect 442144 520494 442464 527258
rect 442144 520258 442186 520494
rect 442422 520258 442464 520494
rect 442144 513494 442464 520258
rect 442144 513258 442186 513494
rect 442422 513258 442464 513494
rect 442144 506494 442464 513258
rect 442144 506258 442186 506494
rect 442422 506258 442464 506494
rect 442144 499494 442464 506258
rect 442144 499258 442186 499494
rect 442422 499258 442464 499494
rect 442144 492494 442464 499258
rect 442144 492258 442186 492494
rect 442422 492258 442464 492494
rect 442144 485494 442464 492258
rect 442144 485258 442186 485494
rect 442422 485258 442464 485494
rect 442144 478494 442464 485258
rect 442144 478258 442186 478494
rect 442422 478258 442464 478494
rect 442144 471494 442464 478258
rect 442144 471258 442186 471494
rect 442422 471258 442464 471494
rect 442144 464494 442464 471258
rect 442144 464258 442186 464494
rect 442422 464258 442464 464494
rect 442144 457494 442464 464258
rect 442144 457258 442186 457494
rect 442422 457258 442464 457494
rect 442144 450494 442464 457258
rect 442144 450258 442186 450494
rect 442422 450258 442464 450494
rect 442144 443494 442464 450258
rect 442144 443258 442186 443494
rect 442422 443258 442464 443494
rect 442144 436494 442464 443258
rect 442144 436258 442186 436494
rect 442422 436258 442464 436494
rect 442144 429494 442464 436258
rect 442144 429258 442186 429494
rect 442422 429258 442464 429494
rect 442144 422494 442464 429258
rect 442144 422258 442186 422494
rect 442422 422258 442464 422494
rect 442144 415494 442464 422258
rect 442144 415258 442186 415494
rect 442422 415258 442464 415494
rect 442144 408494 442464 415258
rect 442144 408258 442186 408494
rect 442422 408258 442464 408494
rect 442144 401494 442464 408258
rect 442144 401258 442186 401494
rect 442422 401258 442464 401494
rect 442144 394494 442464 401258
rect 442144 394258 442186 394494
rect 442422 394258 442464 394494
rect 442144 387494 442464 394258
rect 442144 387258 442186 387494
rect 442422 387258 442464 387494
rect 442144 380494 442464 387258
rect 442144 380258 442186 380494
rect 442422 380258 442464 380494
rect 442144 373494 442464 380258
rect 442144 373258 442186 373494
rect 442422 373258 442464 373494
rect 442144 366494 442464 373258
rect 442144 366258 442186 366494
rect 442422 366258 442464 366494
rect 442144 359494 442464 366258
rect 442144 359258 442186 359494
rect 442422 359258 442464 359494
rect 442144 352494 442464 359258
rect 442144 352258 442186 352494
rect 442422 352258 442464 352494
rect 442144 345494 442464 352258
rect 442144 345258 442186 345494
rect 442422 345258 442464 345494
rect 442144 338494 442464 345258
rect 442144 338258 442186 338494
rect 442422 338258 442464 338494
rect 442144 331494 442464 338258
rect 442144 331258 442186 331494
rect 442422 331258 442464 331494
rect 442144 324494 442464 331258
rect 442144 324258 442186 324494
rect 442422 324258 442464 324494
rect 442144 317494 442464 324258
rect 442144 317258 442186 317494
rect 442422 317258 442464 317494
rect 442144 310494 442464 317258
rect 442144 310258 442186 310494
rect 442422 310258 442464 310494
rect 442144 303494 442464 310258
rect 442144 303258 442186 303494
rect 442422 303258 442464 303494
rect 442144 296494 442464 303258
rect 442144 296258 442186 296494
rect 442422 296258 442464 296494
rect 442144 289494 442464 296258
rect 442144 289258 442186 289494
rect 442422 289258 442464 289494
rect 442144 282494 442464 289258
rect 442144 282258 442186 282494
rect 442422 282258 442464 282494
rect 442144 275494 442464 282258
rect 442144 275258 442186 275494
rect 442422 275258 442464 275494
rect 442144 268494 442464 275258
rect 442144 268258 442186 268494
rect 442422 268258 442464 268494
rect 442144 261494 442464 268258
rect 442144 261258 442186 261494
rect 442422 261258 442464 261494
rect 442144 254494 442464 261258
rect 442144 254258 442186 254494
rect 442422 254258 442464 254494
rect 442144 247494 442464 254258
rect 442144 247258 442186 247494
rect 442422 247258 442464 247494
rect 442144 240494 442464 247258
rect 442144 240258 442186 240494
rect 442422 240258 442464 240494
rect 442144 233494 442464 240258
rect 442144 233258 442186 233494
rect 442422 233258 442464 233494
rect 442144 226494 442464 233258
rect 442144 226258 442186 226494
rect 442422 226258 442464 226494
rect 442144 219494 442464 226258
rect 442144 219258 442186 219494
rect 442422 219258 442464 219494
rect 442144 212494 442464 219258
rect 442144 212258 442186 212494
rect 442422 212258 442464 212494
rect 442144 205494 442464 212258
rect 442144 205258 442186 205494
rect 442422 205258 442464 205494
rect 442144 198494 442464 205258
rect 442144 198258 442186 198494
rect 442422 198258 442464 198494
rect 442144 191494 442464 198258
rect 442144 191258 442186 191494
rect 442422 191258 442464 191494
rect 442144 184494 442464 191258
rect 442144 184258 442186 184494
rect 442422 184258 442464 184494
rect 442144 177494 442464 184258
rect 442144 177258 442186 177494
rect 442422 177258 442464 177494
rect 442144 170494 442464 177258
rect 442144 170258 442186 170494
rect 442422 170258 442464 170494
rect 442144 163494 442464 170258
rect 442144 163258 442186 163494
rect 442422 163258 442464 163494
rect 442144 156494 442464 163258
rect 442144 156258 442186 156494
rect 442422 156258 442464 156494
rect 442144 149494 442464 156258
rect 442144 149258 442186 149494
rect 442422 149258 442464 149494
rect 442144 142494 442464 149258
rect 442144 142258 442186 142494
rect 442422 142258 442464 142494
rect 442144 135494 442464 142258
rect 442144 135258 442186 135494
rect 442422 135258 442464 135494
rect 442144 128494 442464 135258
rect 442144 128258 442186 128494
rect 442422 128258 442464 128494
rect 442144 121494 442464 128258
rect 442144 121258 442186 121494
rect 442422 121258 442464 121494
rect 442144 114494 442464 121258
rect 442144 114258 442186 114494
rect 442422 114258 442464 114494
rect 442144 107494 442464 114258
rect 442144 107258 442186 107494
rect 442422 107258 442464 107494
rect 442144 100494 442464 107258
rect 442144 100258 442186 100494
rect 442422 100258 442464 100494
rect 442144 93494 442464 100258
rect 442144 93258 442186 93494
rect 442422 93258 442464 93494
rect 442144 86494 442464 93258
rect 442144 86258 442186 86494
rect 442422 86258 442464 86494
rect 442144 79494 442464 86258
rect 442144 79258 442186 79494
rect 442422 79258 442464 79494
rect 442144 72494 442464 79258
rect 442144 72258 442186 72494
rect 442422 72258 442464 72494
rect 442144 65494 442464 72258
rect 442144 65258 442186 65494
rect 442422 65258 442464 65494
rect 442144 58494 442464 65258
rect 442144 58258 442186 58494
rect 442422 58258 442464 58494
rect 442144 51494 442464 58258
rect 442144 51258 442186 51494
rect 442422 51258 442464 51494
rect 442144 44494 442464 51258
rect 442144 44258 442186 44494
rect 442422 44258 442464 44494
rect 442144 37494 442464 44258
rect 442144 37258 442186 37494
rect 442422 37258 442464 37494
rect 442144 30494 442464 37258
rect 442144 30258 442186 30494
rect 442422 30258 442464 30494
rect 442144 23494 442464 30258
rect 442144 23258 442186 23494
rect 442422 23258 442464 23494
rect 442144 16494 442464 23258
rect 442144 16258 442186 16494
rect 442422 16258 442464 16494
rect 442144 9494 442464 16258
rect 442144 9258 442186 9494
rect 442422 9258 442464 9494
rect 442144 2494 442464 9258
rect 442144 2258 442186 2494
rect 442422 2258 442464 2494
rect 442144 -746 442464 2258
rect 442144 -982 442186 -746
rect 442422 -982 442464 -746
rect 442144 -1066 442464 -982
rect 442144 -1302 442186 -1066
rect 442422 -1302 442464 -1066
rect 442144 -2294 442464 -1302
rect 443876 706198 444196 706230
rect 443876 705962 443918 706198
rect 444154 705962 444196 706198
rect 443876 705878 444196 705962
rect 443876 705642 443918 705878
rect 444154 705642 444196 705878
rect 443876 696434 444196 705642
rect 443876 696198 443918 696434
rect 444154 696198 444196 696434
rect 443876 689434 444196 696198
rect 443876 689198 443918 689434
rect 444154 689198 444196 689434
rect 443876 682434 444196 689198
rect 443876 682198 443918 682434
rect 444154 682198 444196 682434
rect 443876 675434 444196 682198
rect 443876 675198 443918 675434
rect 444154 675198 444196 675434
rect 443876 668434 444196 675198
rect 443876 668198 443918 668434
rect 444154 668198 444196 668434
rect 443876 661434 444196 668198
rect 443876 661198 443918 661434
rect 444154 661198 444196 661434
rect 443876 654434 444196 661198
rect 443876 654198 443918 654434
rect 444154 654198 444196 654434
rect 443876 647434 444196 654198
rect 443876 647198 443918 647434
rect 444154 647198 444196 647434
rect 443876 640434 444196 647198
rect 443876 640198 443918 640434
rect 444154 640198 444196 640434
rect 443876 633434 444196 640198
rect 443876 633198 443918 633434
rect 444154 633198 444196 633434
rect 443876 626434 444196 633198
rect 443876 626198 443918 626434
rect 444154 626198 444196 626434
rect 443876 619434 444196 626198
rect 443876 619198 443918 619434
rect 444154 619198 444196 619434
rect 443876 612434 444196 619198
rect 443876 612198 443918 612434
rect 444154 612198 444196 612434
rect 443876 605434 444196 612198
rect 443876 605198 443918 605434
rect 444154 605198 444196 605434
rect 443876 598434 444196 605198
rect 443876 598198 443918 598434
rect 444154 598198 444196 598434
rect 443876 591434 444196 598198
rect 443876 591198 443918 591434
rect 444154 591198 444196 591434
rect 443876 584434 444196 591198
rect 443876 584198 443918 584434
rect 444154 584198 444196 584434
rect 443876 577434 444196 584198
rect 443876 577198 443918 577434
rect 444154 577198 444196 577434
rect 443876 570434 444196 577198
rect 443876 570198 443918 570434
rect 444154 570198 444196 570434
rect 443876 563434 444196 570198
rect 443876 563198 443918 563434
rect 444154 563198 444196 563434
rect 443876 556434 444196 563198
rect 443876 556198 443918 556434
rect 444154 556198 444196 556434
rect 443876 549434 444196 556198
rect 443876 549198 443918 549434
rect 444154 549198 444196 549434
rect 443876 542434 444196 549198
rect 443876 542198 443918 542434
rect 444154 542198 444196 542434
rect 443876 535434 444196 542198
rect 443876 535198 443918 535434
rect 444154 535198 444196 535434
rect 443876 528434 444196 535198
rect 443876 528198 443918 528434
rect 444154 528198 444196 528434
rect 443876 521434 444196 528198
rect 443876 521198 443918 521434
rect 444154 521198 444196 521434
rect 443876 514434 444196 521198
rect 443876 514198 443918 514434
rect 444154 514198 444196 514434
rect 443876 507434 444196 514198
rect 443876 507198 443918 507434
rect 444154 507198 444196 507434
rect 443876 500434 444196 507198
rect 443876 500198 443918 500434
rect 444154 500198 444196 500434
rect 443876 493434 444196 500198
rect 443876 493198 443918 493434
rect 444154 493198 444196 493434
rect 443876 486434 444196 493198
rect 443876 486198 443918 486434
rect 444154 486198 444196 486434
rect 443876 479434 444196 486198
rect 443876 479198 443918 479434
rect 444154 479198 444196 479434
rect 443876 472434 444196 479198
rect 443876 472198 443918 472434
rect 444154 472198 444196 472434
rect 443876 465434 444196 472198
rect 443876 465198 443918 465434
rect 444154 465198 444196 465434
rect 443876 458434 444196 465198
rect 443876 458198 443918 458434
rect 444154 458198 444196 458434
rect 443876 451434 444196 458198
rect 443876 451198 443918 451434
rect 444154 451198 444196 451434
rect 443876 444434 444196 451198
rect 443876 444198 443918 444434
rect 444154 444198 444196 444434
rect 443876 437434 444196 444198
rect 443876 437198 443918 437434
rect 444154 437198 444196 437434
rect 443876 430434 444196 437198
rect 443876 430198 443918 430434
rect 444154 430198 444196 430434
rect 443876 423434 444196 430198
rect 443876 423198 443918 423434
rect 444154 423198 444196 423434
rect 443876 416434 444196 423198
rect 443876 416198 443918 416434
rect 444154 416198 444196 416434
rect 443876 409434 444196 416198
rect 443876 409198 443918 409434
rect 444154 409198 444196 409434
rect 443876 402434 444196 409198
rect 443876 402198 443918 402434
rect 444154 402198 444196 402434
rect 443876 395434 444196 402198
rect 443876 395198 443918 395434
rect 444154 395198 444196 395434
rect 443876 388434 444196 395198
rect 443876 388198 443918 388434
rect 444154 388198 444196 388434
rect 443876 381434 444196 388198
rect 443876 381198 443918 381434
rect 444154 381198 444196 381434
rect 443876 374434 444196 381198
rect 443876 374198 443918 374434
rect 444154 374198 444196 374434
rect 443876 367434 444196 374198
rect 443876 367198 443918 367434
rect 444154 367198 444196 367434
rect 443876 360434 444196 367198
rect 443876 360198 443918 360434
rect 444154 360198 444196 360434
rect 443876 353434 444196 360198
rect 443876 353198 443918 353434
rect 444154 353198 444196 353434
rect 443876 346434 444196 353198
rect 443876 346198 443918 346434
rect 444154 346198 444196 346434
rect 443876 339434 444196 346198
rect 443876 339198 443918 339434
rect 444154 339198 444196 339434
rect 443876 332434 444196 339198
rect 443876 332198 443918 332434
rect 444154 332198 444196 332434
rect 443876 325434 444196 332198
rect 443876 325198 443918 325434
rect 444154 325198 444196 325434
rect 443876 318434 444196 325198
rect 443876 318198 443918 318434
rect 444154 318198 444196 318434
rect 443876 311434 444196 318198
rect 443876 311198 443918 311434
rect 444154 311198 444196 311434
rect 443876 304434 444196 311198
rect 443876 304198 443918 304434
rect 444154 304198 444196 304434
rect 443876 297434 444196 304198
rect 443876 297198 443918 297434
rect 444154 297198 444196 297434
rect 443876 290434 444196 297198
rect 443876 290198 443918 290434
rect 444154 290198 444196 290434
rect 443876 283434 444196 290198
rect 443876 283198 443918 283434
rect 444154 283198 444196 283434
rect 443876 276434 444196 283198
rect 443876 276198 443918 276434
rect 444154 276198 444196 276434
rect 443876 269434 444196 276198
rect 443876 269198 443918 269434
rect 444154 269198 444196 269434
rect 443876 262434 444196 269198
rect 443876 262198 443918 262434
rect 444154 262198 444196 262434
rect 443876 255434 444196 262198
rect 443876 255198 443918 255434
rect 444154 255198 444196 255434
rect 443876 248434 444196 255198
rect 443876 248198 443918 248434
rect 444154 248198 444196 248434
rect 443876 241434 444196 248198
rect 443876 241198 443918 241434
rect 444154 241198 444196 241434
rect 443876 234434 444196 241198
rect 443876 234198 443918 234434
rect 444154 234198 444196 234434
rect 443876 227434 444196 234198
rect 443876 227198 443918 227434
rect 444154 227198 444196 227434
rect 443876 220434 444196 227198
rect 443876 220198 443918 220434
rect 444154 220198 444196 220434
rect 443876 213434 444196 220198
rect 443876 213198 443918 213434
rect 444154 213198 444196 213434
rect 443876 206434 444196 213198
rect 443876 206198 443918 206434
rect 444154 206198 444196 206434
rect 443876 199434 444196 206198
rect 443876 199198 443918 199434
rect 444154 199198 444196 199434
rect 443876 192434 444196 199198
rect 443876 192198 443918 192434
rect 444154 192198 444196 192434
rect 443876 185434 444196 192198
rect 443876 185198 443918 185434
rect 444154 185198 444196 185434
rect 443876 178434 444196 185198
rect 443876 178198 443918 178434
rect 444154 178198 444196 178434
rect 443876 171434 444196 178198
rect 443876 171198 443918 171434
rect 444154 171198 444196 171434
rect 443876 164434 444196 171198
rect 443876 164198 443918 164434
rect 444154 164198 444196 164434
rect 443876 157434 444196 164198
rect 443876 157198 443918 157434
rect 444154 157198 444196 157434
rect 443876 150434 444196 157198
rect 443876 150198 443918 150434
rect 444154 150198 444196 150434
rect 443876 143434 444196 150198
rect 443876 143198 443918 143434
rect 444154 143198 444196 143434
rect 443876 136434 444196 143198
rect 443876 136198 443918 136434
rect 444154 136198 444196 136434
rect 443876 129434 444196 136198
rect 443876 129198 443918 129434
rect 444154 129198 444196 129434
rect 443876 122434 444196 129198
rect 443876 122198 443918 122434
rect 444154 122198 444196 122434
rect 443876 115434 444196 122198
rect 443876 115198 443918 115434
rect 444154 115198 444196 115434
rect 443876 108434 444196 115198
rect 443876 108198 443918 108434
rect 444154 108198 444196 108434
rect 443876 101434 444196 108198
rect 443876 101198 443918 101434
rect 444154 101198 444196 101434
rect 443876 94434 444196 101198
rect 443876 94198 443918 94434
rect 444154 94198 444196 94434
rect 443876 87434 444196 94198
rect 443876 87198 443918 87434
rect 444154 87198 444196 87434
rect 443876 80434 444196 87198
rect 443876 80198 443918 80434
rect 444154 80198 444196 80434
rect 443876 73434 444196 80198
rect 443876 73198 443918 73434
rect 444154 73198 444196 73434
rect 443876 66434 444196 73198
rect 443876 66198 443918 66434
rect 444154 66198 444196 66434
rect 443876 59434 444196 66198
rect 443876 59198 443918 59434
rect 444154 59198 444196 59434
rect 443876 52434 444196 59198
rect 443876 52198 443918 52434
rect 444154 52198 444196 52434
rect 443876 45434 444196 52198
rect 443876 45198 443918 45434
rect 444154 45198 444196 45434
rect 443876 38434 444196 45198
rect 443876 38198 443918 38434
rect 444154 38198 444196 38434
rect 443876 31434 444196 38198
rect 443876 31198 443918 31434
rect 444154 31198 444196 31434
rect 443876 24434 444196 31198
rect 443876 24198 443918 24434
rect 444154 24198 444196 24434
rect 443876 17434 444196 24198
rect 443876 17198 443918 17434
rect 444154 17198 444196 17434
rect 443876 10434 444196 17198
rect 443876 10198 443918 10434
rect 444154 10198 444196 10434
rect 443876 3434 444196 10198
rect 443876 3198 443918 3434
rect 444154 3198 444196 3434
rect 443876 -1706 444196 3198
rect 443876 -1942 443918 -1706
rect 444154 -1942 444196 -1706
rect 443876 -2026 444196 -1942
rect 443876 -2262 443918 -2026
rect 444154 -2262 444196 -2026
rect 443876 -2294 444196 -2262
rect 449144 705238 449464 706230
rect 449144 705002 449186 705238
rect 449422 705002 449464 705238
rect 449144 704918 449464 705002
rect 449144 704682 449186 704918
rect 449422 704682 449464 704918
rect 449144 695494 449464 704682
rect 449144 695258 449186 695494
rect 449422 695258 449464 695494
rect 449144 688494 449464 695258
rect 449144 688258 449186 688494
rect 449422 688258 449464 688494
rect 449144 681494 449464 688258
rect 449144 681258 449186 681494
rect 449422 681258 449464 681494
rect 449144 674494 449464 681258
rect 449144 674258 449186 674494
rect 449422 674258 449464 674494
rect 449144 667494 449464 674258
rect 449144 667258 449186 667494
rect 449422 667258 449464 667494
rect 449144 660494 449464 667258
rect 449144 660258 449186 660494
rect 449422 660258 449464 660494
rect 449144 653494 449464 660258
rect 449144 653258 449186 653494
rect 449422 653258 449464 653494
rect 449144 646494 449464 653258
rect 449144 646258 449186 646494
rect 449422 646258 449464 646494
rect 449144 639494 449464 646258
rect 449144 639258 449186 639494
rect 449422 639258 449464 639494
rect 449144 632494 449464 639258
rect 449144 632258 449186 632494
rect 449422 632258 449464 632494
rect 449144 625494 449464 632258
rect 449144 625258 449186 625494
rect 449422 625258 449464 625494
rect 449144 618494 449464 625258
rect 449144 618258 449186 618494
rect 449422 618258 449464 618494
rect 449144 611494 449464 618258
rect 449144 611258 449186 611494
rect 449422 611258 449464 611494
rect 449144 604494 449464 611258
rect 449144 604258 449186 604494
rect 449422 604258 449464 604494
rect 449144 597494 449464 604258
rect 449144 597258 449186 597494
rect 449422 597258 449464 597494
rect 449144 590494 449464 597258
rect 449144 590258 449186 590494
rect 449422 590258 449464 590494
rect 449144 583494 449464 590258
rect 449144 583258 449186 583494
rect 449422 583258 449464 583494
rect 449144 576494 449464 583258
rect 449144 576258 449186 576494
rect 449422 576258 449464 576494
rect 449144 569494 449464 576258
rect 449144 569258 449186 569494
rect 449422 569258 449464 569494
rect 449144 562494 449464 569258
rect 449144 562258 449186 562494
rect 449422 562258 449464 562494
rect 449144 555494 449464 562258
rect 449144 555258 449186 555494
rect 449422 555258 449464 555494
rect 449144 548494 449464 555258
rect 449144 548258 449186 548494
rect 449422 548258 449464 548494
rect 449144 541494 449464 548258
rect 449144 541258 449186 541494
rect 449422 541258 449464 541494
rect 449144 534494 449464 541258
rect 449144 534258 449186 534494
rect 449422 534258 449464 534494
rect 449144 527494 449464 534258
rect 449144 527258 449186 527494
rect 449422 527258 449464 527494
rect 449144 520494 449464 527258
rect 449144 520258 449186 520494
rect 449422 520258 449464 520494
rect 449144 513494 449464 520258
rect 449144 513258 449186 513494
rect 449422 513258 449464 513494
rect 449144 506494 449464 513258
rect 449144 506258 449186 506494
rect 449422 506258 449464 506494
rect 449144 499494 449464 506258
rect 449144 499258 449186 499494
rect 449422 499258 449464 499494
rect 449144 492494 449464 499258
rect 449144 492258 449186 492494
rect 449422 492258 449464 492494
rect 449144 485494 449464 492258
rect 449144 485258 449186 485494
rect 449422 485258 449464 485494
rect 449144 478494 449464 485258
rect 449144 478258 449186 478494
rect 449422 478258 449464 478494
rect 449144 471494 449464 478258
rect 449144 471258 449186 471494
rect 449422 471258 449464 471494
rect 449144 464494 449464 471258
rect 449144 464258 449186 464494
rect 449422 464258 449464 464494
rect 449144 457494 449464 464258
rect 449144 457258 449186 457494
rect 449422 457258 449464 457494
rect 449144 450494 449464 457258
rect 449144 450258 449186 450494
rect 449422 450258 449464 450494
rect 449144 443494 449464 450258
rect 449144 443258 449186 443494
rect 449422 443258 449464 443494
rect 449144 436494 449464 443258
rect 449144 436258 449186 436494
rect 449422 436258 449464 436494
rect 449144 429494 449464 436258
rect 449144 429258 449186 429494
rect 449422 429258 449464 429494
rect 449144 422494 449464 429258
rect 449144 422258 449186 422494
rect 449422 422258 449464 422494
rect 449144 415494 449464 422258
rect 449144 415258 449186 415494
rect 449422 415258 449464 415494
rect 449144 408494 449464 415258
rect 449144 408258 449186 408494
rect 449422 408258 449464 408494
rect 449144 401494 449464 408258
rect 449144 401258 449186 401494
rect 449422 401258 449464 401494
rect 449144 394494 449464 401258
rect 449144 394258 449186 394494
rect 449422 394258 449464 394494
rect 449144 387494 449464 394258
rect 449144 387258 449186 387494
rect 449422 387258 449464 387494
rect 449144 380494 449464 387258
rect 449144 380258 449186 380494
rect 449422 380258 449464 380494
rect 449144 373494 449464 380258
rect 449144 373258 449186 373494
rect 449422 373258 449464 373494
rect 449144 366494 449464 373258
rect 449144 366258 449186 366494
rect 449422 366258 449464 366494
rect 449144 359494 449464 366258
rect 449144 359258 449186 359494
rect 449422 359258 449464 359494
rect 449144 352494 449464 359258
rect 449144 352258 449186 352494
rect 449422 352258 449464 352494
rect 449144 345494 449464 352258
rect 449144 345258 449186 345494
rect 449422 345258 449464 345494
rect 449144 338494 449464 345258
rect 449144 338258 449186 338494
rect 449422 338258 449464 338494
rect 449144 331494 449464 338258
rect 449144 331258 449186 331494
rect 449422 331258 449464 331494
rect 449144 324494 449464 331258
rect 449144 324258 449186 324494
rect 449422 324258 449464 324494
rect 449144 317494 449464 324258
rect 449144 317258 449186 317494
rect 449422 317258 449464 317494
rect 449144 310494 449464 317258
rect 449144 310258 449186 310494
rect 449422 310258 449464 310494
rect 449144 303494 449464 310258
rect 449144 303258 449186 303494
rect 449422 303258 449464 303494
rect 449144 296494 449464 303258
rect 449144 296258 449186 296494
rect 449422 296258 449464 296494
rect 449144 289494 449464 296258
rect 449144 289258 449186 289494
rect 449422 289258 449464 289494
rect 449144 282494 449464 289258
rect 449144 282258 449186 282494
rect 449422 282258 449464 282494
rect 449144 275494 449464 282258
rect 449144 275258 449186 275494
rect 449422 275258 449464 275494
rect 449144 268494 449464 275258
rect 449144 268258 449186 268494
rect 449422 268258 449464 268494
rect 449144 261494 449464 268258
rect 449144 261258 449186 261494
rect 449422 261258 449464 261494
rect 449144 254494 449464 261258
rect 449144 254258 449186 254494
rect 449422 254258 449464 254494
rect 449144 247494 449464 254258
rect 449144 247258 449186 247494
rect 449422 247258 449464 247494
rect 449144 240494 449464 247258
rect 449144 240258 449186 240494
rect 449422 240258 449464 240494
rect 449144 233494 449464 240258
rect 449144 233258 449186 233494
rect 449422 233258 449464 233494
rect 449144 226494 449464 233258
rect 449144 226258 449186 226494
rect 449422 226258 449464 226494
rect 449144 219494 449464 226258
rect 449144 219258 449186 219494
rect 449422 219258 449464 219494
rect 449144 212494 449464 219258
rect 449144 212258 449186 212494
rect 449422 212258 449464 212494
rect 449144 205494 449464 212258
rect 449144 205258 449186 205494
rect 449422 205258 449464 205494
rect 449144 198494 449464 205258
rect 449144 198258 449186 198494
rect 449422 198258 449464 198494
rect 449144 191494 449464 198258
rect 449144 191258 449186 191494
rect 449422 191258 449464 191494
rect 449144 184494 449464 191258
rect 449144 184258 449186 184494
rect 449422 184258 449464 184494
rect 449144 177494 449464 184258
rect 449144 177258 449186 177494
rect 449422 177258 449464 177494
rect 449144 170494 449464 177258
rect 449144 170258 449186 170494
rect 449422 170258 449464 170494
rect 449144 163494 449464 170258
rect 449144 163258 449186 163494
rect 449422 163258 449464 163494
rect 449144 156494 449464 163258
rect 449144 156258 449186 156494
rect 449422 156258 449464 156494
rect 449144 149494 449464 156258
rect 449144 149258 449186 149494
rect 449422 149258 449464 149494
rect 449144 142494 449464 149258
rect 449144 142258 449186 142494
rect 449422 142258 449464 142494
rect 449144 135494 449464 142258
rect 449144 135258 449186 135494
rect 449422 135258 449464 135494
rect 449144 128494 449464 135258
rect 449144 128258 449186 128494
rect 449422 128258 449464 128494
rect 449144 121494 449464 128258
rect 449144 121258 449186 121494
rect 449422 121258 449464 121494
rect 449144 114494 449464 121258
rect 449144 114258 449186 114494
rect 449422 114258 449464 114494
rect 449144 107494 449464 114258
rect 449144 107258 449186 107494
rect 449422 107258 449464 107494
rect 449144 100494 449464 107258
rect 449144 100258 449186 100494
rect 449422 100258 449464 100494
rect 449144 93494 449464 100258
rect 449144 93258 449186 93494
rect 449422 93258 449464 93494
rect 449144 86494 449464 93258
rect 449144 86258 449186 86494
rect 449422 86258 449464 86494
rect 449144 79494 449464 86258
rect 449144 79258 449186 79494
rect 449422 79258 449464 79494
rect 449144 72494 449464 79258
rect 449144 72258 449186 72494
rect 449422 72258 449464 72494
rect 449144 65494 449464 72258
rect 449144 65258 449186 65494
rect 449422 65258 449464 65494
rect 449144 58494 449464 65258
rect 449144 58258 449186 58494
rect 449422 58258 449464 58494
rect 449144 51494 449464 58258
rect 449144 51258 449186 51494
rect 449422 51258 449464 51494
rect 449144 44494 449464 51258
rect 449144 44258 449186 44494
rect 449422 44258 449464 44494
rect 449144 37494 449464 44258
rect 449144 37258 449186 37494
rect 449422 37258 449464 37494
rect 449144 30494 449464 37258
rect 449144 30258 449186 30494
rect 449422 30258 449464 30494
rect 449144 23494 449464 30258
rect 449144 23258 449186 23494
rect 449422 23258 449464 23494
rect 449144 16494 449464 23258
rect 449144 16258 449186 16494
rect 449422 16258 449464 16494
rect 449144 9494 449464 16258
rect 449144 9258 449186 9494
rect 449422 9258 449464 9494
rect 449144 2494 449464 9258
rect 449144 2258 449186 2494
rect 449422 2258 449464 2494
rect 449144 -746 449464 2258
rect 449144 -982 449186 -746
rect 449422 -982 449464 -746
rect 449144 -1066 449464 -982
rect 449144 -1302 449186 -1066
rect 449422 -1302 449464 -1066
rect 449144 -2294 449464 -1302
rect 450876 706198 451196 706230
rect 450876 705962 450918 706198
rect 451154 705962 451196 706198
rect 450876 705878 451196 705962
rect 450876 705642 450918 705878
rect 451154 705642 451196 705878
rect 450876 696434 451196 705642
rect 450876 696198 450918 696434
rect 451154 696198 451196 696434
rect 450876 689434 451196 696198
rect 450876 689198 450918 689434
rect 451154 689198 451196 689434
rect 450876 682434 451196 689198
rect 450876 682198 450918 682434
rect 451154 682198 451196 682434
rect 450876 675434 451196 682198
rect 450876 675198 450918 675434
rect 451154 675198 451196 675434
rect 450876 668434 451196 675198
rect 450876 668198 450918 668434
rect 451154 668198 451196 668434
rect 450876 661434 451196 668198
rect 450876 661198 450918 661434
rect 451154 661198 451196 661434
rect 450876 654434 451196 661198
rect 450876 654198 450918 654434
rect 451154 654198 451196 654434
rect 450876 647434 451196 654198
rect 450876 647198 450918 647434
rect 451154 647198 451196 647434
rect 450876 640434 451196 647198
rect 450876 640198 450918 640434
rect 451154 640198 451196 640434
rect 450876 633434 451196 640198
rect 450876 633198 450918 633434
rect 451154 633198 451196 633434
rect 450876 626434 451196 633198
rect 450876 626198 450918 626434
rect 451154 626198 451196 626434
rect 450876 619434 451196 626198
rect 450876 619198 450918 619434
rect 451154 619198 451196 619434
rect 450876 612434 451196 619198
rect 450876 612198 450918 612434
rect 451154 612198 451196 612434
rect 450876 605434 451196 612198
rect 450876 605198 450918 605434
rect 451154 605198 451196 605434
rect 450876 598434 451196 605198
rect 450876 598198 450918 598434
rect 451154 598198 451196 598434
rect 450876 591434 451196 598198
rect 450876 591198 450918 591434
rect 451154 591198 451196 591434
rect 450876 584434 451196 591198
rect 450876 584198 450918 584434
rect 451154 584198 451196 584434
rect 450876 577434 451196 584198
rect 450876 577198 450918 577434
rect 451154 577198 451196 577434
rect 450876 570434 451196 577198
rect 450876 570198 450918 570434
rect 451154 570198 451196 570434
rect 450876 563434 451196 570198
rect 450876 563198 450918 563434
rect 451154 563198 451196 563434
rect 450876 556434 451196 563198
rect 450876 556198 450918 556434
rect 451154 556198 451196 556434
rect 450876 549434 451196 556198
rect 450876 549198 450918 549434
rect 451154 549198 451196 549434
rect 450876 542434 451196 549198
rect 450876 542198 450918 542434
rect 451154 542198 451196 542434
rect 450876 535434 451196 542198
rect 450876 535198 450918 535434
rect 451154 535198 451196 535434
rect 450876 528434 451196 535198
rect 450876 528198 450918 528434
rect 451154 528198 451196 528434
rect 450876 521434 451196 528198
rect 450876 521198 450918 521434
rect 451154 521198 451196 521434
rect 450876 514434 451196 521198
rect 450876 514198 450918 514434
rect 451154 514198 451196 514434
rect 450876 507434 451196 514198
rect 450876 507198 450918 507434
rect 451154 507198 451196 507434
rect 450876 500434 451196 507198
rect 450876 500198 450918 500434
rect 451154 500198 451196 500434
rect 450876 493434 451196 500198
rect 450876 493198 450918 493434
rect 451154 493198 451196 493434
rect 450876 486434 451196 493198
rect 450876 486198 450918 486434
rect 451154 486198 451196 486434
rect 450876 479434 451196 486198
rect 450876 479198 450918 479434
rect 451154 479198 451196 479434
rect 450876 472434 451196 479198
rect 450876 472198 450918 472434
rect 451154 472198 451196 472434
rect 450876 465434 451196 472198
rect 450876 465198 450918 465434
rect 451154 465198 451196 465434
rect 450876 458434 451196 465198
rect 450876 458198 450918 458434
rect 451154 458198 451196 458434
rect 450876 451434 451196 458198
rect 450876 451198 450918 451434
rect 451154 451198 451196 451434
rect 450876 444434 451196 451198
rect 450876 444198 450918 444434
rect 451154 444198 451196 444434
rect 450876 437434 451196 444198
rect 450876 437198 450918 437434
rect 451154 437198 451196 437434
rect 450876 430434 451196 437198
rect 450876 430198 450918 430434
rect 451154 430198 451196 430434
rect 450876 423434 451196 430198
rect 450876 423198 450918 423434
rect 451154 423198 451196 423434
rect 450876 416434 451196 423198
rect 450876 416198 450918 416434
rect 451154 416198 451196 416434
rect 450876 409434 451196 416198
rect 450876 409198 450918 409434
rect 451154 409198 451196 409434
rect 450876 402434 451196 409198
rect 450876 402198 450918 402434
rect 451154 402198 451196 402434
rect 450876 395434 451196 402198
rect 450876 395198 450918 395434
rect 451154 395198 451196 395434
rect 450876 388434 451196 395198
rect 450876 388198 450918 388434
rect 451154 388198 451196 388434
rect 450876 381434 451196 388198
rect 450876 381198 450918 381434
rect 451154 381198 451196 381434
rect 450876 374434 451196 381198
rect 450876 374198 450918 374434
rect 451154 374198 451196 374434
rect 450876 367434 451196 374198
rect 450876 367198 450918 367434
rect 451154 367198 451196 367434
rect 450876 360434 451196 367198
rect 450876 360198 450918 360434
rect 451154 360198 451196 360434
rect 450876 353434 451196 360198
rect 450876 353198 450918 353434
rect 451154 353198 451196 353434
rect 450876 346434 451196 353198
rect 450876 346198 450918 346434
rect 451154 346198 451196 346434
rect 450876 339434 451196 346198
rect 450876 339198 450918 339434
rect 451154 339198 451196 339434
rect 450876 332434 451196 339198
rect 450876 332198 450918 332434
rect 451154 332198 451196 332434
rect 450876 325434 451196 332198
rect 450876 325198 450918 325434
rect 451154 325198 451196 325434
rect 450876 318434 451196 325198
rect 450876 318198 450918 318434
rect 451154 318198 451196 318434
rect 450876 311434 451196 318198
rect 450876 311198 450918 311434
rect 451154 311198 451196 311434
rect 450876 304434 451196 311198
rect 450876 304198 450918 304434
rect 451154 304198 451196 304434
rect 450876 297434 451196 304198
rect 450876 297198 450918 297434
rect 451154 297198 451196 297434
rect 450876 290434 451196 297198
rect 450876 290198 450918 290434
rect 451154 290198 451196 290434
rect 450876 283434 451196 290198
rect 450876 283198 450918 283434
rect 451154 283198 451196 283434
rect 450876 276434 451196 283198
rect 450876 276198 450918 276434
rect 451154 276198 451196 276434
rect 450876 269434 451196 276198
rect 450876 269198 450918 269434
rect 451154 269198 451196 269434
rect 450876 262434 451196 269198
rect 450876 262198 450918 262434
rect 451154 262198 451196 262434
rect 450876 255434 451196 262198
rect 450876 255198 450918 255434
rect 451154 255198 451196 255434
rect 450876 248434 451196 255198
rect 450876 248198 450918 248434
rect 451154 248198 451196 248434
rect 450876 241434 451196 248198
rect 450876 241198 450918 241434
rect 451154 241198 451196 241434
rect 450876 234434 451196 241198
rect 450876 234198 450918 234434
rect 451154 234198 451196 234434
rect 450876 227434 451196 234198
rect 450876 227198 450918 227434
rect 451154 227198 451196 227434
rect 450876 220434 451196 227198
rect 450876 220198 450918 220434
rect 451154 220198 451196 220434
rect 450876 213434 451196 220198
rect 450876 213198 450918 213434
rect 451154 213198 451196 213434
rect 450876 206434 451196 213198
rect 450876 206198 450918 206434
rect 451154 206198 451196 206434
rect 450876 199434 451196 206198
rect 450876 199198 450918 199434
rect 451154 199198 451196 199434
rect 450876 192434 451196 199198
rect 450876 192198 450918 192434
rect 451154 192198 451196 192434
rect 450876 185434 451196 192198
rect 450876 185198 450918 185434
rect 451154 185198 451196 185434
rect 450876 178434 451196 185198
rect 450876 178198 450918 178434
rect 451154 178198 451196 178434
rect 450876 171434 451196 178198
rect 450876 171198 450918 171434
rect 451154 171198 451196 171434
rect 450876 164434 451196 171198
rect 450876 164198 450918 164434
rect 451154 164198 451196 164434
rect 450876 157434 451196 164198
rect 450876 157198 450918 157434
rect 451154 157198 451196 157434
rect 450876 150434 451196 157198
rect 450876 150198 450918 150434
rect 451154 150198 451196 150434
rect 450876 143434 451196 150198
rect 450876 143198 450918 143434
rect 451154 143198 451196 143434
rect 450876 136434 451196 143198
rect 450876 136198 450918 136434
rect 451154 136198 451196 136434
rect 450876 129434 451196 136198
rect 450876 129198 450918 129434
rect 451154 129198 451196 129434
rect 450876 122434 451196 129198
rect 450876 122198 450918 122434
rect 451154 122198 451196 122434
rect 450876 115434 451196 122198
rect 450876 115198 450918 115434
rect 451154 115198 451196 115434
rect 450876 108434 451196 115198
rect 450876 108198 450918 108434
rect 451154 108198 451196 108434
rect 450876 101434 451196 108198
rect 450876 101198 450918 101434
rect 451154 101198 451196 101434
rect 450876 94434 451196 101198
rect 450876 94198 450918 94434
rect 451154 94198 451196 94434
rect 450876 87434 451196 94198
rect 450876 87198 450918 87434
rect 451154 87198 451196 87434
rect 450876 80434 451196 87198
rect 450876 80198 450918 80434
rect 451154 80198 451196 80434
rect 450876 73434 451196 80198
rect 450876 73198 450918 73434
rect 451154 73198 451196 73434
rect 450876 66434 451196 73198
rect 450876 66198 450918 66434
rect 451154 66198 451196 66434
rect 450876 59434 451196 66198
rect 450876 59198 450918 59434
rect 451154 59198 451196 59434
rect 450876 52434 451196 59198
rect 450876 52198 450918 52434
rect 451154 52198 451196 52434
rect 450876 45434 451196 52198
rect 450876 45198 450918 45434
rect 451154 45198 451196 45434
rect 450876 38434 451196 45198
rect 450876 38198 450918 38434
rect 451154 38198 451196 38434
rect 450876 31434 451196 38198
rect 450876 31198 450918 31434
rect 451154 31198 451196 31434
rect 450876 24434 451196 31198
rect 450876 24198 450918 24434
rect 451154 24198 451196 24434
rect 450876 17434 451196 24198
rect 450876 17198 450918 17434
rect 451154 17198 451196 17434
rect 450876 10434 451196 17198
rect 450876 10198 450918 10434
rect 451154 10198 451196 10434
rect 450876 3434 451196 10198
rect 450876 3198 450918 3434
rect 451154 3198 451196 3434
rect 450876 -1706 451196 3198
rect 450876 -1942 450918 -1706
rect 451154 -1942 451196 -1706
rect 450876 -2026 451196 -1942
rect 450876 -2262 450918 -2026
rect 451154 -2262 451196 -2026
rect 450876 -2294 451196 -2262
rect 456144 705238 456464 706230
rect 456144 705002 456186 705238
rect 456422 705002 456464 705238
rect 456144 704918 456464 705002
rect 456144 704682 456186 704918
rect 456422 704682 456464 704918
rect 456144 695494 456464 704682
rect 456144 695258 456186 695494
rect 456422 695258 456464 695494
rect 456144 688494 456464 695258
rect 456144 688258 456186 688494
rect 456422 688258 456464 688494
rect 456144 681494 456464 688258
rect 456144 681258 456186 681494
rect 456422 681258 456464 681494
rect 456144 674494 456464 681258
rect 456144 674258 456186 674494
rect 456422 674258 456464 674494
rect 456144 667494 456464 674258
rect 456144 667258 456186 667494
rect 456422 667258 456464 667494
rect 456144 660494 456464 667258
rect 456144 660258 456186 660494
rect 456422 660258 456464 660494
rect 456144 653494 456464 660258
rect 456144 653258 456186 653494
rect 456422 653258 456464 653494
rect 456144 646494 456464 653258
rect 456144 646258 456186 646494
rect 456422 646258 456464 646494
rect 456144 639494 456464 646258
rect 456144 639258 456186 639494
rect 456422 639258 456464 639494
rect 456144 632494 456464 639258
rect 456144 632258 456186 632494
rect 456422 632258 456464 632494
rect 456144 625494 456464 632258
rect 456144 625258 456186 625494
rect 456422 625258 456464 625494
rect 456144 618494 456464 625258
rect 456144 618258 456186 618494
rect 456422 618258 456464 618494
rect 456144 611494 456464 618258
rect 456144 611258 456186 611494
rect 456422 611258 456464 611494
rect 456144 604494 456464 611258
rect 456144 604258 456186 604494
rect 456422 604258 456464 604494
rect 456144 597494 456464 604258
rect 456144 597258 456186 597494
rect 456422 597258 456464 597494
rect 456144 590494 456464 597258
rect 456144 590258 456186 590494
rect 456422 590258 456464 590494
rect 456144 583494 456464 590258
rect 456144 583258 456186 583494
rect 456422 583258 456464 583494
rect 456144 576494 456464 583258
rect 456144 576258 456186 576494
rect 456422 576258 456464 576494
rect 456144 569494 456464 576258
rect 456144 569258 456186 569494
rect 456422 569258 456464 569494
rect 456144 562494 456464 569258
rect 456144 562258 456186 562494
rect 456422 562258 456464 562494
rect 456144 555494 456464 562258
rect 456144 555258 456186 555494
rect 456422 555258 456464 555494
rect 456144 548494 456464 555258
rect 456144 548258 456186 548494
rect 456422 548258 456464 548494
rect 456144 541494 456464 548258
rect 456144 541258 456186 541494
rect 456422 541258 456464 541494
rect 456144 534494 456464 541258
rect 456144 534258 456186 534494
rect 456422 534258 456464 534494
rect 456144 527494 456464 534258
rect 456144 527258 456186 527494
rect 456422 527258 456464 527494
rect 456144 520494 456464 527258
rect 456144 520258 456186 520494
rect 456422 520258 456464 520494
rect 456144 513494 456464 520258
rect 456144 513258 456186 513494
rect 456422 513258 456464 513494
rect 456144 506494 456464 513258
rect 456144 506258 456186 506494
rect 456422 506258 456464 506494
rect 456144 499494 456464 506258
rect 456144 499258 456186 499494
rect 456422 499258 456464 499494
rect 456144 492494 456464 499258
rect 456144 492258 456186 492494
rect 456422 492258 456464 492494
rect 456144 485494 456464 492258
rect 456144 485258 456186 485494
rect 456422 485258 456464 485494
rect 456144 478494 456464 485258
rect 456144 478258 456186 478494
rect 456422 478258 456464 478494
rect 456144 471494 456464 478258
rect 456144 471258 456186 471494
rect 456422 471258 456464 471494
rect 456144 464494 456464 471258
rect 456144 464258 456186 464494
rect 456422 464258 456464 464494
rect 456144 457494 456464 464258
rect 456144 457258 456186 457494
rect 456422 457258 456464 457494
rect 456144 450494 456464 457258
rect 456144 450258 456186 450494
rect 456422 450258 456464 450494
rect 456144 443494 456464 450258
rect 456144 443258 456186 443494
rect 456422 443258 456464 443494
rect 456144 436494 456464 443258
rect 456144 436258 456186 436494
rect 456422 436258 456464 436494
rect 456144 429494 456464 436258
rect 456144 429258 456186 429494
rect 456422 429258 456464 429494
rect 456144 422494 456464 429258
rect 456144 422258 456186 422494
rect 456422 422258 456464 422494
rect 456144 415494 456464 422258
rect 456144 415258 456186 415494
rect 456422 415258 456464 415494
rect 456144 408494 456464 415258
rect 456144 408258 456186 408494
rect 456422 408258 456464 408494
rect 456144 401494 456464 408258
rect 456144 401258 456186 401494
rect 456422 401258 456464 401494
rect 456144 394494 456464 401258
rect 456144 394258 456186 394494
rect 456422 394258 456464 394494
rect 456144 387494 456464 394258
rect 456144 387258 456186 387494
rect 456422 387258 456464 387494
rect 456144 380494 456464 387258
rect 456144 380258 456186 380494
rect 456422 380258 456464 380494
rect 456144 373494 456464 380258
rect 456144 373258 456186 373494
rect 456422 373258 456464 373494
rect 456144 366494 456464 373258
rect 456144 366258 456186 366494
rect 456422 366258 456464 366494
rect 456144 359494 456464 366258
rect 456144 359258 456186 359494
rect 456422 359258 456464 359494
rect 456144 352494 456464 359258
rect 456144 352258 456186 352494
rect 456422 352258 456464 352494
rect 456144 345494 456464 352258
rect 456144 345258 456186 345494
rect 456422 345258 456464 345494
rect 456144 338494 456464 345258
rect 456144 338258 456186 338494
rect 456422 338258 456464 338494
rect 456144 331494 456464 338258
rect 456144 331258 456186 331494
rect 456422 331258 456464 331494
rect 456144 324494 456464 331258
rect 456144 324258 456186 324494
rect 456422 324258 456464 324494
rect 456144 317494 456464 324258
rect 456144 317258 456186 317494
rect 456422 317258 456464 317494
rect 456144 310494 456464 317258
rect 456144 310258 456186 310494
rect 456422 310258 456464 310494
rect 456144 303494 456464 310258
rect 456144 303258 456186 303494
rect 456422 303258 456464 303494
rect 456144 296494 456464 303258
rect 456144 296258 456186 296494
rect 456422 296258 456464 296494
rect 456144 289494 456464 296258
rect 456144 289258 456186 289494
rect 456422 289258 456464 289494
rect 456144 282494 456464 289258
rect 456144 282258 456186 282494
rect 456422 282258 456464 282494
rect 456144 275494 456464 282258
rect 456144 275258 456186 275494
rect 456422 275258 456464 275494
rect 456144 268494 456464 275258
rect 456144 268258 456186 268494
rect 456422 268258 456464 268494
rect 456144 261494 456464 268258
rect 456144 261258 456186 261494
rect 456422 261258 456464 261494
rect 456144 254494 456464 261258
rect 456144 254258 456186 254494
rect 456422 254258 456464 254494
rect 456144 247494 456464 254258
rect 456144 247258 456186 247494
rect 456422 247258 456464 247494
rect 456144 240494 456464 247258
rect 456144 240258 456186 240494
rect 456422 240258 456464 240494
rect 456144 233494 456464 240258
rect 456144 233258 456186 233494
rect 456422 233258 456464 233494
rect 456144 226494 456464 233258
rect 456144 226258 456186 226494
rect 456422 226258 456464 226494
rect 456144 219494 456464 226258
rect 456144 219258 456186 219494
rect 456422 219258 456464 219494
rect 456144 212494 456464 219258
rect 456144 212258 456186 212494
rect 456422 212258 456464 212494
rect 456144 205494 456464 212258
rect 456144 205258 456186 205494
rect 456422 205258 456464 205494
rect 456144 198494 456464 205258
rect 456144 198258 456186 198494
rect 456422 198258 456464 198494
rect 456144 191494 456464 198258
rect 456144 191258 456186 191494
rect 456422 191258 456464 191494
rect 456144 184494 456464 191258
rect 456144 184258 456186 184494
rect 456422 184258 456464 184494
rect 456144 177494 456464 184258
rect 456144 177258 456186 177494
rect 456422 177258 456464 177494
rect 456144 170494 456464 177258
rect 456144 170258 456186 170494
rect 456422 170258 456464 170494
rect 456144 163494 456464 170258
rect 456144 163258 456186 163494
rect 456422 163258 456464 163494
rect 456144 156494 456464 163258
rect 456144 156258 456186 156494
rect 456422 156258 456464 156494
rect 456144 149494 456464 156258
rect 456144 149258 456186 149494
rect 456422 149258 456464 149494
rect 456144 142494 456464 149258
rect 456144 142258 456186 142494
rect 456422 142258 456464 142494
rect 456144 135494 456464 142258
rect 456144 135258 456186 135494
rect 456422 135258 456464 135494
rect 456144 128494 456464 135258
rect 456144 128258 456186 128494
rect 456422 128258 456464 128494
rect 456144 121494 456464 128258
rect 456144 121258 456186 121494
rect 456422 121258 456464 121494
rect 456144 114494 456464 121258
rect 456144 114258 456186 114494
rect 456422 114258 456464 114494
rect 456144 107494 456464 114258
rect 456144 107258 456186 107494
rect 456422 107258 456464 107494
rect 456144 100494 456464 107258
rect 456144 100258 456186 100494
rect 456422 100258 456464 100494
rect 456144 93494 456464 100258
rect 456144 93258 456186 93494
rect 456422 93258 456464 93494
rect 456144 86494 456464 93258
rect 456144 86258 456186 86494
rect 456422 86258 456464 86494
rect 456144 79494 456464 86258
rect 456144 79258 456186 79494
rect 456422 79258 456464 79494
rect 456144 72494 456464 79258
rect 456144 72258 456186 72494
rect 456422 72258 456464 72494
rect 456144 65494 456464 72258
rect 456144 65258 456186 65494
rect 456422 65258 456464 65494
rect 456144 58494 456464 65258
rect 456144 58258 456186 58494
rect 456422 58258 456464 58494
rect 456144 51494 456464 58258
rect 456144 51258 456186 51494
rect 456422 51258 456464 51494
rect 456144 44494 456464 51258
rect 456144 44258 456186 44494
rect 456422 44258 456464 44494
rect 456144 37494 456464 44258
rect 456144 37258 456186 37494
rect 456422 37258 456464 37494
rect 456144 30494 456464 37258
rect 456144 30258 456186 30494
rect 456422 30258 456464 30494
rect 456144 23494 456464 30258
rect 456144 23258 456186 23494
rect 456422 23258 456464 23494
rect 456144 16494 456464 23258
rect 456144 16258 456186 16494
rect 456422 16258 456464 16494
rect 456144 9494 456464 16258
rect 456144 9258 456186 9494
rect 456422 9258 456464 9494
rect 456144 2494 456464 9258
rect 456144 2258 456186 2494
rect 456422 2258 456464 2494
rect 456144 -746 456464 2258
rect 456144 -982 456186 -746
rect 456422 -982 456464 -746
rect 456144 -1066 456464 -982
rect 456144 -1302 456186 -1066
rect 456422 -1302 456464 -1066
rect 456144 -2294 456464 -1302
rect 457876 706198 458196 706230
rect 457876 705962 457918 706198
rect 458154 705962 458196 706198
rect 457876 705878 458196 705962
rect 457876 705642 457918 705878
rect 458154 705642 458196 705878
rect 457876 696434 458196 705642
rect 457876 696198 457918 696434
rect 458154 696198 458196 696434
rect 457876 689434 458196 696198
rect 457876 689198 457918 689434
rect 458154 689198 458196 689434
rect 457876 682434 458196 689198
rect 457876 682198 457918 682434
rect 458154 682198 458196 682434
rect 457876 675434 458196 682198
rect 457876 675198 457918 675434
rect 458154 675198 458196 675434
rect 457876 668434 458196 675198
rect 457876 668198 457918 668434
rect 458154 668198 458196 668434
rect 457876 661434 458196 668198
rect 457876 661198 457918 661434
rect 458154 661198 458196 661434
rect 457876 654434 458196 661198
rect 457876 654198 457918 654434
rect 458154 654198 458196 654434
rect 457876 647434 458196 654198
rect 457876 647198 457918 647434
rect 458154 647198 458196 647434
rect 457876 640434 458196 647198
rect 457876 640198 457918 640434
rect 458154 640198 458196 640434
rect 457876 633434 458196 640198
rect 457876 633198 457918 633434
rect 458154 633198 458196 633434
rect 457876 626434 458196 633198
rect 457876 626198 457918 626434
rect 458154 626198 458196 626434
rect 457876 619434 458196 626198
rect 457876 619198 457918 619434
rect 458154 619198 458196 619434
rect 457876 612434 458196 619198
rect 457876 612198 457918 612434
rect 458154 612198 458196 612434
rect 457876 605434 458196 612198
rect 457876 605198 457918 605434
rect 458154 605198 458196 605434
rect 457876 598434 458196 605198
rect 457876 598198 457918 598434
rect 458154 598198 458196 598434
rect 457876 591434 458196 598198
rect 457876 591198 457918 591434
rect 458154 591198 458196 591434
rect 457876 584434 458196 591198
rect 457876 584198 457918 584434
rect 458154 584198 458196 584434
rect 457876 577434 458196 584198
rect 457876 577198 457918 577434
rect 458154 577198 458196 577434
rect 457876 570434 458196 577198
rect 457876 570198 457918 570434
rect 458154 570198 458196 570434
rect 457876 563434 458196 570198
rect 457876 563198 457918 563434
rect 458154 563198 458196 563434
rect 457876 556434 458196 563198
rect 457876 556198 457918 556434
rect 458154 556198 458196 556434
rect 457876 549434 458196 556198
rect 457876 549198 457918 549434
rect 458154 549198 458196 549434
rect 457876 542434 458196 549198
rect 457876 542198 457918 542434
rect 458154 542198 458196 542434
rect 457876 535434 458196 542198
rect 457876 535198 457918 535434
rect 458154 535198 458196 535434
rect 457876 528434 458196 535198
rect 457876 528198 457918 528434
rect 458154 528198 458196 528434
rect 457876 521434 458196 528198
rect 457876 521198 457918 521434
rect 458154 521198 458196 521434
rect 457876 514434 458196 521198
rect 457876 514198 457918 514434
rect 458154 514198 458196 514434
rect 457876 507434 458196 514198
rect 457876 507198 457918 507434
rect 458154 507198 458196 507434
rect 457876 500434 458196 507198
rect 457876 500198 457918 500434
rect 458154 500198 458196 500434
rect 457876 493434 458196 500198
rect 457876 493198 457918 493434
rect 458154 493198 458196 493434
rect 457876 486434 458196 493198
rect 457876 486198 457918 486434
rect 458154 486198 458196 486434
rect 457876 479434 458196 486198
rect 457876 479198 457918 479434
rect 458154 479198 458196 479434
rect 457876 472434 458196 479198
rect 457876 472198 457918 472434
rect 458154 472198 458196 472434
rect 457876 465434 458196 472198
rect 457876 465198 457918 465434
rect 458154 465198 458196 465434
rect 457876 458434 458196 465198
rect 457876 458198 457918 458434
rect 458154 458198 458196 458434
rect 457876 451434 458196 458198
rect 457876 451198 457918 451434
rect 458154 451198 458196 451434
rect 457876 444434 458196 451198
rect 457876 444198 457918 444434
rect 458154 444198 458196 444434
rect 457876 437434 458196 444198
rect 457876 437198 457918 437434
rect 458154 437198 458196 437434
rect 457876 430434 458196 437198
rect 457876 430198 457918 430434
rect 458154 430198 458196 430434
rect 457876 423434 458196 430198
rect 457876 423198 457918 423434
rect 458154 423198 458196 423434
rect 457876 416434 458196 423198
rect 457876 416198 457918 416434
rect 458154 416198 458196 416434
rect 457876 409434 458196 416198
rect 457876 409198 457918 409434
rect 458154 409198 458196 409434
rect 457876 402434 458196 409198
rect 457876 402198 457918 402434
rect 458154 402198 458196 402434
rect 457876 395434 458196 402198
rect 457876 395198 457918 395434
rect 458154 395198 458196 395434
rect 457876 388434 458196 395198
rect 457876 388198 457918 388434
rect 458154 388198 458196 388434
rect 457876 381434 458196 388198
rect 457876 381198 457918 381434
rect 458154 381198 458196 381434
rect 457876 374434 458196 381198
rect 457876 374198 457918 374434
rect 458154 374198 458196 374434
rect 457876 367434 458196 374198
rect 457876 367198 457918 367434
rect 458154 367198 458196 367434
rect 457876 360434 458196 367198
rect 457876 360198 457918 360434
rect 458154 360198 458196 360434
rect 457876 353434 458196 360198
rect 457876 353198 457918 353434
rect 458154 353198 458196 353434
rect 457876 346434 458196 353198
rect 457876 346198 457918 346434
rect 458154 346198 458196 346434
rect 457876 339434 458196 346198
rect 457876 339198 457918 339434
rect 458154 339198 458196 339434
rect 457876 332434 458196 339198
rect 457876 332198 457918 332434
rect 458154 332198 458196 332434
rect 457876 325434 458196 332198
rect 457876 325198 457918 325434
rect 458154 325198 458196 325434
rect 457876 318434 458196 325198
rect 457876 318198 457918 318434
rect 458154 318198 458196 318434
rect 457876 311434 458196 318198
rect 457876 311198 457918 311434
rect 458154 311198 458196 311434
rect 457876 304434 458196 311198
rect 457876 304198 457918 304434
rect 458154 304198 458196 304434
rect 457876 297434 458196 304198
rect 457876 297198 457918 297434
rect 458154 297198 458196 297434
rect 457876 290434 458196 297198
rect 457876 290198 457918 290434
rect 458154 290198 458196 290434
rect 457876 283434 458196 290198
rect 457876 283198 457918 283434
rect 458154 283198 458196 283434
rect 457876 276434 458196 283198
rect 457876 276198 457918 276434
rect 458154 276198 458196 276434
rect 457876 269434 458196 276198
rect 457876 269198 457918 269434
rect 458154 269198 458196 269434
rect 457876 262434 458196 269198
rect 457876 262198 457918 262434
rect 458154 262198 458196 262434
rect 457876 255434 458196 262198
rect 457876 255198 457918 255434
rect 458154 255198 458196 255434
rect 457876 248434 458196 255198
rect 457876 248198 457918 248434
rect 458154 248198 458196 248434
rect 457876 241434 458196 248198
rect 457876 241198 457918 241434
rect 458154 241198 458196 241434
rect 457876 234434 458196 241198
rect 457876 234198 457918 234434
rect 458154 234198 458196 234434
rect 457876 227434 458196 234198
rect 457876 227198 457918 227434
rect 458154 227198 458196 227434
rect 457876 220434 458196 227198
rect 457876 220198 457918 220434
rect 458154 220198 458196 220434
rect 457876 213434 458196 220198
rect 457876 213198 457918 213434
rect 458154 213198 458196 213434
rect 457876 206434 458196 213198
rect 457876 206198 457918 206434
rect 458154 206198 458196 206434
rect 457876 199434 458196 206198
rect 457876 199198 457918 199434
rect 458154 199198 458196 199434
rect 457876 192434 458196 199198
rect 457876 192198 457918 192434
rect 458154 192198 458196 192434
rect 457876 185434 458196 192198
rect 457876 185198 457918 185434
rect 458154 185198 458196 185434
rect 457876 178434 458196 185198
rect 457876 178198 457918 178434
rect 458154 178198 458196 178434
rect 457876 171434 458196 178198
rect 457876 171198 457918 171434
rect 458154 171198 458196 171434
rect 457876 164434 458196 171198
rect 457876 164198 457918 164434
rect 458154 164198 458196 164434
rect 457876 157434 458196 164198
rect 457876 157198 457918 157434
rect 458154 157198 458196 157434
rect 457876 150434 458196 157198
rect 457876 150198 457918 150434
rect 458154 150198 458196 150434
rect 457876 143434 458196 150198
rect 457876 143198 457918 143434
rect 458154 143198 458196 143434
rect 457876 136434 458196 143198
rect 457876 136198 457918 136434
rect 458154 136198 458196 136434
rect 457876 129434 458196 136198
rect 457876 129198 457918 129434
rect 458154 129198 458196 129434
rect 457876 122434 458196 129198
rect 457876 122198 457918 122434
rect 458154 122198 458196 122434
rect 457876 115434 458196 122198
rect 457876 115198 457918 115434
rect 458154 115198 458196 115434
rect 457876 108434 458196 115198
rect 457876 108198 457918 108434
rect 458154 108198 458196 108434
rect 457876 101434 458196 108198
rect 457876 101198 457918 101434
rect 458154 101198 458196 101434
rect 457876 94434 458196 101198
rect 457876 94198 457918 94434
rect 458154 94198 458196 94434
rect 457876 87434 458196 94198
rect 457876 87198 457918 87434
rect 458154 87198 458196 87434
rect 457876 80434 458196 87198
rect 457876 80198 457918 80434
rect 458154 80198 458196 80434
rect 457876 73434 458196 80198
rect 457876 73198 457918 73434
rect 458154 73198 458196 73434
rect 457876 66434 458196 73198
rect 457876 66198 457918 66434
rect 458154 66198 458196 66434
rect 457876 59434 458196 66198
rect 457876 59198 457918 59434
rect 458154 59198 458196 59434
rect 457876 52434 458196 59198
rect 457876 52198 457918 52434
rect 458154 52198 458196 52434
rect 457876 45434 458196 52198
rect 457876 45198 457918 45434
rect 458154 45198 458196 45434
rect 457876 38434 458196 45198
rect 457876 38198 457918 38434
rect 458154 38198 458196 38434
rect 457876 31434 458196 38198
rect 457876 31198 457918 31434
rect 458154 31198 458196 31434
rect 457876 24434 458196 31198
rect 457876 24198 457918 24434
rect 458154 24198 458196 24434
rect 457876 17434 458196 24198
rect 457876 17198 457918 17434
rect 458154 17198 458196 17434
rect 457876 10434 458196 17198
rect 457876 10198 457918 10434
rect 458154 10198 458196 10434
rect 457876 3434 458196 10198
rect 457876 3198 457918 3434
rect 458154 3198 458196 3434
rect 457876 -1706 458196 3198
rect 457876 -1942 457918 -1706
rect 458154 -1942 458196 -1706
rect 457876 -2026 458196 -1942
rect 457876 -2262 457918 -2026
rect 458154 -2262 458196 -2026
rect 457876 -2294 458196 -2262
rect 463144 705238 463464 706230
rect 463144 705002 463186 705238
rect 463422 705002 463464 705238
rect 463144 704918 463464 705002
rect 463144 704682 463186 704918
rect 463422 704682 463464 704918
rect 463144 695494 463464 704682
rect 463144 695258 463186 695494
rect 463422 695258 463464 695494
rect 463144 688494 463464 695258
rect 463144 688258 463186 688494
rect 463422 688258 463464 688494
rect 463144 681494 463464 688258
rect 463144 681258 463186 681494
rect 463422 681258 463464 681494
rect 463144 674494 463464 681258
rect 463144 674258 463186 674494
rect 463422 674258 463464 674494
rect 463144 667494 463464 674258
rect 463144 667258 463186 667494
rect 463422 667258 463464 667494
rect 463144 660494 463464 667258
rect 463144 660258 463186 660494
rect 463422 660258 463464 660494
rect 463144 653494 463464 660258
rect 463144 653258 463186 653494
rect 463422 653258 463464 653494
rect 463144 646494 463464 653258
rect 463144 646258 463186 646494
rect 463422 646258 463464 646494
rect 463144 639494 463464 646258
rect 463144 639258 463186 639494
rect 463422 639258 463464 639494
rect 463144 632494 463464 639258
rect 463144 632258 463186 632494
rect 463422 632258 463464 632494
rect 463144 625494 463464 632258
rect 463144 625258 463186 625494
rect 463422 625258 463464 625494
rect 463144 618494 463464 625258
rect 463144 618258 463186 618494
rect 463422 618258 463464 618494
rect 463144 611494 463464 618258
rect 463144 611258 463186 611494
rect 463422 611258 463464 611494
rect 463144 604494 463464 611258
rect 463144 604258 463186 604494
rect 463422 604258 463464 604494
rect 463144 597494 463464 604258
rect 463144 597258 463186 597494
rect 463422 597258 463464 597494
rect 463144 590494 463464 597258
rect 463144 590258 463186 590494
rect 463422 590258 463464 590494
rect 463144 583494 463464 590258
rect 463144 583258 463186 583494
rect 463422 583258 463464 583494
rect 463144 576494 463464 583258
rect 463144 576258 463186 576494
rect 463422 576258 463464 576494
rect 463144 569494 463464 576258
rect 463144 569258 463186 569494
rect 463422 569258 463464 569494
rect 463144 562494 463464 569258
rect 463144 562258 463186 562494
rect 463422 562258 463464 562494
rect 463144 555494 463464 562258
rect 463144 555258 463186 555494
rect 463422 555258 463464 555494
rect 463144 548494 463464 555258
rect 463144 548258 463186 548494
rect 463422 548258 463464 548494
rect 463144 541494 463464 548258
rect 463144 541258 463186 541494
rect 463422 541258 463464 541494
rect 463144 534494 463464 541258
rect 463144 534258 463186 534494
rect 463422 534258 463464 534494
rect 463144 527494 463464 534258
rect 463144 527258 463186 527494
rect 463422 527258 463464 527494
rect 463144 520494 463464 527258
rect 463144 520258 463186 520494
rect 463422 520258 463464 520494
rect 463144 513494 463464 520258
rect 463144 513258 463186 513494
rect 463422 513258 463464 513494
rect 463144 506494 463464 513258
rect 463144 506258 463186 506494
rect 463422 506258 463464 506494
rect 463144 499494 463464 506258
rect 463144 499258 463186 499494
rect 463422 499258 463464 499494
rect 463144 492494 463464 499258
rect 463144 492258 463186 492494
rect 463422 492258 463464 492494
rect 463144 485494 463464 492258
rect 463144 485258 463186 485494
rect 463422 485258 463464 485494
rect 463144 478494 463464 485258
rect 463144 478258 463186 478494
rect 463422 478258 463464 478494
rect 463144 471494 463464 478258
rect 463144 471258 463186 471494
rect 463422 471258 463464 471494
rect 463144 464494 463464 471258
rect 463144 464258 463186 464494
rect 463422 464258 463464 464494
rect 463144 457494 463464 464258
rect 463144 457258 463186 457494
rect 463422 457258 463464 457494
rect 463144 450494 463464 457258
rect 463144 450258 463186 450494
rect 463422 450258 463464 450494
rect 463144 443494 463464 450258
rect 463144 443258 463186 443494
rect 463422 443258 463464 443494
rect 463144 436494 463464 443258
rect 463144 436258 463186 436494
rect 463422 436258 463464 436494
rect 463144 429494 463464 436258
rect 463144 429258 463186 429494
rect 463422 429258 463464 429494
rect 463144 422494 463464 429258
rect 463144 422258 463186 422494
rect 463422 422258 463464 422494
rect 463144 415494 463464 422258
rect 463144 415258 463186 415494
rect 463422 415258 463464 415494
rect 463144 408494 463464 415258
rect 463144 408258 463186 408494
rect 463422 408258 463464 408494
rect 463144 401494 463464 408258
rect 463144 401258 463186 401494
rect 463422 401258 463464 401494
rect 463144 394494 463464 401258
rect 463144 394258 463186 394494
rect 463422 394258 463464 394494
rect 463144 387494 463464 394258
rect 463144 387258 463186 387494
rect 463422 387258 463464 387494
rect 463144 380494 463464 387258
rect 463144 380258 463186 380494
rect 463422 380258 463464 380494
rect 463144 373494 463464 380258
rect 463144 373258 463186 373494
rect 463422 373258 463464 373494
rect 463144 366494 463464 373258
rect 463144 366258 463186 366494
rect 463422 366258 463464 366494
rect 463144 359494 463464 366258
rect 463144 359258 463186 359494
rect 463422 359258 463464 359494
rect 463144 352494 463464 359258
rect 463144 352258 463186 352494
rect 463422 352258 463464 352494
rect 463144 345494 463464 352258
rect 463144 345258 463186 345494
rect 463422 345258 463464 345494
rect 463144 338494 463464 345258
rect 463144 338258 463186 338494
rect 463422 338258 463464 338494
rect 463144 331494 463464 338258
rect 463144 331258 463186 331494
rect 463422 331258 463464 331494
rect 463144 324494 463464 331258
rect 463144 324258 463186 324494
rect 463422 324258 463464 324494
rect 463144 317494 463464 324258
rect 463144 317258 463186 317494
rect 463422 317258 463464 317494
rect 463144 310494 463464 317258
rect 463144 310258 463186 310494
rect 463422 310258 463464 310494
rect 463144 303494 463464 310258
rect 463144 303258 463186 303494
rect 463422 303258 463464 303494
rect 463144 296494 463464 303258
rect 463144 296258 463186 296494
rect 463422 296258 463464 296494
rect 463144 289494 463464 296258
rect 463144 289258 463186 289494
rect 463422 289258 463464 289494
rect 463144 282494 463464 289258
rect 463144 282258 463186 282494
rect 463422 282258 463464 282494
rect 463144 275494 463464 282258
rect 463144 275258 463186 275494
rect 463422 275258 463464 275494
rect 463144 268494 463464 275258
rect 463144 268258 463186 268494
rect 463422 268258 463464 268494
rect 463144 261494 463464 268258
rect 463144 261258 463186 261494
rect 463422 261258 463464 261494
rect 463144 254494 463464 261258
rect 463144 254258 463186 254494
rect 463422 254258 463464 254494
rect 463144 247494 463464 254258
rect 463144 247258 463186 247494
rect 463422 247258 463464 247494
rect 463144 240494 463464 247258
rect 463144 240258 463186 240494
rect 463422 240258 463464 240494
rect 463144 233494 463464 240258
rect 463144 233258 463186 233494
rect 463422 233258 463464 233494
rect 463144 226494 463464 233258
rect 463144 226258 463186 226494
rect 463422 226258 463464 226494
rect 463144 219494 463464 226258
rect 463144 219258 463186 219494
rect 463422 219258 463464 219494
rect 463144 212494 463464 219258
rect 463144 212258 463186 212494
rect 463422 212258 463464 212494
rect 463144 205494 463464 212258
rect 463144 205258 463186 205494
rect 463422 205258 463464 205494
rect 463144 198494 463464 205258
rect 463144 198258 463186 198494
rect 463422 198258 463464 198494
rect 463144 191494 463464 198258
rect 463144 191258 463186 191494
rect 463422 191258 463464 191494
rect 463144 184494 463464 191258
rect 463144 184258 463186 184494
rect 463422 184258 463464 184494
rect 463144 177494 463464 184258
rect 463144 177258 463186 177494
rect 463422 177258 463464 177494
rect 463144 170494 463464 177258
rect 463144 170258 463186 170494
rect 463422 170258 463464 170494
rect 463144 163494 463464 170258
rect 463144 163258 463186 163494
rect 463422 163258 463464 163494
rect 463144 156494 463464 163258
rect 463144 156258 463186 156494
rect 463422 156258 463464 156494
rect 463144 149494 463464 156258
rect 463144 149258 463186 149494
rect 463422 149258 463464 149494
rect 463144 142494 463464 149258
rect 463144 142258 463186 142494
rect 463422 142258 463464 142494
rect 463144 135494 463464 142258
rect 463144 135258 463186 135494
rect 463422 135258 463464 135494
rect 463144 128494 463464 135258
rect 463144 128258 463186 128494
rect 463422 128258 463464 128494
rect 463144 121494 463464 128258
rect 463144 121258 463186 121494
rect 463422 121258 463464 121494
rect 463144 114494 463464 121258
rect 463144 114258 463186 114494
rect 463422 114258 463464 114494
rect 463144 107494 463464 114258
rect 463144 107258 463186 107494
rect 463422 107258 463464 107494
rect 463144 100494 463464 107258
rect 463144 100258 463186 100494
rect 463422 100258 463464 100494
rect 463144 93494 463464 100258
rect 463144 93258 463186 93494
rect 463422 93258 463464 93494
rect 463144 86494 463464 93258
rect 463144 86258 463186 86494
rect 463422 86258 463464 86494
rect 463144 79494 463464 86258
rect 463144 79258 463186 79494
rect 463422 79258 463464 79494
rect 463144 72494 463464 79258
rect 463144 72258 463186 72494
rect 463422 72258 463464 72494
rect 463144 65494 463464 72258
rect 463144 65258 463186 65494
rect 463422 65258 463464 65494
rect 463144 58494 463464 65258
rect 463144 58258 463186 58494
rect 463422 58258 463464 58494
rect 463144 51494 463464 58258
rect 463144 51258 463186 51494
rect 463422 51258 463464 51494
rect 463144 44494 463464 51258
rect 463144 44258 463186 44494
rect 463422 44258 463464 44494
rect 463144 37494 463464 44258
rect 463144 37258 463186 37494
rect 463422 37258 463464 37494
rect 463144 30494 463464 37258
rect 463144 30258 463186 30494
rect 463422 30258 463464 30494
rect 463144 23494 463464 30258
rect 463144 23258 463186 23494
rect 463422 23258 463464 23494
rect 463144 16494 463464 23258
rect 463144 16258 463186 16494
rect 463422 16258 463464 16494
rect 463144 9494 463464 16258
rect 463144 9258 463186 9494
rect 463422 9258 463464 9494
rect 463144 2494 463464 9258
rect 463144 2258 463186 2494
rect 463422 2258 463464 2494
rect 463144 -746 463464 2258
rect 463144 -982 463186 -746
rect 463422 -982 463464 -746
rect 463144 -1066 463464 -982
rect 463144 -1302 463186 -1066
rect 463422 -1302 463464 -1066
rect 463144 -2294 463464 -1302
rect 464876 706198 465196 706230
rect 464876 705962 464918 706198
rect 465154 705962 465196 706198
rect 464876 705878 465196 705962
rect 464876 705642 464918 705878
rect 465154 705642 465196 705878
rect 464876 696434 465196 705642
rect 464876 696198 464918 696434
rect 465154 696198 465196 696434
rect 464876 689434 465196 696198
rect 464876 689198 464918 689434
rect 465154 689198 465196 689434
rect 464876 682434 465196 689198
rect 464876 682198 464918 682434
rect 465154 682198 465196 682434
rect 464876 675434 465196 682198
rect 464876 675198 464918 675434
rect 465154 675198 465196 675434
rect 464876 668434 465196 675198
rect 464876 668198 464918 668434
rect 465154 668198 465196 668434
rect 464876 661434 465196 668198
rect 464876 661198 464918 661434
rect 465154 661198 465196 661434
rect 464876 654434 465196 661198
rect 464876 654198 464918 654434
rect 465154 654198 465196 654434
rect 464876 647434 465196 654198
rect 464876 647198 464918 647434
rect 465154 647198 465196 647434
rect 464876 640434 465196 647198
rect 464876 640198 464918 640434
rect 465154 640198 465196 640434
rect 464876 633434 465196 640198
rect 464876 633198 464918 633434
rect 465154 633198 465196 633434
rect 464876 626434 465196 633198
rect 464876 626198 464918 626434
rect 465154 626198 465196 626434
rect 464876 619434 465196 626198
rect 464876 619198 464918 619434
rect 465154 619198 465196 619434
rect 464876 612434 465196 619198
rect 464876 612198 464918 612434
rect 465154 612198 465196 612434
rect 464876 605434 465196 612198
rect 464876 605198 464918 605434
rect 465154 605198 465196 605434
rect 464876 598434 465196 605198
rect 464876 598198 464918 598434
rect 465154 598198 465196 598434
rect 464876 591434 465196 598198
rect 464876 591198 464918 591434
rect 465154 591198 465196 591434
rect 464876 584434 465196 591198
rect 464876 584198 464918 584434
rect 465154 584198 465196 584434
rect 464876 577434 465196 584198
rect 464876 577198 464918 577434
rect 465154 577198 465196 577434
rect 464876 570434 465196 577198
rect 464876 570198 464918 570434
rect 465154 570198 465196 570434
rect 464876 563434 465196 570198
rect 464876 563198 464918 563434
rect 465154 563198 465196 563434
rect 464876 556434 465196 563198
rect 464876 556198 464918 556434
rect 465154 556198 465196 556434
rect 464876 549434 465196 556198
rect 464876 549198 464918 549434
rect 465154 549198 465196 549434
rect 464876 542434 465196 549198
rect 464876 542198 464918 542434
rect 465154 542198 465196 542434
rect 464876 535434 465196 542198
rect 464876 535198 464918 535434
rect 465154 535198 465196 535434
rect 464876 528434 465196 535198
rect 464876 528198 464918 528434
rect 465154 528198 465196 528434
rect 464876 521434 465196 528198
rect 464876 521198 464918 521434
rect 465154 521198 465196 521434
rect 464876 514434 465196 521198
rect 464876 514198 464918 514434
rect 465154 514198 465196 514434
rect 464876 507434 465196 514198
rect 464876 507198 464918 507434
rect 465154 507198 465196 507434
rect 464876 500434 465196 507198
rect 464876 500198 464918 500434
rect 465154 500198 465196 500434
rect 464876 493434 465196 500198
rect 464876 493198 464918 493434
rect 465154 493198 465196 493434
rect 464876 486434 465196 493198
rect 464876 486198 464918 486434
rect 465154 486198 465196 486434
rect 464876 479434 465196 486198
rect 464876 479198 464918 479434
rect 465154 479198 465196 479434
rect 464876 472434 465196 479198
rect 464876 472198 464918 472434
rect 465154 472198 465196 472434
rect 464876 465434 465196 472198
rect 464876 465198 464918 465434
rect 465154 465198 465196 465434
rect 464876 458434 465196 465198
rect 464876 458198 464918 458434
rect 465154 458198 465196 458434
rect 464876 451434 465196 458198
rect 464876 451198 464918 451434
rect 465154 451198 465196 451434
rect 464876 444434 465196 451198
rect 464876 444198 464918 444434
rect 465154 444198 465196 444434
rect 464876 437434 465196 444198
rect 464876 437198 464918 437434
rect 465154 437198 465196 437434
rect 464876 430434 465196 437198
rect 464876 430198 464918 430434
rect 465154 430198 465196 430434
rect 464876 423434 465196 430198
rect 464876 423198 464918 423434
rect 465154 423198 465196 423434
rect 464876 416434 465196 423198
rect 464876 416198 464918 416434
rect 465154 416198 465196 416434
rect 464876 409434 465196 416198
rect 464876 409198 464918 409434
rect 465154 409198 465196 409434
rect 464876 402434 465196 409198
rect 464876 402198 464918 402434
rect 465154 402198 465196 402434
rect 464876 395434 465196 402198
rect 464876 395198 464918 395434
rect 465154 395198 465196 395434
rect 464876 388434 465196 395198
rect 464876 388198 464918 388434
rect 465154 388198 465196 388434
rect 464876 381434 465196 388198
rect 464876 381198 464918 381434
rect 465154 381198 465196 381434
rect 464876 374434 465196 381198
rect 464876 374198 464918 374434
rect 465154 374198 465196 374434
rect 464876 367434 465196 374198
rect 464876 367198 464918 367434
rect 465154 367198 465196 367434
rect 464876 360434 465196 367198
rect 464876 360198 464918 360434
rect 465154 360198 465196 360434
rect 464876 353434 465196 360198
rect 464876 353198 464918 353434
rect 465154 353198 465196 353434
rect 464876 346434 465196 353198
rect 464876 346198 464918 346434
rect 465154 346198 465196 346434
rect 464876 339434 465196 346198
rect 464876 339198 464918 339434
rect 465154 339198 465196 339434
rect 464876 332434 465196 339198
rect 464876 332198 464918 332434
rect 465154 332198 465196 332434
rect 464876 325434 465196 332198
rect 464876 325198 464918 325434
rect 465154 325198 465196 325434
rect 464876 318434 465196 325198
rect 464876 318198 464918 318434
rect 465154 318198 465196 318434
rect 464876 311434 465196 318198
rect 464876 311198 464918 311434
rect 465154 311198 465196 311434
rect 464876 304434 465196 311198
rect 464876 304198 464918 304434
rect 465154 304198 465196 304434
rect 464876 297434 465196 304198
rect 464876 297198 464918 297434
rect 465154 297198 465196 297434
rect 464876 290434 465196 297198
rect 464876 290198 464918 290434
rect 465154 290198 465196 290434
rect 464876 283434 465196 290198
rect 464876 283198 464918 283434
rect 465154 283198 465196 283434
rect 464876 276434 465196 283198
rect 464876 276198 464918 276434
rect 465154 276198 465196 276434
rect 464876 269434 465196 276198
rect 464876 269198 464918 269434
rect 465154 269198 465196 269434
rect 464876 262434 465196 269198
rect 464876 262198 464918 262434
rect 465154 262198 465196 262434
rect 464876 255434 465196 262198
rect 464876 255198 464918 255434
rect 465154 255198 465196 255434
rect 464876 248434 465196 255198
rect 464876 248198 464918 248434
rect 465154 248198 465196 248434
rect 464876 241434 465196 248198
rect 464876 241198 464918 241434
rect 465154 241198 465196 241434
rect 464876 234434 465196 241198
rect 464876 234198 464918 234434
rect 465154 234198 465196 234434
rect 464876 227434 465196 234198
rect 464876 227198 464918 227434
rect 465154 227198 465196 227434
rect 464876 220434 465196 227198
rect 464876 220198 464918 220434
rect 465154 220198 465196 220434
rect 464876 213434 465196 220198
rect 464876 213198 464918 213434
rect 465154 213198 465196 213434
rect 464876 206434 465196 213198
rect 464876 206198 464918 206434
rect 465154 206198 465196 206434
rect 464876 199434 465196 206198
rect 464876 199198 464918 199434
rect 465154 199198 465196 199434
rect 464876 192434 465196 199198
rect 464876 192198 464918 192434
rect 465154 192198 465196 192434
rect 464876 185434 465196 192198
rect 464876 185198 464918 185434
rect 465154 185198 465196 185434
rect 464876 178434 465196 185198
rect 464876 178198 464918 178434
rect 465154 178198 465196 178434
rect 464876 171434 465196 178198
rect 464876 171198 464918 171434
rect 465154 171198 465196 171434
rect 464876 164434 465196 171198
rect 464876 164198 464918 164434
rect 465154 164198 465196 164434
rect 464876 157434 465196 164198
rect 464876 157198 464918 157434
rect 465154 157198 465196 157434
rect 464876 150434 465196 157198
rect 464876 150198 464918 150434
rect 465154 150198 465196 150434
rect 464876 143434 465196 150198
rect 464876 143198 464918 143434
rect 465154 143198 465196 143434
rect 464876 136434 465196 143198
rect 464876 136198 464918 136434
rect 465154 136198 465196 136434
rect 464876 129434 465196 136198
rect 464876 129198 464918 129434
rect 465154 129198 465196 129434
rect 464876 122434 465196 129198
rect 464876 122198 464918 122434
rect 465154 122198 465196 122434
rect 464876 115434 465196 122198
rect 464876 115198 464918 115434
rect 465154 115198 465196 115434
rect 464876 108434 465196 115198
rect 464876 108198 464918 108434
rect 465154 108198 465196 108434
rect 464876 101434 465196 108198
rect 464876 101198 464918 101434
rect 465154 101198 465196 101434
rect 464876 94434 465196 101198
rect 464876 94198 464918 94434
rect 465154 94198 465196 94434
rect 464876 87434 465196 94198
rect 464876 87198 464918 87434
rect 465154 87198 465196 87434
rect 464876 80434 465196 87198
rect 464876 80198 464918 80434
rect 465154 80198 465196 80434
rect 464876 73434 465196 80198
rect 464876 73198 464918 73434
rect 465154 73198 465196 73434
rect 464876 66434 465196 73198
rect 464876 66198 464918 66434
rect 465154 66198 465196 66434
rect 464876 59434 465196 66198
rect 464876 59198 464918 59434
rect 465154 59198 465196 59434
rect 464876 52434 465196 59198
rect 464876 52198 464918 52434
rect 465154 52198 465196 52434
rect 464876 45434 465196 52198
rect 464876 45198 464918 45434
rect 465154 45198 465196 45434
rect 464876 38434 465196 45198
rect 464876 38198 464918 38434
rect 465154 38198 465196 38434
rect 464876 31434 465196 38198
rect 464876 31198 464918 31434
rect 465154 31198 465196 31434
rect 464876 24434 465196 31198
rect 464876 24198 464918 24434
rect 465154 24198 465196 24434
rect 464876 17434 465196 24198
rect 464876 17198 464918 17434
rect 465154 17198 465196 17434
rect 464876 10434 465196 17198
rect 464876 10198 464918 10434
rect 465154 10198 465196 10434
rect 464876 3434 465196 10198
rect 464876 3198 464918 3434
rect 465154 3198 465196 3434
rect 464876 -1706 465196 3198
rect 464876 -1942 464918 -1706
rect 465154 -1942 465196 -1706
rect 464876 -2026 465196 -1942
rect 464876 -2262 464918 -2026
rect 465154 -2262 465196 -2026
rect 464876 -2294 465196 -2262
rect 470144 705238 470464 706230
rect 470144 705002 470186 705238
rect 470422 705002 470464 705238
rect 470144 704918 470464 705002
rect 470144 704682 470186 704918
rect 470422 704682 470464 704918
rect 470144 695494 470464 704682
rect 470144 695258 470186 695494
rect 470422 695258 470464 695494
rect 470144 688494 470464 695258
rect 470144 688258 470186 688494
rect 470422 688258 470464 688494
rect 470144 681494 470464 688258
rect 470144 681258 470186 681494
rect 470422 681258 470464 681494
rect 470144 674494 470464 681258
rect 470144 674258 470186 674494
rect 470422 674258 470464 674494
rect 470144 667494 470464 674258
rect 470144 667258 470186 667494
rect 470422 667258 470464 667494
rect 470144 660494 470464 667258
rect 470144 660258 470186 660494
rect 470422 660258 470464 660494
rect 470144 653494 470464 660258
rect 470144 653258 470186 653494
rect 470422 653258 470464 653494
rect 470144 646494 470464 653258
rect 470144 646258 470186 646494
rect 470422 646258 470464 646494
rect 470144 639494 470464 646258
rect 470144 639258 470186 639494
rect 470422 639258 470464 639494
rect 470144 632494 470464 639258
rect 470144 632258 470186 632494
rect 470422 632258 470464 632494
rect 470144 625494 470464 632258
rect 470144 625258 470186 625494
rect 470422 625258 470464 625494
rect 470144 618494 470464 625258
rect 470144 618258 470186 618494
rect 470422 618258 470464 618494
rect 470144 611494 470464 618258
rect 470144 611258 470186 611494
rect 470422 611258 470464 611494
rect 470144 604494 470464 611258
rect 470144 604258 470186 604494
rect 470422 604258 470464 604494
rect 470144 597494 470464 604258
rect 470144 597258 470186 597494
rect 470422 597258 470464 597494
rect 470144 590494 470464 597258
rect 470144 590258 470186 590494
rect 470422 590258 470464 590494
rect 470144 583494 470464 590258
rect 470144 583258 470186 583494
rect 470422 583258 470464 583494
rect 470144 576494 470464 583258
rect 470144 576258 470186 576494
rect 470422 576258 470464 576494
rect 470144 569494 470464 576258
rect 470144 569258 470186 569494
rect 470422 569258 470464 569494
rect 470144 562494 470464 569258
rect 470144 562258 470186 562494
rect 470422 562258 470464 562494
rect 470144 555494 470464 562258
rect 470144 555258 470186 555494
rect 470422 555258 470464 555494
rect 470144 548494 470464 555258
rect 470144 548258 470186 548494
rect 470422 548258 470464 548494
rect 470144 541494 470464 548258
rect 470144 541258 470186 541494
rect 470422 541258 470464 541494
rect 470144 534494 470464 541258
rect 470144 534258 470186 534494
rect 470422 534258 470464 534494
rect 470144 527494 470464 534258
rect 470144 527258 470186 527494
rect 470422 527258 470464 527494
rect 470144 520494 470464 527258
rect 470144 520258 470186 520494
rect 470422 520258 470464 520494
rect 470144 513494 470464 520258
rect 470144 513258 470186 513494
rect 470422 513258 470464 513494
rect 470144 506494 470464 513258
rect 470144 506258 470186 506494
rect 470422 506258 470464 506494
rect 470144 499494 470464 506258
rect 470144 499258 470186 499494
rect 470422 499258 470464 499494
rect 470144 492494 470464 499258
rect 470144 492258 470186 492494
rect 470422 492258 470464 492494
rect 470144 485494 470464 492258
rect 470144 485258 470186 485494
rect 470422 485258 470464 485494
rect 470144 478494 470464 485258
rect 470144 478258 470186 478494
rect 470422 478258 470464 478494
rect 470144 471494 470464 478258
rect 470144 471258 470186 471494
rect 470422 471258 470464 471494
rect 470144 464494 470464 471258
rect 470144 464258 470186 464494
rect 470422 464258 470464 464494
rect 470144 457494 470464 464258
rect 470144 457258 470186 457494
rect 470422 457258 470464 457494
rect 470144 450494 470464 457258
rect 470144 450258 470186 450494
rect 470422 450258 470464 450494
rect 470144 443494 470464 450258
rect 470144 443258 470186 443494
rect 470422 443258 470464 443494
rect 470144 436494 470464 443258
rect 470144 436258 470186 436494
rect 470422 436258 470464 436494
rect 470144 429494 470464 436258
rect 470144 429258 470186 429494
rect 470422 429258 470464 429494
rect 470144 422494 470464 429258
rect 470144 422258 470186 422494
rect 470422 422258 470464 422494
rect 470144 415494 470464 422258
rect 470144 415258 470186 415494
rect 470422 415258 470464 415494
rect 470144 408494 470464 415258
rect 470144 408258 470186 408494
rect 470422 408258 470464 408494
rect 470144 401494 470464 408258
rect 470144 401258 470186 401494
rect 470422 401258 470464 401494
rect 470144 394494 470464 401258
rect 470144 394258 470186 394494
rect 470422 394258 470464 394494
rect 470144 387494 470464 394258
rect 470144 387258 470186 387494
rect 470422 387258 470464 387494
rect 470144 380494 470464 387258
rect 470144 380258 470186 380494
rect 470422 380258 470464 380494
rect 470144 373494 470464 380258
rect 470144 373258 470186 373494
rect 470422 373258 470464 373494
rect 470144 366494 470464 373258
rect 470144 366258 470186 366494
rect 470422 366258 470464 366494
rect 470144 359494 470464 366258
rect 470144 359258 470186 359494
rect 470422 359258 470464 359494
rect 470144 352494 470464 359258
rect 470144 352258 470186 352494
rect 470422 352258 470464 352494
rect 470144 345494 470464 352258
rect 470144 345258 470186 345494
rect 470422 345258 470464 345494
rect 470144 338494 470464 345258
rect 470144 338258 470186 338494
rect 470422 338258 470464 338494
rect 470144 331494 470464 338258
rect 470144 331258 470186 331494
rect 470422 331258 470464 331494
rect 470144 324494 470464 331258
rect 470144 324258 470186 324494
rect 470422 324258 470464 324494
rect 470144 317494 470464 324258
rect 470144 317258 470186 317494
rect 470422 317258 470464 317494
rect 470144 310494 470464 317258
rect 470144 310258 470186 310494
rect 470422 310258 470464 310494
rect 470144 303494 470464 310258
rect 470144 303258 470186 303494
rect 470422 303258 470464 303494
rect 470144 296494 470464 303258
rect 470144 296258 470186 296494
rect 470422 296258 470464 296494
rect 470144 289494 470464 296258
rect 470144 289258 470186 289494
rect 470422 289258 470464 289494
rect 470144 282494 470464 289258
rect 470144 282258 470186 282494
rect 470422 282258 470464 282494
rect 470144 275494 470464 282258
rect 470144 275258 470186 275494
rect 470422 275258 470464 275494
rect 470144 268494 470464 275258
rect 470144 268258 470186 268494
rect 470422 268258 470464 268494
rect 470144 261494 470464 268258
rect 470144 261258 470186 261494
rect 470422 261258 470464 261494
rect 470144 254494 470464 261258
rect 470144 254258 470186 254494
rect 470422 254258 470464 254494
rect 470144 247494 470464 254258
rect 470144 247258 470186 247494
rect 470422 247258 470464 247494
rect 470144 240494 470464 247258
rect 470144 240258 470186 240494
rect 470422 240258 470464 240494
rect 470144 233494 470464 240258
rect 470144 233258 470186 233494
rect 470422 233258 470464 233494
rect 470144 226494 470464 233258
rect 470144 226258 470186 226494
rect 470422 226258 470464 226494
rect 470144 219494 470464 226258
rect 470144 219258 470186 219494
rect 470422 219258 470464 219494
rect 470144 212494 470464 219258
rect 470144 212258 470186 212494
rect 470422 212258 470464 212494
rect 470144 205494 470464 212258
rect 470144 205258 470186 205494
rect 470422 205258 470464 205494
rect 470144 198494 470464 205258
rect 470144 198258 470186 198494
rect 470422 198258 470464 198494
rect 470144 191494 470464 198258
rect 470144 191258 470186 191494
rect 470422 191258 470464 191494
rect 470144 184494 470464 191258
rect 470144 184258 470186 184494
rect 470422 184258 470464 184494
rect 470144 177494 470464 184258
rect 470144 177258 470186 177494
rect 470422 177258 470464 177494
rect 470144 170494 470464 177258
rect 470144 170258 470186 170494
rect 470422 170258 470464 170494
rect 470144 163494 470464 170258
rect 470144 163258 470186 163494
rect 470422 163258 470464 163494
rect 470144 156494 470464 163258
rect 470144 156258 470186 156494
rect 470422 156258 470464 156494
rect 470144 149494 470464 156258
rect 470144 149258 470186 149494
rect 470422 149258 470464 149494
rect 470144 142494 470464 149258
rect 470144 142258 470186 142494
rect 470422 142258 470464 142494
rect 470144 135494 470464 142258
rect 470144 135258 470186 135494
rect 470422 135258 470464 135494
rect 470144 128494 470464 135258
rect 470144 128258 470186 128494
rect 470422 128258 470464 128494
rect 470144 121494 470464 128258
rect 470144 121258 470186 121494
rect 470422 121258 470464 121494
rect 470144 114494 470464 121258
rect 470144 114258 470186 114494
rect 470422 114258 470464 114494
rect 470144 107494 470464 114258
rect 470144 107258 470186 107494
rect 470422 107258 470464 107494
rect 470144 100494 470464 107258
rect 470144 100258 470186 100494
rect 470422 100258 470464 100494
rect 470144 93494 470464 100258
rect 470144 93258 470186 93494
rect 470422 93258 470464 93494
rect 470144 86494 470464 93258
rect 470144 86258 470186 86494
rect 470422 86258 470464 86494
rect 470144 79494 470464 86258
rect 470144 79258 470186 79494
rect 470422 79258 470464 79494
rect 470144 72494 470464 79258
rect 470144 72258 470186 72494
rect 470422 72258 470464 72494
rect 470144 65494 470464 72258
rect 470144 65258 470186 65494
rect 470422 65258 470464 65494
rect 470144 58494 470464 65258
rect 470144 58258 470186 58494
rect 470422 58258 470464 58494
rect 470144 51494 470464 58258
rect 470144 51258 470186 51494
rect 470422 51258 470464 51494
rect 470144 44494 470464 51258
rect 470144 44258 470186 44494
rect 470422 44258 470464 44494
rect 470144 37494 470464 44258
rect 470144 37258 470186 37494
rect 470422 37258 470464 37494
rect 470144 30494 470464 37258
rect 470144 30258 470186 30494
rect 470422 30258 470464 30494
rect 470144 23494 470464 30258
rect 470144 23258 470186 23494
rect 470422 23258 470464 23494
rect 470144 16494 470464 23258
rect 470144 16258 470186 16494
rect 470422 16258 470464 16494
rect 470144 9494 470464 16258
rect 470144 9258 470186 9494
rect 470422 9258 470464 9494
rect 470144 2494 470464 9258
rect 470144 2258 470186 2494
rect 470422 2258 470464 2494
rect 470144 -746 470464 2258
rect 470144 -982 470186 -746
rect 470422 -982 470464 -746
rect 470144 -1066 470464 -982
rect 470144 -1302 470186 -1066
rect 470422 -1302 470464 -1066
rect 470144 -2294 470464 -1302
rect 471876 706198 472196 706230
rect 471876 705962 471918 706198
rect 472154 705962 472196 706198
rect 471876 705878 472196 705962
rect 471876 705642 471918 705878
rect 472154 705642 472196 705878
rect 471876 696434 472196 705642
rect 471876 696198 471918 696434
rect 472154 696198 472196 696434
rect 471876 689434 472196 696198
rect 471876 689198 471918 689434
rect 472154 689198 472196 689434
rect 471876 682434 472196 689198
rect 471876 682198 471918 682434
rect 472154 682198 472196 682434
rect 471876 675434 472196 682198
rect 471876 675198 471918 675434
rect 472154 675198 472196 675434
rect 471876 668434 472196 675198
rect 471876 668198 471918 668434
rect 472154 668198 472196 668434
rect 471876 661434 472196 668198
rect 471876 661198 471918 661434
rect 472154 661198 472196 661434
rect 471876 654434 472196 661198
rect 471876 654198 471918 654434
rect 472154 654198 472196 654434
rect 471876 647434 472196 654198
rect 471876 647198 471918 647434
rect 472154 647198 472196 647434
rect 471876 640434 472196 647198
rect 471876 640198 471918 640434
rect 472154 640198 472196 640434
rect 471876 633434 472196 640198
rect 471876 633198 471918 633434
rect 472154 633198 472196 633434
rect 471876 626434 472196 633198
rect 471876 626198 471918 626434
rect 472154 626198 472196 626434
rect 471876 619434 472196 626198
rect 471876 619198 471918 619434
rect 472154 619198 472196 619434
rect 471876 612434 472196 619198
rect 471876 612198 471918 612434
rect 472154 612198 472196 612434
rect 471876 605434 472196 612198
rect 471876 605198 471918 605434
rect 472154 605198 472196 605434
rect 471876 598434 472196 605198
rect 471876 598198 471918 598434
rect 472154 598198 472196 598434
rect 471876 591434 472196 598198
rect 471876 591198 471918 591434
rect 472154 591198 472196 591434
rect 471876 584434 472196 591198
rect 471876 584198 471918 584434
rect 472154 584198 472196 584434
rect 471876 577434 472196 584198
rect 471876 577198 471918 577434
rect 472154 577198 472196 577434
rect 471876 570434 472196 577198
rect 471876 570198 471918 570434
rect 472154 570198 472196 570434
rect 471876 563434 472196 570198
rect 471876 563198 471918 563434
rect 472154 563198 472196 563434
rect 471876 556434 472196 563198
rect 471876 556198 471918 556434
rect 472154 556198 472196 556434
rect 471876 549434 472196 556198
rect 471876 549198 471918 549434
rect 472154 549198 472196 549434
rect 471876 542434 472196 549198
rect 471876 542198 471918 542434
rect 472154 542198 472196 542434
rect 471876 535434 472196 542198
rect 471876 535198 471918 535434
rect 472154 535198 472196 535434
rect 471876 528434 472196 535198
rect 471876 528198 471918 528434
rect 472154 528198 472196 528434
rect 471876 521434 472196 528198
rect 471876 521198 471918 521434
rect 472154 521198 472196 521434
rect 471876 514434 472196 521198
rect 471876 514198 471918 514434
rect 472154 514198 472196 514434
rect 471876 507434 472196 514198
rect 471876 507198 471918 507434
rect 472154 507198 472196 507434
rect 471876 500434 472196 507198
rect 471876 500198 471918 500434
rect 472154 500198 472196 500434
rect 471876 493434 472196 500198
rect 471876 493198 471918 493434
rect 472154 493198 472196 493434
rect 471876 486434 472196 493198
rect 471876 486198 471918 486434
rect 472154 486198 472196 486434
rect 471876 479434 472196 486198
rect 471876 479198 471918 479434
rect 472154 479198 472196 479434
rect 471876 472434 472196 479198
rect 471876 472198 471918 472434
rect 472154 472198 472196 472434
rect 471876 465434 472196 472198
rect 471876 465198 471918 465434
rect 472154 465198 472196 465434
rect 471876 458434 472196 465198
rect 471876 458198 471918 458434
rect 472154 458198 472196 458434
rect 471876 451434 472196 458198
rect 471876 451198 471918 451434
rect 472154 451198 472196 451434
rect 471876 444434 472196 451198
rect 471876 444198 471918 444434
rect 472154 444198 472196 444434
rect 471876 437434 472196 444198
rect 471876 437198 471918 437434
rect 472154 437198 472196 437434
rect 471876 430434 472196 437198
rect 471876 430198 471918 430434
rect 472154 430198 472196 430434
rect 471876 423434 472196 430198
rect 471876 423198 471918 423434
rect 472154 423198 472196 423434
rect 471876 416434 472196 423198
rect 471876 416198 471918 416434
rect 472154 416198 472196 416434
rect 471876 409434 472196 416198
rect 471876 409198 471918 409434
rect 472154 409198 472196 409434
rect 471876 402434 472196 409198
rect 471876 402198 471918 402434
rect 472154 402198 472196 402434
rect 471876 395434 472196 402198
rect 471876 395198 471918 395434
rect 472154 395198 472196 395434
rect 471876 388434 472196 395198
rect 471876 388198 471918 388434
rect 472154 388198 472196 388434
rect 471876 381434 472196 388198
rect 471876 381198 471918 381434
rect 472154 381198 472196 381434
rect 471876 374434 472196 381198
rect 471876 374198 471918 374434
rect 472154 374198 472196 374434
rect 471876 367434 472196 374198
rect 471876 367198 471918 367434
rect 472154 367198 472196 367434
rect 471876 360434 472196 367198
rect 471876 360198 471918 360434
rect 472154 360198 472196 360434
rect 471876 353434 472196 360198
rect 471876 353198 471918 353434
rect 472154 353198 472196 353434
rect 471876 346434 472196 353198
rect 471876 346198 471918 346434
rect 472154 346198 472196 346434
rect 471876 339434 472196 346198
rect 471876 339198 471918 339434
rect 472154 339198 472196 339434
rect 471876 332434 472196 339198
rect 471876 332198 471918 332434
rect 472154 332198 472196 332434
rect 471876 325434 472196 332198
rect 471876 325198 471918 325434
rect 472154 325198 472196 325434
rect 471876 318434 472196 325198
rect 471876 318198 471918 318434
rect 472154 318198 472196 318434
rect 471876 311434 472196 318198
rect 471876 311198 471918 311434
rect 472154 311198 472196 311434
rect 471876 304434 472196 311198
rect 471876 304198 471918 304434
rect 472154 304198 472196 304434
rect 471876 297434 472196 304198
rect 471876 297198 471918 297434
rect 472154 297198 472196 297434
rect 471876 290434 472196 297198
rect 471876 290198 471918 290434
rect 472154 290198 472196 290434
rect 471876 283434 472196 290198
rect 471876 283198 471918 283434
rect 472154 283198 472196 283434
rect 471876 276434 472196 283198
rect 471876 276198 471918 276434
rect 472154 276198 472196 276434
rect 471876 269434 472196 276198
rect 471876 269198 471918 269434
rect 472154 269198 472196 269434
rect 471876 262434 472196 269198
rect 471876 262198 471918 262434
rect 472154 262198 472196 262434
rect 471876 255434 472196 262198
rect 471876 255198 471918 255434
rect 472154 255198 472196 255434
rect 471876 248434 472196 255198
rect 471876 248198 471918 248434
rect 472154 248198 472196 248434
rect 471876 241434 472196 248198
rect 471876 241198 471918 241434
rect 472154 241198 472196 241434
rect 471876 234434 472196 241198
rect 471876 234198 471918 234434
rect 472154 234198 472196 234434
rect 471876 227434 472196 234198
rect 471876 227198 471918 227434
rect 472154 227198 472196 227434
rect 471876 220434 472196 227198
rect 471876 220198 471918 220434
rect 472154 220198 472196 220434
rect 471876 213434 472196 220198
rect 471876 213198 471918 213434
rect 472154 213198 472196 213434
rect 471876 206434 472196 213198
rect 471876 206198 471918 206434
rect 472154 206198 472196 206434
rect 471876 199434 472196 206198
rect 471876 199198 471918 199434
rect 472154 199198 472196 199434
rect 471876 192434 472196 199198
rect 471876 192198 471918 192434
rect 472154 192198 472196 192434
rect 471876 185434 472196 192198
rect 471876 185198 471918 185434
rect 472154 185198 472196 185434
rect 471876 178434 472196 185198
rect 471876 178198 471918 178434
rect 472154 178198 472196 178434
rect 471876 171434 472196 178198
rect 471876 171198 471918 171434
rect 472154 171198 472196 171434
rect 471876 164434 472196 171198
rect 471876 164198 471918 164434
rect 472154 164198 472196 164434
rect 471876 157434 472196 164198
rect 471876 157198 471918 157434
rect 472154 157198 472196 157434
rect 471876 150434 472196 157198
rect 471876 150198 471918 150434
rect 472154 150198 472196 150434
rect 471876 143434 472196 150198
rect 471876 143198 471918 143434
rect 472154 143198 472196 143434
rect 471876 136434 472196 143198
rect 471876 136198 471918 136434
rect 472154 136198 472196 136434
rect 471876 129434 472196 136198
rect 471876 129198 471918 129434
rect 472154 129198 472196 129434
rect 471876 122434 472196 129198
rect 471876 122198 471918 122434
rect 472154 122198 472196 122434
rect 471876 115434 472196 122198
rect 471876 115198 471918 115434
rect 472154 115198 472196 115434
rect 471876 108434 472196 115198
rect 471876 108198 471918 108434
rect 472154 108198 472196 108434
rect 471876 101434 472196 108198
rect 471876 101198 471918 101434
rect 472154 101198 472196 101434
rect 471876 94434 472196 101198
rect 471876 94198 471918 94434
rect 472154 94198 472196 94434
rect 471876 87434 472196 94198
rect 471876 87198 471918 87434
rect 472154 87198 472196 87434
rect 471876 80434 472196 87198
rect 471876 80198 471918 80434
rect 472154 80198 472196 80434
rect 471876 73434 472196 80198
rect 471876 73198 471918 73434
rect 472154 73198 472196 73434
rect 471876 66434 472196 73198
rect 471876 66198 471918 66434
rect 472154 66198 472196 66434
rect 471876 59434 472196 66198
rect 471876 59198 471918 59434
rect 472154 59198 472196 59434
rect 471876 52434 472196 59198
rect 471876 52198 471918 52434
rect 472154 52198 472196 52434
rect 471876 45434 472196 52198
rect 471876 45198 471918 45434
rect 472154 45198 472196 45434
rect 471876 38434 472196 45198
rect 471876 38198 471918 38434
rect 472154 38198 472196 38434
rect 471876 31434 472196 38198
rect 471876 31198 471918 31434
rect 472154 31198 472196 31434
rect 471876 24434 472196 31198
rect 471876 24198 471918 24434
rect 472154 24198 472196 24434
rect 471876 17434 472196 24198
rect 471876 17198 471918 17434
rect 472154 17198 472196 17434
rect 471876 10434 472196 17198
rect 471876 10198 471918 10434
rect 472154 10198 472196 10434
rect 471876 3434 472196 10198
rect 471876 3198 471918 3434
rect 472154 3198 472196 3434
rect 471876 -1706 472196 3198
rect 471876 -1942 471918 -1706
rect 472154 -1942 472196 -1706
rect 471876 -2026 472196 -1942
rect 471876 -2262 471918 -2026
rect 472154 -2262 472196 -2026
rect 471876 -2294 472196 -2262
rect 477144 705238 477464 706230
rect 477144 705002 477186 705238
rect 477422 705002 477464 705238
rect 477144 704918 477464 705002
rect 477144 704682 477186 704918
rect 477422 704682 477464 704918
rect 477144 695494 477464 704682
rect 477144 695258 477186 695494
rect 477422 695258 477464 695494
rect 477144 688494 477464 695258
rect 477144 688258 477186 688494
rect 477422 688258 477464 688494
rect 477144 681494 477464 688258
rect 477144 681258 477186 681494
rect 477422 681258 477464 681494
rect 477144 674494 477464 681258
rect 477144 674258 477186 674494
rect 477422 674258 477464 674494
rect 477144 667494 477464 674258
rect 477144 667258 477186 667494
rect 477422 667258 477464 667494
rect 477144 660494 477464 667258
rect 477144 660258 477186 660494
rect 477422 660258 477464 660494
rect 477144 653494 477464 660258
rect 477144 653258 477186 653494
rect 477422 653258 477464 653494
rect 477144 646494 477464 653258
rect 477144 646258 477186 646494
rect 477422 646258 477464 646494
rect 477144 639494 477464 646258
rect 477144 639258 477186 639494
rect 477422 639258 477464 639494
rect 477144 632494 477464 639258
rect 477144 632258 477186 632494
rect 477422 632258 477464 632494
rect 477144 625494 477464 632258
rect 477144 625258 477186 625494
rect 477422 625258 477464 625494
rect 477144 618494 477464 625258
rect 477144 618258 477186 618494
rect 477422 618258 477464 618494
rect 477144 611494 477464 618258
rect 477144 611258 477186 611494
rect 477422 611258 477464 611494
rect 477144 604494 477464 611258
rect 477144 604258 477186 604494
rect 477422 604258 477464 604494
rect 477144 597494 477464 604258
rect 477144 597258 477186 597494
rect 477422 597258 477464 597494
rect 477144 590494 477464 597258
rect 477144 590258 477186 590494
rect 477422 590258 477464 590494
rect 477144 583494 477464 590258
rect 477144 583258 477186 583494
rect 477422 583258 477464 583494
rect 477144 576494 477464 583258
rect 477144 576258 477186 576494
rect 477422 576258 477464 576494
rect 477144 569494 477464 576258
rect 477144 569258 477186 569494
rect 477422 569258 477464 569494
rect 477144 562494 477464 569258
rect 477144 562258 477186 562494
rect 477422 562258 477464 562494
rect 477144 555494 477464 562258
rect 477144 555258 477186 555494
rect 477422 555258 477464 555494
rect 477144 548494 477464 555258
rect 477144 548258 477186 548494
rect 477422 548258 477464 548494
rect 477144 541494 477464 548258
rect 477144 541258 477186 541494
rect 477422 541258 477464 541494
rect 477144 534494 477464 541258
rect 477144 534258 477186 534494
rect 477422 534258 477464 534494
rect 477144 527494 477464 534258
rect 477144 527258 477186 527494
rect 477422 527258 477464 527494
rect 477144 520494 477464 527258
rect 477144 520258 477186 520494
rect 477422 520258 477464 520494
rect 477144 513494 477464 520258
rect 477144 513258 477186 513494
rect 477422 513258 477464 513494
rect 477144 506494 477464 513258
rect 477144 506258 477186 506494
rect 477422 506258 477464 506494
rect 477144 499494 477464 506258
rect 477144 499258 477186 499494
rect 477422 499258 477464 499494
rect 477144 492494 477464 499258
rect 477144 492258 477186 492494
rect 477422 492258 477464 492494
rect 477144 485494 477464 492258
rect 477144 485258 477186 485494
rect 477422 485258 477464 485494
rect 477144 478494 477464 485258
rect 477144 478258 477186 478494
rect 477422 478258 477464 478494
rect 477144 471494 477464 478258
rect 477144 471258 477186 471494
rect 477422 471258 477464 471494
rect 477144 464494 477464 471258
rect 477144 464258 477186 464494
rect 477422 464258 477464 464494
rect 477144 457494 477464 464258
rect 477144 457258 477186 457494
rect 477422 457258 477464 457494
rect 477144 450494 477464 457258
rect 477144 450258 477186 450494
rect 477422 450258 477464 450494
rect 477144 443494 477464 450258
rect 477144 443258 477186 443494
rect 477422 443258 477464 443494
rect 477144 436494 477464 443258
rect 477144 436258 477186 436494
rect 477422 436258 477464 436494
rect 477144 429494 477464 436258
rect 477144 429258 477186 429494
rect 477422 429258 477464 429494
rect 477144 422494 477464 429258
rect 477144 422258 477186 422494
rect 477422 422258 477464 422494
rect 477144 415494 477464 422258
rect 477144 415258 477186 415494
rect 477422 415258 477464 415494
rect 477144 408494 477464 415258
rect 477144 408258 477186 408494
rect 477422 408258 477464 408494
rect 477144 401494 477464 408258
rect 477144 401258 477186 401494
rect 477422 401258 477464 401494
rect 477144 394494 477464 401258
rect 477144 394258 477186 394494
rect 477422 394258 477464 394494
rect 477144 387494 477464 394258
rect 477144 387258 477186 387494
rect 477422 387258 477464 387494
rect 477144 380494 477464 387258
rect 477144 380258 477186 380494
rect 477422 380258 477464 380494
rect 477144 373494 477464 380258
rect 477144 373258 477186 373494
rect 477422 373258 477464 373494
rect 477144 366494 477464 373258
rect 477144 366258 477186 366494
rect 477422 366258 477464 366494
rect 477144 359494 477464 366258
rect 477144 359258 477186 359494
rect 477422 359258 477464 359494
rect 477144 352494 477464 359258
rect 477144 352258 477186 352494
rect 477422 352258 477464 352494
rect 477144 345494 477464 352258
rect 477144 345258 477186 345494
rect 477422 345258 477464 345494
rect 477144 338494 477464 345258
rect 477144 338258 477186 338494
rect 477422 338258 477464 338494
rect 477144 331494 477464 338258
rect 477144 331258 477186 331494
rect 477422 331258 477464 331494
rect 477144 324494 477464 331258
rect 477144 324258 477186 324494
rect 477422 324258 477464 324494
rect 477144 317494 477464 324258
rect 477144 317258 477186 317494
rect 477422 317258 477464 317494
rect 477144 310494 477464 317258
rect 477144 310258 477186 310494
rect 477422 310258 477464 310494
rect 477144 303494 477464 310258
rect 477144 303258 477186 303494
rect 477422 303258 477464 303494
rect 477144 296494 477464 303258
rect 477144 296258 477186 296494
rect 477422 296258 477464 296494
rect 477144 289494 477464 296258
rect 477144 289258 477186 289494
rect 477422 289258 477464 289494
rect 477144 282494 477464 289258
rect 477144 282258 477186 282494
rect 477422 282258 477464 282494
rect 477144 275494 477464 282258
rect 477144 275258 477186 275494
rect 477422 275258 477464 275494
rect 477144 268494 477464 275258
rect 477144 268258 477186 268494
rect 477422 268258 477464 268494
rect 477144 261494 477464 268258
rect 477144 261258 477186 261494
rect 477422 261258 477464 261494
rect 477144 254494 477464 261258
rect 477144 254258 477186 254494
rect 477422 254258 477464 254494
rect 477144 247494 477464 254258
rect 477144 247258 477186 247494
rect 477422 247258 477464 247494
rect 477144 240494 477464 247258
rect 477144 240258 477186 240494
rect 477422 240258 477464 240494
rect 477144 233494 477464 240258
rect 477144 233258 477186 233494
rect 477422 233258 477464 233494
rect 477144 226494 477464 233258
rect 477144 226258 477186 226494
rect 477422 226258 477464 226494
rect 477144 219494 477464 226258
rect 477144 219258 477186 219494
rect 477422 219258 477464 219494
rect 477144 212494 477464 219258
rect 477144 212258 477186 212494
rect 477422 212258 477464 212494
rect 477144 205494 477464 212258
rect 477144 205258 477186 205494
rect 477422 205258 477464 205494
rect 477144 198494 477464 205258
rect 477144 198258 477186 198494
rect 477422 198258 477464 198494
rect 477144 191494 477464 198258
rect 477144 191258 477186 191494
rect 477422 191258 477464 191494
rect 477144 184494 477464 191258
rect 477144 184258 477186 184494
rect 477422 184258 477464 184494
rect 477144 177494 477464 184258
rect 477144 177258 477186 177494
rect 477422 177258 477464 177494
rect 477144 170494 477464 177258
rect 477144 170258 477186 170494
rect 477422 170258 477464 170494
rect 477144 163494 477464 170258
rect 477144 163258 477186 163494
rect 477422 163258 477464 163494
rect 477144 156494 477464 163258
rect 477144 156258 477186 156494
rect 477422 156258 477464 156494
rect 477144 149494 477464 156258
rect 477144 149258 477186 149494
rect 477422 149258 477464 149494
rect 477144 142494 477464 149258
rect 477144 142258 477186 142494
rect 477422 142258 477464 142494
rect 477144 135494 477464 142258
rect 477144 135258 477186 135494
rect 477422 135258 477464 135494
rect 477144 128494 477464 135258
rect 477144 128258 477186 128494
rect 477422 128258 477464 128494
rect 477144 121494 477464 128258
rect 477144 121258 477186 121494
rect 477422 121258 477464 121494
rect 477144 114494 477464 121258
rect 477144 114258 477186 114494
rect 477422 114258 477464 114494
rect 477144 107494 477464 114258
rect 477144 107258 477186 107494
rect 477422 107258 477464 107494
rect 477144 100494 477464 107258
rect 477144 100258 477186 100494
rect 477422 100258 477464 100494
rect 477144 93494 477464 100258
rect 477144 93258 477186 93494
rect 477422 93258 477464 93494
rect 477144 86494 477464 93258
rect 477144 86258 477186 86494
rect 477422 86258 477464 86494
rect 477144 79494 477464 86258
rect 477144 79258 477186 79494
rect 477422 79258 477464 79494
rect 477144 72494 477464 79258
rect 477144 72258 477186 72494
rect 477422 72258 477464 72494
rect 477144 65494 477464 72258
rect 477144 65258 477186 65494
rect 477422 65258 477464 65494
rect 477144 58494 477464 65258
rect 477144 58258 477186 58494
rect 477422 58258 477464 58494
rect 477144 51494 477464 58258
rect 477144 51258 477186 51494
rect 477422 51258 477464 51494
rect 477144 44494 477464 51258
rect 477144 44258 477186 44494
rect 477422 44258 477464 44494
rect 477144 37494 477464 44258
rect 477144 37258 477186 37494
rect 477422 37258 477464 37494
rect 477144 30494 477464 37258
rect 477144 30258 477186 30494
rect 477422 30258 477464 30494
rect 477144 23494 477464 30258
rect 477144 23258 477186 23494
rect 477422 23258 477464 23494
rect 477144 16494 477464 23258
rect 477144 16258 477186 16494
rect 477422 16258 477464 16494
rect 477144 9494 477464 16258
rect 477144 9258 477186 9494
rect 477422 9258 477464 9494
rect 477144 2494 477464 9258
rect 477144 2258 477186 2494
rect 477422 2258 477464 2494
rect 477144 -746 477464 2258
rect 477144 -982 477186 -746
rect 477422 -982 477464 -746
rect 477144 -1066 477464 -982
rect 477144 -1302 477186 -1066
rect 477422 -1302 477464 -1066
rect 477144 -2294 477464 -1302
rect 478876 706198 479196 706230
rect 478876 705962 478918 706198
rect 479154 705962 479196 706198
rect 478876 705878 479196 705962
rect 478876 705642 478918 705878
rect 479154 705642 479196 705878
rect 478876 696434 479196 705642
rect 478876 696198 478918 696434
rect 479154 696198 479196 696434
rect 478876 689434 479196 696198
rect 478876 689198 478918 689434
rect 479154 689198 479196 689434
rect 478876 682434 479196 689198
rect 478876 682198 478918 682434
rect 479154 682198 479196 682434
rect 478876 675434 479196 682198
rect 478876 675198 478918 675434
rect 479154 675198 479196 675434
rect 478876 668434 479196 675198
rect 478876 668198 478918 668434
rect 479154 668198 479196 668434
rect 478876 661434 479196 668198
rect 478876 661198 478918 661434
rect 479154 661198 479196 661434
rect 478876 654434 479196 661198
rect 478876 654198 478918 654434
rect 479154 654198 479196 654434
rect 478876 647434 479196 654198
rect 478876 647198 478918 647434
rect 479154 647198 479196 647434
rect 478876 640434 479196 647198
rect 478876 640198 478918 640434
rect 479154 640198 479196 640434
rect 478876 633434 479196 640198
rect 478876 633198 478918 633434
rect 479154 633198 479196 633434
rect 478876 626434 479196 633198
rect 478876 626198 478918 626434
rect 479154 626198 479196 626434
rect 478876 619434 479196 626198
rect 478876 619198 478918 619434
rect 479154 619198 479196 619434
rect 478876 612434 479196 619198
rect 478876 612198 478918 612434
rect 479154 612198 479196 612434
rect 478876 605434 479196 612198
rect 478876 605198 478918 605434
rect 479154 605198 479196 605434
rect 478876 598434 479196 605198
rect 478876 598198 478918 598434
rect 479154 598198 479196 598434
rect 478876 591434 479196 598198
rect 478876 591198 478918 591434
rect 479154 591198 479196 591434
rect 478876 584434 479196 591198
rect 478876 584198 478918 584434
rect 479154 584198 479196 584434
rect 478876 577434 479196 584198
rect 478876 577198 478918 577434
rect 479154 577198 479196 577434
rect 478876 570434 479196 577198
rect 478876 570198 478918 570434
rect 479154 570198 479196 570434
rect 478876 563434 479196 570198
rect 478876 563198 478918 563434
rect 479154 563198 479196 563434
rect 478876 556434 479196 563198
rect 478876 556198 478918 556434
rect 479154 556198 479196 556434
rect 478876 549434 479196 556198
rect 478876 549198 478918 549434
rect 479154 549198 479196 549434
rect 478876 542434 479196 549198
rect 478876 542198 478918 542434
rect 479154 542198 479196 542434
rect 478876 535434 479196 542198
rect 478876 535198 478918 535434
rect 479154 535198 479196 535434
rect 478876 528434 479196 535198
rect 478876 528198 478918 528434
rect 479154 528198 479196 528434
rect 478876 521434 479196 528198
rect 478876 521198 478918 521434
rect 479154 521198 479196 521434
rect 478876 514434 479196 521198
rect 478876 514198 478918 514434
rect 479154 514198 479196 514434
rect 478876 507434 479196 514198
rect 478876 507198 478918 507434
rect 479154 507198 479196 507434
rect 478876 500434 479196 507198
rect 478876 500198 478918 500434
rect 479154 500198 479196 500434
rect 478876 493434 479196 500198
rect 478876 493198 478918 493434
rect 479154 493198 479196 493434
rect 478876 486434 479196 493198
rect 478876 486198 478918 486434
rect 479154 486198 479196 486434
rect 478876 479434 479196 486198
rect 478876 479198 478918 479434
rect 479154 479198 479196 479434
rect 478876 472434 479196 479198
rect 478876 472198 478918 472434
rect 479154 472198 479196 472434
rect 478876 465434 479196 472198
rect 478876 465198 478918 465434
rect 479154 465198 479196 465434
rect 478876 458434 479196 465198
rect 478876 458198 478918 458434
rect 479154 458198 479196 458434
rect 478876 451434 479196 458198
rect 478876 451198 478918 451434
rect 479154 451198 479196 451434
rect 478876 444434 479196 451198
rect 478876 444198 478918 444434
rect 479154 444198 479196 444434
rect 478876 437434 479196 444198
rect 478876 437198 478918 437434
rect 479154 437198 479196 437434
rect 478876 430434 479196 437198
rect 478876 430198 478918 430434
rect 479154 430198 479196 430434
rect 478876 423434 479196 430198
rect 478876 423198 478918 423434
rect 479154 423198 479196 423434
rect 478876 416434 479196 423198
rect 478876 416198 478918 416434
rect 479154 416198 479196 416434
rect 478876 409434 479196 416198
rect 478876 409198 478918 409434
rect 479154 409198 479196 409434
rect 478876 402434 479196 409198
rect 478876 402198 478918 402434
rect 479154 402198 479196 402434
rect 478876 395434 479196 402198
rect 478876 395198 478918 395434
rect 479154 395198 479196 395434
rect 478876 388434 479196 395198
rect 478876 388198 478918 388434
rect 479154 388198 479196 388434
rect 478876 381434 479196 388198
rect 478876 381198 478918 381434
rect 479154 381198 479196 381434
rect 478876 374434 479196 381198
rect 478876 374198 478918 374434
rect 479154 374198 479196 374434
rect 478876 367434 479196 374198
rect 478876 367198 478918 367434
rect 479154 367198 479196 367434
rect 478876 360434 479196 367198
rect 478876 360198 478918 360434
rect 479154 360198 479196 360434
rect 478876 353434 479196 360198
rect 478876 353198 478918 353434
rect 479154 353198 479196 353434
rect 478876 346434 479196 353198
rect 478876 346198 478918 346434
rect 479154 346198 479196 346434
rect 478876 339434 479196 346198
rect 478876 339198 478918 339434
rect 479154 339198 479196 339434
rect 478876 332434 479196 339198
rect 478876 332198 478918 332434
rect 479154 332198 479196 332434
rect 478876 325434 479196 332198
rect 478876 325198 478918 325434
rect 479154 325198 479196 325434
rect 478876 318434 479196 325198
rect 478876 318198 478918 318434
rect 479154 318198 479196 318434
rect 478876 311434 479196 318198
rect 478876 311198 478918 311434
rect 479154 311198 479196 311434
rect 478876 304434 479196 311198
rect 478876 304198 478918 304434
rect 479154 304198 479196 304434
rect 478876 297434 479196 304198
rect 478876 297198 478918 297434
rect 479154 297198 479196 297434
rect 478876 290434 479196 297198
rect 478876 290198 478918 290434
rect 479154 290198 479196 290434
rect 478876 283434 479196 290198
rect 478876 283198 478918 283434
rect 479154 283198 479196 283434
rect 478876 276434 479196 283198
rect 478876 276198 478918 276434
rect 479154 276198 479196 276434
rect 478876 269434 479196 276198
rect 478876 269198 478918 269434
rect 479154 269198 479196 269434
rect 478876 262434 479196 269198
rect 478876 262198 478918 262434
rect 479154 262198 479196 262434
rect 478876 255434 479196 262198
rect 478876 255198 478918 255434
rect 479154 255198 479196 255434
rect 478876 248434 479196 255198
rect 478876 248198 478918 248434
rect 479154 248198 479196 248434
rect 478876 241434 479196 248198
rect 478876 241198 478918 241434
rect 479154 241198 479196 241434
rect 478876 234434 479196 241198
rect 478876 234198 478918 234434
rect 479154 234198 479196 234434
rect 478876 227434 479196 234198
rect 478876 227198 478918 227434
rect 479154 227198 479196 227434
rect 478876 220434 479196 227198
rect 478876 220198 478918 220434
rect 479154 220198 479196 220434
rect 478876 213434 479196 220198
rect 478876 213198 478918 213434
rect 479154 213198 479196 213434
rect 478876 206434 479196 213198
rect 478876 206198 478918 206434
rect 479154 206198 479196 206434
rect 478876 199434 479196 206198
rect 478876 199198 478918 199434
rect 479154 199198 479196 199434
rect 478876 192434 479196 199198
rect 478876 192198 478918 192434
rect 479154 192198 479196 192434
rect 478876 185434 479196 192198
rect 478876 185198 478918 185434
rect 479154 185198 479196 185434
rect 478876 178434 479196 185198
rect 478876 178198 478918 178434
rect 479154 178198 479196 178434
rect 478876 171434 479196 178198
rect 478876 171198 478918 171434
rect 479154 171198 479196 171434
rect 478876 164434 479196 171198
rect 478876 164198 478918 164434
rect 479154 164198 479196 164434
rect 478876 157434 479196 164198
rect 478876 157198 478918 157434
rect 479154 157198 479196 157434
rect 478876 150434 479196 157198
rect 478876 150198 478918 150434
rect 479154 150198 479196 150434
rect 478876 143434 479196 150198
rect 478876 143198 478918 143434
rect 479154 143198 479196 143434
rect 478876 136434 479196 143198
rect 478876 136198 478918 136434
rect 479154 136198 479196 136434
rect 478876 129434 479196 136198
rect 478876 129198 478918 129434
rect 479154 129198 479196 129434
rect 478876 122434 479196 129198
rect 478876 122198 478918 122434
rect 479154 122198 479196 122434
rect 478876 115434 479196 122198
rect 478876 115198 478918 115434
rect 479154 115198 479196 115434
rect 478876 108434 479196 115198
rect 478876 108198 478918 108434
rect 479154 108198 479196 108434
rect 478876 101434 479196 108198
rect 478876 101198 478918 101434
rect 479154 101198 479196 101434
rect 478876 94434 479196 101198
rect 478876 94198 478918 94434
rect 479154 94198 479196 94434
rect 478876 87434 479196 94198
rect 478876 87198 478918 87434
rect 479154 87198 479196 87434
rect 478876 80434 479196 87198
rect 478876 80198 478918 80434
rect 479154 80198 479196 80434
rect 478876 73434 479196 80198
rect 478876 73198 478918 73434
rect 479154 73198 479196 73434
rect 478876 66434 479196 73198
rect 478876 66198 478918 66434
rect 479154 66198 479196 66434
rect 478876 59434 479196 66198
rect 478876 59198 478918 59434
rect 479154 59198 479196 59434
rect 478876 52434 479196 59198
rect 478876 52198 478918 52434
rect 479154 52198 479196 52434
rect 478876 45434 479196 52198
rect 478876 45198 478918 45434
rect 479154 45198 479196 45434
rect 478876 38434 479196 45198
rect 478876 38198 478918 38434
rect 479154 38198 479196 38434
rect 478876 31434 479196 38198
rect 478876 31198 478918 31434
rect 479154 31198 479196 31434
rect 478876 24434 479196 31198
rect 478876 24198 478918 24434
rect 479154 24198 479196 24434
rect 478876 17434 479196 24198
rect 478876 17198 478918 17434
rect 479154 17198 479196 17434
rect 478876 10434 479196 17198
rect 478876 10198 478918 10434
rect 479154 10198 479196 10434
rect 478876 3434 479196 10198
rect 478876 3198 478918 3434
rect 479154 3198 479196 3434
rect 478876 -1706 479196 3198
rect 478876 -1942 478918 -1706
rect 479154 -1942 479196 -1706
rect 478876 -2026 479196 -1942
rect 478876 -2262 478918 -2026
rect 479154 -2262 479196 -2026
rect 478876 -2294 479196 -2262
rect 484144 705238 484464 706230
rect 484144 705002 484186 705238
rect 484422 705002 484464 705238
rect 484144 704918 484464 705002
rect 484144 704682 484186 704918
rect 484422 704682 484464 704918
rect 484144 695494 484464 704682
rect 484144 695258 484186 695494
rect 484422 695258 484464 695494
rect 484144 688494 484464 695258
rect 484144 688258 484186 688494
rect 484422 688258 484464 688494
rect 484144 681494 484464 688258
rect 484144 681258 484186 681494
rect 484422 681258 484464 681494
rect 484144 674494 484464 681258
rect 484144 674258 484186 674494
rect 484422 674258 484464 674494
rect 484144 667494 484464 674258
rect 484144 667258 484186 667494
rect 484422 667258 484464 667494
rect 484144 660494 484464 667258
rect 484144 660258 484186 660494
rect 484422 660258 484464 660494
rect 484144 653494 484464 660258
rect 484144 653258 484186 653494
rect 484422 653258 484464 653494
rect 484144 646494 484464 653258
rect 484144 646258 484186 646494
rect 484422 646258 484464 646494
rect 484144 639494 484464 646258
rect 484144 639258 484186 639494
rect 484422 639258 484464 639494
rect 484144 632494 484464 639258
rect 484144 632258 484186 632494
rect 484422 632258 484464 632494
rect 484144 625494 484464 632258
rect 484144 625258 484186 625494
rect 484422 625258 484464 625494
rect 484144 618494 484464 625258
rect 484144 618258 484186 618494
rect 484422 618258 484464 618494
rect 484144 611494 484464 618258
rect 484144 611258 484186 611494
rect 484422 611258 484464 611494
rect 484144 604494 484464 611258
rect 484144 604258 484186 604494
rect 484422 604258 484464 604494
rect 484144 597494 484464 604258
rect 484144 597258 484186 597494
rect 484422 597258 484464 597494
rect 484144 590494 484464 597258
rect 484144 590258 484186 590494
rect 484422 590258 484464 590494
rect 484144 583494 484464 590258
rect 484144 583258 484186 583494
rect 484422 583258 484464 583494
rect 484144 576494 484464 583258
rect 484144 576258 484186 576494
rect 484422 576258 484464 576494
rect 484144 569494 484464 576258
rect 484144 569258 484186 569494
rect 484422 569258 484464 569494
rect 484144 562494 484464 569258
rect 484144 562258 484186 562494
rect 484422 562258 484464 562494
rect 484144 555494 484464 562258
rect 484144 555258 484186 555494
rect 484422 555258 484464 555494
rect 484144 548494 484464 555258
rect 484144 548258 484186 548494
rect 484422 548258 484464 548494
rect 484144 541494 484464 548258
rect 484144 541258 484186 541494
rect 484422 541258 484464 541494
rect 484144 534494 484464 541258
rect 484144 534258 484186 534494
rect 484422 534258 484464 534494
rect 484144 527494 484464 534258
rect 484144 527258 484186 527494
rect 484422 527258 484464 527494
rect 484144 520494 484464 527258
rect 484144 520258 484186 520494
rect 484422 520258 484464 520494
rect 484144 513494 484464 520258
rect 484144 513258 484186 513494
rect 484422 513258 484464 513494
rect 484144 506494 484464 513258
rect 484144 506258 484186 506494
rect 484422 506258 484464 506494
rect 484144 499494 484464 506258
rect 484144 499258 484186 499494
rect 484422 499258 484464 499494
rect 484144 492494 484464 499258
rect 484144 492258 484186 492494
rect 484422 492258 484464 492494
rect 484144 485494 484464 492258
rect 484144 485258 484186 485494
rect 484422 485258 484464 485494
rect 484144 478494 484464 485258
rect 484144 478258 484186 478494
rect 484422 478258 484464 478494
rect 484144 471494 484464 478258
rect 484144 471258 484186 471494
rect 484422 471258 484464 471494
rect 484144 464494 484464 471258
rect 484144 464258 484186 464494
rect 484422 464258 484464 464494
rect 484144 457494 484464 464258
rect 484144 457258 484186 457494
rect 484422 457258 484464 457494
rect 484144 450494 484464 457258
rect 484144 450258 484186 450494
rect 484422 450258 484464 450494
rect 484144 443494 484464 450258
rect 484144 443258 484186 443494
rect 484422 443258 484464 443494
rect 484144 436494 484464 443258
rect 484144 436258 484186 436494
rect 484422 436258 484464 436494
rect 484144 429494 484464 436258
rect 484144 429258 484186 429494
rect 484422 429258 484464 429494
rect 484144 422494 484464 429258
rect 484144 422258 484186 422494
rect 484422 422258 484464 422494
rect 484144 415494 484464 422258
rect 484144 415258 484186 415494
rect 484422 415258 484464 415494
rect 484144 408494 484464 415258
rect 484144 408258 484186 408494
rect 484422 408258 484464 408494
rect 484144 401494 484464 408258
rect 484144 401258 484186 401494
rect 484422 401258 484464 401494
rect 484144 394494 484464 401258
rect 484144 394258 484186 394494
rect 484422 394258 484464 394494
rect 484144 387494 484464 394258
rect 484144 387258 484186 387494
rect 484422 387258 484464 387494
rect 484144 380494 484464 387258
rect 484144 380258 484186 380494
rect 484422 380258 484464 380494
rect 484144 373494 484464 380258
rect 484144 373258 484186 373494
rect 484422 373258 484464 373494
rect 484144 366494 484464 373258
rect 484144 366258 484186 366494
rect 484422 366258 484464 366494
rect 484144 359494 484464 366258
rect 484144 359258 484186 359494
rect 484422 359258 484464 359494
rect 484144 352494 484464 359258
rect 484144 352258 484186 352494
rect 484422 352258 484464 352494
rect 484144 345494 484464 352258
rect 484144 345258 484186 345494
rect 484422 345258 484464 345494
rect 484144 338494 484464 345258
rect 484144 338258 484186 338494
rect 484422 338258 484464 338494
rect 484144 331494 484464 338258
rect 484144 331258 484186 331494
rect 484422 331258 484464 331494
rect 484144 324494 484464 331258
rect 484144 324258 484186 324494
rect 484422 324258 484464 324494
rect 484144 317494 484464 324258
rect 484144 317258 484186 317494
rect 484422 317258 484464 317494
rect 484144 310494 484464 317258
rect 484144 310258 484186 310494
rect 484422 310258 484464 310494
rect 484144 303494 484464 310258
rect 484144 303258 484186 303494
rect 484422 303258 484464 303494
rect 484144 296494 484464 303258
rect 484144 296258 484186 296494
rect 484422 296258 484464 296494
rect 484144 289494 484464 296258
rect 484144 289258 484186 289494
rect 484422 289258 484464 289494
rect 484144 282494 484464 289258
rect 484144 282258 484186 282494
rect 484422 282258 484464 282494
rect 484144 275494 484464 282258
rect 484144 275258 484186 275494
rect 484422 275258 484464 275494
rect 484144 268494 484464 275258
rect 484144 268258 484186 268494
rect 484422 268258 484464 268494
rect 484144 261494 484464 268258
rect 484144 261258 484186 261494
rect 484422 261258 484464 261494
rect 484144 254494 484464 261258
rect 484144 254258 484186 254494
rect 484422 254258 484464 254494
rect 484144 247494 484464 254258
rect 484144 247258 484186 247494
rect 484422 247258 484464 247494
rect 484144 240494 484464 247258
rect 484144 240258 484186 240494
rect 484422 240258 484464 240494
rect 484144 233494 484464 240258
rect 484144 233258 484186 233494
rect 484422 233258 484464 233494
rect 484144 226494 484464 233258
rect 484144 226258 484186 226494
rect 484422 226258 484464 226494
rect 484144 219494 484464 226258
rect 484144 219258 484186 219494
rect 484422 219258 484464 219494
rect 484144 212494 484464 219258
rect 484144 212258 484186 212494
rect 484422 212258 484464 212494
rect 484144 205494 484464 212258
rect 484144 205258 484186 205494
rect 484422 205258 484464 205494
rect 484144 198494 484464 205258
rect 484144 198258 484186 198494
rect 484422 198258 484464 198494
rect 484144 191494 484464 198258
rect 484144 191258 484186 191494
rect 484422 191258 484464 191494
rect 484144 184494 484464 191258
rect 484144 184258 484186 184494
rect 484422 184258 484464 184494
rect 484144 177494 484464 184258
rect 484144 177258 484186 177494
rect 484422 177258 484464 177494
rect 484144 170494 484464 177258
rect 484144 170258 484186 170494
rect 484422 170258 484464 170494
rect 484144 163494 484464 170258
rect 484144 163258 484186 163494
rect 484422 163258 484464 163494
rect 484144 156494 484464 163258
rect 484144 156258 484186 156494
rect 484422 156258 484464 156494
rect 484144 149494 484464 156258
rect 484144 149258 484186 149494
rect 484422 149258 484464 149494
rect 484144 142494 484464 149258
rect 484144 142258 484186 142494
rect 484422 142258 484464 142494
rect 484144 135494 484464 142258
rect 484144 135258 484186 135494
rect 484422 135258 484464 135494
rect 484144 128494 484464 135258
rect 484144 128258 484186 128494
rect 484422 128258 484464 128494
rect 484144 121494 484464 128258
rect 484144 121258 484186 121494
rect 484422 121258 484464 121494
rect 484144 114494 484464 121258
rect 484144 114258 484186 114494
rect 484422 114258 484464 114494
rect 484144 107494 484464 114258
rect 484144 107258 484186 107494
rect 484422 107258 484464 107494
rect 484144 100494 484464 107258
rect 484144 100258 484186 100494
rect 484422 100258 484464 100494
rect 484144 93494 484464 100258
rect 484144 93258 484186 93494
rect 484422 93258 484464 93494
rect 484144 86494 484464 93258
rect 484144 86258 484186 86494
rect 484422 86258 484464 86494
rect 484144 79494 484464 86258
rect 484144 79258 484186 79494
rect 484422 79258 484464 79494
rect 484144 72494 484464 79258
rect 484144 72258 484186 72494
rect 484422 72258 484464 72494
rect 484144 65494 484464 72258
rect 484144 65258 484186 65494
rect 484422 65258 484464 65494
rect 484144 58494 484464 65258
rect 484144 58258 484186 58494
rect 484422 58258 484464 58494
rect 484144 51494 484464 58258
rect 484144 51258 484186 51494
rect 484422 51258 484464 51494
rect 484144 44494 484464 51258
rect 484144 44258 484186 44494
rect 484422 44258 484464 44494
rect 484144 37494 484464 44258
rect 484144 37258 484186 37494
rect 484422 37258 484464 37494
rect 484144 30494 484464 37258
rect 484144 30258 484186 30494
rect 484422 30258 484464 30494
rect 484144 23494 484464 30258
rect 484144 23258 484186 23494
rect 484422 23258 484464 23494
rect 484144 16494 484464 23258
rect 484144 16258 484186 16494
rect 484422 16258 484464 16494
rect 484144 9494 484464 16258
rect 484144 9258 484186 9494
rect 484422 9258 484464 9494
rect 484144 2494 484464 9258
rect 484144 2258 484186 2494
rect 484422 2258 484464 2494
rect 484144 -746 484464 2258
rect 484144 -982 484186 -746
rect 484422 -982 484464 -746
rect 484144 -1066 484464 -982
rect 484144 -1302 484186 -1066
rect 484422 -1302 484464 -1066
rect 484144 -2294 484464 -1302
rect 485876 706198 486196 706230
rect 485876 705962 485918 706198
rect 486154 705962 486196 706198
rect 485876 705878 486196 705962
rect 485876 705642 485918 705878
rect 486154 705642 486196 705878
rect 485876 696434 486196 705642
rect 485876 696198 485918 696434
rect 486154 696198 486196 696434
rect 485876 689434 486196 696198
rect 485876 689198 485918 689434
rect 486154 689198 486196 689434
rect 485876 682434 486196 689198
rect 485876 682198 485918 682434
rect 486154 682198 486196 682434
rect 485876 675434 486196 682198
rect 485876 675198 485918 675434
rect 486154 675198 486196 675434
rect 485876 668434 486196 675198
rect 485876 668198 485918 668434
rect 486154 668198 486196 668434
rect 485876 661434 486196 668198
rect 485876 661198 485918 661434
rect 486154 661198 486196 661434
rect 485876 654434 486196 661198
rect 485876 654198 485918 654434
rect 486154 654198 486196 654434
rect 485876 647434 486196 654198
rect 485876 647198 485918 647434
rect 486154 647198 486196 647434
rect 485876 640434 486196 647198
rect 485876 640198 485918 640434
rect 486154 640198 486196 640434
rect 485876 633434 486196 640198
rect 485876 633198 485918 633434
rect 486154 633198 486196 633434
rect 485876 626434 486196 633198
rect 485876 626198 485918 626434
rect 486154 626198 486196 626434
rect 485876 619434 486196 626198
rect 485876 619198 485918 619434
rect 486154 619198 486196 619434
rect 485876 612434 486196 619198
rect 485876 612198 485918 612434
rect 486154 612198 486196 612434
rect 485876 605434 486196 612198
rect 485876 605198 485918 605434
rect 486154 605198 486196 605434
rect 485876 598434 486196 605198
rect 485876 598198 485918 598434
rect 486154 598198 486196 598434
rect 485876 591434 486196 598198
rect 485876 591198 485918 591434
rect 486154 591198 486196 591434
rect 485876 584434 486196 591198
rect 485876 584198 485918 584434
rect 486154 584198 486196 584434
rect 485876 577434 486196 584198
rect 485876 577198 485918 577434
rect 486154 577198 486196 577434
rect 485876 570434 486196 577198
rect 485876 570198 485918 570434
rect 486154 570198 486196 570434
rect 485876 563434 486196 570198
rect 485876 563198 485918 563434
rect 486154 563198 486196 563434
rect 485876 556434 486196 563198
rect 485876 556198 485918 556434
rect 486154 556198 486196 556434
rect 485876 549434 486196 556198
rect 485876 549198 485918 549434
rect 486154 549198 486196 549434
rect 485876 542434 486196 549198
rect 485876 542198 485918 542434
rect 486154 542198 486196 542434
rect 485876 535434 486196 542198
rect 485876 535198 485918 535434
rect 486154 535198 486196 535434
rect 485876 528434 486196 535198
rect 485876 528198 485918 528434
rect 486154 528198 486196 528434
rect 485876 521434 486196 528198
rect 485876 521198 485918 521434
rect 486154 521198 486196 521434
rect 485876 514434 486196 521198
rect 485876 514198 485918 514434
rect 486154 514198 486196 514434
rect 485876 507434 486196 514198
rect 485876 507198 485918 507434
rect 486154 507198 486196 507434
rect 485876 500434 486196 507198
rect 485876 500198 485918 500434
rect 486154 500198 486196 500434
rect 485876 493434 486196 500198
rect 485876 493198 485918 493434
rect 486154 493198 486196 493434
rect 485876 486434 486196 493198
rect 485876 486198 485918 486434
rect 486154 486198 486196 486434
rect 485876 479434 486196 486198
rect 485876 479198 485918 479434
rect 486154 479198 486196 479434
rect 485876 472434 486196 479198
rect 485876 472198 485918 472434
rect 486154 472198 486196 472434
rect 485876 465434 486196 472198
rect 485876 465198 485918 465434
rect 486154 465198 486196 465434
rect 485876 458434 486196 465198
rect 485876 458198 485918 458434
rect 486154 458198 486196 458434
rect 485876 451434 486196 458198
rect 485876 451198 485918 451434
rect 486154 451198 486196 451434
rect 485876 444434 486196 451198
rect 485876 444198 485918 444434
rect 486154 444198 486196 444434
rect 485876 437434 486196 444198
rect 485876 437198 485918 437434
rect 486154 437198 486196 437434
rect 485876 430434 486196 437198
rect 485876 430198 485918 430434
rect 486154 430198 486196 430434
rect 485876 423434 486196 430198
rect 485876 423198 485918 423434
rect 486154 423198 486196 423434
rect 485876 416434 486196 423198
rect 485876 416198 485918 416434
rect 486154 416198 486196 416434
rect 485876 409434 486196 416198
rect 485876 409198 485918 409434
rect 486154 409198 486196 409434
rect 485876 402434 486196 409198
rect 485876 402198 485918 402434
rect 486154 402198 486196 402434
rect 485876 395434 486196 402198
rect 485876 395198 485918 395434
rect 486154 395198 486196 395434
rect 485876 388434 486196 395198
rect 485876 388198 485918 388434
rect 486154 388198 486196 388434
rect 485876 381434 486196 388198
rect 485876 381198 485918 381434
rect 486154 381198 486196 381434
rect 485876 374434 486196 381198
rect 485876 374198 485918 374434
rect 486154 374198 486196 374434
rect 485876 367434 486196 374198
rect 485876 367198 485918 367434
rect 486154 367198 486196 367434
rect 485876 360434 486196 367198
rect 485876 360198 485918 360434
rect 486154 360198 486196 360434
rect 485876 353434 486196 360198
rect 485876 353198 485918 353434
rect 486154 353198 486196 353434
rect 485876 346434 486196 353198
rect 485876 346198 485918 346434
rect 486154 346198 486196 346434
rect 485876 339434 486196 346198
rect 485876 339198 485918 339434
rect 486154 339198 486196 339434
rect 485876 332434 486196 339198
rect 485876 332198 485918 332434
rect 486154 332198 486196 332434
rect 485876 325434 486196 332198
rect 485876 325198 485918 325434
rect 486154 325198 486196 325434
rect 485876 318434 486196 325198
rect 485876 318198 485918 318434
rect 486154 318198 486196 318434
rect 485876 311434 486196 318198
rect 485876 311198 485918 311434
rect 486154 311198 486196 311434
rect 485876 304434 486196 311198
rect 485876 304198 485918 304434
rect 486154 304198 486196 304434
rect 485876 297434 486196 304198
rect 485876 297198 485918 297434
rect 486154 297198 486196 297434
rect 485876 290434 486196 297198
rect 485876 290198 485918 290434
rect 486154 290198 486196 290434
rect 485876 283434 486196 290198
rect 485876 283198 485918 283434
rect 486154 283198 486196 283434
rect 485876 276434 486196 283198
rect 485876 276198 485918 276434
rect 486154 276198 486196 276434
rect 485876 269434 486196 276198
rect 485876 269198 485918 269434
rect 486154 269198 486196 269434
rect 485876 262434 486196 269198
rect 485876 262198 485918 262434
rect 486154 262198 486196 262434
rect 485876 255434 486196 262198
rect 485876 255198 485918 255434
rect 486154 255198 486196 255434
rect 485876 248434 486196 255198
rect 485876 248198 485918 248434
rect 486154 248198 486196 248434
rect 485876 241434 486196 248198
rect 485876 241198 485918 241434
rect 486154 241198 486196 241434
rect 485876 234434 486196 241198
rect 485876 234198 485918 234434
rect 486154 234198 486196 234434
rect 485876 227434 486196 234198
rect 485876 227198 485918 227434
rect 486154 227198 486196 227434
rect 485876 220434 486196 227198
rect 485876 220198 485918 220434
rect 486154 220198 486196 220434
rect 485876 213434 486196 220198
rect 485876 213198 485918 213434
rect 486154 213198 486196 213434
rect 485876 206434 486196 213198
rect 485876 206198 485918 206434
rect 486154 206198 486196 206434
rect 485876 199434 486196 206198
rect 485876 199198 485918 199434
rect 486154 199198 486196 199434
rect 485876 192434 486196 199198
rect 485876 192198 485918 192434
rect 486154 192198 486196 192434
rect 485876 185434 486196 192198
rect 485876 185198 485918 185434
rect 486154 185198 486196 185434
rect 485876 178434 486196 185198
rect 485876 178198 485918 178434
rect 486154 178198 486196 178434
rect 485876 171434 486196 178198
rect 485876 171198 485918 171434
rect 486154 171198 486196 171434
rect 485876 164434 486196 171198
rect 485876 164198 485918 164434
rect 486154 164198 486196 164434
rect 485876 157434 486196 164198
rect 485876 157198 485918 157434
rect 486154 157198 486196 157434
rect 485876 150434 486196 157198
rect 485876 150198 485918 150434
rect 486154 150198 486196 150434
rect 485876 143434 486196 150198
rect 485876 143198 485918 143434
rect 486154 143198 486196 143434
rect 485876 136434 486196 143198
rect 485876 136198 485918 136434
rect 486154 136198 486196 136434
rect 485876 129434 486196 136198
rect 485876 129198 485918 129434
rect 486154 129198 486196 129434
rect 485876 122434 486196 129198
rect 485876 122198 485918 122434
rect 486154 122198 486196 122434
rect 485876 115434 486196 122198
rect 485876 115198 485918 115434
rect 486154 115198 486196 115434
rect 485876 108434 486196 115198
rect 485876 108198 485918 108434
rect 486154 108198 486196 108434
rect 485876 101434 486196 108198
rect 485876 101198 485918 101434
rect 486154 101198 486196 101434
rect 485876 94434 486196 101198
rect 485876 94198 485918 94434
rect 486154 94198 486196 94434
rect 485876 87434 486196 94198
rect 485876 87198 485918 87434
rect 486154 87198 486196 87434
rect 485876 80434 486196 87198
rect 485876 80198 485918 80434
rect 486154 80198 486196 80434
rect 485876 73434 486196 80198
rect 485876 73198 485918 73434
rect 486154 73198 486196 73434
rect 485876 66434 486196 73198
rect 485876 66198 485918 66434
rect 486154 66198 486196 66434
rect 485876 59434 486196 66198
rect 485876 59198 485918 59434
rect 486154 59198 486196 59434
rect 485876 52434 486196 59198
rect 485876 52198 485918 52434
rect 486154 52198 486196 52434
rect 485876 45434 486196 52198
rect 485876 45198 485918 45434
rect 486154 45198 486196 45434
rect 485876 38434 486196 45198
rect 485876 38198 485918 38434
rect 486154 38198 486196 38434
rect 485876 31434 486196 38198
rect 485876 31198 485918 31434
rect 486154 31198 486196 31434
rect 485876 24434 486196 31198
rect 485876 24198 485918 24434
rect 486154 24198 486196 24434
rect 485876 17434 486196 24198
rect 485876 17198 485918 17434
rect 486154 17198 486196 17434
rect 485876 10434 486196 17198
rect 485876 10198 485918 10434
rect 486154 10198 486196 10434
rect 485876 3434 486196 10198
rect 485876 3198 485918 3434
rect 486154 3198 486196 3434
rect 485876 -1706 486196 3198
rect 485876 -1942 485918 -1706
rect 486154 -1942 486196 -1706
rect 485876 -2026 486196 -1942
rect 485876 -2262 485918 -2026
rect 486154 -2262 486196 -2026
rect 485876 -2294 486196 -2262
rect 491144 705238 491464 706230
rect 491144 705002 491186 705238
rect 491422 705002 491464 705238
rect 491144 704918 491464 705002
rect 491144 704682 491186 704918
rect 491422 704682 491464 704918
rect 491144 695494 491464 704682
rect 491144 695258 491186 695494
rect 491422 695258 491464 695494
rect 491144 688494 491464 695258
rect 491144 688258 491186 688494
rect 491422 688258 491464 688494
rect 491144 681494 491464 688258
rect 491144 681258 491186 681494
rect 491422 681258 491464 681494
rect 491144 674494 491464 681258
rect 491144 674258 491186 674494
rect 491422 674258 491464 674494
rect 491144 667494 491464 674258
rect 491144 667258 491186 667494
rect 491422 667258 491464 667494
rect 491144 660494 491464 667258
rect 491144 660258 491186 660494
rect 491422 660258 491464 660494
rect 491144 653494 491464 660258
rect 491144 653258 491186 653494
rect 491422 653258 491464 653494
rect 491144 646494 491464 653258
rect 491144 646258 491186 646494
rect 491422 646258 491464 646494
rect 491144 639494 491464 646258
rect 491144 639258 491186 639494
rect 491422 639258 491464 639494
rect 491144 632494 491464 639258
rect 491144 632258 491186 632494
rect 491422 632258 491464 632494
rect 491144 625494 491464 632258
rect 491144 625258 491186 625494
rect 491422 625258 491464 625494
rect 491144 618494 491464 625258
rect 491144 618258 491186 618494
rect 491422 618258 491464 618494
rect 491144 611494 491464 618258
rect 491144 611258 491186 611494
rect 491422 611258 491464 611494
rect 491144 604494 491464 611258
rect 491144 604258 491186 604494
rect 491422 604258 491464 604494
rect 491144 597494 491464 604258
rect 491144 597258 491186 597494
rect 491422 597258 491464 597494
rect 491144 590494 491464 597258
rect 491144 590258 491186 590494
rect 491422 590258 491464 590494
rect 491144 583494 491464 590258
rect 491144 583258 491186 583494
rect 491422 583258 491464 583494
rect 491144 576494 491464 583258
rect 491144 576258 491186 576494
rect 491422 576258 491464 576494
rect 491144 569494 491464 576258
rect 491144 569258 491186 569494
rect 491422 569258 491464 569494
rect 491144 562494 491464 569258
rect 491144 562258 491186 562494
rect 491422 562258 491464 562494
rect 491144 555494 491464 562258
rect 491144 555258 491186 555494
rect 491422 555258 491464 555494
rect 491144 548494 491464 555258
rect 491144 548258 491186 548494
rect 491422 548258 491464 548494
rect 491144 541494 491464 548258
rect 491144 541258 491186 541494
rect 491422 541258 491464 541494
rect 491144 534494 491464 541258
rect 491144 534258 491186 534494
rect 491422 534258 491464 534494
rect 491144 527494 491464 534258
rect 491144 527258 491186 527494
rect 491422 527258 491464 527494
rect 491144 520494 491464 527258
rect 491144 520258 491186 520494
rect 491422 520258 491464 520494
rect 491144 513494 491464 520258
rect 491144 513258 491186 513494
rect 491422 513258 491464 513494
rect 491144 506494 491464 513258
rect 491144 506258 491186 506494
rect 491422 506258 491464 506494
rect 491144 499494 491464 506258
rect 491144 499258 491186 499494
rect 491422 499258 491464 499494
rect 491144 492494 491464 499258
rect 491144 492258 491186 492494
rect 491422 492258 491464 492494
rect 491144 485494 491464 492258
rect 491144 485258 491186 485494
rect 491422 485258 491464 485494
rect 491144 478494 491464 485258
rect 491144 478258 491186 478494
rect 491422 478258 491464 478494
rect 491144 471494 491464 478258
rect 491144 471258 491186 471494
rect 491422 471258 491464 471494
rect 491144 464494 491464 471258
rect 491144 464258 491186 464494
rect 491422 464258 491464 464494
rect 491144 457494 491464 464258
rect 491144 457258 491186 457494
rect 491422 457258 491464 457494
rect 491144 450494 491464 457258
rect 491144 450258 491186 450494
rect 491422 450258 491464 450494
rect 491144 443494 491464 450258
rect 491144 443258 491186 443494
rect 491422 443258 491464 443494
rect 491144 436494 491464 443258
rect 491144 436258 491186 436494
rect 491422 436258 491464 436494
rect 491144 429494 491464 436258
rect 491144 429258 491186 429494
rect 491422 429258 491464 429494
rect 491144 422494 491464 429258
rect 491144 422258 491186 422494
rect 491422 422258 491464 422494
rect 491144 415494 491464 422258
rect 491144 415258 491186 415494
rect 491422 415258 491464 415494
rect 491144 408494 491464 415258
rect 491144 408258 491186 408494
rect 491422 408258 491464 408494
rect 491144 401494 491464 408258
rect 491144 401258 491186 401494
rect 491422 401258 491464 401494
rect 491144 394494 491464 401258
rect 491144 394258 491186 394494
rect 491422 394258 491464 394494
rect 491144 387494 491464 394258
rect 491144 387258 491186 387494
rect 491422 387258 491464 387494
rect 491144 380494 491464 387258
rect 491144 380258 491186 380494
rect 491422 380258 491464 380494
rect 491144 373494 491464 380258
rect 491144 373258 491186 373494
rect 491422 373258 491464 373494
rect 491144 366494 491464 373258
rect 491144 366258 491186 366494
rect 491422 366258 491464 366494
rect 491144 359494 491464 366258
rect 491144 359258 491186 359494
rect 491422 359258 491464 359494
rect 491144 352494 491464 359258
rect 491144 352258 491186 352494
rect 491422 352258 491464 352494
rect 491144 345494 491464 352258
rect 491144 345258 491186 345494
rect 491422 345258 491464 345494
rect 491144 338494 491464 345258
rect 491144 338258 491186 338494
rect 491422 338258 491464 338494
rect 491144 331494 491464 338258
rect 491144 331258 491186 331494
rect 491422 331258 491464 331494
rect 491144 324494 491464 331258
rect 491144 324258 491186 324494
rect 491422 324258 491464 324494
rect 491144 317494 491464 324258
rect 491144 317258 491186 317494
rect 491422 317258 491464 317494
rect 491144 310494 491464 317258
rect 491144 310258 491186 310494
rect 491422 310258 491464 310494
rect 491144 303494 491464 310258
rect 491144 303258 491186 303494
rect 491422 303258 491464 303494
rect 491144 296494 491464 303258
rect 491144 296258 491186 296494
rect 491422 296258 491464 296494
rect 491144 289494 491464 296258
rect 491144 289258 491186 289494
rect 491422 289258 491464 289494
rect 491144 282494 491464 289258
rect 491144 282258 491186 282494
rect 491422 282258 491464 282494
rect 491144 275494 491464 282258
rect 491144 275258 491186 275494
rect 491422 275258 491464 275494
rect 491144 268494 491464 275258
rect 491144 268258 491186 268494
rect 491422 268258 491464 268494
rect 491144 261494 491464 268258
rect 491144 261258 491186 261494
rect 491422 261258 491464 261494
rect 491144 254494 491464 261258
rect 491144 254258 491186 254494
rect 491422 254258 491464 254494
rect 491144 247494 491464 254258
rect 491144 247258 491186 247494
rect 491422 247258 491464 247494
rect 491144 240494 491464 247258
rect 491144 240258 491186 240494
rect 491422 240258 491464 240494
rect 491144 233494 491464 240258
rect 491144 233258 491186 233494
rect 491422 233258 491464 233494
rect 491144 226494 491464 233258
rect 491144 226258 491186 226494
rect 491422 226258 491464 226494
rect 491144 219494 491464 226258
rect 491144 219258 491186 219494
rect 491422 219258 491464 219494
rect 491144 212494 491464 219258
rect 491144 212258 491186 212494
rect 491422 212258 491464 212494
rect 491144 205494 491464 212258
rect 491144 205258 491186 205494
rect 491422 205258 491464 205494
rect 491144 198494 491464 205258
rect 491144 198258 491186 198494
rect 491422 198258 491464 198494
rect 491144 191494 491464 198258
rect 491144 191258 491186 191494
rect 491422 191258 491464 191494
rect 491144 184494 491464 191258
rect 491144 184258 491186 184494
rect 491422 184258 491464 184494
rect 491144 177494 491464 184258
rect 491144 177258 491186 177494
rect 491422 177258 491464 177494
rect 491144 170494 491464 177258
rect 491144 170258 491186 170494
rect 491422 170258 491464 170494
rect 491144 163494 491464 170258
rect 491144 163258 491186 163494
rect 491422 163258 491464 163494
rect 491144 156494 491464 163258
rect 491144 156258 491186 156494
rect 491422 156258 491464 156494
rect 491144 149494 491464 156258
rect 491144 149258 491186 149494
rect 491422 149258 491464 149494
rect 491144 142494 491464 149258
rect 491144 142258 491186 142494
rect 491422 142258 491464 142494
rect 491144 135494 491464 142258
rect 491144 135258 491186 135494
rect 491422 135258 491464 135494
rect 491144 128494 491464 135258
rect 491144 128258 491186 128494
rect 491422 128258 491464 128494
rect 491144 121494 491464 128258
rect 491144 121258 491186 121494
rect 491422 121258 491464 121494
rect 491144 114494 491464 121258
rect 491144 114258 491186 114494
rect 491422 114258 491464 114494
rect 491144 107494 491464 114258
rect 491144 107258 491186 107494
rect 491422 107258 491464 107494
rect 491144 100494 491464 107258
rect 491144 100258 491186 100494
rect 491422 100258 491464 100494
rect 491144 93494 491464 100258
rect 491144 93258 491186 93494
rect 491422 93258 491464 93494
rect 491144 86494 491464 93258
rect 491144 86258 491186 86494
rect 491422 86258 491464 86494
rect 491144 79494 491464 86258
rect 491144 79258 491186 79494
rect 491422 79258 491464 79494
rect 491144 72494 491464 79258
rect 491144 72258 491186 72494
rect 491422 72258 491464 72494
rect 491144 65494 491464 72258
rect 491144 65258 491186 65494
rect 491422 65258 491464 65494
rect 491144 58494 491464 65258
rect 491144 58258 491186 58494
rect 491422 58258 491464 58494
rect 491144 51494 491464 58258
rect 491144 51258 491186 51494
rect 491422 51258 491464 51494
rect 491144 44494 491464 51258
rect 491144 44258 491186 44494
rect 491422 44258 491464 44494
rect 491144 37494 491464 44258
rect 491144 37258 491186 37494
rect 491422 37258 491464 37494
rect 491144 30494 491464 37258
rect 491144 30258 491186 30494
rect 491422 30258 491464 30494
rect 491144 23494 491464 30258
rect 491144 23258 491186 23494
rect 491422 23258 491464 23494
rect 491144 16494 491464 23258
rect 491144 16258 491186 16494
rect 491422 16258 491464 16494
rect 491144 9494 491464 16258
rect 491144 9258 491186 9494
rect 491422 9258 491464 9494
rect 491144 2494 491464 9258
rect 491144 2258 491186 2494
rect 491422 2258 491464 2494
rect 491144 -746 491464 2258
rect 491144 -982 491186 -746
rect 491422 -982 491464 -746
rect 491144 -1066 491464 -982
rect 491144 -1302 491186 -1066
rect 491422 -1302 491464 -1066
rect 491144 -2294 491464 -1302
rect 492876 706198 493196 706230
rect 492876 705962 492918 706198
rect 493154 705962 493196 706198
rect 492876 705878 493196 705962
rect 492876 705642 492918 705878
rect 493154 705642 493196 705878
rect 492876 696434 493196 705642
rect 492876 696198 492918 696434
rect 493154 696198 493196 696434
rect 492876 689434 493196 696198
rect 492876 689198 492918 689434
rect 493154 689198 493196 689434
rect 492876 682434 493196 689198
rect 492876 682198 492918 682434
rect 493154 682198 493196 682434
rect 492876 675434 493196 682198
rect 492876 675198 492918 675434
rect 493154 675198 493196 675434
rect 492876 668434 493196 675198
rect 492876 668198 492918 668434
rect 493154 668198 493196 668434
rect 492876 661434 493196 668198
rect 492876 661198 492918 661434
rect 493154 661198 493196 661434
rect 492876 654434 493196 661198
rect 492876 654198 492918 654434
rect 493154 654198 493196 654434
rect 492876 647434 493196 654198
rect 492876 647198 492918 647434
rect 493154 647198 493196 647434
rect 492876 640434 493196 647198
rect 492876 640198 492918 640434
rect 493154 640198 493196 640434
rect 492876 633434 493196 640198
rect 492876 633198 492918 633434
rect 493154 633198 493196 633434
rect 492876 626434 493196 633198
rect 492876 626198 492918 626434
rect 493154 626198 493196 626434
rect 492876 619434 493196 626198
rect 492876 619198 492918 619434
rect 493154 619198 493196 619434
rect 492876 612434 493196 619198
rect 492876 612198 492918 612434
rect 493154 612198 493196 612434
rect 492876 605434 493196 612198
rect 492876 605198 492918 605434
rect 493154 605198 493196 605434
rect 492876 598434 493196 605198
rect 492876 598198 492918 598434
rect 493154 598198 493196 598434
rect 492876 591434 493196 598198
rect 492876 591198 492918 591434
rect 493154 591198 493196 591434
rect 492876 584434 493196 591198
rect 492876 584198 492918 584434
rect 493154 584198 493196 584434
rect 492876 577434 493196 584198
rect 492876 577198 492918 577434
rect 493154 577198 493196 577434
rect 492876 570434 493196 577198
rect 492876 570198 492918 570434
rect 493154 570198 493196 570434
rect 492876 563434 493196 570198
rect 492876 563198 492918 563434
rect 493154 563198 493196 563434
rect 492876 556434 493196 563198
rect 492876 556198 492918 556434
rect 493154 556198 493196 556434
rect 492876 549434 493196 556198
rect 492876 549198 492918 549434
rect 493154 549198 493196 549434
rect 492876 542434 493196 549198
rect 492876 542198 492918 542434
rect 493154 542198 493196 542434
rect 492876 535434 493196 542198
rect 492876 535198 492918 535434
rect 493154 535198 493196 535434
rect 492876 528434 493196 535198
rect 492876 528198 492918 528434
rect 493154 528198 493196 528434
rect 492876 521434 493196 528198
rect 492876 521198 492918 521434
rect 493154 521198 493196 521434
rect 492876 514434 493196 521198
rect 492876 514198 492918 514434
rect 493154 514198 493196 514434
rect 492876 507434 493196 514198
rect 492876 507198 492918 507434
rect 493154 507198 493196 507434
rect 492876 500434 493196 507198
rect 492876 500198 492918 500434
rect 493154 500198 493196 500434
rect 492876 493434 493196 500198
rect 492876 493198 492918 493434
rect 493154 493198 493196 493434
rect 492876 486434 493196 493198
rect 492876 486198 492918 486434
rect 493154 486198 493196 486434
rect 492876 479434 493196 486198
rect 492876 479198 492918 479434
rect 493154 479198 493196 479434
rect 492876 472434 493196 479198
rect 492876 472198 492918 472434
rect 493154 472198 493196 472434
rect 492876 465434 493196 472198
rect 492876 465198 492918 465434
rect 493154 465198 493196 465434
rect 492876 458434 493196 465198
rect 492876 458198 492918 458434
rect 493154 458198 493196 458434
rect 492876 451434 493196 458198
rect 492876 451198 492918 451434
rect 493154 451198 493196 451434
rect 492876 444434 493196 451198
rect 492876 444198 492918 444434
rect 493154 444198 493196 444434
rect 492876 437434 493196 444198
rect 492876 437198 492918 437434
rect 493154 437198 493196 437434
rect 492876 430434 493196 437198
rect 492876 430198 492918 430434
rect 493154 430198 493196 430434
rect 492876 423434 493196 430198
rect 492876 423198 492918 423434
rect 493154 423198 493196 423434
rect 492876 416434 493196 423198
rect 492876 416198 492918 416434
rect 493154 416198 493196 416434
rect 492876 409434 493196 416198
rect 492876 409198 492918 409434
rect 493154 409198 493196 409434
rect 492876 402434 493196 409198
rect 492876 402198 492918 402434
rect 493154 402198 493196 402434
rect 492876 395434 493196 402198
rect 492876 395198 492918 395434
rect 493154 395198 493196 395434
rect 492876 388434 493196 395198
rect 492876 388198 492918 388434
rect 493154 388198 493196 388434
rect 492876 381434 493196 388198
rect 492876 381198 492918 381434
rect 493154 381198 493196 381434
rect 492876 374434 493196 381198
rect 492876 374198 492918 374434
rect 493154 374198 493196 374434
rect 492876 367434 493196 374198
rect 492876 367198 492918 367434
rect 493154 367198 493196 367434
rect 492876 360434 493196 367198
rect 492876 360198 492918 360434
rect 493154 360198 493196 360434
rect 492876 353434 493196 360198
rect 492876 353198 492918 353434
rect 493154 353198 493196 353434
rect 492876 346434 493196 353198
rect 492876 346198 492918 346434
rect 493154 346198 493196 346434
rect 492876 339434 493196 346198
rect 492876 339198 492918 339434
rect 493154 339198 493196 339434
rect 492876 332434 493196 339198
rect 492876 332198 492918 332434
rect 493154 332198 493196 332434
rect 492876 325434 493196 332198
rect 492876 325198 492918 325434
rect 493154 325198 493196 325434
rect 492876 318434 493196 325198
rect 492876 318198 492918 318434
rect 493154 318198 493196 318434
rect 492876 311434 493196 318198
rect 492876 311198 492918 311434
rect 493154 311198 493196 311434
rect 492876 304434 493196 311198
rect 492876 304198 492918 304434
rect 493154 304198 493196 304434
rect 492876 297434 493196 304198
rect 492876 297198 492918 297434
rect 493154 297198 493196 297434
rect 492876 290434 493196 297198
rect 492876 290198 492918 290434
rect 493154 290198 493196 290434
rect 492876 283434 493196 290198
rect 492876 283198 492918 283434
rect 493154 283198 493196 283434
rect 492876 276434 493196 283198
rect 492876 276198 492918 276434
rect 493154 276198 493196 276434
rect 492876 269434 493196 276198
rect 492876 269198 492918 269434
rect 493154 269198 493196 269434
rect 492876 262434 493196 269198
rect 492876 262198 492918 262434
rect 493154 262198 493196 262434
rect 492876 255434 493196 262198
rect 492876 255198 492918 255434
rect 493154 255198 493196 255434
rect 492876 248434 493196 255198
rect 492876 248198 492918 248434
rect 493154 248198 493196 248434
rect 492876 241434 493196 248198
rect 492876 241198 492918 241434
rect 493154 241198 493196 241434
rect 492876 234434 493196 241198
rect 492876 234198 492918 234434
rect 493154 234198 493196 234434
rect 492876 227434 493196 234198
rect 492876 227198 492918 227434
rect 493154 227198 493196 227434
rect 492876 220434 493196 227198
rect 492876 220198 492918 220434
rect 493154 220198 493196 220434
rect 492876 213434 493196 220198
rect 492876 213198 492918 213434
rect 493154 213198 493196 213434
rect 492876 206434 493196 213198
rect 492876 206198 492918 206434
rect 493154 206198 493196 206434
rect 492876 199434 493196 206198
rect 492876 199198 492918 199434
rect 493154 199198 493196 199434
rect 492876 192434 493196 199198
rect 492876 192198 492918 192434
rect 493154 192198 493196 192434
rect 492876 185434 493196 192198
rect 492876 185198 492918 185434
rect 493154 185198 493196 185434
rect 492876 178434 493196 185198
rect 492876 178198 492918 178434
rect 493154 178198 493196 178434
rect 492876 171434 493196 178198
rect 492876 171198 492918 171434
rect 493154 171198 493196 171434
rect 492876 164434 493196 171198
rect 492876 164198 492918 164434
rect 493154 164198 493196 164434
rect 492876 157434 493196 164198
rect 492876 157198 492918 157434
rect 493154 157198 493196 157434
rect 492876 150434 493196 157198
rect 492876 150198 492918 150434
rect 493154 150198 493196 150434
rect 492876 143434 493196 150198
rect 492876 143198 492918 143434
rect 493154 143198 493196 143434
rect 492876 136434 493196 143198
rect 492876 136198 492918 136434
rect 493154 136198 493196 136434
rect 492876 129434 493196 136198
rect 492876 129198 492918 129434
rect 493154 129198 493196 129434
rect 492876 122434 493196 129198
rect 492876 122198 492918 122434
rect 493154 122198 493196 122434
rect 492876 115434 493196 122198
rect 492876 115198 492918 115434
rect 493154 115198 493196 115434
rect 492876 108434 493196 115198
rect 492876 108198 492918 108434
rect 493154 108198 493196 108434
rect 492876 101434 493196 108198
rect 492876 101198 492918 101434
rect 493154 101198 493196 101434
rect 492876 94434 493196 101198
rect 492876 94198 492918 94434
rect 493154 94198 493196 94434
rect 492876 87434 493196 94198
rect 492876 87198 492918 87434
rect 493154 87198 493196 87434
rect 492876 80434 493196 87198
rect 492876 80198 492918 80434
rect 493154 80198 493196 80434
rect 492876 73434 493196 80198
rect 492876 73198 492918 73434
rect 493154 73198 493196 73434
rect 492876 66434 493196 73198
rect 492876 66198 492918 66434
rect 493154 66198 493196 66434
rect 492876 59434 493196 66198
rect 492876 59198 492918 59434
rect 493154 59198 493196 59434
rect 492876 52434 493196 59198
rect 492876 52198 492918 52434
rect 493154 52198 493196 52434
rect 492876 45434 493196 52198
rect 492876 45198 492918 45434
rect 493154 45198 493196 45434
rect 492876 38434 493196 45198
rect 492876 38198 492918 38434
rect 493154 38198 493196 38434
rect 492876 31434 493196 38198
rect 492876 31198 492918 31434
rect 493154 31198 493196 31434
rect 492876 24434 493196 31198
rect 492876 24198 492918 24434
rect 493154 24198 493196 24434
rect 492876 17434 493196 24198
rect 492876 17198 492918 17434
rect 493154 17198 493196 17434
rect 492876 10434 493196 17198
rect 492876 10198 492918 10434
rect 493154 10198 493196 10434
rect 492876 3434 493196 10198
rect 492876 3198 492918 3434
rect 493154 3198 493196 3434
rect 492876 -1706 493196 3198
rect 492876 -1942 492918 -1706
rect 493154 -1942 493196 -1706
rect 492876 -2026 493196 -1942
rect 492876 -2262 492918 -2026
rect 493154 -2262 493196 -2026
rect 492876 -2294 493196 -2262
rect 498144 705238 498464 706230
rect 498144 705002 498186 705238
rect 498422 705002 498464 705238
rect 498144 704918 498464 705002
rect 498144 704682 498186 704918
rect 498422 704682 498464 704918
rect 498144 695494 498464 704682
rect 498144 695258 498186 695494
rect 498422 695258 498464 695494
rect 498144 688494 498464 695258
rect 498144 688258 498186 688494
rect 498422 688258 498464 688494
rect 498144 681494 498464 688258
rect 498144 681258 498186 681494
rect 498422 681258 498464 681494
rect 498144 674494 498464 681258
rect 498144 674258 498186 674494
rect 498422 674258 498464 674494
rect 498144 667494 498464 674258
rect 498144 667258 498186 667494
rect 498422 667258 498464 667494
rect 498144 660494 498464 667258
rect 498144 660258 498186 660494
rect 498422 660258 498464 660494
rect 498144 653494 498464 660258
rect 498144 653258 498186 653494
rect 498422 653258 498464 653494
rect 498144 646494 498464 653258
rect 498144 646258 498186 646494
rect 498422 646258 498464 646494
rect 498144 639494 498464 646258
rect 498144 639258 498186 639494
rect 498422 639258 498464 639494
rect 498144 632494 498464 639258
rect 498144 632258 498186 632494
rect 498422 632258 498464 632494
rect 498144 625494 498464 632258
rect 498144 625258 498186 625494
rect 498422 625258 498464 625494
rect 498144 618494 498464 625258
rect 498144 618258 498186 618494
rect 498422 618258 498464 618494
rect 498144 611494 498464 618258
rect 498144 611258 498186 611494
rect 498422 611258 498464 611494
rect 498144 604494 498464 611258
rect 498144 604258 498186 604494
rect 498422 604258 498464 604494
rect 498144 597494 498464 604258
rect 498144 597258 498186 597494
rect 498422 597258 498464 597494
rect 498144 590494 498464 597258
rect 498144 590258 498186 590494
rect 498422 590258 498464 590494
rect 498144 583494 498464 590258
rect 498144 583258 498186 583494
rect 498422 583258 498464 583494
rect 498144 576494 498464 583258
rect 498144 576258 498186 576494
rect 498422 576258 498464 576494
rect 498144 569494 498464 576258
rect 498144 569258 498186 569494
rect 498422 569258 498464 569494
rect 498144 562494 498464 569258
rect 498144 562258 498186 562494
rect 498422 562258 498464 562494
rect 498144 555494 498464 562258
rect 498144 555258 498186 555494
rect 498422 555258 498464 555494
rect 498144 548494 498464 555258
rect 498144 548258 498186 548494
rect 498422 548258 498464 548494
rect 498144 541494 498464 548258
rect 498144 541258 498186 541494
rect 498422 541258 498464 541494
rect 498144 534494 498464 541258
rect 498144 534258 498186 534494
rect 498422 534258 498464 534494
rect 498144 527494 498464 534258
rect 498144 527258 498186 527494
rect 498422 527258 498464 527494
rect 498144 520494 498464 527258
rect 498144 520258 498186 520494
rect 498422 520258 498464 520494
rect 498144 513494 498464 520258
rect 498144 513258 498186 513494
rect 498422 513258 498464 513494
rect 498144 506494 498464 513258
rect 498144 506258 498186 506494
rect 498422 506258 498464 506494
rect 498144 499494 498464 506258
rect 498144 499258 498186 499494
rect 498422 499258 498464 499494
rect 498144 492494 498464 499258
rect 498144 492258 498186 492494
rect 498422 492258 498464 492494
rect 498144 485494 498464 492258
rect 498144 485258 498186 485494
rect 498422 485258 498464 485494
rect 498144 478494 498464 485258
rect 498144 478258 498186 478494
rect 498422 478258 498464 478494
rect 498144 471494 498464 478258
rect 498144 471258 498186 471494
rect 498422 471258 498464 471494
rect 498144 464494 498464 471258
rect 498144 464258 498186 464494
rect 498422 464258 498464 464494
rect 498144 457494 498464 464258
rect 498144 457258 498186 457494
rect 498422 457258 498464 457494
rect 498144 450494 498464 457258
rect 498144 450258 498186 450494
rect 498422 450258 498464 450494
rect 498144 443494 498464 450258
rect 498144 443258 498186 443494
rect 498422 443258 498464 443494
rect 498144 436494 498464 443258
rect 498144 436258 498186 436494
rect 498422 436258 498464 436494
rect 498144 429494 498464 436258
rect 498144 429258 498186 429494
rect 498422 429258 498464 429494
rect 498144 422494 498464 429258
rect 498144 422258 498186 422494
rect 498422 422258 498464 422494
rect 498144 415494 498464 422258
rect 498144 415258 498186 415494
rect 498422 415258 498464 415494
rect 498144 408494 498464 415258
rect 498144 408258 498186 408494
rect 498422 408258 498464 408494
rect 498144 401494 498464 408258
rect 498144 401258 498186 401494
rect 498422 401258 498464 401494
rect 498144 394494 498464 401258
rect 498144 394258 498186 394494
rect 498422 394258 498464 394494
rect 498144 387494 498464 394258
rect 498144 387258 498186 387494
rect 498422 387258 498464 387494
rect 498144 380494 498464 387258
rect 498144 380258 498186 380494
rect 498422 380258 498464 380494
rect 498144 373494 498464 380258
rect 498144 373258 498186 373494
rect 498422 373258 498464 373494
rect 498144 366494 498464 373258
rect 498144 366258 498186 366494
rect 498422 366258 498464 366494
rect 498144 359494 498464 366258
rect 498144 359258 498186 359494
rect 498422 359258 498464 359494
rect 498144 352494 498464 359258
rect 498144 352258 498186 352494
rect 498422 352258 498464 352494
rect 498144 345494 498464 352258
rect 498144 345258 498186 345494
rect 498422 345258 498464 345494
rect 498144 338494 498464 345258
rect 498144 338258 498186 338494
rect 498422 338258 498464 338494
rect 498144 331494 498464 338258
rect 498144 331258 498186 331494
rect 498422 331258 498464 331494
rect 498144 324494 498464 331258
rect 498144 324258 498186 324494
rect 498422 324258 498464 324494
rect 498144 317494 498464 324258
rect 498144 317258 498186 317494
rect 498422 317258 498464 317494
rect 498144 310494 498464 317258
rect 498144 310258 498186 310494
rect 498422 310258 498464 310494
rect 498144 303494 498464 310258
rect 498144 303258 498186 303494
rect 498422 303258 498464 303494
rect 498144 296494 498464 303258
rect 498144 296258 498186 296494
rect 498422 296258 498464 296494
rect 498144 289494 498464 296258
rect 498144 289258 498186 289494
rect 498422 289258 498464 289494
rect 498144 282494 498464 289258
rect 498144 282258 498186 282494
rect 498422 282258 498464 282494
rect 498144 275494 498464 282258
rect 498144 275258 498186 275494
rect 498422 275258 498464 275494
rect 498144 268494 498464 275258
rect 498144 268258 498186 268494
rect 498422 268258 498464 268494
rect 498144 261494 498464 268258
rect 498144 261258 498186 261494
rect 498422 261258 498464 261494
rect 498144 254494 498464 261258
rect 498144 254258 498186 254494
rect 498422 254258 498464 254494
rect 498144 247494 498464 254258
rect 498144 247258 498186 247494
rect 498422 247258 498464 247494
rect 498144 240494 498464 247258
rect 498144 240258 498186 240494
rect 498422 240258 498464 240494
rect 498144 233494 498464 240258
rect 498144 233258 498186 233494
rect 498422 233258 498464 233494
rect 498144 226494 498464 233258
rect 498144 226258 498186 226494
rect 498422 226258 498464 226494
rect 498144 219494 498464 226258
rect 498144 219258 498186 219494
rect 498422 219258 498464 219494
rect 498144 212494 498464 219258
rect 498144 212258 498186 212494
rect 498422 212258 498464 212494
rect 498144 205494 498464 212258
rect 498144 205258 498186 205494
rect 498422 205258 498464 205494
rect 498144 198494 498464 205258
rect 498144 198258 498186 198494
rect 498422 198258 498464 198494
rect 498144 191494 498464 198258
rect 498144 191258 498186 191494
rect 498422 191258 498464 191494
rect 498144 184494 498464 191258
rect 498144 184258 498186 184494
rect 498422 184258 498464 184494
rect 498144 177494 498464 184258
rect 498144 177258 498186 177494
rect 498422 177258 498464 177494
rect 498144 170494 498464 177258
rect 498144 170258 498186 170494
rect 498422 170258 498464 170494
rect 498144 163494 498464 170258
rect 498144 163258 498186 163494
rect 498422 163258 498464 163494
rect 498144 156494 498464 163258
rect 498144 156258 498186 156494
rect 498422 156258 498464 156494
rect 498144 149494 498464 156258
rect 498144 149258 498186 149494
rect 498422 149258 498464 149494
rect 498144 142494 498464 149258
rect 498144 142258 498186 142494
rect 498422 142258 498464 142494
rect 498144 135494 498464 142258
rect 498144 135258 498186 135494
rect 498422 135258 498464 135494
rect 498144 128494 498464 135258
rect 498144 128258 498186 128494
rect 498422 128258 498464 128494
rect 498144 121494 498464 128258
rect 498144 121258 498186 121494
rect 498422 121258 498464 121494
rect 498144 114494 498464 121258
rect 498144 114258 498186 114494
rect 498422 114258 498464 114494
rect 498144 107494 498464 114258
rect 498144 107258 498186 107494
rect 498422 107258 498464 107494
rect 498144 100494 498464 107258
rect 498144 100258 498186 100494
rect 498422 100258 498464 100494
rect 498144 93494 498464 100258
rect 498144 93258 498186 93494
rect 498422 93258 498464 93494
rect 498144 86494 498464 93258
rect 498144 86258 498186 86494
rect 498422 86258 498464 86494
rect 498144 79494 498464 86258
rect 498144 79258 498186 79494
rect 498422 79258 498464 79494
rect 498144 72494 498464 79258
rect 498144 72258 498186 72494
rect 498422 72258 498464 72494
rect 498144 65494 498464 72258
rect 498144 65258 498186 65494
rect 498422 65258 498464 65494
rect 498144 58494 498464 65258
rect 498144 58258 498186 58494
rect 498422 58258 498464 58494
rect 498144 51494 498464 58258
rect 498144 51258 498186 51494
rect 498422 51258 498464 51494
rect 498144 44494 498464 51258
rect 498144 44258 498186 44494
rect 498422 44258 498464 44494
rect 498144 37494 498464 44258
rect 498144 37258 498186 37494
rect 498422 37258 498464 37494
rect 498144 30494 498464 37258
rect 498144 30258 498186 30494
rect 498422 30258 498464 30494
rect 498144 23494 498464 30258
rect 498144 23258 498186 23494
rect 498422 23258 498464 23494
rect 498144 16494 498464 23258
rect 498144 16258 498186 16494
rect 498422 16258 498464 16494
rect 498144 9494 498464 16258
rect 498144 9258 498186 9494
rect 498422 9258 498464 9494
rect 498144 2494 498464 9258
rect 498144 2258 498186 2494
rect 498422 2258 498464 2494
rect 498144 -746 498464 2258
rect 498144 -982 498186 -746
rect 498422 -982 498464 -746
rect 498144 -1066 498464 -982
rect 498144 -1302 498186 -1066
rect 498422 -1302 498464 -1066
rect 498144 -2294 498464 -1302
rect 499876 706198 500196 706230
rect 499876 705962 499918 706198
rect 500154 705962 500196 706198
rect 499876 705878 500196 705962
rect 499876 705642 499918 705878
rect 500154 705642 500196 705878
rect 499876 696434 500196 705642
rect 499876 696198 499918 696434
rect 500154 696198 500196 696434
rect 499876 689434 500196 696198
rect 499876 689198 499918 689434
rect 500154 689198 500196 689434
rect 499876 682434 500196 689198
rect 499876 682198 499918 682434
rect 500154 682198 500196 682434
rect 499876 675434 500196 682198
rect 499876 675198 499918 675434
rect 500154 675198 500196 675434
rect 499876 668434 500196 675198
rect 499876 668198 499918 668434
rect 500154 668198 500196 668434
rect 499876 661434 500196 668198
rect 499876 661198 499918 661434
rect 500154 661198 500196 661434
rect 499876 654434 500196 661198
rect 499876 654198 499918 654434
rect 500154 654198 500196 654434
rect 499876 647434 500196 654198
rect 499876 647198 499918 647434
rect 500154 647198 500196 647434
rect 499876 640434 500196 647198
rect 499876 640198 499918 640434
rect 500154 640198 500196 640434
rect 499876 633434 500196 640198
rect 499876 633198 499918 633434
rect 500154 633198 500196 633434
rect 499876 626434 500196 633198
rect 499876 626198 499918 626434
rect 500154 626198 500196 626434
rect 499876 619434 500196 626198
rect 499876 619198 499918 619434
rect 500154 619198 500196 619434
rect 499876 612434 500196 619198
rect 499876 612198 499918 612434
rect 500154 612198 500196 612434
rect 499876 605434 500196 612198
rect 499876 605198 499918 605434
rect 500154 605198 500196 605434
rect 499876 598434 500196 605198
rect 499876 598198 499918 598434
rect 500154 598198 500196 598434
rect 499876 591434 500196 598198
rect 499876 591198 499918 591434
rect 500154 591198 500196 591434
rect 499876 584434 500196 591198
rect 499876 584198 499918 584434
rect 500154 584198 500196 584434
rect 499876 577434 500196 584198
rect 499876 577198 499918 577434
rect 500154 577198 500196 577434
rect 499876 570434 500196 577198
rect 499876 570198 499918 570434
rect 500154 570198 500196 570434
rect 499876 563434 500196 570198
rect 499876 563198 499918 563434
rect 500154 563198 500196 563434
rect 499876 556434 500196 563198
rect 499876 556198 499918 556434
rect 500154 556198 500196 556434
rect 499876 549434 500196 556198
rect 499876 549198 499918 549434
rect 500154 549198 500196 549434
rect 499876 542434 500196 549198
rect 499876 542198 499918 542434
rect 500154 542198 500196 542434
rect 499876 535434 500196 542198
rect 499876 535198 499918 535434
rect 500154 535198 500196 535434
rect 499876 528434 500196 535198
rect 499876 528198 499918 528434
rect 500154 528198 500196 528434
rect 499876 521434 500196 528198
rect 499876 521198 499918 521434
rect 500154 521198 500196 521434
rect 499876 514434 500196 521198
rect 499876 514198 499918 514434
rect 500154 514198 500196 514434
rect 499876 507434 500196 514198
rect 499876 507198 499918 507434
rect 500154 507198 500196 507434
rect 499876 500434 500196 507198
rect 499876 500198 499918 500434
rect 500154 500198 500196 500434
rect 499876 493434 500196 500198
rect 499876 493198 499918 493434
rect 500154 493198 500196 493434
rect 499876 486434 500196 493198
rect 499876 486198 499918 486434
rect 500154 486198 500196 486434
rect 499876 479434 500196 486198
rect 499876 479198 499918 479434
rect 500154 479198 500196 479434
rect 499876 472434 500196 479198
rect 499876 472198 499918 472434
rect 500154 472198 500196 472434
rect 499876 465434 500196 472198
rect 499876 465198 499918 465434
rect 500154 465198 500196 465434
rect 499876 458434 500196 465198
rect 499876 458198 499918 458434
rect 500154 458198 500196 458434
rect 499876 451434 500196 458198
rect 499876 451198 499918 451434
rect 500154 451198 500196 451434
rect 499876 444434 500196 451198
rect 499876 444198 499918 444434
rect 500154 444198 500196 444434
rect 499876 437434 500196 444198
rect 499876 437198 499918 437434
rect 500154 437198 500196 437434
rect 499876 430434 500196 437198
rect 499876 430198 499918 430434
rect 500154 430198 500196 430434
rect 499876 423434 500196 430198
rect 499876 423198 499918 423434
rect 500154 423198 500196 423434
rect 499876 416434 500196 423198
rect 499876 416198 499918 416434
rect 500154 416198 500196 416434
rect 499876 409434 500196 416198
rect 499876 409198 499918 409434
rect 500154 409198 500196 409434
rect 499876 402434 500196 409198
rect 499876 402198 499918 402434
rect 500154 402198 500196 402434
rect 499876 395434 500196 402198
rect 499876 395198 499918 395434
rect 500154 395198 500196 395434
rect 499876 388434 500196 395198
rect 499876 388198 499918 388434
rect 500154 388198 500196 388434
rect 499876 381434 500196 388198
rect 499876 381198 499918 381434
rect 500154 381198 500196 381434
rect 499876 374434 500196 381198
rect 499876 374198 499918 374434
rect 500154 374198 500196 374434
rect 499876 367434 500196 374198
rect 499876 367198 499918 367434
rect 500154 367198 500196 367434
rect 499876 360434 500196 367198
rect 499876 360198 499918 360434
rect 500154 360198 500196 360434
rect 499876 353434 500196 360198
rect 499876 353198 499918 353434
rect 500154 353198 500196 353434
rect 499876 346434 500196 353198
rect 499876 346198 499918 346434
rect 500154 346198 500196 346434
rect 499876 339434 500196 346198
rect 499876 339198 499918 339434
rect 500154 339198 500196 339434
rect 499876 332434 500196 339198
rect 499876 332198 499918 332434
rect 500154 332198 500196 332434
rect 499876 325434 500196 332198
rect 499876 325198 499918 325434
rect 500154 325198 500196 325434
rect 499876 318434 500196 325198
rect 499876 318198 499918 318434
rect 500154 318198 500196 318434
rect 499876 311434 500196 318198
rect 499876 311198 499918 311434
rect 500154 311198 500196 311434
rect 499876 304434 500196 311198
rect 499876 304198 499918 304434
rect 500154 304198 500196 304434
rect 499876 297434 500196 304198
rect 499876 297198 499918 297434
rect 500154 297198 500196 297434
rect 499876 290434 500196 297198
rect 499876 290198 499918 290434
rect 500154 290198 500196 290434
rect 499876 283434 500196 290198
rect 499876 283198 499918 283434
rect 500154 283198 500196 283434
rect 499876 276434 500196 283198
rect 499876 276198 499918 276434
rect 500154 276198 500196 276434
rect 499876 269434 500196 276198
rect 499876 269198 499918 269434
rect 500154 269198 500196 269434
rect 499876 262434 500196 269198
rect 499876 262198 499918 262434
rect 500154 262198 500196 262434
rect 499876 255434 500196 262198
rect 499876 255198 499918 255434
rect 500154 255198 500196 255434
rect 499876 248434 500196 255198
rect 499876 248198 499918 248434
rect 500154 248198 500196 248434
rect 499876 241434 500196 248198
rect 499876 241198 499918 241434
rect 500154 241198 500196 241434
rect 499876 234434 500196 241198
rect 499876 234198 499918 234434
rect 500154 234198 500196 234434
rect 499876 227434 500196 234198
rect 499876 227198 499918 227434
rect 500154 227198 500196 227434
rect 499876 220434 500196 227198
rect 499876 220198 499918 220434
rect 500154 220198 500196 220434
rect 499876 213434 500196 220198
rect 499876 213198 499918 213434
rect 500154 213198 500196 213434
rect 499876 206434 500196 213198
rect 499876 206198 499918 206434
rect 500154 206198 500196 206434
rect 499876 199434 500196 206198
rect 499876 199198 499918 199434
rect 500154 199198 500196 199434
rect 499876 192434 500196 199198
rect 499876 192198 499918 192434
rect 500154 192198 500196 192434
rect 499876 185434 500196 192198
rect 499876 185198 499918 185434
rect 500154 185198 500196 185434
rect 499876 178434 500196 185198
rect 499876 178198 499918 178434
rect 500154 178198 500196 178434
rect 499876 171434 500196 178198
rect 499876 171198 499918 171434
rect 500154 171198 500196 171434
rect 499876 164434 500196 171198
rect 499876 164198 499918 164434
rect 500154 164198 500196 164434
rect 499876 157434 500196 164198
rect 499876 157198 499918 157434
rect 500154 157198 500196 157434
rect 499876 150434 500196 157198
rect 499876 150198 499918 150434
rect 500154 150198 500196 150434
rect 499876 143434 500196 150198
rect 499876 143198 499918 143434
rect 500154 143198 500196 143434
rect 499876 136434 500196 143198
rect 499876 136198 499918 136434
rect 500154 136198 500196 136434
rect 499876 129434 500196 136198
rect 499876 129198 499918 129434
rect 500154 129198 500196 129434
rect 499876 122434 500196 129198
rect 499876 122198 499918 122434
rect 500154 122198 500196 122434
rect 499876 115434 500196 122198
rect 499876 115198 499918 115434
rect 500154 115198 500196 115434
rect 499876 108434 500196 115198
rect 499876 108198 499918 108434
rect 500154 108198 500196 108434
rect 499876 101434 500196 108198
rect 499876 101198 499918 101434
rect 500154 101198 500196 101434
rect 499876 94434 500196 101198
rect 499876 94198 499918 94434
rect 500154 94198 500196 94434
rect 499876 87434 500196 94198
rect 499876 87198 499918 87434
rect 500154 87198 500196 87434
rect 499876 80434 500196 87198
rect 499876 80198 499918 80434
rect 500154 80198 500196 80434
rect 499876 73434 500196 80198
rect 499876 73198 499918 73434
rect 500154 73198 500196 73434
rect 499876 66434 500196 73198
rect 499876 66198 499918 66434
rect 500154 66198 500196 66434
rect 499876 59434 500196 66198
rect 499876 59198 499918 59434
rect 500154 59198 500196 59434
rect 499876 52434 500196 59198
rect 499876 52198 499918 52434
rect 500154 52198 500196 52434
rect 499876 45434 500196 52198
rect 499876 45198 499918 45434
rect 500154 45198 500196 45434
rect 499876 38434 500196 45198
rect 499876 38198 499918 38434
rect 500154 38198 500196 38434
rect 499876 31434 500196 38198
rect 499876 31198 499918 31434
rect 500154 31198 500196 31434
rect 499876 24434 500196 31198
rect 499876 24198 499918 24434
rect 500154 24198 500196 24434
rect 499876 17434 500196 24198
rect 499876 17198 499918 17434
rect 500154 17198 500196 17434
rect 499876 10434 500196 17198
rect 499876 10198 499918 10434
rect 500154 10198 500196 10434
rect 499876 3434 500196 10198
rect 499876 3198 499918 3434
rect 500154 3198 500196 3434
rect 499876 -1706 500196 3198
rect 499876 -1942 499918 -1706
rect 500154 -1942 500196 -1706
rect 499876 -2026 500196 -1942
rect 499876 -2262 499918 -2026
rect 500154 -2262 500196 -2026
rect 499876 -2294 500196 -2262
rect 505144 705238 505464 706230
rect 505144 705002 505186 705238
rect 505422 705002 505464 705238
rect 505144 704918 505464 705002
rect 505144 704682 505186 704918
rect 505422 704682 505464 704918
rect 505144 695494 505464 704682
rect 505144 695258 505186 695494
rect 505422 695258 505464 695494
rect 505144 688494 505464 695258
rect 505144 688258 505186 688494
rect 505422 688258 505464 688494
rect 505144 681494 505464 688258
rect 505144 681258 505186 681494
rect 505422 681258 505464 681494
rect 505144 674494 505464 681258
rect 505144 674258 505186 674494
rect 505422 674258 505464 674494
rect 505144 667494 505464 674258
rect 505144 667258 505186 667494
rect 505422 667258 505464 667494
rect 505144 660494 505464 667258
rect 505144 660258 505186 660494
rect 505422 660258 505464 660494
rect 505144 653494 505464 660258
rect 505144 653258 505186 653494
rect 505422 653258 505464 653494
rect 505144 646494 505464 653258
rect 505144 646258 505186 646494
rect 505422 646258 505464 646494
rect 505144 639494 505464 646258
rect 505144 639258 505186 639494
rect 505422 639258 505464 639494
rect 505144 632494 505464 639258
rect 505144 632258 505186 632494
rect 505422 632258 505464 632494
rect 505144 625494 505464 632258
rect 505144 625258 505186 625494
rect 505422 625258 505464 625494
rect 505144 618494 505464 625258
rect 505144 618258 505186 618494
rect 505422 618258 505464 618494
rect 505144 611494 505464 618258
rect 505144 611258 505186 611494
rect 505422 611258 505464 611494
rect 505144 604494 505464 611258
rect 505144 604258 505186 604494
rect 505422 604258 505464 604494
rect 505144 597494 505464 604258
rect 505144 597258 505186 597494
rect 505422 597258 505464 597494
rect 505144 590494 505464 597258
rect 505144 590258 505186 590494
rect 505422 590258 505464 590494
rect 505144 583494 505464 590258
rect 505144 583258 505186 583494
rect 505422 583258 505464 583494
rect 505144 576494 505464 583258
rect 505144 576258 505186 576494
rect 505422 576258 505464 576494
rect 505144 569494 505464 576258
rect 505144 569258 505186 569494
rect 505422 569258 505464 569494
rect 505144 562494 505464 569258
rect 505144 562258 505186 562494
rect 505422 562258 505464 562494
rect 505144 555494 505464 562258
rect 505144 555258 505186 555494
rect 505422 555258 505464 555494
rect 505144 548494 505464 555258
rect 505144 548258 505186 548494
rect 505422 548258 505464 548494
rect 505144 541494 505464 548258
rect 505144 541258 505186 541494
rect 505422 541258 505464 541494
rect 505144 534494 505464 541258
rect 505144 534258 505186 534494
rect 505422 534258 505464 534494
rect 505144 527494 505464 534258
rect 505144 527258 505186 527494
rect 505422 527258 505464 527494
rect 505144 520494 505464 527258
rect 505144 520258 505186 520494
rect 505422 520258 505464 520494
rect 505144 513494 505464 520258
rect 505144 513258 505186 513494
rect 505422 513258 505464 513494
rect 505144 506494 505464 513258
rect 505144 506258 505186 506494
rect 505422 506258 505464 506494
rect 505144 499494 505464 506258
rect 505144 499258 505186 499494
rect 505422 499258 505464 499494
rect 505144 492494 505464 499258
rect 505144 492258 505186 492494
rect 505422 492258 505464 492494
rect 505144 485494 505464 492258
rect 505144 485258 505186 485494
rect 505422 485258 505464 485494
rect 505144 478494 505464 485258
rect 505144 478258 505186 478494
rect 505422 478258 505464 478494
rect 505144 471494 505464 478258
rect 505144 471258 505186 471494
rect 505422 471258 505464 471494
rect 505144 464494 505464 471258
rect 505144 464258 505186 464494
rect 505422 464258 505464 464494
rect 505144 457494 505464 464258
rect 505144 457258 505186 457494
rect 505422 457258 505464 457494
rect 505144 450494 505464 457258
rect 505144 450258 505186 450494
rect 505422 450258 505464 450494
rect 505144 443494 505464 450258
rect 505144 443258 505186 443494
rect 505422 443258 505464 443494
rect 505144 436494 505464 443258
rect 505144 436258 505186 436494
rect 505422 436258 505464 436494
rect 505144 429494 505464 436258
rect 505144 429258 505186 429494
rect 505422 429258 505464 429494
rect 505144 422494 505464 429258
rect 505144 422258 505186 422494
rect 505422 422258 505464 422494
rect 505144 415494 505464 422258
rect 505144 415258 505186 415494
rect 505422 415258 505464 415494
rect 505144 408494 505464 415258
rect 505144 408258 505186 408494
rect 505422 408258 505464 408494
rect 505144 401494 505464 408258
rect 505144 401258 505186 401494
rect 505422 401258 505464 401494
rect 505144 394494 505464 401258
rect 505144 394258 505186 394494
rect 505422 394258 505464 394494
rect 505144 387494 505464 394258
rect 505144 387258 505186 387494
rect 505422 387258 505464 387494
rect 505144 380494 505464 387258
rect 505144 380258 505186 380494
rect 505422 380258 505464 380494
rect 505144 373494 505464 380258
rect 505144 373258 505186 373494
rect 505422 373258 505464 373494
rect 505144 366494 505464 373258
rect 505144 366258 505186 366494
rect 505422 366258 505464 366494
rect 505144 359494 505464 366258
rect 505144 359258 505186 359494
rect 505422 359258 505464 359494
rect 505144 352494 505464 359258
rect 505144 352258 505186 352494
rect 505422 352258 505464 352494
rect 505144 345494 505464 352258
rect 505144 345258 505186 345494
rect 505422 345258 505464 345494
rect 505144 338494 505464 345258
rect 505144 338258 505186 338494
rect 505422 338258 505464 338494
rect 505144 331494 505464 338258
rect 505144 331258 505186 331494
rect 505422 331258 505464 331494
rect 505144 324494 505464 331258
rect 505144 324258 505186 324494
rect 505422 324258 505464 324494
rect 505144 317494 505464 324258
rect 505144 317258 505186 317494
rect 505422 317258 505464 317494
rect 505144 310494 505464 317258
rect 505144 310258 505186 310494
rect 505422 310258 505464 310494
rect 505144 303494 505464 310258
rect 505144 303258 505186 303494
rect 505422 303258 505464 303494
rect 505144 296494 505464 303258
rect 505144 296258 505186 296494
rect 505422 296258 505464 296494
rect 505144 289494 505464 296258
rect 505144 289258 505186 289494
rect 505422 289258 505464 289494
rect 505144 282494 505464 289258
rect 505144 282258 505186 282494
rect 505422 282258 505464 282494
rect 505144 275494 505464 282258
rect 505144 275258 505186 275494
rect 505422 275258 505464 275494
rect 505144 268494 505464 275258
rect 505144 268258 505186 268494
rect 505422 268258 505464 268494
rect 505144 261494 505464 268258
rect 505144 261258 505186 261494
rect 505422 261258 505464 261494
rect 505144 254494 505464 261258
rect 505144 254258 505186 254494
rect 505422 254258 505464 254494
rect 505144 247494 505464 254258
rect 505144 247258 505186 247494
rect 505422 247258 505464 247494
rect 505144 240494 505464 247258
rect 505144 240258 505186 240494
rect 505422 240258 505464 240494
rect 505144 233494 505464 240258
rect 505144 233258 505186 233494
rect 505422 233258 505464 233494
rect 505144 226494 505464 233258
rect 505144 226258 505186 226494
rect 505422 226258 505464 226494
rect 505144 219494 505464 226258
rect 505144 219258 505186 219494
rect 505422 219258 505464 219494
rect 505144 212494 505464 219258
rect 505144 212258 505186 212494
rect 505422 212258 505464 212494
rect 505144 205494 505464 212258
rect 505144 205258 505186 205494
rect 505422 205258 505464 205494
rect 505144 198494 505464 205258
rect 505144 198258 505186 198494
rect 505422 198258 505464 198494
rect 505144 191494 505464 198258
rect 505144 191258 505186 191494
rect 505422 191258 505464 191494
rect 505144 184494 505464 191258
rect 505144 184258 505186 184494
rect 505422 184258 505464 184494
rect 505144 177494 505464 184258
rect 505144 177258 505186 177494
rect 505422 177258 505464 177494
rect 505144 170494 505464 177258
rect 505144 170258 505186 170494
rect 505422 170258 505464 170494
rect 505144 163494 505464 170258
rect 505144 163258 505186 163494
rect 505422 163258 505464 163494
rect 505144 156494 505464 163258
rect 505144 156258 505186 156494
rect 505422 156258 505464 156494
rect 505144 149494 505464 156258
rect 505144 149258 505186 149494
rect 505422 149258 505464 149494
rect 505144 142494 505464 149258
rect 505144 142258 505186 142494
rect 505422 142258 505464 142494
rect 505144 135494 505464 142258
rect 505144 135258 505186 135494
rect 505422 135258 505464 135494
rect 505144 128494 505464 135258
rect 505144 128258 505186 128494
rect 505422 128258 505464 128494
rect 505144 121494 505464 128258
rect 505144 121258 505186 121494
rect 505422 121258 505464 121494
rect 505144 114494 505464 121258
rect 505144 114258 505186 114494
rect 505422 114258 505464 114494
rect 505144 107494 505464 114258
rect 505144 107258 505186 107494
rect 505422 107258 505464 107494
rect 505144 100494 505464 107258
rect 505144 100258 505186 100494
rect 505422 100258 505464 100494
rect 505144 93494 505464 100258
rect 505144 93258 505186 93494
rect 505422 93258 505464 93494
rect 505144 86494 505464 93258
rect 505144 86258 505186 86494
rect 505422 86258 505464 86494
rect 505144 79494 505464 86258
rect 505144 79258 505186 79494
rect 505422 79258 505464 79494
rect 505144 72494 505464 79258
rect 505144 72258 505186 72494
rect 505422 72258 505464 72494
rect 505144 65494 505464 72258
rect 505144 65258 505186 65494
rect 505422 65258 505464 65494
rect 505144 58494 505464 65258
rect 505144 58258 505186 58494
rect 505422 58258 505464 58494
rect 505144 51494 505464 58258
rect 505144 51258 505186 51494
rect 505422 51258 505464 51494
rect 505144 44494 505464 51258
rect 505144 44258 505186 44494
rect 505422 44258 505464 44494
rect 505144 37494 505464 44258
rect 505144 37258 505186 37494
rect 505422 37258 505464 37494
rect 505144 30494 505464 37258
rect 505144 30258 505186 30494
rect 505422 30258 505464 30494
rect 505144 23494 505464 30258
rect 505144 23258 505186 23494
rect 505422 23258 505464 23494
rect 505144 16494 505464 23258
rect 505144 16258 505186 16494
rect 505422 16258 505464 16494
rect 505144 9494 505464 16258
rect 505144 9258 505186 9494
rect 505422 9258 505464 9494
rect 505144 2494 505464 9258
rect 505144 2258 505186 2494
rect 505422 2258 505464 2494
rect 505144 -746 505464 2258
rect 505144 -982 505186 -746
rect 505422 -982 505464 -746
rect 505144 -1066 505464 -982
rect 505144 -1302 505186 -1066
rect 505422 -1302 505464 -1066
rect 505144 -2294 505464 -1302
rect 506876 706198 507196 706230
rect 506876 705962 506918 706198
rect 507154 705962 507196 706198
rect 506876 705878 507196 705962
rect 506876 705642 506918 705878
rect 507154 705642 507196 705878
rect 506876 696434 507196 705642
rect 506876 696198 506918 696434
rect 507154 696198 507196 696434
rect 506876 689434 507196 696198
rect 506876 689198 506918 689434
rect 507154 689198 507196 689434
rect 506876 682434 507196 689198
rect 506876 682198 506918 682434
rect 507154 682198 507196 682434
rect 506876 675434 507196 682198
rect 506876 675198 506918 675434
rect 507154 675198 507196 675434
rect 506876 668434 507196 675198
rect 506876 668198 506918 668434
rect 507154 668198 507196 668434
rect 506876 661434 507196 668198
rect 506876 661198 506918 661434
rect 507154 661198 507196 661434
rect 506876 654434 507196 661198
rect 506876 654198 506918 654434
rect 507154 654198 507196 654434
rect 506876 647434 507196 654198
rect 506876 647198 506918 647434
rect 507154 647198 507196 647434
rect 506876 640434 507196 647198
rect 506876 640198 506918 640434
rect 507154 640198 507196 640434
rect 506876 633434 507196 640198
rect 506876 633198 506918 633434
rect 507154 633198 507196 633434
rect 506876 626434 507196 633198
rect 506876 626198 506918 626434
rect 507154 626198 507196 626434
rect 506876 619434 507196 626198
rect 506876 619198 506918 619434
rect 507154 619198 507196 619434
rect 506876 612434 507196 619198
rect 506876 612198 506918 612434
rect 507154 612198 507196 612434
rect 506876 605434 507196 612198
rect 506876 605198 506918 605434
rect 507154 605198 507196 605434
rect 506876 598434 507196 605198
rect 506876 598198 506918 598434
rect 507154 598198 507196 598434
rect 506876 591434 507196 598198
rect 506876 591198 506918 591434
rect 507154 591198 507196 591434
rect 506876 584434 507196 591198
rect 506876 584198 506918 584434
rect 507154 584198 507196 584434
rect 506876 577434 507196 584198
rect 506876 577198 506918 577434
rect 507154 577198 507196 577434
rect 506876 570434 507196 577198
rect 506876 570198 506918 570434
rect 507154 570198 507196 570434
rect 506876 563434 507196 570198
rect 506876 563198 506918 563434
rect 507154 563198 507196 563434
rect 506876 556434 507196 563198
rect 506876 556198 506918 556434
rect 507154 556198 507196 556434
rect 506876 549434 507196 556198
rect 506876 549198 506918 549434
rect 507154 549198 507196 549434
rect 506876 542434 507196 549198
rect 506876 542198 506918 542434
rect 507154 542198 507196 542434
rect 506876 535434 507196 542198
rect 506876 535198 506918 535434
rect 507154 535198 507196 535434
rect 506876 528434 507196 535198
rect 506876 528198 506918 528434
rect 507154 528198 507196 528434
rect 506876 521434 507196 528198
rect 506876 521198 506918 521434
rect 507154 521198 507196 521434
rect 506876 514434 507196 521198
rect 506876 514198 506918 514434
rect 507154 514198 507196 514434
rect 506876 507434 507196 514198
rect 506876 507198 506918 507434
rect 507154 507198 507196 507434
rect 506876 500434 507196 507198
rect 506876 500198 506918 500434
rect 507154 500198 507196 500434
rect 506876 493434 507196 500198
rect 506876 493198 506918 493434
rect 507154 493198 507196 493434
rect 506876 486434 507196 493198
rect 506876 486198 506918 486434
rect 507154 486198 507196 486434
rect 506876 479434 507196 486198
rect 506876 479198 506918 479434
rect 507154 479198 507196 479434
rect 506876 472434 507196 479198
rect 506876 472198 506918 472434
rect 507154 472198 507196 472434
rect 506876 465434 507196 472198
rect 506876 465198 506918 465434
rect 507154 465198 507196 465434
rect 506876 458434 507196 465198
rect 506876 458198 506918 458434
rect 507154 458198 507196 458434
rect 506876 451434 507196 458198
rect 506876 451198 506918 451434
rect 507154 451198 507196 451434
rect 506876 444434 507196 451198
rect 506876 444198 506918 444434
rect 507154 444198 507196 444434
rect 506876 437434 507196 444198
rect 506876 437198 506918 437434
rect 507154 437198 507196 437434
rect 506876 430434 507196 437198
rect 506876 430198 506918 430434
rect 507154 430198 507196 430434
rect 506876 423434 507196 430198
rect 506876 423198 506918 423434
rect 507154 423198 507196 423434
rect 506876 416434 507196 423198
rect 506876 416198 506918 416434
rect 507154 416198 507196 416434
rect 506876 409434 507196 416198
rect 506876 409198 506918 409434
rect 507154 409198 507196 409434
rect 506876 402434 507196 409198
rect 506876 402198 506918 402434
rect 507154 402198 507196 402434
rect 506876 395434 507196 402198
rect 506876 395198 506918 395434
rect 507154 395198 507196 395434
rect 506876 388434 507196 395198
rect 506876 388198 506918 388434
rect 507154 388198 507196 388434
rect 506876 381434 507196 388198
rect 506876 381198 506918 381434
rect 507154 381198 507196 381434
rect 506876 374434 507196 381198
rect 506876 374198 506918 374434
rect 507154 374198 507196 374434
rect 506876 367434 507196 374198
rect 506876 367198 506918 367434
rect 507154 367198 507196 367434
rect 506876 360434 507196 367198
rect 506876 360198 506918 360434
rect 507154 360198 507196 360434
rect 506876 353434 507196 360198
rect 506876 353198 506918 353434
rect 507154 353198 507196 353434
rect 506876 346434 507196 353198
rect 506876 346198 506918 346434
rect 507154 346198 507196 346434
rect 506876 339434 507196 346198
rect 506876 339198 506918 339434
rect 507154 339198 507196 339434
rect 506876 332434 507196 339198
rect 506876 332198 506918 332434
rect 507154 332198 507196 332434
rect 506876 325434 507196 332198
rect 506876 325198 506918 325434
rect 507154 325198 507196 325434
rect 506876 318434 507196 325198
rect 506876 318198 506918 318434
rect 507154 318198 507196 318434
rect 506876 311434 507196 318198
rect 506876 311198 506918 311434
rect 507154 311198 507196 311434
rect 506876 304434 507196 311198
rect 506876 304198 506918 304434
rect 507154 304198 507196 304434
rect 506876 297434 507196 304198
rect 506876 297198 506918 297434
rect 507154 297198 507196 297434
rect 506876 290434 507196 297198
rect 506876 290198 506918 290434
rect 507154 290198 507196 290434
rect 506876 283434 507196 290198
rect 506876 283198 506918 283434
rect 507154 283198 507196 283434
rect 506876 276434 507196 283198
rect 506876 276198 506918 276434
rect 507154 276198 507196 276434
rect 506876 269434 507196 276198
rect 506876 269198 506918 269434
rect 507154 269198 507196 269434
rect 506876 262434 507196 269198
rect 506876 262198 506918 262434
rect 507154 262198 507196 262434
rect 506876 255434 507196 262198
rect 506876 255198 506918 255434
rect 507154 255198 507196 255434
rect 506876 248434 507196 255198
rect 506876 248198 506918 248434
rect 507154 248198 507196 248434
rect 506876 241434 507196 248198
rect 506876 241198 506918 241434
rect 507154 241198 507196 241434
rect 506876 234434 507196 241198
rect 506876 234198 506918 234434
rect 507154 234198 507196 234434
rect 506876 227434 507196 234198
rect 506876 227198 506918 227434
rect 507154 227198 507196 227434
rect 506876 220434 507196 227198
rect 506876 220198 506918 220434
rect 507154 220198 507196 220434
rect 506876 213434 507196 220198
rect 506876 213198 506918 213434
rect 507154 213198 507196 213434
rect 506876 206434 507196 213198
rect 506876 206198 506918 206434
rect 507154 206198 507196 206434
rect 506876 199434 507196 206198
rect 506876 199198 506918 199434
rect 507154 199198 507196 199434
rect 506876 192434 507196 199198
rect 506876 192198 506918 192434
rect 507154 192198 507196 192434
rect 506876 185434 507196 192198
rect 506876 185198 506918 185434
rect 507154 185198 507196 185434
rect 506876 178434 507196 185198
rect 506876 178198 506918 178434
rect 507154 178198 507196 178434
rect 506876 171434 507196 178198
rect 506876 171198 506918 171434
rect 507154 171198 507196 171434
rect 506876 164434 507196 171198
rect 506876 164198 506918 164434
rect 507154 164198 507196 164434
rect 506876 157434 507196 164198
rect 506876 157198 506918 157434
rect 507154 157198 507196 157434
rect 506876 150434 507196 157198
rect 506876 150198 506918 150434
rect 507154 150198 507196 150434
rect 506876 143434 507196 150198
rect 506876 143198 506918 143434
rect 507154 143198 507196 143434
rect 506876 136434 507196 143198
rect 506876 136198 506918 136434
rect 507154 136198 507196 136434
rect 506876 129434 507196 136198
rect 506876 129198 506918 129434
rect 507154 129198 507196 129434
rect 506876 122434 507196 129198
rect 506876 122198 506918 122434
rect 507154 122198 507196 122434
rect 506876 115434 507196 122198
rect 506876 115198 506918 115434
rect 507154 115198 507196 115434
rect 506876 108434 507196 115198
rect 506876 108198 506918 108434
rect 507154 108198 507196 108434
rect 506876 101434 507196 108198
rect 506876 101198 506918 101434
rect 507154 101198 507196 101434
rect 506876 94434 507196 101198
rect 506876 94198 506918 94434
rect 507154 94198 507196 94434
rect 506876 87434 507196 94198
rect 506876 87198 506918 87434
rect 507154 87198 507196 87434
rect 506876 80434 507196 87198
rect 506876 80198 506918 80434
rect 507154 80198 507196 80434
rect 506876 73434 507196 80198
rect 506876 73198 506918 73434
rect 507154 73198 507196 73434
rect 506876 66434 507196 73198
rect 506876 66198 506918 66434
rect 507154 66198 507196 66434
rect 506876 59434 507196 66198
rect 506876 59198 506918 59434
rect 507154 59198 507196 59434
rect 506876 52434 507196 59198
rect 506876 52198 506918 52434
rect 507154 52198 507196 52434
rect 506876 45434 507196 52198
rect 506876 45198 506918 45434
rect 507154 45198 507196 45434
rect 506876 38434 507196 45198
rect 506876 38198 506918 38434
rect 507154 38198 507196 38434
rect 506876 31434 507196 38198
rect 506876 31198 506918 31434
rect 507154 31198 507196 31434
rect 506876 24434 507196 31198
rect 506876 24198 506918 24434
rect 507154 24198 507196 24434
rect 506876 17434 507196 24198
rect 506876 17198 506918 17434
rect 507154 17198 507196 17434
rect 506876 10434 507196 17198
rect 506876 10198 506918 10434
rect 507154 10198 507196 10434
rect 506876 3434 507196 10198
rect 506876 3198 506918 3434
rect 507154 3198 507196 3434
rect 506876 -1706 507196 3198
rect 506876 -1942 506918 -1706
rect 507154 -1942 507196 -1706
rect 506876 -2026 507196 -1942
rect 506876 -2262 506918 -2026
rect 507154 -2262 507196 -2026
rect 506876 -2294 507196 -2262
rect 512144 705238 512464 706230
rect 512144 705002 512186 705238
rect 512422 705002 512464 705238
rect 512144 704918 512464 705002
rect 512144 704682 512186 704918
rect 512422 704682 512464 704918
rect 512144 695494 512464 704682
rect 512144 695258 512186 695494
rect 512422 695258 512464 695494
rect 512144 688494 512464 695258
rect 512144 688258 512186 688494
rect 512422 688258 512464 688494
rect 512144 681494 512464 688258
rect 512144 681258 512186 681494
rect 512422 681258 512464 681494
rect 512144 674494 512464 681258
rect 512144 674258 512186 674494
rect 512422 674258 512464 674494
rect 512144 667494 512464 674258
rect 512144 667258 512186 667494
rect 512422 667258 512464 667494
rect 512144 660494 512464 667258
rect 512144 660258 512186 660494
rect 512422 660258 512464 660494
rect 512144 653494 512464 660258
rect 512144 653258 512186 653494
rect 512422 653258 512464 653494
rect 512144 646494 512464 653258
rect 512144 646258 512186 646494
rect 512422 646258 512464 646494
rect 512144 639494 512464 646258
rect 512144 639258 512186 639494
rect 512422 639258 512464 639494
rect 512144 632494 512464 639258
rect 512144 632258 512186 632494
rect 512422 632258 512464 632494
rect 512144 625494 512464 632258
rect 512144 625258 512186 625494
rect 512422 625258 512464 625494
rect 512144 618494 512464 625258
rect 512144 618258 512186 618494
rect 512422 618258 512464 618494
rect 512144 611494 512464 618258
rect 512144 611258 512186 611494
rect 512422 611258 512464 611494
rect 512144 604494 512464 611258
rect 512144 604258 512186 604494
rect 512422 604258 512464 604494
rect 512144 597494 512464 604258
rect 512144 597258 512186 597494
rect 512422 597258 512464 597494
rect 512144 590494 512464 597258
rect 512144 590258 512186 590494
rect 512422 590258 512464 590494
rect 512144 583494 512464 590258
rect 512144 583258 512186 583494
rect 512422 583258 512464 583494
rect 512144 576494 512464 583258
rect 512144 576258 512186 576494
rect 512422 576258 512464 576494
rect 512144 569494 512464 576258
rect 512144 569258 512186 569494
rect 512422 569258 512464 569494
rect 512144 562494 512464 569258
rect 512144 562258 512186 562494
rect 512422 562258 512464 562494
rect 512144 555494 512464 562258
rect 512144 555258 512186 555494
rect 512422 555258 512464 555494
rect 512144 548494 512464 555258
rect 512144 548258 512186 548494
rect 512422 548258 512464 548494
rect 512144 541494 512464 548258
rect 512144 541258 512186 541494
rect 512422 541258 512464 541494
rect 512144 534494 512464 541258
rect 512144 534258 512186 534494
rect 512422 534258 512464 534494
rect 512144 527494 512464 534258
rect 512144 527258 512186 527494
rect 512422 527258 512464 527494
rect 512144 520494 512464 527258
rect 512144 520258 512186 520494
rect 512422 520258 512464 520494
rect 512144 513494 512464 520258
rect 512144 513258 512186 513494
rect 512422 513258 512464 513494
rect 512144 506494 512464 513258
rect 512144 506258 512186 506494
rect 512422 506258 512464 506494
rect 512144 499494 512464 506258
rect 512144 499258 512186 499494
rect 512422 499258 512464 499494
rect 512144 492494 512464 499258
rect 512144 492258 512186 492494
rect 512422 492258 512464 492494
rect 512144 485494 512464 492258
rect 512144 485258 512186 485494
rect 512422 485258 512464 485494
rect 512144 478494 512464 485258
rect 512144 478258 512186 478494
rect 512422 478258 512464 478494
rect 512144 471494 512464 478258
rect 512144 471258 512186 471494
rect 512422 471258 512464 471494
rect 512144 464494 512464 471258
rect 512144 464258 512186 464494
rect 512422 464258 512464 464494
rect 512144 457494 512464 464258
rect 512144 457258 512186 457494
rect 512422 457258 512464 457494
rect 512144 450494 512464 457258
rect 512144 450258 512186 450494
rect 512422 450258 512464 450494
rect 512144 443494 512464 450258
rect 512144 443258 512186 443494
rect 512422 443258 512464 443494
rect 512144 436494 512464 443258
rect 512144 436258 512186 436494
rect 512422 436258 512464 436494
rect 512144 429494 512464 436258
rect 512144 429258 512186 429494
rect 512422 429258 512464 429494
rect 512144 422494 512464 429258
rect 512144 422258 512186 422494
rect 512422 422258 512464 422494
rect 512144 415494 512464 422258
rect 512144 415258 512186 415494
rect 512422 415258 512464 415494
rect 512144 408494 512464 415258
rect 512144 408258 512186 408494
rect 512422 408258 512464 408494
rect 512144 401494 512464 408258
rect 512144 401258 512186 401494
rect 512422 401258 512464 401494
rect 512144 394494 512464 401258
rect 512144 394258 512186 394494
rect 512422 394258 512464 394494
rect 512144 387494 512464 394258
rect 512144 387258 512186 387494
rect 512422 387258 512464 387494
rect 512144 380494 512464 387258
rect 512144 380258 512186 380494
rect 512422 380258 512464 380494
rect 512144 373494 512464 380258
rect 512144 373258 512186 373494
rect 512422 373258 512464 373494
rect 512144 366494 512464 373258
rect 512144 366258 512186 366494
rect 512422 366258 512464 366494
rect 512144 359494 512464 366258
rect 512144 359258 512186 359494
rect 512422 359258 512464 359494
rect 512144 352494 512464 359258
rect 512144 352258 512186 352494
rect 512422 352258 512464 352494
rect 512144 345494 512464 352258
rect 512144 345258 512186 345494
rect 512422 345258 512464 345494
rect 512144 338494 512464 345258
rect 512144 338258 512186 338494
rect 512422 338258 512464 338494
rect 512144 331494 512464 338258
rect 512144 331258 512186 331494
rect 512422 331258 512464 331494
rect 512144 324494 512464 331258
rect 512144 324258 512186 324494
rect 512422 324258 512464 324494
rect 512144 317494 512464 324258
rect 512144 317258 512186 317494
rect 512422 317258 512464 317494
rect 512144 310494 512464 317258
rect 512144 310258 512186 310494
rect 512422 310258 512464 310494
rect 512144 303494 512464 310258
rect 512144 303258 512186 303494
rect 512422 303258 512464 303494
rect 512144 296494 512464 303258
rect 512144 296258 512186 296494
rect 512422 296258 512464 296494
rect 512144 289494 512464 296258
rect 512144 289258 512186 289494
rect 512422 289258 512464 289494
rect 512144 282494 512464 289258
rect 512144 282258 512186 282494
rect 512422 282258 512464 282494
rect 512144 275494 512464 282258
rect 512144 275258 512186 275494
rect 512422 275258 512464 275494
rect 512144 268494 512464 275258
rect 512144 268258 512186 268494
rect 512422 268258 512464 268494
rect 512144 261494 512464 268258
rect 512144 261258 512186 261494
rect 512422 261258 512464 261494
rect 512144 254494 512464 261258
rect 512144 254258 512186 254494
rect 512422 254258 512464 254494
rect 512144 247494 512464 254258
rect 512144 247258 512186 247494
rect 512422 247258 512464 247494
rect 512144 240494 512464 247258
rect 512144 240258 512186 240494
rect 512422 240258 512464 240494
rect 512144 233494 512464 240258
rect 512144 233258 512186 233494
rect 512422 233258 512464 233494
rect 512144 226494 512464 233258
rect 512144 226258 512186 226494
rect 512422 226258 512464 226494
rect 512144 219494 512464 226258
rect 512144 219258 512186 219494
rect 512422 219258 512464 219494
rect 512144 212494 512464 219258
rect 512144 212258 512186 212494
rect 512422 212258 512464 212494
rect 512144 205494 512464 212258
rect 512144 205258 512186 205494
rect 512422 205258 512464 205494
rect 512144 198494 512464 205258
rect 512144 198258 512186 198494
rect 512422 198258 512464 198494
rect 512144 191494 512464 198258
rect 512144 191258 512186 191494
rect 512422 191258 512464 191494
rect 512144 184494 512464 191258
rect 512144 184258 512186 184494
rect 512422 184258 512464 184494
rect 512144 177494 512464 184258
rect 512144 177258 512186 177494
rect 512422 177258 512464 177494
rect 512144 170494 512464 177258
rect 512144 170258 512186 170494
rect 512422 170258 512464 170494
rect 512144 163494 512464 170258
rect 512144 163258 512186 163494
rect 512422 163258 512464 163494
rect 512144 156494 512464 163258
rect 512144 156258 512186 156494
rect 512422 156258 512464 156494
rect 512144 149494 512464 156258
rect 512144 149258 512186 149494
rect 512422 149258 512464 149494
rect 512144 142494 512464 149258
rect 512144 142258 512186 142494
rect 512422 142258 512464 142494
rect 512144 135494 512464 142258
rect 512144 135258 512186 135494
rect 512422 135258 512464 135494
rect 512144 128494 512464 135258
rect 512144 128258 512186 128494
rect 512422 128258 512464 128494
rect 512144 121494 512464 128258
rect 512144 121258 512186 121494
rect 512422 121258 512464 121494
rect 512144 114494 512464 121258
rect 512144 114258 512186 114494
rect 512422 114258 512464 114494
rect 512144 107494 512464 114258
rect 512144 107258 512186 107494
rect 512422 107258 512464 107494
rect 512144 100494 512464 107258
rect 512144 100258 512186 100494
rect 512422 100258 512464 100494
rect 512144 93494 512464 100258
rect 512144 93258 512186 93494
rect 512422 93258 512464 93494
rect 512144 86494 512464 93258
rect 512144 86258 512186 86494
rect 512422 86258 512464 86494
rect 512144 79494 512464 86258
rect 512144 79258 512186 79494
rect 512422 79258 512464 79494
rect 512144 72494 512464 79258
rect 512144 72258 512186 72494
rect 512422 72258 512464 72494
rect 512144 65494 512464 72258
rect 512144 65258 512186 65494
rect 512422 65258 512464 65494
rect 512144 58494 512464 65258
rect 512144 58258 512186 58494
rect 512422 58258 512464 58494
rect 512144 51494 512464 58258
rect 512144 51258 512186 51494
rect 512422 51258 512464 51494
rect 512144 44494 512464 51258
rect 512144 44258 512186 44494
rect 512422 44258 512464 44494
rect 512144 37494 512464 44258
rect 512144 37258 512186 37494
rect 512422 37258 512464 37494
rect 512144 30494 512464 37258
rect 512144 30258 512186 30494
rect 512422 30258 512464 30494
rect 512144 23494 512464 30258
rect 512144 23258 512186 23494
rect 512422 23258 512464 23494
rect 512144 16494 512464 23258
rect 512144 16258 512186 16494
rect 512422 16258 512464 16494
rect 512144 9494 512464 16258
rect 512144 9258 512186 9494
rect 512422 9258 512464 9494
rect 512144 2494 512464 9258
rect 512144 2258 512186 2494
rect 512422 2258 512464 2494
rect 512144 -746 512464 2258
rect 512144 -982 512186 -746
rect 512422 -982 512464 -746
rect 512144 -1066 512464 -982
rect 512144 -1302 512186 -1066
rect 512422 -1302 512464 -1066
rect 512144 -2294 512464 -1302
rect 513876 706198 514196 706230
rect 513876 705962 513918 706198
rect 514154 705962 514196 706198
rect 513876 705878 514196 705962
rect 513876 705642 513918 705878
rect 514154 705642 514196 705878
rect 513876 696434 514196 705642
rect 513876 696198 513918 696434
rect 514154 696198 514196 696434
rect 513876 689434 514196 696198
rect 513876 689198 513918 689434
rect 514154 689198 514196 689434
rect 513876 682434 514196 689198
rect 513876 682198 513918 682434
rect 514154 682198 514196 682434
rect 513876 675434 514196 682198
rect 513876 675198 513918 675434
rect 514154 675198 514196 675434
rect 513876 668434 514196 675198
rect 513876 668198 513918 668434
rect 514154 668198 514196 668434
rect 513876 661434 514196 668198
rect 513876 661198 513918 661434
rect 514154 661198 514196 661434
rect 513876 654434 514196 661198
rect 513876 654198 513918 654434
rect 514154 654198 514196 654434
rect 513876 647434 514196 654198
rect 513876 647198 513918 647434
rect 514154 647198 514196 647434
rect 513876 640434 514196 647198
rect 513876 640198 513918 640434
rect 514154 640198 514196 640434
rect 513876 633434 514196 640198
rect 513876 633198 513918 633434
rect 514154 633198 514196 633434
rect 513876 626434 514196 633198
rect 513876 626198 513918 626434
rect 514154 626198 514196 626434
rect 513876 619434 514196 626198
rect 513876 619198 513918 619434
rect 514154 619198 514196 619434
rect 513876 612434 514196 619198
rect 513876 612198 513918 612434
rect 514154 612198 514196 612434
rect 513876 605434 514196 612198
rect 513876 605198 513918 605434
rect 514154 605198 514196 605434
rect 513876 598434 514196 605198
rect 513876 598198 513918 598434
rect 514154 598198 514196 598434
rect 513876 591434 514196 598198
rect 513876 591198 513918 591434
rect 514154 591198 514196 591434
rect 513876 584434 514196 591198
rect 513876 584198 513918 584434
rect 514154 584198 514196 584434
rect 513876 577434 514196 584198
rect 513876 577198 513918 577434
rect 514154 577198 514196 577434
rect 513876 570434 514196 577198
rect 513876 570198 513918 570434
rect 514154 570198 514196 570434
rect 513876 563434 514196 570198
rect 513876 563198 513918 563434
rect 514154 563198 514196 563434
rect 513876 556434 514196 563198
rect 513876 556198 513918 556434
rect 514154 556198 514196 556434
rect 513876 549434 514196 556198
rect 513876 549198 513918 549434
rect 514154 549198 514196 549434
rect 513876 542434 514196 549198
rect 513876 542198 513918 542434
rect 514154 542198 514196 542434
rect 513876 535434 514196 542198
rect 513876 535198 513918 535434
rect 514154 535198 514196 535434
rect 513876 528434 514196 535198
rect 513876 528198 513918 528434
rect 514154 528198 514196 528434
rect 513876 521434 514196 528198
rect 513876 521198 513918 521434
rect 514154 521198 514196 521434
rect 513876 514434 514196 521198
rect 513876 514198 513918 514434
rect 514154 514198 514196 514434
rect 513876 507434 514196 514198
rect 513876 507198 513918 507434
rect 514154 507198 514196 507434
rect 513876 500434 514196 507198
rect 513876 500198 513918 500434
rect 514154 500198 514196 500434
rect 513876 493434 514196 500198
rect 513876 493198 513918 493434
rect 514154 493198 514196 493434
rect 513876 486434 514196 493198
rect 513876 486198 513918 486434
rect 514154 486198 514196 486434
rect 513876 479434 514196 486198
rect 513876 479198 513918 479434
rect 514154 479198 514196 479434
rect 513876 472434 514196 479198
rect 513876 472198 513918 472434
rect 514154 472198 514196 472434
rect 513876 465434 514196 472198
rect 513876 465198 513918 465434
rect 514154 465198 514196 465434
rect 513876 458434 514196 465198
rect 513876 458198 513918 458434
rect 514154 458198 514196 458434
rect 513876 451434 514196 458198
rect 513876 451198 513918 451434
rect 514154 451198 514196 451434
rect 513876 444434 514196 451198
rect 513876 444198 513918 444434
rect 514154 444198 514196 444434
rect 513876 437434 514196 444198
rect 513876 437198 513918 437434
rect 514154 437198 514196 437434
rect 513876 430434 514196 437198
rect 513876 430198 513918 430434
rect 514154 430198 514196 430434
rect 513876 423434 514196 430198
rect 513876 423198 513918 423434
rect 514154 423198 514196 423434
rect 513876 416434 514196 423198
rect 513876 416198 513918 416434
rect 514154 416198 514196 416434
rect 513876 409434 514196 416198
rect 513876 409198 513918 409434
rect 514154 409198 514196 409434
rect 513876 402434 514196 409198
rect 513876 402198 513918 402434
rect 514154 402198 514196 402434
rect 513876 395434 514196 402198
rect 513876 395198 513918 395434
rect 514154 395198 514196 395434
rect 513876 388434 514196 395198
rect 513876 388198 513918 388434
rect 514154 388198 514196 388434
rect 513876 381434 514196 388198
rect 513876 381198 513918 381434
rect 514154 381198 514196 381434
rect 513876 374434 514196 381198
rect 513876 374198 513918 374434
rect 514154 374198 514196 374434
rect 513876 367434 514196 374198
rect 513876 367198 513918 367434
rect 514154 367198 514196 367434
rect 513876 360434 514196 367198
rect 513876 360198 513918 360434
rect 514154 360198 514196 360434
rect 513876 353434 514196 360198
rect 513876 353198 513918 353434
rect 514154 353198 514196 353434
rect 513876 346434 514196 353198
rect 513876 346198 513918 346434
rect 514154 346198 514196 346434
rect 513876 339434 514196 346198
rect 513876 339198 513918 339434
rect 514154 339198 514196 339434
rect 513876 332434 514196 339198
rect 513876 332198 513918 332434
rect 514154 332198 514196 332434
rect 513876 325434 514196 332198
rect 513876 325198 513918 325434
rect 514154 325198 514196 325434
rect 513876 318434 514196 325198
rect 513876 318198 513918 318434
rect 514154 318198 514196 318434
rect 513876 311434 514196 318198
rect 513876 311198 513918 311434
rect 514154 311198 514196 311434
rect 513876 304434 514196 311198
rect 513876 304198 513918 304434
rect 514154 304198 514196 304434
rect 513876 297434 514196 304198
rect 513876 297198 513918 297434
rect 514154 297198 514196 297434
rect 513876 290434 514196 297198
rect 513876 290198 513918 290434
rect 514154 290198 514196 290434
rect 513876 283434 514196 290198
rect 513876 283198 513918 283434
rect 514154 283198 514196 283434
rect 513876 276434 514196 283198
rect 513876 276198 513918 276434
rect 514154 276198 514196 276434
rect 513876 269434 514196 276198
rect 513876 269198 513918 269434
rect 514154 269198 514196 269434
rect 513876 262434 514196 269198
rect 513876 262198 513918 262434
rect 514154 262198 514196 262434
rect 513876 255434 514196 262198
rect 513876 255198 513918 255434
rect 514154 255198 514196 255434
rect 513876 248434 514196 255198
rect 513876 248198 513918 248434
rect 514154 248198 514196 248434
rect 513876 241434 514196 248198
rect 513876 241198 513918 241434
rect 514154 241198 514196 241434
rect 513876 234434 514196 241198
rect 513876 234198 513918 234434
rect 514154 234198 514196 234434
rect 513876 227434 514196 234198
rect 513876 227198 513918 227434
rect 514154 227198 514196 227434
rect 513876 220434 514196 227198
rect 513876 220198 513918 220434
rect 514154 220198 514196 220434
rect 513876 213434 514196 220198
rect 513876 213198 513918 213434
rect 514154 213198 514196 213434
rect 513876 206434 514196 213198
rect 513876 206198 513918 206434
rect 514154 206198 514196 206434
rect 513876 199434 514196 206198
rect 513876 199198 513918 199434
rect 514154 199198 514196 199434
rect 513876 192434 514196 199198
rect 513876 192198 513918 192434
rect 514154 192198 514196 192434
rect 513876 185434 514196 192198
rect 513876 185198 513918 185434
rect 514154 185198 514196 185434
rect 513876 178434 514196 185198
rect 513876 178198 513918 178434
rect 514154 178198 514196 178434
rect 513876 171434 514196 178198
rect 513876 171198 513918 171434
rect 514154 171198 514196 171434
rect 513876 164434 514196 171198
rect 513876 164198 513918 164434
rect 514154 164198 514196 164434
rect 513876 157434 514196 164198
rect 513876 157198 513918 157434
rect 514154 157198 514196 157434
rect 513876 150434 514196 157198
rect 513876 150198 513918 150434
rect 514154 150198 514196 150434
rect 513876 143434 514196 150198
rect 513876 143198 513918 143434
rect 514154 143198 514196 143434
rect 513876 136434 514196 143198
rect 513876 136198 513918 136434
rect 514154 136198 514196 136434
rect 513876 129434 514196 136198
rect 513876 129198 513918 129434
rect 514154 129198 514196 129434
rect 513876 122434 514196 129198
rect 513876 122198 513918 122434
rect 514154 122198 514196 122434
rect 513876 115434 514196 122198
rect 513876 115198 513918 115434
rect 514154 115198 514196 115434
rect 513876 108434 514196 115198
rect 513876 108198 513918 108434
rect 514154 108198 514196 108434
rect 513876 101434 514196 108198
rect 513876 101198 513918 101434
rect 514154 101198 514196 101434
rect 513876 94434 514196 101198
rect 513876 94198 513918 94434
rect 514154 94198 514196 94434
rect 513876 87434 514196 94198
rect 513876 87198 513918 87434
rect 514154 87198 514196 87434
rect 513876 80434 514196 87198
rect 513876 80198 513918 80434
rect 514154 80198 514196 80434
rect 513876 73434 514196 80198
rect 513876 73198 513918 73434
rect 514154 73198 514196 73434
rect 513876 66434 514196 73198
rect 513876 66198 513918 66434
rect 514154 66198 514196 66434
rect 513876 59434 514196 66198
rect 513876 59198 513918 59434
rect 514154 59198 514196 59434
rect 513876 52434 514196 59198
rect 513876 52198 513918 52434
rect 514154 52198 514196 52434
rect 513876 45434 514196 52198
rect 513876 45198 513918 45434
rect 514154 45198 514196 45434
rect 513876 38434 514196 45198
rect 513876 38198 513918 38434
rect 514154 38198 514196 38434
rect 513876 31434 514196 38198
rect 513876 31198 513918 31434
rect 514154 31198 514196 31434
rect 513876 24434 514196 31198
rect 513876 24198 513918 24434
rect 514154 24198 514196 24434
rect 513876 17434 514196 24198
rect 513876 17198 513918 17434
rect 514154 17198 514196 17434
rect 513876 10434 514196 17198
rect 513876 10198 513918 10434
rect 514154 10198 514196 10434
rect 513876 3434 514196 10198
rect 513876 3198 513918 3434
rect 514154 3198 514196 3434
rect 513876 -1706 514196 3198
rect 513876 -1942 513918 -1706
rect 514154 -1942 514196 -1706
rect 513876 -2026 514196 -1942
rect 513876 -2262 513918 -2026
rect 514154 -2262 514196 -2026
rect 513876 -2294 514196 -2262
rect 519144 705238 519464 706230
rect 519144 705002 519186 705238
rect 519422 705002 519464 705238
rect 519144 704918 519464 705002
rect 519144 704682 519186 704918
rect 519422 704682 519464 704918
rect 519144 695494 519464 704682
rect 519144 695258 519186 695494
rect 519422 695258 519464 695494
rect 519144 688494 519464 695258
rect 519144 688258 519186 688494
rect 519422 688258 519464 688494
rect 519144 681494 519464 688258
rect 519144 681258 519186 681494
rect 519422 681258 519464 681494
rect 519144 674494 519464 681258
rect 519144 674258 519186 674494
rect 519422 674258 519464 674494
rect 519144 667494 519464 674258
rect 519144 667258 519186 667494
rect 519422 667258 519464 667494
rect 519144 660494 519464 667258
rect 519144 660258 519186 660494
rect 519422 660258 519464 660494
rect 519144 653494 519464 660258
rect 519144 653258 519186 653494
rect 519422 653258 519464 653494
rect 519144 646494 519464 653258
rect 519144 646258 519186 646494
rect 519422 646258 519464 646494
rect 519144 639494 519464 646258
rect 519144 639258 519186 639494
rect 519422 639258 519464 639494
rect 519144 632494 519464 639258
rect 519144 632258 519186 632494
rect 519422 632258 519464 632494
rect 519144 625494 519464 632258
rect 519144 625258 519186 625494
rect 519422 625258 519464 625494
rect 519144 618494 519464 625258
rect 519144 618258 519186 618494
rect 519422 618258 519464 618494
rect 519144 611494 519464 618258
rect 519144 611258 519186 611494
rect 519422 611258 519464 611494
rect 519144 604494 519464 611258
rect 519144 604258 519186 604494
rect 519422 604258 519464 604494
rect 519144 597494 519464 604258
rect 519144 597258 519186 597494
rect 519422 597258 519464 597494
rect 519144 590494 519464 597258
rect 519144 590258 519186 590494
rect 519422 590258 519464 590494
rect 519144 583494 519464 590258
rect 519144 583258 519186 583494
rect 519422 583258 519464 583494
rect 519144 576494 519464 583258
rect 519144 576258 519186 576494
rect 519422 576258 519464 576494
rect 519144 569494 519464 576258
rect 519144 569258 519186 569494
rect 519422 569258 519464 569494
rect 519144 562494 519464 569258
rect 519144 562258 519186 562494
rect 519422 562258 519464 562494
rect 519144 555494 519464 562258
rect 519144 555258 519186 555494
rect 519422 555258 519464 555494
rect 519144 548494 519464 555258
rect 519144 548258 519186 548494
rect 519422 548258 519464 548494
rect 519144 541494 519464 548258
rect 519144 541258 519186 541494
rect 519422 541258 519464 541494
rect 519144 534494 519464 541258
rect 519144 534258 519186 534494
rect 519422 534258 519464 534494
rect 519144 527494 519464 534258
rect 519144 527258 519186 527494
rect 519422 527258 519464 527494
rect 519144 520494 519464 527258
rect 519144 520258 519186 520494
rect 519422 520258 519464 520494
rect 519144 513494 519464 520258
rect 519144 513258 519186 513494
rect 519422 513258 519464 513494
rect 519144 506494 519464 513258
rect 519144 506258 519186 506494
rect 519422 506258 519464 506494
rect 519144 499494 519464 506258
rect 519144 499258 519186 499494
rect 519422 499258 519464 499494
rect 519144 492494 519464 499258
rect 519144 492258 519186 492494
rect 519422 492258 519464 492494
rect 519144 485494 519464 492258
rect 519144 485258 519186 485494
rect 519422 485258 519464 485494
rect 519144 478494 519464 485258
rect 519144 478258 519186 478494
rect 519422 478258 519464 478494
rect 519144 471494 519464 478258
rect 519144 471258 519186 471494
rect 519422 471258 519464 471494
rect 519144 464494 519464 471258
rect 519144 464258 519186 464494
rect 519422 464258 519464 464494
rect 519144 457494 519464 464258
rect 519144 457258 519186 457494
rect 519422 457258 519464 457494
rect 519144 450494 519464 457258
rect 519144 450258 519186 450494
rect 519422 450258 519464 450494
rect 519144 443494 519464 450258
rect 519144 443258 519186 443494
rect 519422 443258 519464 443494
rect 519144 436494 519464 443258
rect 519144 436258 519186 436494
rect 519422 436258 519464 436494
rect 519144 429494 519464 436258
rect 519144 429258 519186 429494
rect 519422 429258 519464 429494
rect 519144 422494 519464 429258
rect 519144 422258 519186 422494
rect 519422 422258 519464 422494
rect 519144 415494 519464 422258
rect 520876 706198 521196 706230
rect 520876 705962 520918 706198
rect 521154 705962 521196 706198
rect 520876 705878 521196 705962
rect 520876 705642 520918 705878
rect 521154 705642 521196 705878
rect 520876 696434 521196 705642
rect 520876 696198 520918 696434
rect 521154 696198 521196 696434
rect 520876 689434 521196 696198
rect 520876 689198 520918 689434
rect 521154 689198 521196 689434
rect 520876 682434 521196 689198
rect 520876 682198 520918 682434
rect 521154 682198 521196 682434
rect 520876 675434 521196 682198
rect 520876 675198 520918 675434
rect 521154 675198 521196 675434
rect 520876 668434 521196 675198
rect 520876 668198 520918 668434
rect 521154 668198 521196 668434
rect 520876 661434 521196 668198
rect 520876 661198 520918 661434
rect 521154 661198 521196 661434
rect 520876 654434 521196 661198
rect 520876 654198 520918 654434
rect 521154 654198 521196 654434
rect 520876 647434 521196 654198
rect 520876 647198 520918 647434
rect 521154 647198 521196 647434
rect 520876 640434 521196 647198
rect 520876 640198 520918 640434
rect 521154 640198 521196 640434
rect 520876 633434 521196 640198
rect 520876 633198 520918 633434
rect 521154 633198 521196 633434
rect 520876 626434 521196 633198
rect 520876 626198 520918 626434
rect 521154 626198 521196 626434
rect 520876 619434 521196 626198
rect 520876 619198 520918 619434
rect 521154 619198 521196 619434
rect 520876 612434 521196 619198
rect 520876 612198 520918 612434
rect 521154 612198 521196 612434
rect 520876 605434 521196 612198
rect 520876 605198 520918 605434
rect 521154 605198 521196 605434
rect 520876 598434 521196 605198
rect 520876 598198 520918 598434
rect 521154 598198 521196 598434
rect 520876 591434 521196 598198
rect 520876 591198 520918 591434
rect 521154 591198 521196 591434
rect 520876 584434 521196 591198
rect 520876 584198 520918 584434
rect 521154 584198 521196 584434
rect 520876 577434 521196 584198
rect 520876 577198 520918 577434
rect 521154 577198 521196 577434
rect 520876 570434 521196 577198
rect 520876 570198 520918 570434
rect 521154 570198 521196 570434
rect 520876 563434 521196 570198
rect 520876 563198 520918 563434
rect 521154 563198 521196 563434
rect 520876 556434 521196 563198
rect 520876 556198 520918 556434
rect 521154 556198 521196 556434
rect 520876 549434 521196 556198
rect 520876 549198 520918 549434
rect 521154 549198 521196 549434
rect 520876 542434 521196 549198
rect 520876 542198 520918 542434
rect 521154 542198 521196 542434
rect 520876 535434 521196 542198
rect 520876 535198 520918 535434
rect 521154 535198 521196 535434
rect 520876 528434 521196 535198
rect 520876 528198 520918 528434
rect 521154 528198 521196 528434
rect 520876 521434 521196 528198
rect 520876 521198 520918 521434
rect 521154 521198 521196 521434
rect 520876 514434 521196 521198
rect 520876 514198 520918 514434
rect 521154 514198 521196 514434
rect 520876 507434 521196 514198
rect 520876 507198 520918 507434
rect 521154 507198 521196 507434
rect 520876 500434 521196 507198
rect 520876 500198 520918 500434
rect 521154 500198 521196 500434
rect 520876 493434 521196 500198
rect 520876 493198 520918 493434
rect 521154 493198 521196 493434
rect 520876 486434 521196 493198
rect 520876 486198 520918 486434
rect 521154 486198 521196 486434
rect 520876 479434 521196 486198
rect 520876 479198 520918 479434
rect 521154 479198 521196 479434
rect 520876 472434 521196 479198
rect 520876 472198 520918 472434
rect 521154 472198 521196 472434
rect 520876 465434 521196 472198
rect 520876 465198 520918 465434
rect 521154 465198 521196 465434
rect 520876 458434 521196 465198
rect 520876 458198 520918 458434
rect 521154 458198 521196 458434
rect 520876 451434 521196 458198
rect 520876 451198 520918 451434
rect 521154 451198 521196 451434
rect 520876 444434 521196 451198
rect 520876 444198 520918 444434
rect 521154 444198 521196 444434
rect 520876 437434 521196 444198
rect 520876 437198 520918 437434
rect 521154 437198 521196 437434
rect 520876 430434 521196 437198
rect 520876 430198 520918 430434
rect 521154 430198 521196 430434
rect 520876 423434 521196 430198
rect 520876 423198 520918 423434
rect 521154 423198 521196 423434
rect 520876 421752 521196 423198
rect 526144 705238 526464 706230
rect 526144 705002 526186 705238
rect 526422 705002 526464 705238
rect 526144 704918 526464 705002
rect 526144 704682 526186 704918
rect 526422 704682 526464 704918
rect 526144 695494 526464 704682
rect 526144 695258 526186 695494
rect 526422 695258 526464 695494
rect 526144 688494 526464 695258
rect 526144 688258 526186 688494
rect 526422 688258 526464 688494
rect 526144 681494 526464 688258
rect 526144 681258 526186 681494
rect 526422 681258 526464 681494
rect 526144 674494 526464 681258
rect 526144 674258 526186 674494
rect 526422 674258 526464 674494
rect 526144 667494 526464 674258
rect 526144 667258 526186 667494
rect 526422 667258 526464 667494
rect 526144 660494 526464 667258
rect 526144 660258 526186 660494
rect 526422 660258 526464 660494
rect 526144 653494 526464 660258
rect 526144 653258 526186 653494
rect 526422 653258 526464 653494
rect 526144 646494 526464 653258
rect 526144 646258 526186 646494
rect 526422 646258 526464 646494
rect 526144 639494 526464 646258
rect 526144 639258 526186 639494
rect 526422 639258 526464 639494
rect 526144 632494 526464 639258
rect 526144 632258 526186 632494
rect 526422 632258 526464 632494
rect 526144 625494 526464 632258
rect 526144 625258 526186 625494
rect 526422 625258 526464 625494
rect 526144 618494 526464 625258
rect 526144 618258 526186 618494
rect 526422 618258 526464 618494
rect 526144 611494 526464 618258
rect 526144 611258 526186 611494
rect 526422 611258 526464 611494
rect 526144 604494 526464 611258
rect 526144 604258 526186 604494
rect 526422 604258 526464 604494
rect 526144 597494 526464 604258
rect 526144 597258 526186 597494
rect 526422 597258 526464 597494
rect 526144 590494 526464 597258
rect 526144 590258 526186 590494
rect 526422 590258 526464 590494
rect 526144 583494 526464 590258
rect 526144 583258 526186 583494
rect 526422 583258 526464 583494
rect 526144 576494 526464 583258
rect 526144 576258 526186 576494
rect 526422 576258 526464 576494
rect 526144 569494 526464 576258
rect 526144 569258 526186 569494
rect 526422 569258 526464 569494
rect 526144 562494 526464 569258
rect 526144 562258 526186 562494
rect 526422 562258 526464 562494
rect 526144 555494 526464 562258
rect 526144 555258 526186 555494
rect 526422 555258 526464 555494
rect 526144 548494 526464 555258
rect 526144 548258 526186 548494
rect 526422 548258 526464 548494
rect 526144 541494 526464 548258
rect 526144 541258 526186 541494
rect 526422 541258 526464 541494
rect 526144 534494 526464 541258
rect 526144 534258 526186 534494
rect 526422 534258 526464 534494
rect 526144 527494 526464 534258
rect 526144 527258 526186 527494
rect 526422 527258 526464 527494
rect 526144 520494 526464 527258
rect 526144 520258 526186 520494
rect 526422 520258 526464 520494
rect 526144 513494 526464 520258
rect 526144 513258 526186 513494
rect 526422 513258 526464 513494
rect 526144 506494 526464 513258
rect 526144 506258 526186 506494
rect 526422 506258 526464 506494
rect 526144 499494 526464 506258
rect 526144 499258 526186 499494
rect 526422 499258 526464 499494
rect 526144 492494 526464 499258
rect 526144 492258 526186 492494
rect 526422 492258 526464 492494
rect 526144 485494 526464 492258
rect 526144 485258 526186 485494
rect 526422 485258 526464 485494
rect 526144 478494 526464 485258
rect 526144 478258 526186 478494
rect 526422 478258 526464 478494
rect 526144 471494 526464 478258
rect 526144 471258 526186 471494
rect 526422 471258 526464 471494
rect 526144 464494 526464 471258
rect 526144 464258 526186 464494
rect 526422 464258 526464 464494
rect 526144 457494 526464 464258
rect 526144 457258 526186 457494
rect 526422 457258 526464 457494
rect 526144 450494 526464 457258
rect 526144 450258 526186 450494
rect 526422 450258 526464 450494
rect 526144 443494 526464 450258
rect 526144 443258 526186 443494
rect 526422 443258 526464 443494
rect 526144 436494 526464 443258
rect 526144 436258 526186 436494
rect 526422 436258 526464 436494
rect 526144 429494 526464 436258
rect 526144 429258 526186 429494
rect 526422 429258 526464 429494
rect 526144 422494 526464 429258
rect 526144 422258 526186 422494
rect 526422 422258 526464 422494
rect 526144 421752 526464 422258
rect 527876 706198 528196 706230
rect 527876 705962 527918 706198
rect 528154 705962 528196 706198
rect 527876 705878 528196 705962
rect 527876 705642 527918 705878
rect 528154 705642 528196 705878
rect 527876 696434 528196 705642
rect 527876 696198 527918 696434
rect 528154 696198 528196 696434
rect 527876 689434 528196 696198
rect 527876 689198 527918 689434
rect 528154 689198 528196 689434
rect 527876 682434 528196 689198
rect 527876 682198 527918 682434
rect 528154 682198 528196 682434
rect 527876 675434 528196 682198
rect 527876 675198 527918 675434
rect 528154 675198 528196 675434
rect 527876 668434 528196 675198
rect 527876 668198 527918 668434
rect 528154 668198 528196 668434
rect 527876 661434 528196 668198
rect 527876 661198 527918 661434
rect 528154 661198 528196 661434
rect 527876 654434 528196 661198
rect 527876 654198 527918 654434
rect 528154 654198 528196 654434
rect 527876 647434 528196 654198
rect 527876 647198 527918 647434
rect 528154 647198 528196 647434
rect 527876 640434 528196 647198
rect 527876 640198 527918 640434
rect 528154 640198 528196 640434
rect 527876 633434 528196 640198
rect 527876 633198 527918 633434
rect 528154 633198 528196 633434
rect 527876 626434 528196 633198
rect 527876 626198 527918 626434
rect 528154 626198 528196 626434
rect 527876 619434 528196 626198
rect 527876 619198 527918 619434
rect 528154 619198 528196 619434
rect 527876 612434 528196 619198
rect 527876 612198 527918 612434
rect 528154 612198 528196 612434
rect 527876 605434 528196 612198
rect 527876 605198 527918 605434
rect 528154 605198 528196 605434
rect 527876 598434 528196 605198
rect 527876 598198 527918 598434
rect 528154 598198 528196 598434
rect 527876 591434 528196 598198
rect 527876 591198 527918 591434
rect 528154 591198 528196 591434
rect 527876 584434 528196 591198
rect 527876 584198 527918 584434
rect 528154 584198 528196 584434
rect 527876 577434 528196 584198
rect 527876 577198 527918 577434
rect 528154 577198 528196 577434
rect 527876 570434 528196 577198
rect 527876 570198 527918 570434
rect 528154 570198 528196 570434
rect 527876 563434 528196 570198
rect 527876 563198 527918 563434
rect 528154 563198 528196 563434
rect 527876 556434 528196 563198
rect 527876 556198 527918 556434
rect 528154 556198 528196 556434
rect 527876 549434 528196 556198
rect 527876 549198 527918 549434
rect 528154 549198 528196 549434
rect 527876 542434 528196 549198
rect 527876 542198 527918 542434
rect 528154 542198 528196 542434
rect 527876 535434 528196 542198
rect 527876 535198 527918 535434
rect 528154 535198 528196 535434
rect 527876 528434 528196 535198
rect 527876 528198 527918 528434
rect 528154 528198 528196 528434
rect 527876 521434 528196 528198
rect 527876 521198 527918 521434
rect 528154 521198 528196 521434
rect 527876 514434 528196 521198
rect 527876 514198 527918 514434
rect 528154 514198 528196 514434
rect 527876 507434 528196 514198
rect 527876 507198 527918 507434
rect 528154 507198 528196 507434
rect 527876 500434 528196 507198
rect 527876 500198 527918 500434
rect 528154 500198 528196 500434
rect 527876 493434 528196 500198
rect 527876 493198 527918 493434
rect 528154 493198 528196 493434
rect 527876 486434 528196 493198
rect 527876 486198 527918 486434
rect 528154 486198 528196 486434
rect 527876 479434 528196 486198
rect 527876 479198 527918 479434
rect 528154 479198 528196 479434
rect 527876 472434 528196 479198
rect 527876 472198 527918 472434
rect 528154 472198 528196 472434
rect 527876 465434 528196 472198
rect 527876 465198 527918 465434
rect 528154 465198 528196 465434
rect 527876 458434 528196 465198
rect 527876 458198 527918 458434
rect 528154 458198 528196 458434
rect 527876 451434 528196 458198
rect 527876 451198 527918 451434
rect 528154 451198 528196 451434
rect 527876 444434 528196 451198
rect 527876 444198 527918 444434
rect 528154 444198 528196 444434
rect 527876 437434 528196 444198
rect 527876 437198 527918 437434
rect 528154 437198 528196 437434
rect 527876 430434 528196 437198
rect 527876 430198 527918 430434
rect 528154 430198 528196 430434
rect 527876 423434 528196 430198
rect 527876 423198 527918 423434
rect 528154 423198 528196 423434
rect 527876 416434 528196 423198
rect 520876 416198 520918 416434
rect 521154 416198 521196 416434
rect 522808 416198 522850 416434
rect 523086 416198 523128 416434
rect 524740 416198 524782 416434
rect 525018 416198 525060 416434
rect 526672 416198 526714 416434
rect 526950 416198 526992 416434
rect 527876 416198 527918 416434
rect 528154 416198 528196 416434
rect 519144 415258 519186 415494
rect 519422 415258 519464 415494
rect 519910 415258 519952 415494
rect 520188 415258 520230 415494
rect 521842 415258 521884 415494
rect 522120 415258 522162 415494
rect 523774 415258 523816 415494
rect 524052 415258 524094 415494
rect 525706 415258 525748 415494
rect 525984 415258 526026 415494
rect 519144 408494 519464 415258
rect 527876 409434 528196 416198
rect 520876 409198 520918 409434
rect 521154 409198 521196 409434
rect 522808 409198 522850 409434
rect 523086 409198 523128 409434
rect 524740 409198 524782 409434
rect 525018 409198 525060 409434
rect 526672 409198 526714 409434
rect 526950 409198 526992 409434
rect 527876 409198 527918 409434
rect 528154 409198 528196 409434
rect 519144 408258 519186 408494
rect 519422 408258 519464 408494
rect 519910 408258 519952 408494
rect 520188 408258 520230 408494
rect 521842 408258 521884 408494
rect 522120 408258 522162 408494
rect 523774 408258 523816 408494
rect 524052 408258 524094 408494
rect 525706 408258 525748 408494
rect 525984 408258 526026 408494
rect 519144 401494 519464 408258
rect 527876 402434 528196 409198
rect 520876 402198 520918 402434
rect 521154 402198 521196 402434
rect 522808 402198 522850 402434
rect 523086 402198 523128 402434
rect 524740 402198 524782 402434
rect 525018 402198 525060 402434
rect 526672 402198 526714 402434
rect 526950 402198 526992 402434
rect 527876 402198 527918 402434
rect 528154 402198 528196 402434
rect 519144 401258 519186 401494
rect 519422 401258 519464 401494
rect 519144 394494 519464 401258
rect 519144 394258 519186 394494
rect 519422 394258 519464 394494
rect 519144 387494 519464 394258
rect 519144 387258 519186 387494
rect 519422 387258 519464 387494
rect 519144 380494 519464 387258
rect 520876 395434 521196 400008
rect 520876 395198 520918 395434
rect 521154 395198 521196 395434
rect 520876 388434 521196 395198
rect 520876 388198 520918 388434
rect 521154 388198 521196 388434
rect 520876 381752 521196 388198
rect 526144 394494 526464 400008
rect 526144 394258 526186 394494
rect 526422 394258 526464 394494
rect 526144 387494 526464 394258
rect 526144 387258 526186 387494
rect 526422 387258 526464 387494
rect 526144 381752 526464 387258
rect 527876 395434 528196 402198
rect 527876 395198 527918 395434
rect 528154 395198 528196 395434
rect 527876 388434 528196 395198
rect 527876 388198 527918 388434
rect 528154 388198 528196 388434
rect 519144 380258 519186 380494
rect 519422 380258 519464 380494
rect 519144 373494 519464 380258
rect 527876 381434 528196 388198
rect 527876 381198 527918 381434
rect 528154 381198 528196 381434
rect 527876 374434 528196 381198
rect 520876 374198 520918 374434
rect 521154 374198 521196 374434
rect 522808 374198 522850 374434
rect 523086 374198 523128 374434
rect 524740 374198 524782 374434
rect 525018 374198 525060 374434
rect 526672 374198 526714 374434
rect 526950 374198 526992 374434
rect 527876 374198 527918 374434
rect 528154 374198 528196 374434
rect 519144 373258 519186 373494
rect 519422 373258 519464 373494
rect 519910 373258 519952 373494
rect 520188 373258 520230 373494
rect 521842 373258 521884 373494
rect 522120 373258 522162 373494
rect 523774 373258 523816 373494
rect 524052 373258 524094 373494
rect 525706 373258 525748 373494
rect 525984 373258 526026 373494
rect 519144 366494 519464 373258
rect 527876 367434 528196 374198
rect 520876 367198 520918 367434
rect 521154 367198 521196 367434
rect 522808 367198 522850 367434
rect 523086 367198 523128 367434
rect 524740 367198 524782 367434
rect 525018 367198 525060 367434
rect 526672 367198 526714 367434
rect 526950 367198 526992 367434
rect 527876 367198 527918 367434
rect 528154 367198 528196 367434
rect 519144 366258 519186 366494
rect 519422 366258 519464 366494
rect 519910 366258 519952 366494
rect 520188 366258 520230 366494
rect 521842 366258 521884 366494
rect 522120 366258 522162 366494
rect 523774 366258 523816 366494
rect 524052 366258 524094 366494
rect 525706 366258 525748 366494
rect 525984 366258 526026 366494
rect 519144 359494 519464 366258
rect 527876 360434 528196 367198
rect 527876 360198 527918 360434
rect 528154 360198 528196 360434
rect 519144 359258 519186 359494
rect 519422 359258 519464 359494
rect 519144 352494 519464 359258
rect 519144 352258 519186 352494
rect 519422 352258 519464 352494
rect 519144 345494 519464 352258
rect 519144 345258 519186 345494
rect 519422 345258 519464 345494
rect 519144 338494 519464 345258
rect 520876 353434 521196 360008
rect 520876 353198 520918 353434
rect 521154 353198 521196 353434
rect 520876 346434 521196 353198
rect 520876 346198 520918 346434
rect 521154 346198 521196 346434
rect 520876 341752 521196 346198
rect 526144 359494 526464 360008
rect 526144 359258 526186 359494
rect 526422 359258 526464 359494
rect 526144 352494 526464 359258
rect 526144 352258 526186 352494
rect 526422 352258 526464 352494
rect 526144 345494 526464 352258
rect 526144 345258 526186 345494
rect 526422 345258 526464 345494
rect 526144 341752 526464 345258
rect 527876 353434 528196 360198
rect 527876 353198 527918 353434
rect 528154 353198 528196 353434
rect 527876 346434 528196 353198
rect 527876 346198 527918 346434
rect 528154 346198 528196 346434
rect 527876 339434 528196 346198
rect 520876 339198 520918 339434
rect 521154 339198 521196 339434
rect 522808 339198 522850 339434
rect 523086 339198 523128 339434
rect 524740 339198 524782 339434
rect 525018 339198 525060 339434
rect 526672 339198 526714 339434
rect 526950 339198 526992 339434
rect 527876 339198 527918 339434
rect 528154 339198 528196 339434
rect 519144 338258 519186 338494
rect 519422 338258 519464 338494
rect 519910 338258 519952 338494
rect 520188 338258 520230 338494
rect 521842 338258 521884 338494
rect 522120 338258 522162 338494
rect 523774 338258 523816 338494
rect 524052 338258 524094 338494
rect 525706 338258 525748 338494
rect 525984 338258 526026 338494
rect 519144 331494 519464 338258
rect 527876 332434 528196 339198
rect 520876 332198 520918 332434
rect 521154 332198 521196 332434
rect 522808 332198 522850 332434
rect 523086 332198 523128 332434
rect 524740 332198 524782 332434
rect 525018 332198 525060 332434
rect 526672 332198 526714 332434
rect 526950 332198 526992 332434
rect 527876 332198 527918 332434
rect 528154 332198 528196 332434
rect 519144 331258 519186 331494
rect 519422 331258 519464 331494
rect 519910 331258 519952 331494
rect 520188 331258 520230 331494
rect 521842 331258 521884 331494
rect 522120 331258 522162 331494
rect 523774 331258 523816 331494
rect 524052 331258 524094 331494
rect 525706 331258 525748 331494
rect 525984 331258 526026 331494
rect 519144 324494 519464 331258
rect 527876 325434 528196 332198
rect 520876 325198 520918 325434
rect 521154 325198 521196 325434
rect 522808 325198 522850 325434
rect 523086 325198 523128 325434
rect 524740 325198 524782 325434
rect 525018 325198 525060 325434
rect 526672 325198 526714 325434
rect 526950 325198 526992 325434
rect 527876 325198 527918 325434
rect 528154 325198 528196 325434
rect 519144 324258 519186 324494
rect 519422 324258 519464 324494
rect 519910 324258 519952 324494
rect 520188 324258 520230 324494
rect 521842 324258 521884 324494
rect 522120 324258 522162 324494
rect 523774 324258 523816 324494
rect 524052 324258 524094 324494
rect 525706 324258 525748 324494
rect 525984 324258 526026 324494
rect 519144 317494 519464 324258
rect 519144 317258 519186 317494
rect 519422 317258 519464 317494
rect 519144 310494 519464 317258
rect 519144 310258 519186 310494
rect 519422 310258 519464 310494
rect 519144 303494 519464 310258
rect 519144 303258 519186 303494
rect 519422 303258 519464 303494
rect 519144 296494 519464 303258
rect 520876 318434 521196 320008
rect 520876 318198 520918 318434
rect 521154 318198 521196 318434
rect 520876 311434 521196 318198
rect 520876 311198 520918 311434
rect 521154 311198 521196 311434
rect 520876 304434 521196 311198
rect 520876 304198 520918 304434
rect 521154 304198 521196 304434
rect 520876 301752 521196 304198
rect 526144 317494 526464 320008
rect 526144 317258 526186 317494
rect 526422 317258 526464 317494
rect 526144 310494 526464 317258
rect 526144 310258 526186 310494
rect 526422 310258 526464 310494
rect 526144 303494 526464 310258
rect 526144 303258 526186 303494
rect 526422 303258 526464 303494
rect 526144 301752 526464 303258
rect 527876 318434 528196 325198
rect 527876 318198 527918 318434
rect 528154 318198 528196 318434
rect 527876 311434 528196 318198
rect 527876 311198 527918 311434
rect 528154 311198 528196 311434
rect 527876 304434 528196 311198
rect 527876 304198 527918 304434
rect 528154 304198 528196 304434
rect 527876 297434 528196 304198
rect 520876 297198 520918 297434
rect 521154 297198 521196 297434
rect 522808 297198 522850 297434
rect 523086 297198 523128 297434
rect 524740 297198 524782 297434
rect 525018 297198 525060 297434
rect 526672 297198 526714 297434
rect 526950 297198 526992 297434
rect 527876 297198 527918 297434
rect 528154 297198 528196 297434
rect 519144 296258 519186 296494
rect 519422 296258 519464 296494
rect 519910 296258 519952 296494
rect 520188 296258 520230 296494
rect 521842 296258 521884 296494
rect 522120 296258 522162 296494
rect 523774 296258 523816 296494
rect 524052 296258 524094 296494
rect 525706 296258 525748 296494
rect 525984 296258 526026 296494
rect 519144 289494 519464 296258
rect 527876 290434 528196 297198
rect 520876 290198 520918 290434
rect 521154 290198 521196 290434
rect 522808 290198 522850 290434
rect 523086 290198 523128 290434
rect 524740 290198 524782 290434
rect 525018 290198 525060 290434
rect 526672 290198 526714 290434
rect 526950 290198 526992 290434
rect 527876 290198 527918 290434
rect 528154 290198 528196 290434
rect 519144 289258 519186 289494
rect 519422 289258 519464 289494
rect 519910 289258 519952 289494
rect 520188 289258 520230 289494
rect 521842 289258 521884 289494
rect 522120 289258 522162 289494
rect 523774 289258 523816 289494
rect 524052 289258 524094 289494
rect 525706 289258 525748 289494
rect 525984 289258 526026 289494
rect 519144 282494 519464 289258
rect 527876 283434 528196 290198
rect 520876 283198 520918 283434
rect 521154 283198 521196 283434
rect 522808 283198 522850 283434
rect 523086 283198 523128 283434
rect 524740 283198 524782 283434
rect 525018 283198 525060 283434
rect 526672 283198 526714 283434
rect 526950 283198 526992 283434
rect 527876 283198 527918 283434
rect 528154 283198 528196 283434
rect 519144 282258 519186 282494
rect 519422 282258 519464 282494
rect 519910 282258 519952 282494
rect 520188 282258 520230 282494
rect 521842 282258 521884 282494
rect 522120 282258 522162 282494
rect 523774 282258 523816 282494
rect 524052 282258 524094 282494
rect 525706 282258 525748 282494
rect 525984 282258 526026 282494
rect 519144 275494 519464 282258
rect 519144 275258 519186 275494
rect 519422 275258 519464 275494
rect 519144 268494 519464 275258
rect 519144 268258 519186 268494
rect 519422 268258 519464 268494
rect 519144 261494 519464 268258
rect 520876 276434 521196 280008
rect 520876 276198 520918 276434
rect 521154 276198 521196 276434
rect 520876 269434 521196 276198
rect 520876 269198 520918 269434
rect 521154 269198 521196 269434
rect 520876 262434 521196 269198
rect 520876 262198 520918 262434
rect 521154 262198 521196 262434
rect 520876 261752 521196 262198
rect 526144 275494 526464 280008
rect 526144 275258 526186 275494
rect 526422 275258 526464 275494
rect 526144 268494 526464 275258
rect 526144 268258 526186 268494
rect 526422 268258 526464 268494
rect 526144 261752 526464 268258
rect 527876 276434 528196 283198
rect 527876 276198 527918 276434
rect 528154 276198 528196 276434
rect 527876 269434 528196 276198
rect 527876 269198 527918 269434
rect 528154 269198 528196 269434
rect 527876 262434 528196 269198
rect 527876 262198 527918 262434
rect 528154 262198 528196 262434
rect 519144 261258 519186 261494
rect 519422 261258 519464 261494
rect 519144 254494 519464 261258
rect 527876 255434 528196 262198
rect 520876 255198 520918 255434
rect 521154 255198 521196 255434
rect 522808 255198 522850 255434
rect 523086 255198 523128 255434
rect 524740 255198 524782 255434
rect 525018 255198 525060 255434
rect 526672 255198 526714 255434
rect 526950 255198 526992 255434
rect 527876 255198 527918 255434
rect 528154 255198 528196 255434
rect 519144 254258 519186 254494
rect 519422 254258 519464 254494
rect 519910 254258 519952 254494
rect 520188 254258 520230 254494
rect 521842 254258 521884 254494
rect 522120 254258 522162 254494
rect 523774 254258 523816 254494
rect 524052 254258 524094 254494
rect 525706 254258 525748 254494
rect 525984 254258 526026 254494
rect 519144 247494 519464 254258
rect 527876 248434 528196 255198
rect 520876 248198 520918 248434
rect 521154 248198 521196 248434
rect 522808 248198 522850 248434
rect 523086 248198 523128 248434
rect 524740 248198 524782 248434
rect 525018 248198 525060 248434
rect 526672 248198 526714 248434
rect 526950 248198 526992 248434
rect 527876 248198 527918 248434
rect 528154 248198 528196 248434
rect 519144 247258 519186 247494
rect 519422 247258 519464 247494
rect 519910 247258 519952 247494
rect 520188 247258 520230 247494
rect 521842 247258 521884 247494
rect 522120 247258 522162 247494
rect 523774 247258 523816 247494
rect 524052 247258 524094 247494
rect 525706 247258 525748 247494
rect 525984 247258 526026 247494
rect 519144 240494 519464 247258
rect 519144 240258 519186 240494
rect 519422 240258 519464 240494
rect 519144 233494 519464 240258
rect 527876 241434 528196 248198
rect 527876 241198 527918 241434
rect 528154 241198 528196 241434
rect 519144 233258 519186 233494
rect 519422 233258 519464 233494
rect 519144 226494 519464 233258
rect 519144 226258 519186 226494
rect 519422 226258 519464 226494
rect 519144 219494 519464 226258
rect 519144 219258 519186 219494
rect 519422 219258 519464 219494
rect 519144 212494 519464 219258
rect 519144 212258 519186 212494
rect 519422 212258 519464 212494
rect 519144 205494 519464 212258
rect 519144 205258 519186 205494
rect 519422 205258 519464 205494
rect 519144 198494 519464 205258
rect 519144 198258 519186 198494
rect 519422 198258 519464 198494
rect 519144 191494 519464 198258
rect 519144 191258 519186 191494
rect 519422 191258 519464 191494
rect 519144 184494 519464 191258
rect 519144 184258 519186 184494
rect 519422 184258 519464 184494
rect 519144 177494 519464 184258
rect 519144 177258 519186 177494
rect 519422 177258 519464 177494
rect 519144 170494 519464 177258
rect 519144 170258 519186 170494
rect 519422 170258 519464 170494
rect 519144 163494 519464 170258
rect 519144 163258 519186 163494
rect 519422 163258 519464 163494
rect 519144 156494 519464 163258
rect 519144 156258 519186 156494
rect 519422 156258 519464 156494
rect 519144 149494 519464 156258
rect 519144 149258 519186 149494
rect 519422 149258 519464 149494
rect 519144 142494 519464 149258
rect 519144 142258 519186 142494
rect 519422 142258 519464 142494
rect 519144 135494 519464 142258
rect 519144 135258 519186 135494
rect 519422 135258 519464 135494
rect 519144 128494 519464 135258
rect 519144 128258 519186 128494
rect 519422 128258 519464 128494
rect 519144 121494 519464 128258
rect 519144 121258 519186 121494
rect 519422 121258 519464 121494
rect 519144 114494 519464 121258
rect 519144 114258 519186 114494
rect 519422 114258 519464 114494
rect 519144 107494 519464 114258
rect 519144 107258 519186 107494
rect 519422 107258 519464 107494
rect 519144 100494 519464 107258
rect 519144 100258 519186 100494
rect 519422 100258 519464 100494
rect 519144 93494 519464 100258
rect 519144 93258 519186 93494
rect 519422 93258 519464 93494
rect 519144 86494 519464 93258
rect 519144 86258 519186 86494
rect 519422 86258 519464 86494
rect 519144 79494 519464 86258
rect 519144 79258 519186 79494
rect 519422 79258 519464 79494
rect 519144 72494 519464 79258
rect 519144 72258 519186 72494
rect 519422 72258 519464 72494
rect 519144 65494 519464 72258
rect 519144 65258 519186 65494
rect 519422 65258 519464 65494
rect 519144 58494 519464 65258
rect 519144 58258 519186 58494
rect 519422 58258 519464 58494
rect 519144 51494 519464 58258
rect 519144 51258 519186 51494
rect 519422 51258 519464 51494
rect 519144 44494 519464 51258
rect 519144 44258 519186 44494
rect 519422 44258 519464 44494
rect 519144 37494 519464 44258
rect 519144 37258 519186 37494
rect 519422 37258 519464 37494
rect 519144 30494 519464 37258
rect 519144 30258 519186 30494
rect 519422 30258 519464 30494
rect 519144 23494 519464 30258
rect 519144 23258 519186 23494
rect 519422 23258 519464 23494
rect 519144 16494 519464 23258
rect 519144 16258 519186 16494
rect 519422 16258 519464 16494
rect 519144 9494 519464 16258
rect 519144 9258 519186 9494
rect 519422 9258 519464 9494
rect 519144 2494 519464 9258
rect 519144 2258 519186 2494
rect 519422 2258 519464 2494
rect 519144 -746 519464 2258
rect 519144 -982 519186 -746
rect 519422 -982 519464 -746
rect 519144 -1066 519464 -982
rect 519144 -1302 519186 -1066
rect 519422 -1302 519464 -1066
rect 519144 -2294 519464 -1302
rect 520876 234434 521196 240008
rect 520876 234198 520918 234434
rect 521154 234198 521196 234434
rect 520876 227434 521196 234198
rect 520876 227198 520918 227434
rect 521154 227198 521196 227434
rect 520876 220434 521196 227198
rect 520876 220198 520918 220434
rect 521154 220198 521196 220434
rect 520876 213434 521196 220198
rect 520876 213198 520918 213434
rect 521154 213198 521196 213434
rect 520876 206434 521196 213198
rect 520876 206198 520918 206434
rect 521154 206198 521196 206434
rect 520876 199434 521196 206198
rect 520876 199198 520918 199434
rect 521154 199198 521196 199434
rect 520876 192434 521196 199198
rect 520876 192198 520918 192434
rect 521154 192198 521196 192434
rect 520876 185434 521196 192198
rect 520876 185198 520918 185434
rect 521154 185198 521196 185434
rect 520876 178434 521196 185198
rect 520876 178198 520918 178434
rect 521154 178198 521196 178434
rect 520876 171434 521196 178198
rect 520876 171198 520918 171434
rect 521154 171198 521196 171434
rect 520876 164434 521196 171198
rect 520876 164198 520918 164434
rect 521154 164198 521196 164434
rect 520876 157434 521196 164198
rect 520876 157198 520918 157434
rect 521154 157198 521196 157434
rect 520876 150434 521196 157198
rect 520876 150198 520918 150434
rect 521154 150198 521196 150434
rect 520876 143434 521196 150198
rect 520876 143198 520918 143434
rect 521154 143198 521196 143434
rect 520876 136434 521196 143198
rect 520876 136198 520918 136434
rect 521154 136198 521196 136434
rect 520876 129434 521196 136198
rect 520876 129198 520918 129434
rect 521154 129198 521196 129434
rect 520876 122434 521196 129198
rect 520876 122198 520918 122434
rect 521154 122198 521196 122434
rect 520876 115434 521196 122198
rect 520876 115198 520918 115434
rect 521154 115198 521196 115434
rect 520876 108434 521196 115198
rect 520876 108198 520918 108434
rect 521154 108198 521196 108434
rect 520876 101434 521196 108198
rect 520876 101198 520918 101434
rect 521154 101198 521196 101434
rect 520876 94434 521196 101198
rect 520876 94198 520918 94434
rect 521154 94198 521196 94434
rect 520876 87434 521196 94198
rect 520876 87198 520918 87434
rect 521154 87198 521196 87434
rect 520876 80434 521196 87198
rect 520876 80198 520918 80434
rect 521154 80198 521196 80434
rect 520876 73434 521196 80198
rect 520876 73198 520918 73434
rect 521154 73198 521196 73434
rect 520876 66434 521196 73198
rect 520876 66198 520918 66434
rect 521154 66198 521196 66434
rect 520876 59434 521196 66198
rect 520876 59198 520918 59434
rect 521154 59198 521196 59434
rect 520876 52434 521196 59198
rect 520876 52198 520918 52434
rect 521154 52198 521196 52434
rect 520876 45434 521196 52198
rect 520876 45198 520918 45434
rect 521154 45198 521196 45434
rect 520876 38434 521196 45198
rect 520876 38198 520918 38434
rect 521154 38198 521196 38434
rect 520876 31434 521196 38198
rect 520876 31198 520918 31434
rect 521154 31198 521196 31434
rect 520876 24434 521196 31198
rect 520876 24198 520918 24434
rect 521154 24198 521196 24434
rect 520876 17434 521196 24198
rect 520876 17198 520918 17434
rect 521154 17198 521196 17434
rect 520876 10434 521196 17198
rect 520876 10198 520918 10434
rect 521154 10198 521196 10434
rect 520876 3434 521196 10198
rect 520876 3198 520918 3434
rect 521154 3198 521196 3434
rect 520876 -1706 521196 3198
rect 520876 -1942 520918 -1706
rect 521154 -1942 521196 -1706
rect 520876 -2026 521196 -1942
rect 520876 -2262 520918 -2026
rect 521154 -2262 521196 -2026
rect 520876 -2294 521196 -2262
rect 526144 233494 526464 240008
rect 526144 233258 526186 233494
rect 526422 233258 526464 233494
rect 526144 226494 526464 233258
rect 526144 226258 526186 226494
rect 526422 226258 526464 226494
rect 526144 219494 526464 226258
rect 526144 219258 526186 219494
rect 526422 219258 526464 219494
rect 526144 212494 526464 219258
rect 526144 212258 526186 212494
rect 526422 212258 526464 212494
rect 526144 205494 526464 212258
rect 526144 205258 526186 205494
rect 526422 205258 526464 205494
rect 526144 198494 526464 205258
rect 526144 198258 526186 198494
rect 526422 198258 526464 198494
rect 526144 191494 526464 198258
rect 526144 191258 526186 191494
rect 526422 191258 526464 191494
rect 526144 184494 526464 191258
rect 526144 184258 526186 184494
rect 526422 184258 526464 184494
rect 526144 177494 526464 184258
rect 526144 177258 526186 177494
rect 526422 177258 526464 177494
rect 526144 170494 526464 177258
rect 526144 170258 526186 170494
rect 526422 170258 526464 170494
rect 526144 163494 526464 170258
rect 526144 163258 526186 163494
rect 526422 163258 526464 163494
rect 526144 156494 526464 163258
rect 526144 156258 526186 156494
rect 526422 156258 526464 156494
rect 526144 149494 526464 156258
rect 526144 149258 526186 149494
rect 526422 149258 526464 149494
rect 526144 142494 526464 149258
rect 526144 142258 526186 142494
rect 526422 142258 526464 142494
rect 526144 135494 526464 142258
rect 526144 135258 526186 135494
rect 526422 135258 526464 135494
rect 526144 128494 526464 135258
rect 526144 128258 526186 128494
rect 526422 128258 526464 128494
rect 526144 121494 526464 128258
rect 526144 121258 526186 121494
rect 526422 121258 526464 121494
rect 526144 114494 526464 121258
rect 526144 114258 526186 114494
rect 526422 114258 526464 114494
rect 526144 107494 526464 114258
rect 526144 107258 526186 107494
rect 526422 107258 526464 107494
rect 526144 100494 526464 107258
rect 526144 100258 526186 100494
rect 526422 100258 526464 100494
rect 526144 93494 526464 100258
rect 526144 93258 526186 93494
rect 526422 93258 526464 93494
rect 526144 86494 526464 93258
rect 526144 86258 526186 86494
rect 526422 86258 526464 86494
rect 526144 79494 526464 86258
rect 526144 79258 526186 79494
rect 526422 79258 526464 79494
rect 526144 72494 526464 79258
rect 526144 72258 526186 72494
rect 526422 72258 526464 72494
rect 526144 65494 526464 72258
rect 526144 65258 526186 65494
rect 526422 65258 526464 65494
rect 526144 58494 526464 65258
rect 526144 58258 526186 58494
rect 526422 58258 526464 58494
rect 526144 51494 526464 58258
rect 526144 51258 526186 51494
rect 526422 51258 526464 51494
rect 526144 44494 526464 51258
rect 526144 44258 526186 44494
rect 526422 44258 526464 44494
rect 526144 37494 526464 44258
rect 526144 37258 526186 37494
rect 526422 37258 526464 37494
rect 526144 30494 526464 37258
rect 526144 30258 526186 30494
rect 526422 30258 526464 30494
rect 526144 23494 526464 30258
rect 526144 23258 526186 23494
rect 526422 23258 526464 23494
rect 526144 16494 526464 23258
rect 526144 16258 526186 16494
rect 526422 16258 526464 16494
rect 526144 9494 526464 16258
rect 526144 9258 526186 9494
rect 526422 9258 526464 9494
rect 526144 2494 526464 9258
rect 526144 2258 526186 2494
rect 526422 2258 526464 2494
rect 526144 -746 526464 2258
rect 526144 -982 526186 -746
rect 526422 -982 526464 -746
rect 526144 -1066 526464 -982
rect 526144 -1302 526186 -1066
rect 526422 -1302 526464 -1066
rect 526144 -2294 526464 -1302
rect 527876 234434 528196 241198
rect 527876 234198 527918 234434
rect 528154 234198 528196 234434
rect 527876 227434 528196 234198
rect 527876 227198 527918 227434
rect 528154 227198 528196 227434
rect 527876 220434 528196 227198
rect 527876 220198 527918 220434
rect 528154 220198 528196 220434
rect 527876 213434 528196 220198
rect 527876 213198 527918 213434
rect 528154 213198 528196 213434
rect 527876 206434 528196 213198
rect 527876 206198 527918 206434
rect 528154 206198 528196 206434
rect 527876 199434 528196 206198
rect 527876 199198 527918 199434
rect 528154 199198 528196 199434
rect 527876 192434 528196 199198
rect 527876 192198 527918 192434
rect 528154 192198 528196 192434
rect 527876 185434 528196 192198
rect 527876 185198 527918 185434
rect 528154 185198 528196 185434
rect 527876 178434 528196 185198
rect 527876 178198 527918 178434
rect 528154 178198 528196 178434
rect 527876 171434 528196 178198
rect 527876 171198 527918 171434
rect 528154 171198 528196 171434
rect 527876 164434 528196 171198
rect 527876 164198 527918 164434
rect 528154 164198 528196 164434
rect 527876 157434 528196 164198
rect 527876 157198 527918 157434
rect 528154 157198 528196 157434
rect 527876 150434 528196 157198
rect 527876 150198 527918 150434
rect 528154 150198 528196 150434
rect 527876 143434 528196 150198
rect 527876 143198 527918 143434
rect 528154 143198 528196 143434
rect 527876 136434 528196 143198
rect 527876 136198 527918 136434
rect 528154 136198 528196 136434
rect 527876 129434 528196 136198
rect 527876 129198 527918 129434
rect 528154 129198 528196 129434
rect 527876 122434 528196 129198
rect 527876 122198 527918 122434
rect 528154 122198 528196 122434
rect 527876 115434 528196 122198
rect 527876 115198 527918 115434
rect 528154 115198 528196 115434
rect 527876 108434 528196 115198
rect 527876 108198 527918 108434
rect 528154 108198 528196 108434
rect 527876 101434 528196 108198
rect 527876 101198 527918 101434
rect 528154 101198 528196 101434
rect 527876 94434 528196 101198
rect 527876 94198 527918 94434
rect 528154 94198 528196 94434
rect 527876 87434 528196 94198
rect 527876 87198 527918 87434
rect 528154 87198 528196 87434
rect 527876 80434 528196 87198
rect 527876 80198 527918 80434
rect 528154 80198 528196 80434
rect 527876 73434 528196 80198
rect 527876 73198 527918 73434
rect 528154 73198 528196 73434
rect 527876 66434 528196 73198
rect 527876 66198 527918 66434
rect 528154 66198 528196 66434
rect 527876 59434 528196 66198
rect 527876 59198 527918 59434
rect 528154 59198 528196 59434
rect 527876 52434 528196 59198
rect 527876 52198 527918 52434
rect 528154 52198 528196 52434
rect 527876 45434 528196 52198
rect 527876 45198 527918 45434
rect 528154 45198 528196 45434
rect 527876 38434 528196 45198
rect 527876 38198 527918 38434
rect 528154 38198 528196 38434
rect 527876 31434 528196 38198
rect 527876 31198 527918 31434
rect 528154 31198 528196 31434
rect 527876 24434 528196 31198
rect 527876 24198 527918 24434
rect 528154 24198 528196 24434
rect 527876 17434 528196 24198
rect 527876 17198 527918 17434
rect 528154 17198 528196 17434
rect 527876 10434 528196 17198
rect 527876 10198 527918 10434
rect 528154 10198 528196 10434
rect 527876 3434 528196 10198
rect 527876 3198 527918 3434
rect 528154 3198 528196 3434
rect 527876 -1706 528196 3198
rect 527876 -1942 527918 -1706
rect 528154 -1942 528196 -1706
rect 527876 -2026 528196 -1942
rect 527876 -2262 527918 -2026
rect 528154 -2262 528196 -2026
rect 527876 -2294 528196 -2262
rect 533144 705238 533464 706230
rect 533144 705002 533186 705238
rect 533422 705002 533464 705238
rect 533144 704918 533464 705002
rect 533144 704682 533186 704918
rect 533422 704682 533464 704918
rect 533144 695494 533464 704682
rect 533144 695258 533186 695494
rect 533422 695258 533464 695494
rect 533144 688494 533464 695258
rect 533144 688258 533186 688494
rect 533422 688258 533464 688494
rect 533144 681494 533464 688258
rect 533144 681258 533186 681494
rect 533422 681258 533464 681494
rect 533144 674494 533464 681258
rect 533144 674258 533186 674494
rect 533422 674258 533464 674494
rect 533144 667494 533464 674258
rect 533144 667258 533186 667494
rect 533422 667258 533464 667494
rect 533144 660494 533464 667258
rect 533144 660258 533186 660494
rect 533422 660258 533464 660494
rect 533144 653494 533464 660258
rect 533144 653258 533186 653494
rect 533422 653258 533464 653494
rect 533144 646494 533464 653258
rect 533144 646258 533186 646494
rect 533422 646258 533464 646494
rect 533144 639494 533464 646258
rect 533144 639258 533186 639494
rect 533422 639258 533464 639494
rect 533144 632494 533464 639258
rect 533144 632258 533186 632494
rect 533422 632258 533464 632494
rect 533144 625494 533464 632258
rect 533144 625258 533186 625494
rect 533422 625258 533464 625494
rect 533144 618494 533464 625258
rect 533144 618258 533186 618494
rect 533422 618258 533464 618494
rect 533144 611494 533464 618258
rect 533144 611258 533186 611494
rect 533422 611258 533464 611494
rect 533144 604494 533464 611258
rect 533144 604258 533186 604494
rect 533422 604258 533464 604494
rect 533144 597494 533464 604258
rect 533144 597258 533186 597494
rect 533422 597258 533464 597494
rect 533144 590494 533464 597258
rect 533144 590258 533186 590494
rect 533422 590258 533464 590494
rect 533144 583494 533464 590258
rect 533144 583258 533186 583494
rect 533422 583258 533464 583494
rect 533144 576494 533464 583258
rect 533144 576258 533186 576494
rect 533422 576258 533464 576494
rect 533144 569494 533464 576258
rect 533144 569258 533186 569494
rect 533422 569258 533464 569494
rect 533144 562494 533464 569258
rect 533144 562258 533186 562494
rect 533422 562258 533464 562494
rect 533144 555494 533464 562258
rect 533144 555258 533186 555494
rect 533422 555258 533464 555494
rect 533144 548494 533464 555258
rect 533144 548258 533186 548494
rect 533422 548258 533464 548494
rect 533144 541494 533464 548258
rect 533144 541258 533186 541494
rect 533422 541258 533464 541494
rect 533144 534494 533464 541258
rect 533144 534258 533186 534494
rect 533422 534258 533464 534494
rect 533144 527494 533464 534258
rect 533144 527258 533186 527494
rect 533422 527258 533464 527494
rect 533144 520494 533464 527258
rect 533144 520258 533186 520494
rect 533422 520258 533464 520494
rect 533144 513494 533464 520258
rect 533144 513258 533186 513494
rect 533422 513258 533464 513494
rect 533144 506494 533464 513258
rect 533144 506258 533186 506494
rect 533422 506258 533464 506494
rect 533144 499494 533464 506258
rect 533144 499258 533186 499494
rect 533422 499258 533464 499494
rect 533144 492494 533464 499258
rect 533144 492258 533186 492494
rect 533422 492258 533464 492494
rect 533144 485494 533464 492258
rect 533144 485258 533186 485494
rect 533422 485258 533464 485494
rect 533144 478494 533464 485258
rect 533144 478258 533186 478494
rect 533422 478258 533464 478494
rect 533144 471494 533464 478258
rect 533144 471258 533186 471494
rect 533422 471258 533464 471494
rect 533144 464494 533464 471258
rect 533144 464258 533186 464494
rect 533422 464258 533464 464494
rect 533144 457494 533464 464258
rect 533144 457258 533186 457494
rect 533422 457258 533464 457494
rect 533144 450494 533464 457258
rect 533144 450258 533186 450494
rect 533422 450258 533464 450494
rect 533144 443494 533464 450258
rect 533144 443258 533186 443494
rect 533422 443258 533464 443494
rect 533144 436494 533464 443258
rect 533144 436258 533186 436494
rect 533422 436258 533464 436494
rect 533144 429494 533464 436258
rect 533144 429258 533186 429494
rect 533422 429258 533464 429494
rect 533144 422494 533464 429258
rect 533144 422258 533186 422494
rect 533422 422258 533464 422494
rect 533144 415494 533464 422258
rect 533144 415258 533186 415494
rect 533422 415258 533464 415494
rect 533144 408494 533464 415258
rect 533144 408258 533186 408494
rect 533422 408258 533464 408494
rect 533144 401494 533464 408258
rect 533144 401258 533186 401494
rect 533422 401258 533464 401494
rect 533144 394494 533464 401258
rect 533144 394258 533186 394494
rect 533422 394258 533464 394494
rect 533144 387494 533464 394258
rect 533144 387258 533186 387494
rect 533422 387258 533464 387494
rect 533144 380494 533464 387258
rect 533144 380258 533186 380494
rect 533422 380258 533464 380494
rect 533144 373494 533464 380258
rect 533144 373258 533186 373494
rect 533422 373258 533464 373494
rect 533144 366494 533464 373258
rect 533144 366258 533186 366494
rect 533422 366258 533464 366494
rect 533144 359494 533464 366258
rect 533144 359258 533186 359494
rect 533422 359258 533464 359494
rect 533144 352494 533464 359258
rect 533144 352258 533186 352494
rect 533422 352258 533464 352494
rect 533144 345494 533464 352258
rect 533144 345258 533186 345494
rect 533422 345258 533464 345494
rect 533144 338494 533464 345258
rect 533144 338258 533186 338494
rect 533422 338258 533464 338494
rect 533144 331494 533464 338258
rect 533144 331258 533186 331494
rect 533422 331258 533464 331494
rect 533144 324494 533464 331258
rect 533144 324258 533186 324494
rect 533422 324258 533464 324494
rect 533144 317494 533464 324258
rect 533144 317258 533186 317494
rect 533422 317258 533464 317494
rect 533144 310494 533464 317258
rect 533144 310258 533186 310494
rect 533422 310258 533464 310494
rect 533144 303494 533464 310258
rect 533144 303258 533186 303494
rect 533422 303258 533464 303494
rect 533144 296494 533464 303258
rect 533144 296258 533186 296494
rect 533422 296258 533464 296494
rect 533144 289494 533464 296258
rect 533144 289258 533186 289494
rect 533422 289258 533464 289494
rect 533144 282494 533464 289258
rect 533144 282258 533186 282494
rect 533422 282258 533464 282494
rect 533144 275494 533464 282258
rect 533144 275258 533186 275494
rect 533422 275258 533464 275494
rect 533144 268494 533464 275258
rect 533144 268258 533186 268494
rect 533422 268258 533464 268494
rect 533144 261494 533464 268258
rect 533144 261258 533186 261494
rect 533422 261258 533464 261494
rect 533144 254494 533464 261258
rect 533144 254258 533186 254494
rect 533422 254258 533464 254494
rect 533144 247494 533464 254258
rect 533144 247258 533186 247494
rect 533422 247258 533464 247494
rect 533144 240494 533464 247258
rect 533144 240258 533186 240494
rect 533422 240258 533464 240494
rect 533144 233494 533464 240258
rect 533144 233258 533186 233494
rect 533422 233258 533464 233494
rect 533144 226494 533464 233258
rect 533144 226258 533186 226494
rect 533422 226258 533464 226494
rect 533144 219494 533464 226258
rect 533144 219258 533186 219494
rect 533422 219258 533464 219494
rect 533144 212494 533464 219258
rect 533144 212258 533186 212494
rect 533422 212258 533464 212494
rect 533144 205494 533464 212258
rect 533144 205258 533186 205494
rect 533422 205258 533464 205494
rect 533144 198494 533464 205258
rect 533144 198258 533186 198494
rect 533422 198258 533464 198494
rect 533144 191494 533464 198258
rect 533144 191258 533186 191494
rect 533422 191258 533464 191494
rect 533144 184494 533464 191258
rect 533144 184258 533186 184494
rect 533422 184258 533464 184494
rect 533144 177494 533464 184258
rect 533144 177258 533186 177494
rect 533422 177258 533464 177494
rect 533144 170494 533464 177258
rect 533144 170258 533186 170494
rect 533422 170258 533464 170494
rect 533144 163494 533464 170258
rect 533144 163258 533186 163494
rect 533422 163258 533464 163494
rect 533144 156494 533464 163258
rect 533144 156258 533186 156494
rect 533422 156258 533464 156494
rect 533144 149494 533464 156258
rect 533144 149258 533186 149494
rect 533422 149258 533464 149494
rect 533144 142494 533464 149258
rect 533144 142258 533186 142494
rect 533422 142258 533464 142494
rect 533144 135494 533464 142258
rect 533144 135258 533186 135494
rect 533422 135258 533464 135494
rect 533144 128494 533464 135258
rect 533144 128258 533186 128494
rect 533422 128258 533464 128494
rect 533144 121494 533464 128258
rect 533144 121258 533186 121494
rect 533422 121258 533464 121494
rect 533144 114494 533464 121258
rect 533144 114258 533186 114494
rect 533422 114258 533464 114494
rect 533144 107494 533464 114258
rect 533144 107258 533186 107494
rect 533422 107258 533464 107494
rect 533144 100494 533464 107258
rect 533144 100258 533186 100494
rect 533422 100258 533464 100494
rect 533144 93494 533464 100258
rect 533144 93258 533186 93494
rect 533422 93258 533464 93494
rect 533144 86494 533464 93258
rect 533144 86258 533186 86494
rect 533422 86258 533464 86494
rect 533144 79494 533464 86258
rect 533144 79258 533186 79494
rect 533422 79258 533464 79494
rect 533144 72494 533464 79258
rect 533144 72258 533186 72494
rect 533422 72258 533464 72494
rect 533144 65494 533464 72258
rect 533144 65258 533186 65494
rect 533422 65258 533464 65494
rect 533144 58494 533464 65258
rect 533144 58258 533186 58494
rect 533422 58258 533464 58494
rect 533144 51494 533464 58258
rect 533144 51258 533186 51494
rect 533422 51258 533464 51494
rect 533144 44494 533464 51258
rect 533144 44258 533186 44494
rect 533422 44258 533464 44494
rect 533144 37494 533464 44258
rect 533144 37258 533186 37494
rect 533422 37258 533464 37494
rect 533144 30494 533464 37258
rect 533144 30258 533186 30494
rect 533422 30258 533464 30494
rect 533144 23494 533464 30258
rect 533144 23258 533186 23494
rect 533422 23258 533464 23494
rect 533144 16494 533464 23258
rect 533144 16258 533186 16494
rect 533422 16258 533464 16494
rect 533144 9494 533464 16258
rect 533144 9258 533186 9494
rect 533422 9258 533464 9494
rect 533144 2494 533464 9258
rect 533144 2258 533186 2494
rect 533422 2258 533464 2494
rect 533144 -746 533464 2258
rect 533144 -982 533186 -746
rect 533422 -982 533464 -746
rect 533144 -1066 533464 -982
rect 533144 -1302 533186 -1066
rect 533422 -1302 533464 -1066
rect 533144 -2294 533464 -1302
rect 534876 706198 535196 706230
rect 534876 705962 534918 706198
rect 535154 705962 535196 706198
rect 534876 705878 535196 705962
rect 534876 705642 534918 705878
rect 535154 705642 535196 705878
rect 534876 696434 535196 705642
rect 534876 696198 534918 696434
rect 535154 696198 535196 696434
rect 534876 689434 535196 696198
rect 534876 689198 534918 689434
rect 535154 689198 535196 689434
rect 534876 682434 535196 689198
rect 534876 682198 534918 682434
rect 535154 682198 535196 682434
rect 534876 675434 535196 682198
rect 534876 675198 534918 675434
rect 535154 675198 535196 675434
rect 534876 668434 535196 675198
rect 534876 668198 534918 668434
rect 535154 668198 535196 668434
rect 534876 661434 535196 668198
rect 534876 661198 534918 661434
rect 535154 661198 535196 661434
rect 534876 654434 535196 661198
rect 534876 654198 534918 654434
rect 535154 654198 535196 654434
rect 534876 647434 535196 654198
rect 534876 647198 534918 647434
rect 535154 647198 535196 647434
rect 534876 640434 535196 647198
rect 534876 640198 534918 640434
rect 535154 640198 535196 640434
rect 534876 633434 535196 640198
rect 534876 633198 534918 633434
rect 535154 633198 535196 633434
rect 534876 626434 535196 633198
rect 534876 626198 534918 626434
rect 535154 626198 535196 626434
rect 534876 619434 535196 626198
rect 534876 619198 534918 619434
rect 535154 619198 535196 619434
rect 534876 612434 535196 619198
rect 534876 612198 534918 612434
rect 535154 612198 535196 612434
rect 534876 605434 535196 612198
rect 534876 605198 534918 605434
rect 535154 605198 535196 605434
rect 534876 598434 535196 605198
rect 534876 598198 534918 598434
rect 535154 598198 535196 598434
rect 534876 591434 535196 598198
rect 534876 591198 534918 591434
rect 535154 591198 535196 591434
rect 534876 584434 535196 591198
rect 534876 584198 534918 584434
rect 535154 584198 535196 584434
rect 534876 577434 535196 584198
rect 534876 577198 534918 577434
rect 535154 577198 535196 577434
rect 534876 570434 535196 577198
rect 534876 570198 534918 570434
rect 535154 570198 535196 570434
rect 534876 563434 535196 570198
rect 534876 563198 534918 563434
rect 535154 563198 535196 563434
rect 534876 556434 535196 563198
rect 534876 556198 534918 556434
rect 535154 556198 535196 556434
rect 534876 549434 535196 556198
rect 534876 549198 534918 549434
rect 535154 549198 535196 549434
rect 534876 542434 535196 549198
rect 534876 542198 534918 542434
rect 535154 542198 535196 542434
rect 534876 535434 535196 542198
rect 534876 535198 534918 535434
rect 535154 535198 535196 535434
rect 534876 528434 535196 535198
rect 534876 528198 534918 528434
rect 535154 528198 535196 528434
rect 534876 521434 535196 528198
rect 534876 521198 534918 521434
rect 535154 521198 535196 521434
rect 534876 514434 535196 521198
rect 534876 514198 534918 514434
rect 535154 514198 535196 514434
rect 534876 507434 535196 514198
rect 534876 507198 534918 507434
rect 535154 507198 535196 507434
rect 534876 500434 535196 507198
rect 534876 500198 534918 500434
rect 535154 500198 535196 500434
rect 534876 493434 535196 500198
rect 534876 493198 534918 493434
rect 535154 493198 535196 493434
rect 534876 486434 535196 493198
rect 534876 486198 534918 486434
rect 535154 486198 535196 486434
rect 534876 479434 535196 486198
rect 534876 479198 534918 479434
rect 535154 479198 535196 479434
rect 534876 472434 535196 479198
rect 534876 472198 534918 472434
rect 535154 472198 535196 472434
rect 534876 465434 535196 472198
rect 534876 465198 534918 465434
rect 535154 465198 535196 465434
rect 534876 458434 535196 465198
rect 534876 458198 534918 458434
rect 535154 458198 535196 458434
rect 534876 451434 535196 458198
rect 534876 451198 534918 451434
rect 535154 451198 535196 451434
rect 534876 444434 535196 451198
rect 534876 444198 534918 444434
rect 535154 444198 535196 444434
rect 534876 437434 535196 444198
rect 534876 437198 534918 437434
rect 535154 437198 535196 437434
rect 534876 430434 535196 437198
rect 534876 430198 534918 430434
rect 535154 430198 535196 430434
rect 534876 423434 535196 430198
rect 534876 423198 534918 423434
rect 535154 423198 535196 423434
rect 534876 416434 535196 423198
rect 534876 416198 534918 416434
rect 535154 416198 535196 416434
rect 534876 409434 535196 416198
rect 534876 409198 534918 409434
rect 535154 409198 535196 409434
rect 534876 402434 535196 409198
rect 534876 402198 534918 402434
rect 535154 402198 535196 402434
rect 534876 395434 535196 402198
rect 534876 395198 534918 395434
rect 535154 395198 535196 395434
rect 534876 388434 535196 395198
rect 534876 388198 534918 388434
rect 535154 388198 535196 388434
rect 534876 381434 535196 388198
rect 534876 381198 534918 381434
rect 535154 381198 535196 381434
rect 534876 374434 535196 381198
rect 534876 374198 534918 374434
rect 535154 374198 535196 374434
rect 534876 367434 535196 374198
rect 534876 367198 534918 367434
rect 535154 367198 535196 367434
rect 534876 360434 535196 367198
rect 534876 360198 534918 360434
rect 535154 360198 535196 360434
rect 534876 353434 535196 360198
rect 534876 353198 534918 353434
rect 535154 353198 535196 353434
rect 534876 346434 535196 353198
rect 534876 346198 534918 346434
rect 535154 346198 535196 346434
rect 534876 339434 535196 346198
rect 534876 339198 534918 339434
rect 535154 339198 535196 339434
rect 534876 332434 535196 339198
rect 534876 332198 534918 332434
rect 535154 332198 535196 332434
rect 534876 325434 535196 332198
rect 534876 325198 534918 325434
rect 535154 325198 535196 325434
rect 534876 318434 535196 325198
rect 534876 318198 534918 318434
rect 535154 318198 535196 318434
rect 534876 311434 535196 318198
rect 534876 311198 534918 311434
rect 535154 311198 535196 311434
rect 534876 304434 535196 311198
rect 534876 304198 534918 304434
rect 535154 304198 535196 304434
rect 534876 297434 535196 304198
rect 534876 297198 534918 297434
rect 535154 297198 535196 297434
rect 534876 290434 535196 297198
rect 534876 290198 534918 290434
rect 535154 290198 535196 290434
rect 534876 283434 535196 290198
rect 534876 283198 534918 283434
rect 535154 283198 535196 283434
rect 534876 276434 535196 283198
rect 534876 276198 534918 276434
rect 535154 276198 535196 276434
rect 534876 269434 535196 276198
rect 534876 269198 534918 269434
rect 535154 269198 535196 269434
rect 534876 262434 535196 269198
rect 534876 262198 534918 262434
rect 535154 262198 535196 262434
rect 534876 255434 535196 262198
rect 534876 255198 534918 255434
rect 535154 255198 535196 255434
rect 534876 248434 535196 255198
rect 534876 248198 534918 248434
rect 535154 248198 535196 248434
rect 534876 241434 535196 248198
rect 534876 241198 534918 241434
rect 535154 241198 535196 241434
rect 534876 234434 535196 241198
rect 534876 234198 534918 234434
rect 535154 234198 535196 234434
rect 534876 227434 535196 234198
rect 534876 227198 534918 227434
rect 535154 227198 535196 227434
rect 534876 220434 535196 227198
rect 534876 220198 534918 220434
rect 535154 220198 535196 220434
rect 534876 213434 535196 220198
rect 534876 213198 534918 213434
rect 535154 213198 535196 213434
rect 534876 206434 535196 213198
rect 534876 206198 534918 206434
rect 535154 206198 535196 206434
rect 534876 199434 535196 206198
rect 534876 199198 534918 199434
rect 535154 199198 535196 199434
rect 534876 192434 535196 199198
rect 534876 192198 534918 192434
rect 535154 192198 535196 192434
rect 534876 185434 535196 192198
rect 534876 185198 534918 185434
rect 535154 185198 535196 185434
rect 534876 178434 535196 185198
rect 534876 178198 534918 178434
rect 535154 178198 535196 178434
rect 534876 171434 535196 178198
rect 534876 171198 534918 171434
rect 535154 171198 535196 171434
rect 534876 164434 535196 171198
rect 534876 164198 534918 164434
rect 535154 164198 535196 164434
rect 534876 157434 535196 164198
rect 534876 157198 534918 157434
rect 535154 157198 535196 157434
rect 534876 150434 535196 157198
rect 534876 150198 534918 150434
rect 535154 150198 535196 150434
rect 534876 143434 535196 150198
rect 534876 143198 534918 143434
rect 535154 143198 535196 143434
rect 534876 136434 535196 143198
rect 534876 136198 534918 136434
rect 535154 136198 535196 136434
rect 534876 129434 535196 136198
rect 534876 129198 534918 129434
rect 535154 129198 535196 129434
rect 534876 122434 535196 129198
rect 534876 122198 534918 122434
rect 535154 122198 535196 122434
rect 534876 115434 535196 122198
rect 534876 115198 534918 115434
rect 535154 115198 535196 115434
rect 534876 108434 535196 115198
rect 534876 108198 534918 108434
rect 535154 108198 535196 108434
rect 534876 101434 535196 108198
rect 534876 101198 534918 101434
rect 535154 101198 535196 101434
rect 534876 94434 535196 101198
rect 534876 94198 534918 94434
rect 535154 94198 535196 94434
rect 534876 87434 535196 94198
rect 534876 87198 534918 87434
rect 535154 87198 535196 87434
rect 534876 80434 535196 87198
rect 534876 80198 534918 80434
rect 535154 80198 535196 80434
rect 534876 73434 535196 80198
rect 534876 73198 534918 73434
rect 535154 73198 535196 73434
rect 534876 66434 535196 73198
rect 534876 66198 534918 66434
rect 535154 66198 535196 66434
rect 534876 59434 535196 66198
rect 534876 59198 534918 59434
rect 535154 59198 535196 59434
rect 534876 52434 535196 59198
rect 534876 52198 534918 52434
rect 535154 52198 535196 52434
rect 534876 45434 535196 52198
rect 534876 45198 534918 45434
rect 535154 45198 535196 45434
rect 534876 38434 535196 45198
rect 534876 38198 534918 38434
rect 535154 38198 535196 38434
rect 534876 31434 535196 38198
rect 534876 31198 534918 31434
rect 535154 31198 535196 31434
rect 534876 24434 535196 31198
rect 534876 24198 534918 24434
rect 535154 24198 535196 24434
rect 534876 17434 535196 24198
rect 534876 17198 534918 17434
rect 535154 17198 535196 17434
rect 534876 10434 535196 17198
rect 534876 10198 534918 10434
rect 535154 10198 535196 10434
rect 534876 3434 535196 10198
rect 534876 3198 534918 3434
rect 535154 3198 535196 3434
rect 534876 -1706 535196 3198
rect 534876 -1942 534918 -1706
rect 535154 -1942 535196 -1706
rect 534876 -2026 535196 -1942
rect 534876 -2262 534918 -2026
rect 535154 -2262 535196 -2026
rect 534876 -2294 535196 -2262
rect 540144 705238 540464 706230
rect 540144 705002 540186 705238
rect 540422 705002 540464 705238
rect 540144 704918 540464 705002
rect 540144 704682 540186 704918
rect 540422 704682 540464 704918
rect 540144 695494 540464 704682
rect 540144 695258 540186 695494
rect 540422 695258 540464 695494
rect 540144 688494 540464 695258
rect 540144 688258 540186 688494
rect 540422 688258 540464 688494
rect 540144 681494 540464 688258
rect 540144 681258 540186 681494
rect 540422 681258 540464 681494
rect 540144 674494 540464 681258
rect 540144 674258 540186 674494
rect 540422 674258 540464 674494
rect 540144 667494 540464 674258
rect 540144 667258 540186 667494
rect 540422 667258 540464 667494
rect 540144 660494 540464 667258
rect 540144 660258 540186 660494
rect 540422 660258 540464 660494
rect 540144 653494 540464 660258
rect 540144 653258 540186 653494
rect 540422 653258 540464 653494
rect 540144 646494 540464 653258
rect 540144 646258 540186 646494
rect 540422 646258 540464 646494
rect 540144 639494 540464 646258
rect 540144 639258 540186 639494
rect 540422 639258 540464 639494
rect 540144 632494 540464 639258
rect 540144 632258 540186 632494
rect 540422 632258 540464 632494
rect 540144 625494 540464 632258
rect 540144 625258 540186 625494
rect 540422 625258 540464 625494
rect 540144 618494 540464 625258
rect 540144 618258 540186 618494
rect 540422 618258 540464 618494
rect 540144 611494 540464 618258
rect 540144 611258 540186 611494
rect 540422 611258 540464 611494
rect 540144 604494 540464 611258
rect 540144 604258 540186 604494
rect 540422 604258 540464 604494
rect 540144 597494 540464 604258
rect 540144 597258 540186 597494
rect 540422 597258 540464 597494
rect 540144 590494 540464 597258
rect 540144 590258 540186 590494
rect 540422 590258 540464 590494
rect 540144 583494 540464 590258
rect 540144 583258 540186 583494
rect 540422 583258 540464 583494
rect 540144 576494 540464 583258
rect 540144 576258 540186 576494
rect 540422 576258 540464 576494
rect 540144 569494 540464 576258
rect 540144 569258 540186 569494
rect 540422 569258 540464 569494
rect 540144 562494 540464 569258
rect 540144 562258 540186 562494
rect 540422 562258 540464 562494
rect 540144 555494 540464 562258
rect 540144 555258 540186 555494
rect 540422 555258 540464 555494
rect 540144 548494 540464 555258
rect 540144 548258 540186 548494
rect 540422 548258 540464 548494
rect 540144 541494 540464 548258
rect 540144 541258 540186 541494
rect 540422 541258 540464 541494
rect 540144 534494 540464 541258
rect 540144 534258 540186 534494
rect 540422 534258 540464 534494
rect 540144 527494 540464 534258
rect 540144 527258 540186 527494
rect 540422 527258 540464 527494
rect 540144 520494 540464 527258
rect 540144 520258 540186 520494
rect 540422 520258 540464 520494
rect 540144 513494 540464 520258
rect 540144 513258 540186 513494
rect 540422 513258 540464 513494
rect 540144 506494 540464 513258
rect 540144 506258 540186 506494
rect 540422 506258 540464 506494
rect 540144 499494 540464 506258
rect 540144 499258 540186 499494
rect 540422 499258 540464 499494
rect 540144 492494 540464 499258
rect 540144 492258 540186 492494
rect 540422 492258 540464 492494
rect 540144 485494 540464 492258
rect 540144 485258 540186 485494
rect 540422 485258 540464 485494
rect 540144 478494 540464 485258
rect 540144 478258 540186 478494
rect 540422 478258 540464 478494
rect 540144 471494 540464 478258
rect 540144 471258 540186 471494
rect 540422 471258 540464 471494
rect 540144 464494 540464 471258
rect 540144 464258 540186 464494
rect 540422 464258 540464 464494
rect 540144 457494 540464 464258
rect 540144 457258 540186 457494
rect 540422 457258 540464 457494
rect 540144 450494 540464 457258
rect 540144 450258 540186 450494
rect 540422 450258 540464 450494
rect 540144 443494 540464 450258
rect 540144 443258 540186 443494
rect 540422 443258 540464 443494
rect 540144 436494 540464 443258
rect 540144 436258 540186 436494
rect 540422 436258 540464 436494
rect 540144 429494 540464 436258
rect 540144 429258 540186 429494
rect 540422 429258 540464 429494
rect 540144 422494 540464 429258
rect 540144 422258 540186 422494
rect 540422 422258 540464 422494
rect 540144 415494 540464 422258
rect 540144 415258 540186 415494
rect 540422 415258 540464 415494
rect 540144 408494 540464 415258
rect 540144 408258 540186 408494
rect 540422 408258 540464 408494
rect 540144 401494 540464 408258
rect 540144 401258 540186 401494
rect 540422 401258 540464 401494
rect 540144 394494 540464 401258
rect 540144 394258 540186 394494
rect 540422 394258 540464 394494
rect 540144 387494 540464 394258
rect 540144 387258 540186 387494
rect 540422 387258 540464 387494
rect 540144 380494 540464 387258
rect 540144 380258 540186 380494
rect 540422 380258 540464 380494
rect 540144 373494 540464 380258
rect 540144 373258 540186 373494
rect 540422 373258 540464 373494
rect 540144 366494 540464 373258
rect 540144 366258 540186 366494
rect 540422 366258 540464 366494
rect 540144 359494 540464 366258
rect 540144 359258 540186 359494
rect 540422 359258 540464 359494
rect 540144 352494 540464 359258
rect 540144 352258 540186 352494
rect 540422 352258 540464 352494
rect 540144 345494 540464 352258
rect 540144 345258 540186 345494
rect 540422 345258 540464 345494
rect 540144 338494 540464 345258
rect 540144 338258 540186 338494
rect 540422 338258 540464 338494
rect 540144 331494 540464 338258
rect 540144 331258 540186 331494
rect 540422 331258 540464 331494
rect 540144 324494 540464 331258
rect 540144 324258 540186 324494
rect 540422 324258 540464 324494
rect 540144 317494 540464 324258
rect 540144 317258 540186 317494
rect 540422 317258 540464 317494
rect 540144 310494 540464 317258
rect 540144 310258 540186 310494
rect 540422 310258 540464 310494
rect 540144 303494 540464 310258
rect 540144 303258 540186 303494
rect 540422 303258 540464 303494
rect 540144 296494 540464 303258
rect 540144 296258 540186 296494
rect 540422 296258 540464 296494
rect 540144 289494 540464 296258
rect 540144 289258 540186 289494
rect 540422 289258 540464 289494
rect 540144 282494 540464 289258
rect 540144 282258 540186 282494
rect 540422 282258 540464 282494
rect 540144 275494 540464 282258
rect 540144 275258 540186 275494
rect 540422 275258 540464 275494
rect 540144 268494 540464 275258
rect 540144 268258 540186 268494
rect 540422 268258 540464 268494
rect 540144 261494 540464 268258
rect 540144 261258 540186 261494
rect 540422 261258 540464 261494
rect 540144 254494 540464 261258
rect 540144 254258 540186 254494
rect 540422 254258 540464 254494
rect 540144 247494 540464 254258
rect 540144 247258 540186 247494
rect 540422 247258 540464 247494
rect 540144 240494 540464 247258
rect 540144 240258 540186 240494
rect 540422 240258 540464 240494
rect 540144 233494 540464 240258
rect 540144 233258 540186 233494
rect 540422 233258 540464 233494
rect 540144 226494 540464 233258
rect 540144 226258 540186 226494
rect 540422 226258 540464 226494
rect 540144 219494 540464 226258
rect 540144 219258 540186 219494
rect 540422 219258 540464 219494
rect 540144 212494 540464 219258
rect 540144 212258 540186 212494
rect 540422 212258 540464 212494
rect 540144 205494 540464 212258
rect 540144 205258 540186 205494
rect 540422 205258 540464 205494
rect 540144 198494 540464 205258
rect 540144 198258 540186 198494
rect 540422 198258 540464 198494
rect 540144 191494 540464 198258
rect 540144 191258 540186 191494
rect 540422 191258 540464 191494
rect 540144 184494 540464 191258
rect 540144 184258 540186 184494
rect 540422 184258 540464 184494
rect 540144 177494 540464 184258
rect 540144 177258 540186 177494
rect 540422 177258 540464 177494
rect 540144 170494 540464 177258
rect 540144 170258 540186 170494
rect 540422 170258 540464 170494
rect 540144 163494 540464 170258
rect 540144 163258 540186 163494
rect 540422 163258 540464 163494
rect 540144 156494 540464 163258
rect 540144 156258 540186 156494
rect 540422 156258 540464 156494
rect 540144 149494 540464 156258
rect 540144 149258 540186 149494
rect 540422 149258 540464 149494
rect 540144 142494 540464 149258
rect 540144 142258 540186 142494
rect 540422 142258 540464 142494
rect 540144 135494 540464 142258
rect 540144 135258 540186 135494
rect 540422 135258 540464 135494
rect 540144 128494 540464 135258
rect 540144 128258 540186 128494
rect 540422 128258 540464 128494
rect 540144 121494 540464 128258
rect 540144 121258 540186 121494
rect 540422 121258 540464 121494
rect 540144 114494 540464 121258
rect 540144 114258 540186 114494
rect 540422 114258 540464 114494
rect 540144 107494 540464 114258
rect 540144 107258 540186 107494
rect 540422 107258 540464 107494
rect 540144 100494 540464 107258
rect 540144 100258 540186 100494
rect 540422 100258 540464 100494
rect 540144 93494 540464 100258
rect 540144 93258 540186 93494
rect 540422 93258 540464 93494
rect 540144 86494 540464 93258
rect 540144 86258 540186 86494
rect 540422 86258 540464 86494
rect 540144 79494 540464 86258
rect 540144 79258 540186 79494
rect 540422 79258 540464 79494
rect 540144 72494 540464 79258
rect 540144 72258 540186 72494
rect 540422 72258 540464 72494
rect 540144 65494 540464 72258
rect 540144 65258 540186 65494
rect 540422 65258 540464 65494
rect 540144 58494 540464 65258
rect 540144 58258 540186 58494
rect 540422 58258 540464 58494
rect 540144 51494 540464 58258
rect 540144 51258 540186 51494
rect 540422 51258 540464 51494
rect 540144 44494 540464 51258
rect 540144 44258 540186 44494
rect 540422 44258 540464 44494
rect 540144 37494 540464 44258
rect 540144 37258 540186 37494
rect 540422 37258 540464 37494
rect 540144 30494 540464 37258
rect 540144 30258 540186 30494
rect 540422 30258 540464 30494
rect 540144 23494 540464 30258
rect 540144 23258 540186 23494
rect 540422 23258 540464 23494
rect 540144 16494 540464 23258
rect 540144 16258 540186 16494
rect 540422 16258 540464 16494
rect 540144 9494 540464 16258
rect 540144 9258 540186 9494
rect 540422 9258 540464 9494
rect 540144 2494 540464 9258
rect 540144 2258 540186 2494
rect 540422 2258 540464 2494
rect 540144 -746 540464 2258
rect 540144 -982 540186 -746
rect 540422 -982 540464 -746
rect 540144 -1066 540464 -982
rect 540144 -1302 540186 -1066
rect 540422 -1302 540464 -1066
rect 540144 -2294 540464 -1302
rect 541876 706198 542196 706230
rect 541876 705962 541918 706198
rect 542154 705962 542196 706198
rect 541876 705878 542196 705962
rect 541876 705642 541918 705878
rect 542154 705642 542196 705878
rect 541876 696434 542196 705642
rect 541876 696198 541918 696434
rect 542154 696198 542196 696434
rect 541876 689434 542196 696198
rect 541876 689198 541918 689434
rect 542154 689198 542196 689434
rect 541876 682434 542196 689198
rect 541876 682198 541918 682434
rect 542154 682198 542196 682434
rect 541876 675434 542196 682198
rect 541876 675198 541918 675434
rect 542154 675198 542196 675434
rect 541876 668434 542196 675198
rect 541876 668198 541918 668434
rect 542154 668198 542196 668434
rect 541876 661434 542196 668198
rect 541876 661198 541918 661434
rect 542154 661198 542196 661434
rect 541876 654434 542196 661198
rect 541876 654198 541918 654434
rect 542154 654198 542196 654434
rect 541876 647434 542196 654198
rect 541876 647198 541918 647434
rect 542154 647198 542196 647434
rect 541876 640434 542196 647198
rect 541876 640198 541918 640434
rect 542154 640198 542196 640434
rect 541876 633434 542196 640198
rect 541876 633198 541918 633434
rect 542154 633198 542196 633434
rect 541876 626434 542196 633198
rect 541876 626198 541918 626434
rect 542154 626198 542196 626434
rect 541876 619434 542196 626198
rect 541876 619198 541918 619434
rect 542154 619198 542196 619434
rect 541876 612434 542196 619198
rect 541876 612198 541918 612434
rect 542154 612198 542196 612434
rect 541876 605434 542196 612198
rect 541876 605198 541918 605434
rect 542154 605198 542196 605434
rect 541876 598434 542196 605198
rect 541876 598198 541918 598434
rect 542154 598198 542196 598434
rect 541876 591434 542196 598198
rect 541876 591198 541918 591434
rect 542154 591198 542196 591434
rect 541876 584434 542196 591198
rect 541876 584198 541918 584434
rect 542154 584198 542196 584434
rect 541876 577434 542196 584198
rect 541876 577198 541918 577434
rect 542154 577198 542196 577434
rect 541876 570434 542196 577198
rect 541876 570198 541918 570434
rect 542154 570198 542196 570434
rect 541876 563434 542196 570198
rect 541876 563198 541918 563434
rect 542154 563198 542196 563434
rect 541876 556434 542196 563198
rect 541876 556198 541918 556434
rect 542154 556198 542196 556434
rect 541876 549434 542196 556198
rect 541876 549198 541918 549434
rect 542154 549198 542196 549434
rect 541876 542434 542196 549198
rect 541876 542198 541918 542434
rect 542154 542198 542196 542434
rect 541876 535434 542196 542198
rect 541876 535198 541918 535434
rect 542154 535198 542196 535434
rect 541876 528434 542196 535198
rect 541876 528198 541918 528434
rect 542154 528198 542196 528434
rect 541876 521434 542196 528198
rect 541876 521198 541918 521434
rect 542154 521198 542196 521434
rect 541876 514434 542196 521198
rect 541876 514198 541918 514434
rect 542154 514198 542196 514434
rect 541876 507434 542196 514198
rect 541876 507198 541918 507434
rect 542154 507198 542196 507434
rect 541876 500434 542196 507198
rect 541876 500198 541918 500434
rect 542154 500198 542196 500434
rect 541876 493434 542196 500198
rect 541876 493198 541918 493434
rect 542154 493198 542196 493434
rect 541876 486434 542196 493198
rect 541876 486198 541918 486434
rect 542154 486198 542196 486434
rect 541876 479434 542196 486198
rect 541876 479198 541918 479434
rect 542154 479198 542196 479434
rect 541876 472434 542196 479198
rect 541876 472198 541918 472434
rect 542154 472198 542196 472434
rect 541876 465434 542196 472198
rect 541876 465198 541918 465434
rect 542154 465198 542196 465434
rect 541876 458434 542196 465198
rect 541876 458198 541918 458434
rect 542154 458198 542196 458434
rect 541876 451434 542196 458198
rect 541876 451198 541918 451434
rect 542154 451198 542196 451434
rect 541876 444434 542196 451198
rect 541876 444198 541918 444434
rect 542154 444198 542196 444434
rect 541876 437434 542196 444198
rect 541876 437198 541918 437434
rect 542154 437198 542196 437434
rect 541876 430434 542196 437198
rect 541876 430198 541918 430434
rect 542154 430198 542196 430434
rect 541876 423434 542196 430198
rect 541876 423198 541918 423434
rect 542154 423198 542196 423434
rect 541876 416434 542196 423198
rect 541876 416198 541918 416434
rect 542154 416198 542196 416434
rect 541876 409434 542196 416198
rect 541876 409198 541918 409434
rect 542154 409198 542196 409434
rect 541876 402434 542196 409198
rect 541876 402198 541918 402434
rect 542154 402198 542196 402434
rect 541876 395434 542196 402198
rect 541876 395198 541918 395434
rect 542154 395198 542196 395434
rect 541876 388434 542196 395198
rect 541876 388198 541918 388434
rect 542154 388198 542196 388434
rect 541876 381434 542196 388198
rect 541876 381198 541918 381434
rect 542154 381198 542196 381434
rect 541876 374434 542196 381198
rect 541876 374198 541918 374434
rect 542154 374198 542196 374434
rect 541876 367434 542196 374198
rect 541876 367198 541918 367434
rect 542154 367198 542196 367434
rect 541876 360434 542196 367198
rect 541876 360198 541918 360434
rect 542154 360198 542196 360434
rect 541876 353434 542196 360198
rect 541876 353198 541918 353434
rect 542154 353198 542196 353434
rect 541876 346434 542196 353198
rect 541876 346198 541918 346434
rect 542154 346198 542196 346434
rect 541876 339434 542196 346198
rect 541876 339198 541918 339434
rect 542154 339198 542196 339434
rect 541876 332434 542196 339198
rect 541876 332198 541918 332434
rect 542154 332198 542196 332434
rect 541876 325434 542196 332198
rect 541876 325198 541918 325434
rect 542154 325198 542196 325434
rect 541876 318434 542196 325198
rect 541876 318198 541918 318434
rect 542154 318198 542196 318434
rect 541876 311434 542196 318198
rect 541876 311198 541918 311434
rect 542154 311198 542196 311434
rect 541876 304434 542196 311198
rect 541876 304198 541918 304434
rect 542154 304198 542196 304434
rect 541876 297434 542196 304198
rect 541876 297198 541918 297434
rect 542154 297198 542196 297434
rect 541876 290434 542196 297198
rect 541876 290198 541918 290434
rect 542154 290198 542196 290434
rect 541876 283434 542196 290198
rect 541876 283198 541918 283434
rect 542154 283198 542196 283434
rect 541876 276434 542196 283198
rect 541876 276198 541918 276434
rect 542154 276198 542196 276434
rect 541876 269434 542196 276198
rect 541876 269198 541918 269434
rect 542154 269198 542196 269434
rect 541876 262434 542196 269198
rect 541876 262198 541918 262434
rect 542154 262198 542196 262434
rect 541876 255434 542196 262198
rect 541876 255198 541918 255434
rect 542154 255198 542196 255434
rect 541876 248434 542196 255198
rect 541876 248198 541918 248434
rect 542154 248198 542196 248434
rect 541876 241434 542196 248198
rect 541876 241198 541918 241434
rect 542154 241198 542196 241434
rect 541876 234434 542196 241198
rect 541876 234198 541918 234434
rect 542154 234198 542196 234434
rect 541876 227434 542196 234198
rect 541876 227198 541918 227434
rect 542154 227198 542196 227434
rect 541876 220434 542196 227198
rect 541876 220198 541918 220434
rect 542154 220198 542196 220434
rect 541876 213434 542196 220198
rect 541876 213198 541918 213434
rect 542154 213198 542196 213434
rect 541876 206434 542196 213198
rect 541876 206198 541918 206434
rect 542154 206198 542196 206434
rect 541876 199434 542196 206198
rect 541876 199198 541918 199434
rect 542154 199198 542196 199434
rect 541876 192434 542196 199198
rect 541876 192198 541918 192434
rect 542154 192198 542196 192434
rect 541876 185434 542196 192198
rect 541876 185198 541918 185434
rect 542154 185198 542196 185434
rect 541876 178434 542196 185198
rect 541876 178198 541918 178434
rect 542154 178198 542196 178434
rect 541876 171434 542196 178198
rect 541876 171198 541918 171434
rect 542154 171198 542196 171434
rect 541876 164434 542196 171198
rect 541876 164198 541918 164434
rect 542154 164198 542196 164434
rect 541876 157434 542196 164198
rect 541876 157198 541918 157434
rect 542154 157198 542196 157434
rect 541876 150434 542196 157198
rect 541876 150198 541918 150434
rect 542154 150198 542196 150434
rect 541876 143434 542196 150198
rect 541876 143198 541918 143434
rect 542154 143198 542196 143434
rect 541876 136434 542196 143198
rect 541876 136198 541918 136434
rect 542154 136198 542196 136434
rect 541876 129434 542196 136198
rect 541876 129198 541918 129434
rect 542154 129198 542196 129434
rect 541876 122434 542196 129198
rect 541876 122198 541918 122434
rect 542154 122198 542196 122434
rect 541876 115434 542196 122198
rect 541876 115198 541918 115434
rect 542154 115198 542196 115434
rect 541876 108434 542196 115198
rect 541876 108198 541918 108434
rect 542154 108198 542196 108434
rect 541876 101434 542196 108198
rect 541876 101198 541918 101434
rect 542154 101198 542196 101434
rect 541876 94434 542196 101198
rect 541876 94198 541918 94434
rect 542154 94198 542196 94434
rect 541876 87434 542196 94198
rect 541876 87198 541918 87434
rect 542154 87198 542196 87434
rect 541876 80434 542196 87198
rect 541876 80198 541918 80434
rect 542154 80198 542196 80434
rect 541876 73434 542196 80198
rect 541876 73198 541918 73434
rect 542154 73198 542196 73434
rect 541876 66434 542196 73198
rect 541876 66198 541918 66434
rect 542154 66198 542196 66434
rect 541876 59434 542196 66198
rect 541876 59198 541918 59434
rect 542154 59198 542196 59434
rect 541876 52434 542196 59198
rect 541876 52198 541918 52434
rect 542154 52198 542196 52434
rect 541876 45434 542196 52198
rect 541876 45198 541918 45434
rect 542154 45198 542196 45434
rect 541876 38434 542196 45198
rect 541876 38198 541918 38434
rect 542154 38198 542196 38434
rect 541876 31434 542196 38198
rect 541876 31198 541918 31434
rect 542154 31198 542196 31434
rect 541876 24434 542196 31198
rect 541876 24198 541918 24434
rect 542154 24198 542196 24434
rect 541876 17434 542196 24198
rect 541876 17198 541918 17434
rect 542154 17198 542196 17434
rect 541876 10434 542196 17198
rect 541876 10198 541918 10434
rect 542154 10198 542196 10434
rect 541876 3434 542196 10198
rect 541876 3198 541918 3434
rect 542154 3198 542196 3434
rect 541876 -1706 542196 3198
rect 541876 -1942 541918 -1706
rect 542154 -1942 542196 -1706
rect 541876 -2026 542196 -1942
rect 541876 -2262 541918 -2026
rect 542154 -2262 542196 -2026
rect 541876 -2294 542196 -2262
rect 547144 705238 547464 706230
rect 547144 705002 547186 705238
rect 547422 705002 547464 705238
rect 547144 704918 547464 705002
rect 547144 704682 547186 704918
rect 547422 704682 547464 704918
rect 547144 695494 547464 704682
rect 547144 695258 547186 695494
rect 547422 695258 547464 695494
rect 547144 688494 547464 695258
rect 547144 688258 547186 688494
rect 547422 688258 547464 688494
rect 547144 681494 547464 688258
rect 547144 681258 547186 681494
rect 547422 681258 547464 681494
rect 547144 674494 547464 681258
rect 547144 674258 547186 674494
rect 547422 674258 547464 674494
rect 547144 667494 547464 674258
rect 547144 667258 547186 667494
rect 547422 667258 547464 667494
rect 547144 660494 547464 667258
rect 547144 660258 547186 660494
rect 547422 660258 547464 660494
rect 547144 653494 547464 660258
rect 547144 653258 547186 653494
rect 547422 653258 547464 653494
rect 547144 646494 547464 653258
rect 547144 646258 547186 646494
rect 547422 646258 547464 646494
rect 547144 639494 547464 646258
rect 547144 639258 547186 639494
rect 547422 639258 547464 639494
rect 547144 632494 547464 639258
rect 547144 632258 547186 632494
rect 547422 632258 547464 632494
rect 547144 625494 547464 632258
rect 547144 625258 547186 625494
rect 547422 625258 547464 625494
rect 547144 618494 547464 625258
rect 547144 618258 547186 618494
rect 547422 618258 547464 618494
rect 547144 611494 547464 618258
rect 547144 611258 547186 611494
rect 547422 611258 547464 611494
rect 547144 604494 547464 611258
rect 547144 604258 547186 604494
rect 547422 604258 547464 604494
rect 547144 597494 547464 604258
rect 547144 597258 547186 597494
rect 547422 597258 547464 597494
rect 547144 590494 547464 597258
rect 547144 590258 547186 590494
rect 547422 590258 547464 590494
rect 547144 583494 547464 590258
rect 547144 583258 547186 583494
rect 547422 583258 547464 583494
rect 547144 576494 547464 583258
rect 547144 576258 547186 576494
rect 547422 576258 547464 576494
rect 547144 569494 547464 576258
rect 547144 569258 547186 569494
rect 547422 569258 547464 569494
rect 547144 562494 547464 569258
rect 547144 562258 547186 562494
rect 547422 562258 547464 562494
rect 547144 555494 547464 562258
rect 547144 555258 547186 555494
rect 547422 555258 547464 555494
rect 547144 548494 547464 555258
rect 547144 548258 547186 548494
rect 547422 548258 547464 548494
rect 547144 541494 547464 548258
rect 547144 541258 547186 541494
rect 547422 541258 547464 541494
rect 547144 534494 547464 541258
rect 547144 534258 547186 534494
rect 547422 534258 547464 534494
rect 547144 527494 547464 534258
rect 547144 527258 547186 527494
rect 547422 527258 547464 527494
rect 547144 520494 547464 527258
rect 547144 520258 547186 520494
rect 547422 520258 547464 520494
rect 547144 513494 547464 520258
rect 547144 513258 547186 513494
rect 547422 513258 547464 513494
rect 547144 506494 547464 513258
rect 547144 506258 547186 506494
rect 547422 506258 547464 506494
rect 547144 499494 547464 506258
rect 547144 499258 547186 499494
rect 547422 499258 547464 499494
rect 547144 492494 547464 499258
rect 547144 492258 547186 492494
rect 547422 492258 547464 492494
rect 547144 485494 547464 492258
rect 547144 485258 547186 485494
rect 547422 485258 547464 485494
rect 547144 478494 547464 485258
rect 547144 478258 547186 478494
rect 547422 478258 547464 478494
rect 547144 471494 547464 478258
rect 547144 471258 547186 471494
rect 547422 471258 547464 471494
rect 547144 464494 547464 471258
rect 547144 464258 547186 464494
rect 547422 464258 547464 464494
rect 547144 457494 547464 464258
rect 547144 457258 547186 457494
rect 547422 457258 547464 457494
rect 547144 450494 547464 457258
rect 547144 450258 547186 450494
rect 547422 450258 547464 450494
rect 547144 443494 547464 450258
rect 547144 443258 547186 443494
rect 547422 443258 547464 443494
rect 547144 436494 547464 443258
rect 547144 436258 547186 436494
rect 547422 436258 547464 436494
rect 547144 429494 547464 436258
rect 547144 429258 547186 429494
rect 547422 429258 547464 429494
rect 547144 422494 547464 429258
rect 547144 422258 547186 422494
rect 547422 422258 547464 422494
rect 547144 415494 547464 422258
rect 547144 415258 547186 415494
rect 547422 415258 547464 415494
rect 547144 408494 547464 415258
rect 547144 408258 547186 408494
rect 547422 408258 547464 408494
rect 547144 401494 547464 408258
rect 547144 401258 547186 401494
rect 547422 401258 547464 401494
rect 547144 394494 547464 401258
rect 547144 394258 547186 394494
rect 547422 394258 547464 394494
rect 547144 387494 547464 394258
rect 547144 387258 547186 387494
rect 547422 387258 547464 387494
rect 547144 380494 547464 387258
rect 547144 380258 547186 380494
rect 547422 380258 547464 380494
rect 547144 373494 547464 380258
rect 547144 373258 547186 373494
rect 547422 373258 547464 373494
rect 547144 366494 547464 373258
rect 547144 366258 547186 366494
rect 547422 366258 547464 366494
rect 547144 359494 547464 366258
rect 547144 359258 547186 359494
rect 547422 359258 547464 359494
rect 547144 352494 547464 359258
rect 547144 352258 547186 352494
rect 547422 352258 547464 352494
rect 547144 345494 547464 352258
rect 547144 345258 547186 345494
rect 547422 345258 547464 345494
rect 547144 338494 547464 345258
rect 547144 338258 547186 338494
rect 547422 338258 547464 338494
rect 547144 331494 547464 338258
rect 547144 331258 547186 331494
rect 547422 331258 547464 331494
rect 547144 324494 547464 331258
rect 547144 324258 547186 324494
rect 547422 324258 547464 324494
rect 547144 317494 547464 324258
rect 547144 317258 547186 317494
rect 547422 317258 547464 317494
rect 547144 310494 547464 317258
rect 547144 310258 547186 310494
rect 547422 310258 547464 310494
rect 547144 303494 547464 310258
rect 547144 303258 547186 303494
rect 547422 303258 547464 303494
rect 547144 296494 547464 303258
rect 547144 296258 547186 296494
rect 547422 296258 547464 296494
rect 547144 289494 547464 296258
rect 547144 289258 547186 289494
rect 547422 289258 547464 289494
rect 547144 282494 547464 289258
rect 547144 282258 547186 282494
rect 547422 282258 547464 282494
rect 547144 275494 547464 282258
rect 547144 275258 547186 275494
rect 547422 275258 547464 275494
rect 547144 268494 547464 275258
rect 547144 268258 547186 268494
rect 547422 268258 547464 268494
rect 547144 261494 547464 268258
rect 547144 261258 547186 261494
rect 547422 261258 547464 261494
rect 547144 254494 547464 261258
rect 547144 254258 547186 254494
rect 547422 254258 547464 254494
rect 547144 247494 547464 254258
rect 547144 247258 547186 247494
rect 547422 247258 547464 247494
rect 547144 240494 547464 247258
rect 547144 240258 547186 240494
rect 547422 240258 547464 240494
rect 547144 233494 547464 240258
rect 547144 233258 547186 233494
rect 547422 233258 547464 233494
rect 547144 226494 547464 233258
rect 547144 226258 547186 226494
rect 547422 226258 547464 226494
rect 547144 219494 547464 226258
rect 547144 219258 547186 219494
rect 547422 219258 547464 219494
rect 547144 212494 547464 219258
rect 547144 212258 547186 212494
rect 547422 212258 547464 212494
rect 547144 205494 547464 212258
rect 547144 205258 547186 205494
rect 547422 205258 547464 205494
rect 547144 198494 547464 205258
rect 547144 198258 547186 198494
rect 547422 198258 547464 198494
rect 547144 191494 547464 198258
rect 547144 191258 547186 191494
rect 547422 191258 547464 191494
rect 547144 184494 547464 191258
rect 547144 184258 547186 184494
rect 547422 184258 547464 184494
rect 547144 177494 547464 184258
rect 547144 177258 547186 177494
rect 547422 177258 547464 177494
rect 547144 170494 547464 177258
rect 547144 170258 547186 170494
rect 547422 170258 547464 170494
rect 547144 163494 547464 170258
rect 547144 163258 547186 163494
rect 547422 163258 547464 163494
rect 547144 156494 547464 163258
rect 547144 156258 547186 156494
rect 547422 156258 547464 156494
rect 547144 149494 547464 156258
rect 547144 149258 547186 149494
rect 547422 149258 547464 149494
rect 547144 142494 547464 149258
rect 547144 142258 547186 142494
rect 547422 142258 547464 142494
rect 547144 135494 547464 142258
rect 547144 135258 547186 135494
rect 547422 135258 547464 135494
rect 547144 128494 547464 135258
rect 547144 128258 547186 128494
rect 547422 128258 547464 128494
rect 547144 121494 547464 128258
rect 547144 121258 547186 121494
rect 547422 121258 547464 121494
rect 547144 114494 547464 121258
rect 547144 114258 547186 114494
rect 547422 114258 547464 114494
rect 547144 107494 547464 114258
rect 547144 107258 547186 107494
rect 547422 107258 547464 107494
rect 547144 100494 547464 107258
rect 547144 100258 547186 100494
rect 547422 100258 547464 100494
rect 547144 93494 547464 100258
rect 547144 93258 547186 93494
rect 547422 93258 547464 93494
rect 547144 86494 547464 93258
rect 547144 86258 547186 86494
rect 547422 86258 547464 86494
rect 547144 79494 547464 86258
rect 547144 79258 547186 79494
rect 547422 79258 547464 79494
rect 547144 72494 547464 79258
rect 547144 72258 547186 72494
rect 547422 72258 547464 72494
rect 547144 65494 547464 72258
rect 547144 65258 547186 65494
rect 547422 65258 547464 65494
rect 547144 58494 547464 65258
rect 547144 58258 547186 58494
rect 547422 58258 547464 58494
rect 547144 51494 547464 58258
rect 547144 51258 547186 51494
rect 547422 51258 547464 51494
rect 547144 44494 547464 51258
rect 547144 44258 547186 44494
rect 547422 44258 547464 44494
rect 547144 37494 547464 44258
rect 547144 37258 547186 37494
rect 547422 37258 547464 37494
rect 547144 30494 547464 37258
rect 547144 30258 547186 30494
rect 547422 30258 547464 30494
rect 547144 23494 547464 30258
rect 547144 23258 547186 23494
rect 547422 23258 547464 23494
rect 547144 16494 547464 23258
rect 547144 16258 547186 16494
rect 547422 16258 547464 16494
rect 547144 9494 547464 16258
rect 547144 9258 547186 9494
rect 547422 9258 547464 9494
rect 547144 2494 547464 9258
rect 547144 2258 547186 2494
rect 547422 2258 547464 2494
rect 547144 -746 547464 2258
rect 547144 -982 547186 -746
rect 547422 -982 547464 -746
rect 547144 -1066 547464 -982
rect 547144 -1302 547186 -1066
rect 547422 -1302 547464 -1066
rect 547144 -2294 547464 -1302
rect 548876 706198 549196 706230
rect 548876 705962 548918 706198
rect 549154 705962 549196 706198
rect 548876 705878 549196 705962
rect 548876 705642 548918 705878
rect 549154 705642 549196 705878
rect 548876 696434 549196 705642
rect 548876 696198 548918 696434
rect 549154 696198 549196 696434
rect 548876 689434 549196 696198
rect 548876 689198 548918 689434
rect 549154 689198 549196 689434
rect 548876 682434 549196 689198
rect 548876 682198 548918 682434
rect 549154 682198 549196 682434
rect 548876 675434 549196 682198
rect 548876 675198 548918 675434
rect 549154 675198 549196 675434
rect 548876 668434 549196 675198
rect 548876 668198 548918 668434
rect 549154 668198 549196 668434
rect 548876 661434 549196 668198
rect 548876 661198 548918 661434
rect 549154 661198 549196 661434
rect 548876 654434 549196 661198
rect 548876 654198 548918 654434
rect 549154 654198 549196 654434
rect 548876 647434 549196 654198
rect 548876 647198 548918 647434
rect 549154 647198 549196 647434
rect 548876 640434 549196 647198
rect 548876 640198 548918 640434
rect 549154 640198 549196 640434
rect 548876 633434 549196 640198
rect 548876 633198 548918 633434
rect 549154 633198 549196 633434
rect 548876 626434 549196 633198
rect 548876 626198 548918 626434
rect 549154 626198 549196 626434
rect 548876 619434 549196 626198
rect 548876 619198 548918 619434
rect 549154 619198 549196 619434
rect 548876 612434 549196 619198
rect 548876 612198 548918 612434
rect 549154 612198 549196 612434
rect 548876 605434 549196 612198
rect 548876 605198 548918 605434
rect 549154 605198 549196 605434
rect 548876 598434 549196 605198
rect 548876 598198 548918 598434
rect 549154 598198 549196 598434
rect 548876 591434 549196 598198
rect 548876 591198 548918 591434
rect 549154 591198 549196 591434
rect 548876 584434 549196 591198
rect 548876 584198 548918 584434
rect 549154 584198 549196 584434
rect 548876 577434 549196 584198
rect 548876 577198 548918 577434
rect 549154 577198 549196 577434
rect 548876 570434 549196 577198
rect 548876 570198 548918 570434
rect 549154 570198 549196 570434
rect 548876 563434 549196 570198
rect 548876 563198 548918 563434
rect 549154 563198 549196 563434
rect 548876 556434 549196 563198
rect 548876 556198 548918 556434
rect 549154 556198 549196 556434
rect 548876 549434 549196 556198
rect 548876 549198 548918 549434
rect 549154 549198 549196 549434
rect 548876 542434 549196 549198
rect 548876 542198 548918 542434
rect 549154 542198 549196 542434
rect 548876 535434 549196 542198
rect 548876 535198 548918 535434
rect 549154 535198 549196 535434
rect 548876 528434 549196 535198
rect 548876 528198 548918 528434
rect 549154 528198 549196 528434
rect 548876 521434 549196 528198
rect 548876 521198 548918 521434
rect 549154 521198 549196 521434
rect 548876 514434 549196 521198
rect 548876 514198 548918 514434
rect 549154 514198 549196 514434
rect 548876 507434 549196 514198
rect 548876 507198 548918 507434
rect 549154 507198 549196 507434
rect 548876 500434 549196 507198
rect 548876 500198 548918 500434
rect 549154 500198 549196 500434
rect 548876 493434 549196 500198
rect 548876 493198 548918 493434
rect 549154 493198 549196 493434
rect 548876 486434 549196 493198
rect 548876 486198 548918 486434
rect 549154 486198 549196 486434
rect 548876 479434 549196 486198
rect 548876 479198 548918 479434
rect 549154 479198 549196 479434
rect 548876 472434 549196 479198
rect 548876 472198 548918 472434
rect 549154 472198 549196 472434
rect 548876 465434 549196 472198
rect 548876 465198 548918 465434
rect 549154 465198 549196 465434
rect 548876 458434 549196 465198
rect 548876 458198 548918 458434
rect 549154 458198 549196 458434
rect 548876 451434 549196 458198
rect 548876 451198 548918 451434
rect 549154 451198 549196 451434
rect 548876 444434 549196 451198
rect 548876 444198 548918 444434
rect 549154 444198 549196 444434
rect 548876 437434 549196 444198
rect 548876 437198 548918 437434
rect 549154 437198 549196 437434
rect 548876 430434 549196 437198
rect 548876 430198 548918 430434
rect 549154 430198 549196 430434
rect 548876 423434 549196 430198
rect 548876 423198 548918 423434
rect 549154 423198 549196 423434
rect 548876 416434 549196 423198
rect 548876 416198 548918 416434
rect 549154 416198 549196 416434
rect 548876 409434 549196 416198
rect 548876 409198 548918 409434
rect 549154 409198 549196 409434
rect 548876 402434 549196 409198
rect 548876 402198 548918 402434
rect 549154 402198 549196 402434
rect 548876 395434 549196 402198
rect 548876 395198 548918 395434
rect 549154 395198 549196 395434
rect 548876 388434 549196 395198
rect 548876 388198 548918 388434
rect 549154 388198 549196 388434
rect 548876 381434 549196 388198
rect 548876 381198 548918 381434
rect 549154 381198 549196 381434
rect 548876 374434 549196 381198
rect 548876 374198 548918 374434
rect 549154 374198 549196 374434
rect 548876 367434 549196 374198
rect 548876 367198 548918 367434
rect 549154 367198 549196 367434
rect 548876 360434 549196 367198
rect 548876 360198 548918 360434
rect 549154 360198 549196 360434
rect 548876 353434 549196 360198
rect 548876 353198 548918 353434
rect 549154 353198 549196 353434
rect 548876 346434 549196 353198
rect 548876 346198 548918 346434
rect 549154 346198 549196 346434
rect 548876 339434 549196 346198
rect 548876 339198 548918 339434
rect 549154 339198 549196 339434
rect 548876 332434 549196 339198
rect 548876 332198 548918 332434
rect 549154 332198 549196 332434
rect 548876 325434 549196 332198
rect 548876 325198 548918 325434
rect 549154 325198 549196 325434
rect 548876 318434 549196 325198
rect 548876 318198 548918 318434
rect 549154 318198 549196 318434
rect 548876 311434 549196 318198
rect 548876 311198 548918 311434
rect 549154 311198 549196 311434
rect 548876 304434 549196 311198
rect 548876 304198 548918 304434
rect 549154 304198 549196 304434
rect 548876 297434 549196 304198
rect 548876 297198 548918 297434
rect 549154 297198 549196 297434
rect 548876 290434 549196 297198
rect 548876 290198 548918 290434
rect 549154 290198 549196 290434
rect 548876 283434 549196 290198
rect 548876 283198 548918 283434
rect 549154 283198 549196 283434
rect 548876 276434 549196 283198
rect 548876 276198 548918 276434
rect 549154 276198 549196 276434
rect 548876 269434 549196 276198
rect 548876 269198 548918 269434
rect 549154 269198 549196 269434
rect 548876 262434 549196 269198
rect 548876 262198 548918 262434
rect 549154 262198 549196 262434
rect 548876 255434 549196 262198
rect 548876 255198 548918 255434
rect 549154 255198 549196 255434
rect 548876 248434 549196 255198
rect 548876 248198 548918 248434
rect 549154 248198 549196 248434
rect 548876 241434 549196 248198
rect 548876 241198 548918 241434
rect 549154 241198 549196 241434
rect 548876 234434 549196 241198
rect 548876 234198 548918 234434
rect 549154 234198 549196 234434
rect 548876 227434 549196 234198
rect 548876 227198 548918 227434
rect 549154 227198 549196 227434
rect 548876 220434 549196 227198
rect 548876 220198 548918 220434
rect 549154 220198 549196 220434
rect 548876 213434 549196 220198
rect 548876 213198 548918 213434
rect 549154 213198 549196 213434
rect 548876 206434 549196 213198
rect 548876 206198 548918 206434
rect 549154 206198 549196 206434
rect 548876 199434 549196 206198
rect 548876 199198 548918 199434
rect 549154 199198 549196 199434
rect 548876 192434 549196 199198
rect 548876 192198 548918 192434
rect 549154 192198 549196 192434
rect 548876 185434 549196 192198
rect 548876 185198 548918 185434
rect 549154 185198 549196 185434
rect 548876 178434 549196 185198
rect 548876 178198 548918 178434
rect 549154 178198 549196 178434
rect 548876 171434 549196 178198
rect 548876 171198 548918 171434
rect 549154 171198 549196 171434
rect 548876 164434 549196 171198
rect 548876 164198 548918 164434
rect 549154 164198 549196 164434
rect 548876 157434 549196 164198
rect 548876 157198 548918 157434
rect 549154 157198 549196 157434
rect 548876 150434 549196 157198
rect 548876 150198 548918 150434
rect 549154 150198 549196 150434
rect 548876 143434 549196 150198
rect 548876 143198 548918 143434
rect 549154 143198 549196 143434
rect 548876 136434 549196 143198
rect 548876 136198 548918 136434
rect 549154 136198 549196 136434
rect 548876 129434 549196 136198
rect 548876 129198 548918 129434
rect 549154 129198 549196 129434
rect 548876 122434 549196 129198
rect 548876 122198 548918 122434
rect 549154 122198 549196 122434
rect 548876 115434 549196 122198
rect 548876 115198 548918 115434
rect 549154 115198 549196 115434
rect 548876 108434 549196 115198
rect 548876 108198 548918 108434
rect 549154 108198 549196 108434
rect 548876 101434 549196 108198
rect 548876 101198 548918 101434
rect 549154 101198 549196 101434
rect 548876 94434 549196 101198
rect 548876 94198 548918 94434
rect 549154 94198 549196 94434
rect 548876 87434 549196 94198
rect 548876 87198 548918 87434
rect 549154 87198 549196 87434
rect 548876 80434 549196 87198
rect 548876 80198 548918 80434
rect 549154 80198 549196 80434
rect 548876 73434 549196 80198
rect 548876 73198 548918 73434
rect 549154 73198 549196 73434
rect 548876 66434 549196 73198
rect 548876 66198 548918 66434
rect 549154 66198 549196 66434
rect 548876 59434 549196 66198
rect 548876 59198 548918 59434
rect 549154 59198 549196 59434
rect 548876 52434 549196 59198
rect 548876 52198 548918 52434
rect 549154 52198 549196 52434
rect 548876 45434 549196 52198
rect 548876 45198 548918 45434
rect 549154 45198 549196 45434
rect 548876 38434 549196 45198
rect 548876 38198 548918 38434
rect 549154 38198 549196 38434
rect 548876 31434 549196 38198
rect 548876 31198 548918 31434
rect 549154 31198 549196 31434
rect 548876 24434 549196 31198
rect 548876 24198 548918 24434
rect 549154 24198 549196 24434
rect 548876 17434 549196 24198
rect 548876 17198 548918 17434
rect 549154 17198 549196 17434
rect 548876 10434 549196 17198
rect 548876 10198 548918 10434
rect 549154 10198 549196 10434
rect 548876 3434 549196 10198
rect 548876 3198 548918 3434
rect 549154 3198 549196 3434
rect 548876 -1706 549196 3198
rect 548876 -1942 548918 -1706
rect 549154 -1942 549196 -1706
rect 548876 -2026 549196 -1942
rect 548876 -2262 548918 -2026
rect 549154 -2262 549196 -2026
rect 548876 -2294 549196 -2262
rect 554144 705238 554464 706230
rect 554144 705002 554186 705238
rect 554422 705002 554464 705238
rect 554144 704918 554464 705002
rect 554144 704682 554186 704918
rect 554422 704682 554464 704918
rect 554144 695494 554464 704682
rect 554144 695258 554186 695494
rect 554422 695258 554464 695494
rect 554144 688494 554464 695258
rect 554144 688258 554186 688494
rect 554422 688258 554464 688494
rect 554144 681494 554464 688258
rect 554144 681258 554186 681494
rect 554422 681258 554464 681494
rect 554144 674494 554464 681258
rect 554144 674258 554186 674494
rect 554422 674258 554464 674494
rect 554144 667494 554464 674258
rect 554144 667258 554186 667494
rect 554422 667258 554464 667494
rect 554144 660494 554464 667258
rect 554144 660258 554186 660494
rect 554422 660258 554464 660494
rect 554144 653494 554464 660258
rect 554144 653258 554186 653494
rect 554422 653258 554464 653494
rect 554144 646494 554464 653258
rect 554144 646258 554186 646494
rect 554422 646258 554464 646494
rect 554144 639494 554464 646258
rect 554144 639258 554186 639494
rect 554422 639258 554464 639494
rect 554144 632494 554464 639258
rect 554144 632258 554186 632494
rect 554422 632258 554464 632494
rect 554144 625494 554464 632258
rect 554144 625258 554186 625494
rect 554422 625258 554464 625494
rect 554144 618494 554464 625258
rect 554144 618258 554186 618494
rect 554422 618258 554464 618494
rect 554144 611494 554464 618258
rect 554144 611258 554186 611494
rect 554422 611258 554464 611494
rect 554144 604494 554464 611258
rect 554144 604258 554186 604494
rect 554422 604258 554464 604494
rect 554144 597494 554464 604258
rect 554144 597258 554186 597494
rect 554422 597258 554464 597494
rect 554144 590494 554464 597258
rect 554144 590258 554186 590494
rect 554422 590258 554464 590494
rect 554144 583494 554464 590258
rect 554144 583258 554186 583494
rect 554422 583258 554464 583494
rect 554144 576494 554464 583258
rect 554144 576258 554186 576494
rect 554422 576258 554464 576494
rect 554144 569494 554464 576258
rect 554144 569258 554186 569494
rect 554422 569258 554464 569494
rect 554144 562494 554464 569258
rect 554144 562258 554186 562494
rect 554422 562258 554464 562494
rect 554144 555494 554464 562258
rect 554144 555258 554186 555494
rect 554422 555258 554464 555494
rect 554144 548494 554464 555258
rect 554144 548258 554186 548494
rect 554422 548258 554464 548494
rect 554144 541494 554464 548258
rect 554144 541258 554186 541494
rect 554422 541258 554464 541494
rect 554144 534494 554464 541258
rect 554144 534258 554186 534494
rect 554422 534258 554464 534494
rect 554144 527494 554464 534258
rect 554144 527258 554186 527494
rect 554422 527258 554464 527494
rect 554144 520494 554464 527258
rect 554144 520258 554186 520494
rect 554422 520258 554464 520494
rect 554144 513494 554464 520258
rect 554144 513258 554186 513494
rect 554422 513258 554464 513494
rect 554144 506494 554464 513258
rect 554144 506258 554186 506494
rect 554422 506258 554464 506494
rect 554144 499494 554464 506258
rect 554144 499258 554186 499494
rect 554422 499258 554464 499494
rect 554144 492494 554464 499258
rect 554144 492258 554186 492494
rect 554422 492258 554464 492494
rect 554144 485494 554464 492258
rect 554144 485258 554186 485494
rect 554422 485258 554464 485494
rect 554144 478494 554464 485258
rect 554144 478258 554186 478494
rect 554422 478258 554464 478494
rect 554144 471494 554464 478258
rect 554144 471258 554186 471494
rect 554422 471258 554464 471494
rect 554144 464494 554464 471258
rect 554144 464258 554186 464494
rect 554422 464258 554464 464494
rect 554144 457494 554464 464258
rect 554144 457258 554186 457494
rect 554422 457258 554464 457494
rect 554144 450494 554464 457258
rect 554144 450258 554186 450494
rect 554422 450258 554464 450494
rect 554144 443494 554464 450258
rect 554144 443258 554186 443494
rect 554422 443258 554464 443494
rect 554144 436494 554464 443258
rect 554144 436258 554186 436494
rect 554422 436258 554464 436494
rect 554144 429494 554464 436258
rect 554144 429258 554186 429494
rect 554422 429258 554464 429494
rect 554144 422494 554464 429258
rect 554144 422258 554186 422494
rect 554422 422258 554464 422494
rect 554144 415494 554464 422258
rect 554144 415258 554186 415494
rect 554422 415258 554464 415494
rect 554144 408494 554464 415258
rect 554144 408258 554186 408494
rect 554422 408258 554464 408494
rect 554144 401494 554464 408258
rect 554144 401258 554186 401494
rect 554422 401258 554464 401494
rect 554144 394494 554464 401258
rect 554144 394258 554186 394494
rect 554422 394258 554464 394494
rect 554144 387494 554464 394258
rect 554144 387258 554186 387494
rect 554422 387258 554464 387494
rect 554144 380494 554464 387258
rect 554144 380258 554186 380494
rect 554422 380258 554464 380494
rect 554144 373494 554464 380258
rect 554144 373258 554186 373494
rect 554422 373258 554464 373494
rect 554144 366494 554464 373258
rect 554144 366258 554186 366494
rect 554422 366258 554464 366494
rect 554144 359494 554464 366258
rect 554144 359258 554186 359494
rect 554422 359258 554464 359494
rect 554144 352494 554464 359258
rect 554144 352258 554186 352494
rect 554422 352258 554464 352494
rect 554144 345494 554464 352258
rect 554144 345258 554186 345494
rect 554422 345258 554464 345494
rect 554144 338494 554464 345258
rect 554144 338258 554186 338494
rect 554422 338258 554464 338494
rect 554144 331494 554464 338258
rect 554144 331258 554186 331494
rect 554422 331258 554464 331494
rect 554144 324494 554464 331258
rect 554144 324258 554186 324494
rect 554422 324258 554464 324494
rect 554144 317494 554464 324258
rect 554144 317258 554186 317494
rect 554422 317258 554464 317494
rect 554144 310494 554464 317258
rect 554144 310258 554186 310494
rect 554422 310258 554464 310494
rect 554144 303494 554464 310258
rect 554144 303258 554186 303494
rect 554422 303258 554464 303494
rect 554144 296494 554464 303258
rect 554144 296258 554186 296494
rect 554422 296258 554464 296494
rect 554144 289494 554464 296258
rect 554144 289258 554186 289494
rect 554422 289258 554464 289494
rect 554144 282494 554464 289258
rect 554144 282258 554186 282494
rect 554422 282258 554464 282494
rect 554144 275494 554464 282258
rect 554144 275258 554186 275494
rect 554422 275258 554464 275494
rect 554144 268494 554464 275258
rect 554144 268258 554186 268494
rect 554422 268258 554464 268494
rect 554144 261494 554464 268258
rect 554144 261258 554186 261494
rect 554422 261258 554464 261494
rect 554144 254494 554464 261258
rect 554144 254258 554186 254494
rect 554422 254258 554464 254494
rect 554144 247494 554464 254258
rect 554144 247258 554186 247494
rect 554422 247258 554464 247494
rect 554144 240494 554464 247258
rect 554144 240258 554186 240494
rect 554422 240258 554464 240494
rect 554144 233494 554464 240258
rect 554144 233258 554186 233494
rect 554422 233258 554464 233494
rect 554144 226494 554464 233258
rect 554144 226258 554186 226494
rect 554422 226258 554464 226494
rect 554144 219494 554464 226258
rect 554144 219258 554186 219494
rect 554422 219258 554464 219494
rect 554144 212494 554464 219258
rect 554144 212258 554186 212494
rect 554422 212258 554464 212494
rect 554144 205494 554464 212258
rect 554144 205258 554186 205494
rect 554422 205258 554464 205494
rect 554144 198494 554464 205258
rect 554144 198258 554186 198494
rect 554422 198258 554464 198494
rect 554144 191494 554464 198258
rect 554144 191258 554186 191494
rect 554422 191258 554464 191494
rect 554144 184494 554464 191258
rect 554144 184258 554186 184494
rect 554422 184258 554464 184494
rect 554144 177494 554464 184258
rect 554144 177258 554186 177494
rect 554422 177258 554464 177494
rect 554144 170494 554464 177258
rect 554144 170258 554186 170494
rect 554422 170258 554464 170494
rect 554144 163494 554464 170258
rect 554144 163258 554186 163494
rect 554422 163258 554464 163494
rect 554144 156494 554464 163258
rect 554144 156258 554186 156494
rect 554422 156258 554464 156494
rect 554144 149494 554464 156258
rect 554144 149258 554186 149494
rect 554422 149258 554464 149494
rect 554144 142494 554464 149258
rect 554144 142258 554186 142494
rect 554422 142258 554464 142494
rect 554144 135494 554464 142258
rect 554144 135258 554186 135494
rect 554422 135258 554464 135494
rect 554144 128494 554464 135258
rect 554144 128258 554186 128494
rect 554422 128258 554464 128494
rect 554144 121494 554464 128258
rect 554144 121258 554186 121494
rect 554422 121258 554464 121494
rect 554144 114494 554464 121258
rect 554144 114258 554186 114494
rect 554422 114258 554464 114494
rect 554144 107494 554464 114258
rect 554144 107258 554186 107494
rect 554422 107258 554464 107494
rect 554144 100494 554464 107258
rect 554144 100258 554186 100494
rect 554422 100258 554464 100494
rect 554144 93494 554464 100258
rect 554144 93258 554186 93494
rect 554422 93258 554464 93494
rect 554144 86494 554464 93258
rect 554144 86258 554186 86494
rect 554422 86258 554464 86494
rect 554144 79494 554464 86258
rect 554144 79258 554186 79494
rect 554422 79258 554464 79494
rect 554144 72494 554464 79258
rect 554144 72258 554186 72494
rect 554422 72258 554464 72494
rect 554144 65494 554464 72258
rect 554144 65258 554186 65494
rect 554422 65258 554464 65494
rect 554144 58494 554464 65258
rect 554144 58258 554186 58494
rect 554422 58258 554464 58494
rect 554144 51494 554464 58258
rect 554144 51258 554186 51494
rect 554422 51258 554464 51494
rect 554144 44494 554464 51258
rect 554144 44258 554186 44494
rect 554422 44258 554464 44494
rect 554144 37494 554464 44258
rect 554144 37258 554186 37494
rect 554422 37258 554464 37494
rect 554144 30494 554464 37258
rect 554144 30258 554186 30494
rect 554422 30258 554464 30494
rect 554144 23494 554464 30258
rect 554144 23258 554186 23494
rect 554422 23258 554464 23494
rect 554144 16494 554464 23258
rect 554144 16258 554186 16494
rect 554422 16258 554464 16494
rect 554144 9494 554464 16258
rect 554144 9258 554186 9494
rect 554422 9258 554464 9494
rect 554144 2494 554464 9258
rect 554144 2258 554186 2494
rect 554422 2258 554464 2494
rect 554144 -746 554464 2258
rect 554144 -982 554186 -746
rect 554422 -982 554464 -746
rect 554144 -1066 554464 -982
rect 554144 -1302 554186 -1066
rect 554422 -1302 554464 -1066
rect 554144 -2294 554464 -1302
rect 555876 706198 556196 706230
rect 555876 705962 555918 706198
rect 556154 705962 556196 706198
rect 555876 705878 556196 705962
rect 555876 705642 555918 705878
rect 556154 705642 556196 705878
rect 555876 696434 556196 705642
rect 555876 696198 555918 696434
rect 556154 696198 556196 696434
rect 555876 689434 556196 696198
rect 555876 689198 555918 689434
rect 556154 689198 556196 689434
rect 555876 682434 556196 689198
rect 555876 682198 555918 682434
rect 556154 682198 556196 682434
rect 555876 675434 556196 682198
rect 555876 675198 555918 675434
rect 556154 675198 556196 675434
rect 555876 668434 556196 675198
rect 555876 668198 555918 668434
rect 556154 668198 556196 668434
rect 555876 661434 556196 668198
rect 555876 661198 555918 661434
rect 556154 661198 556196 661434
rect 555876 654434 556196 661198
rect 555876 654198 555918 654434
rect 556154 654198 556196 654434
rect 555876 647434 556196 654198
rect 555876 647198 555918 647434
rect 556154 647198 556196 647434
rect 555876 640434 556196 647198
rect 555876 640198 555918 640434
rect 556154 640198 556196 640434
rect 555876 633434 556196 640198
rect 555876 633198 555918 633434
rect 556154 633198 556196 633434
rect 555876 626434 556196 633198
rect 555876 626198 555918 626434
rect 556154 626198 556196 626434
rect 555876 619434 556196 626198
rect 555876 619198 555918 619434
rect 556154 619198 556196 619434
rect 555876 612434 556196 619198
rect 555876 612198 555918 612434
rect 556154 612198 556196 612434
rect 555876 605434 556196 612198
rect 555876 605198 555918 605434
rect 556154 605198 556196 605434
rect 555876 598434 556196 605198
rect 555876 598198 555918 598434
rect 556154 598198 556196 598434
rect 555876 591434 556196 598198
rect 555876 591198 555918 591434
rect 556154 591198 556196 591434
rect 555876 584434 556196 591198
rect 555876 584198 555918 584434
rect 556154 584198 556196 584434
rect 555876 577434 556196 584198
rect 555876 577198 555918 577434
rect 556154 577198 556196 577434
rect 555876 570434 556196 577198
rect 555876 570198 555918 570434
rect 556154 570198 556196 570434
rect 555876 563434 556196 570198
rect 555876 563198 555918 563434
rect 556154 563198 556196 563434
rect 555876 556434 556196 563198
rect 555876 556198 555918 556434
rect 556154 556198 556196 556434
rect 555876 549434 556196 556198
rect 555876 549198 555918 549434
rect 556154 549198 556196 549434
rect 555876 542434 556196 549198
rect 555876 542198 555918 542434
rect 556154 542198 556196 542434
rect 555876 535434 556196 542198
rect 555876 535198 555918 535434
rect 556154 535198 556196 535434
rect 555876 528434 556196 535198
rect 555876 528198 555918 528434
rect 556154 528198 556196 528434
rect 555876 521434 556196 528198
rect 555876 521198 555918 521434
rect 556154 521198 556196 521434
rect 555876 514434 556196 521198
rect 555876 514198 555918 514434
rect 556154 514198 556196 514434
rect 555876 507434 556196 514198
rect 555876 507198 555918 507434
rect 556154 507198 556196 507434
rect 555876 500434 556196 507198
rect 555876 500198 555918 500434
rect 556154 500198 556196 500434
rect 555876 493434 556196 500198
rect 555876 493198 555918 493434
rect 556154 493198 556196 493434
rect 555876 486434 556196 493198
rect 555876 486198 555918 486434
rect 556154 486198 556196 486434
rect 555876 479434 556196 486198
rect 555876 479198 555918 479434
rect 556154 479198 556196 479434
rect 555876 472434 556196 479198
rect 555876 472198 555918 472434
rect 556154 472198 556196 472434
rect 555876 465434 556196 472198
rect 555876 465198 555918 465434
rect 556154 465198 556196 465434
rect 555876 458434 556196 465198
rect 555876 458198 555918 458434
rect 556154 458198 556196 458434
rect 555876 451434 556196 458198
rect 555876 451198 555918 451434
rect 556154 451198 556196 451434
rect 555876 444434 556196 451198
rect 555876 444198 555918 444434
rect 556154 444198 556196 444434
rect 555876 437434 556196 444198
rect 555876 437198 555918 437434
rect 556154 437198 556196 437434
rect 555876 430434 556196 437198
rect 555876 430198 555918 430434
rect 556154 430198 556196 430434
rect 555876 423434 556196 430198
rect 555876 423198 555918 423434
rect 556154 423198 556196 423434
rect 555876 416434 556196 423198
rect 555876 416198 555918 416434
rect 556154 416198 556196 416434
rect 555876 409434 556196 416198
rect 555876 409198 555918 409434
rect 556154 409198 556196 409434
rect 555876 402434 556196 409198
rect 555876 402198 555918 402434
rect 556154 402198 556196 402434
rect 555876 395434 556196 402198
rect 555876 395198 555918 395434
rect 556154 395198 556196 395434
rect 555876 388434 556196 395198
rect 555876 388198 555918 388434
rect 556154 388198 556196 388434
rect 555876 381434 556196 388198
rect 555876 381198 555918 381434
rect 556154 381198 556196 381434
rect 555876 374434 556196 381198
rect 555876 374198 555918 374434
rect 556154 374198 556196 374434
rect 555876 367434 556196 374198
rect 555876 367198 555918 367434
rect 556154 367198 556196 367434
rect 555876 360434 556196 367198
rect 555876 360198 555918 360434
rect 556154 360198 556196 360434
rect 555876 353434 556196 360198
rect 555876 353198 555918 353434
rect 556154 353198 556196 353434
rect 555876 346434 556196 353198
rect 555876 346198 555918 346434
rect 556154 346198 556196 346434
rect 555876 339434 556196 346198
rect 555876 339198 555918 339434
rect 556154 339198 556196 339434
rect 555876 332434 556196 339198
rect 555876 332198 555918 332434
rect 556154 332198 556196 332434
rect 555876 325434 556196 332198
rect 555876 325198 555918 325434
rect 556154 325198 556196 325434
rect 555876 318434 556196 325198
rect 555876 318198 555918 318434
rect 556154 318198 556196 318434
rect 555876 311434 556196 318198
rect 555876 311198 555918 311434
rect 556154 311198 556196 311434
rect 555876 304434 556196 311198
rect 555876 304198 555918 304434
rect 556154 304198 556196 304434
rect 555876 297434 556196 304198
rect 555876 297198 555918 297434
rect 556154 297198 556196 297434
rect 555876 290434 556196 297198
rect 555876 290198 555918 290434
rect 556154 290198 556196 290434
rect 555876 283434 556196 290198
rect 555876 283198 555918 283434
rect 556154 283198 556196 283434
rect 555876 276434 556196 283198
rect 555876 276198 555918 276434
rect 556154 276198 556196 276434
rect 555876 269434 556196 276198
rect 555876 269198 555918 269434
rect 556154 269198 556196 269434
rect 555876 262434 556196 269198
rect 555876 262198 555918 262434
rect 556154 262198 556196 262434
rect 555876 255434 556196 262198
rect 555876 255198 555918 255434
rect 556154 255198 556196 255434
rect 555876 248434 556196 255198
rect 555876 248198 555918 248434
rect 556154 248198 556196 248434
rect 555876 241434 556196 248198
rect 555876 241198 555918 241434
rect 556154 241198 556196 241434
rect 555876 234434 556196 241198
rect 555876 234198 555918 234434
rect 556154 234198 556196 234434
rect 555876 227434 556196 234198
rect 555876 227198 555918 227434
rect 556154 227198 556196 227434
rect 555876 220434 556196 227198
rect 555876 220198 555918 220434
rect 556154 220198 556196 220434
rect 555876 213434 556196 220198
rect 555876 213198 555918 213434
rect 556154 213198 556196 213434
rect 555876 206434 556196 213198
rect 555876 206198 555918 206434
rect 556154 206198 556196 206434
rect 555876 199434 556196 206198
rect 555876 199198 555918 199434
rect 556154 199198 556196 199434
rect 555876 192434 556196 199198
rect 555876 192198 555918 192434
rect 556154 192198 556196 192434
rect 555876 185434 556196 192198
rect 555876 185198 555918 185434
rect 556154 185198 556196 185434
rect 555876 178434 556196 185198
rect 555876 178198 555918 178434
rect 556154 178198 556196 178434
rect 555876 171434 556196 178198
rect 555876 171198 555918 171434
rect 556154 171198 556196 171434
rect 555876 164434 556196 171198
rect 555876 164198 555918 164434
rect 556154 164198 556196 164434
rect 555876 157434 556196 164198
rect 555876 157198 555918 157434
rect 556154 157198 556196 157434
rect 555876 150434 556196 157198
rect 555876 150198 555918 150434
rect 556154 150198 556196 150434
rect 555876 143434 556196 150198
rect 555876 143198 555918 143434
rect 556154 143198 556196 143434
rect 555876 136434 556196 143198
rect 555876 136198 555918 136434
rect 556154 136198 556196 136434
rect 555876 129434 556196 136198
rect 555876 129198 555918 129434
rect 556154 129198 556196 129434
rect 555876 122434 556196 129198
rect 555876 122198 555918 122434
rect 556154 122198 556196 122434
rect 555876 115434 556196 122198
rect 555876 115198 555918 115434
rect 556154 115198 556196 115434
rect 555876 108434 556196 115198
rect 555876 108198 555918 108434
rect 556154 108198 556196 108434
rect 555876 101434 556196 108198
rect 555876 101198 555918 101434
rect 556154 101198 556196 101434
rect 555876 94434 556196 101198
rect 555876 94198 555918 94434
rect 556154 94198 556196 94434
rect 555876 87434 556196 94198
rect 555876 87198 555918 87434
rect 556154 87198 556196 87434
rect 555876 80434 556196 87198
rect 555876 80198 555918 80434
rect 556154 80198 556196 80434
rect 555876 73434 556196 80198
rect 555876 73198 555918 73434
rect 556154 73198 556196 73434
rect 555876 66434 556196 73198
rect 555876 66198 555918 66434
rect 556154 66198 556196 66434
rect 555876 59434 556196 66198
rect 555876 59198 555918 59434
rect 556154 59198 556196 59434
rect 555876 52434 556196 59198
rect 555876 52198 555918 52434
rect 556154 52198 556196 52434
rect 555876 45434 556196 52198
rect 555876 45198 555918 45434
rect 556154 45198 556196 45434
rect 555876 38434 556196 45198
rect 555876 38198 555918 38434
rect 556154 38198 556196 38434
rect 555876 31434 556196 38198
rect 555876 31198 555918 31434
rect 556154 31198 556196 31434
rect 555876 24434 556196 31198
rect 555876 24198 555918 24434
rect 556154 24198 556196 24434
rect 555876 17434 556196 24198
rect 555876 17198 555918 17434
rect 556154 17198 556196 17434
rect 555876 10434 556196 17198
rect 555876 10198 555918 10434
rect 556154 10198 556196 10434
rect 555876 3434 556196 10198
rect 555876 3198 555918 3434
rect 556154 3198 556196 3434
rect 555876 -1706 556196 3198
rect 555876 -1942 555918 -1706
rect 556154 -1942 556196 -1706
rect 555876 -2026 556196 -1942
rect 555876 -2262 555918 -2026
rect 556154 -2262 556196 -2026
rect 555876 -2294 556196 -2262
rect 561144 705238 561464 706230
rect 561144 705002 561186 705238
rect 561422 705002 561464 705238
rect 561144 704918 561464 705002
rect 561144 704682 561186 704918
rect 561422 704682 561464 704918
rect 561144 695494 561464 704682
rect 561144 695258 561186 695494
rect 561422 695258 561464 695494
rect 561144 688494 561464 695258
rect 561144 688258 561186 688494
rect 561422 688258 561464 688494
rect 561144 681494 561464 688258
rect 561144 681258 561186 681494
rect 561422 681258 561464 681494
rect 561144 674494 561464 681258
rect 561144 674258 561186 674494
rect 561422 674258 561464 674494
rect 561144 667494 561464 674258
rect 561144 667258 561186 667494
rect 561422 667258 561464 667494
rect 561144 660494 561464 667258
rect 561144 660258 561186 660494
rect 561422 660258 561464 660494
rect 561144 653494 561464 660258
rect 561144 653258 561186 653494
rect 561422 653258 561464 653494
rect 561144 646494 561464 653258
rect 561144 646258 561186 646494
rect 561422 646258 561464 646494
rect 561144 639494 561464 646258
rect 561144 639258 561186 639494
rect 561422 639258 561464 639494
rect 561144 632494 561464 639258
rect 561144 632258 561186 632494
rect 561422 632258 561464 632494
rect 561144 625494 561464 632258
rect 561144 625258 561186 625494
rect 561422 625258 561464 625494
rect 561144 618494 561464 625258
rect 561144 618258 561186 618494
rect 561422 618258 561464 618494
rect 561144 611494 561464 618258
rect 561144 611258 561186 611494
rect 561422 611258 561464 611494
rect 561144 604494 561464 611258
rect 561144 604258 561186 604494
rect 561422 604258 561464 604494
rect 561144 597494 561464 604258
rect 561144 597258 561186 597494
rect 561422 597258 561464 597494
rect 561144 590494 561464 597258
rect 561144 590258 561186 590494
rect 561422 590258 561464 590494
rect 561144 583494 561464 590258
rect 561144 583258 561186 583494
rect 561422 583258 561464 583494
rect 561144 576494 561464 583258
rect 561144 576258 561186 576494
rect 561422 576258 561464 576494
rect 561144 569494 561464 576258
rect 561144 569258 561186 569494
rect 561422 569258 561464 569494
rect 561144 562494 561464 569258
rect 561144 562258 561186 562494
rect 561422 562258 561464 562494
rect 561144 555494 561464 562258
rect 561144 555258 561186 555494
rect 561422 555258 561464 555494
rect 561144 548494 561464 555258
rect 561144 548258 561186 548494
rect 561422 548258 561464 548494
rect 561144 541494 561464 548258
rect 561144 541258 561186 541494
rect 561422 541258 561464 541494
rect 561144 534494 561464 541258
rect 561144 534258 561186 534494
rect 561422 534258 561464 534494
rect 561144 527494 561464 534258
rect 561144 527258 561186 527494
rect 561422 527258 561464 527494
rect 561144 520494 561464 527258
rect 561144 520258 561186 520494
rect 561422 520258 561464 520494
rect 561144 513494 561464 520258
rect 561144 513258 561186 513494
rect 561422 513258 561464 513494
rect 561144 506494 561464 513258
rect 561144 506258 561186 506494
rect 561422 506258 561464 506494
rect 561144 499494 561464 506258
rect 561144 499258 561186 499494
rect 561422 499258 561464 499494
rect 561144 492494 561464 499258
rect 561144 492258 561186 492494
rect 561422 492258 561464 492494
rect 561144 485494 561464 492258
rect 561144 485258 561186 485494
rect 561422 485258 561464 485494
rect 561144 478494 561464 485258
rect 561144 478258 561186 478494
rect 561422 478258 561464 478494
rect 561144 471494 561464 478258
rect 561144 471258 561186 471494
rect 561422 471258 561464 471494
rect 561144 464494 561464 471258
rect 561144 464258 561186 464494
rect 561422 464258 561464 464494
rect 561144 457494 561464 464258
rect 561144 457258 561186 457494
rect 561422 457258 561464 457494
rect 561144 450494 561464 457258
rect 561144 450258 561186 450494
rect 561422 450258 561464 450494
rect 561144 443494 561464 450258
rect 561144 443258 561186 443494
rect 561422 443258 561464 443494
rect 561144 436494 561464 443258
rect 561144 436258 561186 436494
rect 561422 436258 561464 436494
rect 561144 429494 561464 436258
rect 561144 429258 561186 429494
rect 561422 429258 561464 429494
rect 561144 422494 561464 429258
rect 561144 422258 561186 422494
rect 561422 422258 561464 422494
rect 561144 415494 561464 422258
rect 561144 415258 561186 415494
rect 561422 415258 561464 415494
rect 561144 408494 561464 415258
rect 561144 408258 561186 408494
rect 561422 408258 561464 408494
rect 561144 401494 561464 408258
rect 561144 401258 561186 401494
rect 561422 401258 561464 401494
rect 561144 394494 561464 401258
rect 561144 394258 561186 394494
rect 561422 394258 561464 394494
rect 561144 387494 561464 394258
rect 561144 387258 561186 387494
rect 561422 387258 561464 387494
rect 561144 380494 561464 387258
rect 561144 380258 561186 380494
rect 561422 380258 561464 380494
rect 561144 373494 561464 380258
rect 561144 373258 561186 373494
rect 561422 373258 561464 373494
rect 561144 366494 561464 373258
rect 561144 366258 561186 366494
rect 561422 366258 561464 366494
rect 561144 359494 561464 366258
rect 561144 359258 561186 359494
rect 561422 359258 561464 359494
rect 561144 352494 561464 359258
rect 561144 352258 561186 352494
rect 561422 352258 561464 352494
rect 561144 345494 561464 352258
rect 561144 345258 561186 345494
rect 561422 345258 561464 345494
rect 561144 338494 561464 345258
rect 561144 338258 561186 338494
rect 561422 338258 561464 338494
rect 561144 331494 561464 338258
rect 561144 331258 561186 331494
rect 561422 331258 561464 331494
rect 561144 324494 561464 331258
rect 561144 324258 561186 324494
rect 561422 324258 561464 324494
rect 561144 317494 561464 324258
rect 561144 317258 561186 317494
rect 561422 317258 561464 317494
rect 561144 310494 561464 317258
rect 561144 310258 561186 310494
rect 561422 310258 561464 310494
rect 561144 303494 561464 310258
rect 561144 303258 561186 303494
rect 561422 303258 561464 303494
rect 561144 296494 561464 303258
rect 561144 296258 561186 296494
rect 561422 296258 561464 296494
rect 561144 289494 561464 296258
rect 561144 289258 561186 289494
rect 561422 289258 561464 289494
rect 561144 282494 561464 289258
rect 561144 282258 561186 282494
rect 561422 282258 561464 282494
rect 561144 275494 561464 282258
rect 561144 275258 561186 275494
rect 561422 275258 561464 275494
rect 561144 268494 561464 275258
rect 561144 268258 561186 268494
rect 561422 268258 561464 268494
rect 561144 261494 561464 268258
rect 561144 261258 561186 261494
rect 561422 261258 561464 261494
rect 561144 254494 561464 261258
rect 561144 254258 561186 254494
rect 561422 254258 561464 254494
rect 561144 247494 561464 254258
rect 561144 247258 561186 247494
rect 561422 247258 561464 247494
rect 561144 240494 561464 247258
rect 561144 240258 561186 240494
rect 561422 240258 561464 240494
rect 561144 233494 561464 240258
rect 561144 233258 561186 233494
rect 561422 233258 561464 233494
rect 561144 226494 561464 233258
rect 561144 226258 561186 226494
rect 561422 226258 561464 226494
rect 561144 219494 561464 226258
rect 561144 219258 561186 219494
rect 561422 219258 561464 219494
rect 561144 212494 561464 219258
rect 561144 212258 561186 212494
rect 561422 212258 561464 212494
rect 561144 205494 561464 212258
rect 561144 205258 561186 205494
rect 561422 205258 561464 205494
rect 561144 198494 561464 205258
rect 561144 198258 561186 198494
rect 561422 198258 561464 198494
rect 561144 191494 561464 198258
rect 561144 191258 561186 191494
rect 561422 191258 561464 191494
rect 561144 184494 561464 191258
rect 561144 184258 561186 184494
rect 561422 184258 561464 184494
rect 561144 177494 561464 184258
rect 561144 177258 561186 177494
rect 561422 177258 561464 177494
rect 561144 170494 561464 177258
rect 561144 170258 561186 170494
rect 561422 170258 561464 170494
rect 561144 163494 561464 170258
rect 561144 163258 561186 163494
rect 561422 163258 561464 163494
rect 561144 156494 561464 163258
rect 561144 156258 561186 156494
rect 561422 156258 561464 156494
rect 561144 149494 561464 156258
rect 561144 149258 561186 149494
rect 561422 149258 561464 149494
rect 561144 142494 561464 149258
rect 561144 142258 561186 142494
rect 561422 142258 561464 142494
rect 561144 135494 561464 142258
rect 561144 135258 561186 135494
rect 561422 135258 561464 135494
rect 561144 128494 561464 135258
rect 561144 128258 561186 128494
rect 561422 128258 561464 128494
rect 561144 121494 561464 128258
rect 561144 121258 561186 121494
rect 561422 121258 561464 121494
rect 561144 114494 561464 121258
rect 561144 114258 561186 114494
rect 561422 114258 561464 114494
rect 561144 107494 561464 114258
rect 561144 107258 561186 107494
rect 561422 107258 561464 107494
rect 561144 100494 561464 107258
rect 561144 100258 561186 100494
rect 561422 100258 561464 100494
rect 561144 93494 561464 100258
rect 561144 93258 561186 93494
rect 561422 93258 561464 93494
rect 561144 86494 561464 93258
rect 561144 86258 561186 86494
rect 561422 86258 561464 86494
rect 561144 79494 561464 86258
rect 561144 79258 561186 79494
rect 561422 79258 561464 79494
rect 561144 72494 561464 79258
rect 561144 72258 561186 72494
rect 561422 72258 561464 72494
rect 561144 65494 561464 72258
rect 561144 65258 561186 65494
rect 561422 65258 561464 65494
rect 561144 58494 561464 65258
rect 561144 58258 561186 58494
rect 561422 58258 561464 58494
rect 561144 51494 561464 58258
rect 561144 51258 561186 51494
rect 561422 51258 561464 51494
rect 561144 44494 561464 51258
rect 561144 44258 561186 44494
rect 561422 44258 561464 44494
rect 561144 37494 561464 44258
rect 561144 37258 561186 37494
rect 561422 37258 561464 37494
rect 561144 30494 561464 37258
rect 561144 30258 561186 30494
rect 561422 30258 561464 30494
rect 561144 23494 561464 30258
rect 561144 23258 561186 23494
rect 561422 23258 561464 23494
rect 561144 16494 561464 23258
rect 561144 16258 561186 16494
rect 561422 16258 561464 16494
rect 561144 9494 561464 16258
rect 561144 9258 561186 9494
rect 561422 9258 561464 9494
rect 561144 2494 561464 9258
rect 561144 2258 561186 2494
rect 561422 2258 561464 2494
rect 561144 -746 561464 2258
rect 561144 -982 561186 -746
rect 561422 -982 561464 -746
rect 561144 -1066 561464 -982
rect 561144 -1302 561186 -1066
rect 561422 -1302 561464 -1066
rect 561144 -2294 561464 -1302
rect 562876 706198 563196 706230
rect 562876 705962 562918 706198
rect 563154 705962 563196 706198
rect 562876 705878 563196 705962
rect 562876 705642 562918 705878
rect 563154 705642 563196 705878
rect 562876 696434 563196 705642
rect 562876 696198 562918 696434
rect 563154 696198 563196 696434
rect 562876 689434 563196 696198
rect 562876 689198 562918 689434
rect 563154 689198 563196 689434
rect 562876 682434 563196 689198
rect 562876 682198 562918 682434
rect 563154 682198 563196 682434
rect 562876 675434 563196 682198
rect 562876 675198 562918 675434
rect 563154 675198 563196 675434
rect 562876 668434 563196 675198
rect 562876 668198 562918 668434
rect 563154 668198 563196 668434
rect 562876 661434 563196 668198
rect 562876 661198 562918 661434
rect 563154 661198 563196 661434
rect 562876 654434 563196 661198
rect 562876 654198 562918 654434
rect 563154 654198 563196 654434
rect 562876 647434 563196 654198
rect 562876 647198 562918 647434
rect 563154 647198 563196 647434
rect 562876 640434 563196 647198
rect 562876 640198 562918 640434
rect 563154 640198 563196 640434
rect 562876 633434 563196 640198
rect 562876 633198 562918 633434
rect 563154 633198 563196 633434
rect 562876 626434 563196 633198
rect 562876 626198 562918 626434
rect 563154 626198 563196 626434
rect 562876 619434 563196 626198
rect 562876 619198 562918 619434
rect 563154 619198 563196 619434
rect 562876 612434 563196 619198
rect 562876 612198 562918 612434
rect 563154 612198 563196 612434
rect 562876 605434 563196 612198
rect 562876 605198 562918 605434
rect 563154 605198 563196 605434
rect 562876 598434 563196 605198
rect 562876 598198 562918 598434
rect 563154 598198 563196 598434
rect 562876 591434 563196 598198
rect 562876 591198 562918 591434
rect 563154 591198 563196 591434
rect 562876 584434 563196 591198
rect 562876 584198 562918 584434
rect 563154 584198 563196 584434
rect 562876 577434 563196 584198
rect 562876 577198 562918 577434
rect 563154 577198 563196 577434
rect 562876 570434 563196 577198
rect 562876 570198 562918 570434
rect 563154 570198 563196 570434
rect 562876 563434 563196 570198
rect 562876 563198 562918 563434
rect 563154 563198 563196 563434
rect 562876 556434 563196 563198
rect 562876 556198 562918 556434
rect 563154 556198 563196 556434
rect 562876 549434 563196 556198
rect 562876 549198 562918 549434
rect 563154 549198 563196 549434
rect 562876 542434 563196 549198
rect 562876 542198 562918 542434
rect 563154 542198 563196 542434
rect 562876 535434 563196 542198
rect 562876 535198 562918 535434
rect 563154 535198 563196 535434
rect 562876 528434 563196 535198
rect 562876 528198 562918 528434
rect 563154 528198 563196 528434
rect 562876 521434 563196 528198
rect 562876 521198 562918 521434
rect 563154 521198 563196 521434
rect 562876 514434 563196 521198
rect 562876 514198 562918 514434
rect 563154 514198 563196 514434
rect 562876 507434 563196 514198
rect 562876 507198 562918 507434
rect 563154 507198 563196 507434
rect 562876 500434 563196 507198
rect 562876 500198 562918 500434
rect 563154 500198 563196 500434
rect 562876 493434 563196 500198
rect 562876 493198 562918 493434
rect 563154 493198 563196 493434
rect 562876 486434 563196 493198
rect 562876 486198 562918 486434
rect 563154 486198 563196 486434
rect 562876 479434 563196 486198
rect 562876 479198 562918 479434
rect 563154 479198 563196 479434
rect 562876 472434 563196 479198
rect 562876 472198 562918 472434
rect 563154 472198 563196 472434
rect 562876 465434 563196 472198
rect 562876 465198 562918 465434
rect 563154 465198 563196 465434
rect 562876 458434 563196 465198
rect 562876 458198 562918 458434
rect 563154 458198 563196 458434
rect 562876 451434 563196 458198
rect 562876 451198 562918 451434
rect 563154 451198 563196 451434
rect 562876 444434 563196 451198
rect 562876 444198 562918 444434
rect 563154 444198 563196 444434
rect 562876 437434 563196 444198
rect 562876 437198 562918 437434
rect 563154 437198 563196 437434
rect 562876 430434 563196 437198
rect 562876 430198 562918 430434
rect 563154 430198 563196 430434
rect 562876 423434 563196 430198
rect 562876 423198 562918 423434
rect 563154 423198 563196 423434
rect 562876 416434 563196 423198
rect 562876 416198 562918 416434
rect 563154 416198 563196 416434
rect 562876 409434 563196 416198
rect 562876 409198 562918 409434
rect 563154 409198 563196 409434
rect 562876 402434 563196 409198
rect 562876 402198 562918 402434
rect 563154 402198 563196 402434
rect 562876 395434 563196 402198
rect 562876 395198 562918 395434
rect 563154 395198 563196 395434
rect 562876 388434 563196 395198
rect 562876 388198 562918 388434
rect 563154 388198 563196 388434
rect 562876 381434 563196 388198
rect 562876 381198 562918 381434
rect 563154 381198 563196 381434
rect 562876 374434 563196 381198
rect 562876 374198 562918 374434
rect 563154 374198 563196 374434
rect 562876 367434 563196 374198
rect 562876 367198 562918 367434
rect 563154 367198 563196 367434
rect 562876 360434 563196 367198
rect 562876 360198 562918 360434
rect 563154 360198 563196 360434
rect 562876 353434 563196 360198
rect 562876 353198 562918 353434
rect 563154 353198 563196 353434
rect 562876 346434 563196 353198
rect 562876 346198 562918 346434
rect 563154 346198 563196 346434
rect 562876 339434 563196 346198
rect 562876 339198 562918 339434
rect 563154 339198 563196 339434
rect 562876 332434 563196 339198
rect 562876 332198 562918 332434
rect 563154 332198 563196 332434
rect 562876 325434 563196 332198
rect 562876 325198 562918 325434
rect 563154 325198 563196 325434
rect 562876 318434 563196 325198
rect 562876 318198 562918 318434
rect 563154 318198 563196 318434
rect 562876 311434 563196 318198
rect 562876 311198 562918 311434
rect 563154 311198 563196 311434
rect 562876 304434 563196 311198
rect 562876 304198 562918 304434
rect 563154 304198 563196 304434
rect 562876 297434 563196 304198
rect 562876 297198 562918 297434
rect 563154 297198 563196 297434
rect 562876 290434 563196 297198
rect 562876 290198 562918 290434
rect 563154 290198 563196 290434
rect 562876 283434 563196 290198
rect 562876 283198 562918 283434
rect 563154 283198 563196 283434
rect 562876 276434 563196 283198
rect 562876 276198 562918 276434
rect 563154 276198 563196 276434
rect 562876 269434 563196 276198
rect 562876 269198 562918 269434
rect 563154 269198 563196 269434
rect 562876 262434 563196 269198
rect 562876 262198 562918 262434
rect 563154 262198 563196 262434
rect 562876 255434 563196 262198
rect 562876 255198 562918 255434
rect 563154 255198 563196 255434
rect 562876 248434 563196 255198
rect 562876 248198 562918 248434
rect 563154 248198 563196 248434
rect 562876 241434 563196 248198
rect 562876 241198 562918 241434
rect 563154 241198 563196 241434
rect 562876 234434 563196 241198
rect 562876 234198 562918 234434
rect 563154 234198 563196 234434
rect 562876 227434 563196 234198
rect 562876 227198 562918 227434
rect 563154 227198 563196 227434
rect 562876 220434 563196 227198
rect 562876 220198 562918 220434
rect 563154 220198 563196 220434
rect 562876 213434 563196 220198
rect 562876 213198 562918 213434
rect 563154 213198 563196 213434
rect 562876 206434 563196 213198
rect 562876 206198 562918 206434
rect 563154 206198 563196 206434
rect 562876 199434 563196 206198
rect 562876 199198 562918 199434
rect 563154 199198 563196 199434
rect 562876 192434 563196 199198
rect 562876 192198 562918 192434
rect 563154 192198 563196 192434
rect 562876 185434 563196 192198
rect 562876 185198 562918 185434
rect 563154 185198 563196 185434
rect 562876 178434 563196 185198
rect 562876 178198 562918 178434
rect 563154 178198 563196 178434
rect 562876 171434 563196 178198
rect 562876 171198 562918 171434
rect 563154 171198 563196 171434
rect 562876 164434 563196 171198
rect 562876 164198 562918 164434
rect 563154 164198 563196 164434
rect 562876 157434 563196 164198
rect 562876 157198 562918 157434
rect 563154 157198 563196 157434
rect 562876 150434 563196 157198
rect 562876 150198 562918 150434
rect 563154 150198 563196 150434
rect 562876 143434 563196 150198
rect 562876 143198 562918 143434
rect 563154 143198 563196 143434
rect 562876 136434 563196 143198
rect 562876 136198 562918 136434
rect 563154 136198 563196 136434
rect 562876 129434 563196 136198
rect 562876 129198 562918 129434
rect 563154 129198 563196 129434
rect 562876 122434 563196 129198
rect 562876 122198 562918 122434
rect 563154 122198 563196 122434
rect 562876 115434 563196 122198
rect 562876 115198 562918 115434
rect 563154 115198 563196 115434
rect 562876 108434 563196 115198
rect 562876 108198 562918 108434
rect 563154 108198 563196 108434
rect 562876 101434 563196 108198
rect 562876 101198 562918 101434
rect 563154 101198 563196 101434
rect 562876 94434 563196 101198
rect 562876 94198 562918 94434
rect 563154 94198 563196 94434
rect 562876 87434 563196 94198
rect 562876 87198 562918 87434
rect 563154 87198 563196 87434
rect 562876 80434 563196 87198
rect 562876 80198 562918 80434
rect 563154 80198 563196 80434
rect 562876 73434 563196 80198
rect 562876 73198 562918 73434
rect 563154 73198 563196 73434
rect 562876 66434 563196 73198
rect 562876 66198 562918 66434
rect 563154 66198 563196 66434
rect 562876 59434 563196 66198
rect 562876 59198 562918 59434
rect 563154 59198 563196 59434
rect 562876 52434 563196 59198
rect 562876 52198 562918 52434
rect 563154 52198 563196 52434
rect 562876 45434 563196 52198
rect 562876 45198 562918 45434
rect 563154 45198 563196 45434
rect 562876 38434 563196 45198
rect 562876 38198 562918 38434
rect 563154 38198 563196 38434
rect 562876 31434 563196 38198
rect 562876 31198 562918 31434
rect 563154 31198 563196 31434
rect 562876 24434 563196 31198
rect 562876 24198 562918 24434
rect 563154 24198 563196 24434
rect 562876 17434 563196 24198
rect 562876 17198 562918 17434
rect 563154 17198 563196 17434
rect 562876 10434 563196 17198
rect 562876 10198 562918 10434
rect 563154 10198 563196 10434
rect 562876 3434 563196 10198
rect 562876 3198 562918 3434
rect 563154 3198 563196 3434
rect 562876 -1706 563196 3198
rect 562876 -1942 562918 -1706
rect 563154 -1942 563196 -1706
rect 562876 -2026 563196 -1942
rect 562876 -2262 562918 -2026
rect 563154 -2262 563196 -2026
rect 562876 -2294 563196 -2262
rect 568144 705238 568464 706230
rect 568144 705002 568186 705238
rect 568422 705002 568464 705238
rect 568144 704918 568464 705002
rect 568144 704682 568186 704918
rect 568422 704682 568464 704918
rect 568144 695494 568464 704682
rect 568144 695258 568186 695494
rect 568422 695258 568464 695494
rect 568144 688494 568464 695258
rect 568144 688258 568186 688494
rect 568422 688258 568464 688494
rect 568144 681494 568464 688258
rect 568144 681258 568186 681494
rect 568422 681258 568464 681494
rect 568144 674494 568464 681258
rect 568144 674258 568186 674494
rect 568422 674258 568464 674494
rect 568144 667494 568464 674258
rect 568144 667258 568186 667494
rect 568422 667258 568464 667494
rect 568144 660494 568464 667258
rect 568144 660258 568186 660494
rect 568422 660258 568464 660494
rect 568144 653494 568464 660258
rect 568144 653258 568186 653494
rect 568422 653258 568464 653494
rect 568144 646494 568464 653258
rect 568144 646258 568186 646494
rect 568422 646258 568464 646494
rect 568144 639494 568464 646258
rect 568144 639258 568186 639494
rect 568422 639258 568464 639494
rect 568144 632494 568464 639258
rect 568144 632258 568186 632494
rect 568422 632258 568464 632494
rect 568144 625494 568464 632258
rect 568144 625258 568186 625494
rect 568422 625258 568464 625494
rect 568144 618494 568464 625258
rect 568144 618258 568186 618494
rect 568422 618258 568464 618494
rect 568144 611494 568464 618258
rect 568144 611258 568186 611494
rect 568422 611258 568464 611494
rect 568144 604494 568464 611258
rect 568144 604258 568186 604494
rect 568422 604258 568464 604494
rect 568144 597494 568464 604258
rect 568144 597258 568186 597494
rect 568422 597258 568464 597494
rect 568144 590494 568464 597258
rect 568144 590258 568186 590494
rect 568422 590258 568464 590494
rect 568144 583494 568464 590258
rect 568144 583258 568186 583494
rect 568422 583258 568464 583494
rect 568144 576494 568464 583258
rect 568144 576258 568186 576494
rect 568422 576258 568464 576494
rect 568144 569494 568464 576258
rect 568144 569258 568186 569494
rect 568422 569258 568464 569494
rect 568144 562494 568464 569258
rect 568144 562258 568186 562494
rect 568422 562258 568464 562494
rect 568144 555494 568464 562258
rect 568144 555258 568186 555494
rect 568422 555258 568464 555494
rect 568144 548494 568464 555258
rect 568144 548258 568186 548494
rect 568422 548258 568464 548494
rect 568144 541494 568464 548258
rect 568144 541258 568186 541494
rect 568422 541258 568464 541494
rect 568144 534494 568464 541258
rect 568144 534258 568186 534494
rect 568422 534258 568464 534494
rect 568144 527494 568464 534258
rect 568144 527258 568186 527494
rect 568422 527258 568464 527494
rect 568144 520494 568464 527258
rect 568144 520258 568186 520494
rect 568422 520258 568464 520494
rect 568144 513494 568464 520258
rect 568144 513258 568186 513494
rect 568422 513258 568464 513494
rect 568144 506494 568464 513258
rect 568144 506258 568186 506494
rect 568422 506258 568464 506494
rect 568144 499494 568464 506258
rect 568144 499258 568186 499494
rect 568422 499258 568464 499494
rect 568144 492494 568464 499258
rect 568144 492258 568186 492494
rect 568422 492258 568464 492494
rect 568144 485494 568464 492258
rect 568144 485258 568186 485494
rect 568422 485258 568464 485494
rect 568144 478494 568464 485258
rect 568144 478258 568186 478494
rect 568422 478258 568464 478494
rect 568144 471494 568464 478258
rect 568144 471258 568186 471494
rect 568422 471258 568464 471494
rect 568144 464494 568464 471258
rect 568144 464258 568186 464494
rect 568422 464258 568464 464494
rect 568144 457494 568464 464258
rect 568144 457258 568186 457494
rect 568422 457258 568464 457494
rect 568144 450494 568464 457258
rect 568144 450258 568186 450494
rect 568422 450258 568464 450494
rect 568144 443494 568464 450258
rect 568144 443258 568186 443494
rect 568422 443258 568464 443494
rect 568144 436494 568464 443258
rect 568144 436258 568186 436494
rect 568422 436258 568464 436494
rect 568144 429494 568464 436258
rect 568144 429258 568186 429494
rect 568422 429258 568464 429494
rect 568144 422494 568464 429258
rect 568144 422258 568186 422494
rect 568422 422258 568464 422494
rect 568144 415494 568464 422258
rect 568144 415258 568186 415494
rect 568422 415258 568464 415494
rect 568144 408494 568464 415258
rect 568144 408258 568186 408494
rect 568422 408258 568464 408494
rect 568144 401494 568464 408258
rect 568144 401258 568186 401494
rect 568422 401258 568464 401494
rect 568144 394494 568464 401258
rect 568144 394258 568186 394494
rect 568422 394258 568464 394494
rect 568144 387494 568464 394258
rect 568144 387258 568186 387494
rect 568422 387258 568464 387494
rect 568144 380494 568464 387258
rect 568144 380258 568186 380494
rect 568422 380258 568464 380494
rect 568144 373494 568464 380258
rect 568144 373258 568186 373494
rect 568422 373258 568464 373494
rect 568144 366494 568464 373258
rect 568144 366258 568186 366494
rect 568422 366258 568464 366494
rect 568144 359494 568464 366258
rect 568144 359258 568186 359494
rect 568422 359258 568464 359494
rect 568144 352494 568464 359258
rect 568144 352258 568186 352494
rect 568422 352258 568464 352494
rect 568144 345494 568464 352258
rect 568144 345258 568186 345494
rect 568422 345258 568464 345494
rect 568144 338494 568464 345258
rect 568144 338258 568186 338494
rect 568422 338258 568464 338494
rect 568144 331494 568464 338258
rect 568144 331258 568186 331494
rect 568422 331258 568464 331494
rect 568144 324494 568464 331258
rect 568144 324258 568186 324494
rect 568422 324258 568464 324494
rect 568144 317494 568464 324258
rect 568144 317258 568186 317494
rect 568422 317258 568464 317494
rect 568144 310494 568464 317258
rect 568144 310258 568186 310494
rect 568422 310258 568464 310494
rect 568144 303494 568464 310258
rect 568144 303258 568186 303494
rect 568422 303258 568464 303494
rect 568144 296494 568464 303258
rect 568144 296258 568186 296494
rect 568422 296258 568464 296494
rect 568144 289494 568464 296258
rect 568144 289258 568186 289494
rect 568422 289258 568464 289494
rect 568144 282494 568464 289258
rect 568144 282258 568186 282494
rect 568422 282258 568464 282494
rect 568144 275494 568464 282258
rect 568144 275258 568186 275494
rect 568422 275258 568464 275494
rect 568144 268494 568464 275258
rect 568144 268258 568186 268494
rect 568422 268258 568464 268494
rect 568144 261494 568464 268258
rect 568144 261258 568186 261494
rect 568422 261258 568464 261494
rect 568144 254494 568464 261258
rect 568144 254258 568186 254494
rect 568422 254258 568464 254494
rect 568144 247494 568464 254258
rect 568144 247258 568186 247494
rect 568422 247258 568464 247494
rect 568144 240494 568464 247258
rect 568144 240258 568186 240494
rect 568422 240258 568464 240494
rect 568144 233494 568464 240258
rect 568144 233258 568186 233494
rect 568422 233258 568464 233494
rect 568144 226494 568464 233258
rect 568144 226258 568186 226494
rect 568422 226258 568464 226494
rect 568144 219494 568464 226258
rect 568144 219258 568186 219494
rect 568422 219258 568464 219494
rect 568144 212494 568464 219258
rect 568144 212258 568186 212494
rect 568422 212258 568464 212494
rect 568144 205494 568464 212258
rect 568144 205258 568186 205494
rect 568422 205258 568464 205494
rect 568144 198494 568464 205258
rect 568144 198258 568186 198494
rect 568422 198258 568464 198494
rect 568144 191494 568464 198258
rect 568144 191258 568186 191494
rect 568422 191258 568464 191494
rect 568144 184494 568464 191258
rect 568144 184258 568186 184494
rect 568422 184258 568464 184494
rect 568144 177494 568464 184258
rect 568144 177258 568186 177494
rect 568422 177258 568464 177494
rect 568144 170494 568464 177258
rect 568144 170258 568186 170494
rect 568422 170258 568464 170494
rect 568144 163494 568464 170258
rect 568144 163258 568186 163494
rect 568422 163258 568464 163494
rect 568144 156494 568464 163258
rect 568144 156258 568186 156494
rect 568422 156258 568464 156494
rect 568144 149494 568464 156258
rect 568144 149258 568186 149494
rect 568422 149258 568464 149494
rect 568144 142494 568464 149258
rect 568144 142258 568186 142494
rect 568422 142258 568464 142494
rect 568144 135494 568464 142258
rect 568144 135258 568186 135494
rect 568422 135258 568464 135494
rect 568144 128494 568464 135258
rect 568144 128258 568186 128494
rect 568422 128258 568464 128494
rect 568144 121494 568464 128258
rect 568144 121258 568186 121494
rect 568422 121258 568464 121494
rect 568144 114494 568464 121258
rect 568144 114258 568186 114494
rect 568422 114258 568464 114494
rect 568144 107494 568464 114258
rect 568144 107258 568186 107494
rect 568422 107258 568464 107494
rect 568144 100494 568464 107258
rect 568144 100258 568186 100494
rect 568422 100258 568464 100494
rect 568144 93494 568464 100258
rect 568144 93258 568186 93494
rect 568422 93258 568464 93494
rect 568144 86494 568464 93258
rect 568144 86258 568186 86494
rect 568422 86258 568464 86494
rect 568144 79494 568464 86258
rect 568144 79258 568186 79494
rect 568422 79258 568464 79494
rect 568144 72494 568464 79258
rect 568144 72258 568186 72494
rect 568422 72258 568464 72494
rect 568144 65494 568464 72258
rect 568144 65258 568186 65494
rect 568422 65258 568464 65494
rect 568144 58494 568464 65258
rect 568144 58258 568186 58494
rect 568422 58258 568464 58494
rect 568144 51494 568464 58258
rect 568144 51258 568186 51494
rect 568422 51258 568464 51494
rect 568144 44494 568464 51258
rect 568144 44258 568186 44494
rect 568422 44258 568464 44494
rect 568144 37494 568464 44258
rect 568144 37258 568186 37494
rect 568422 37258 568464 37494
rect 568144 30494 568464 37258
rect 568144 30258 568186 30494
rect 568422 30258 568464 30494
rect 568144 23494 568464 30258
rect 568144 23258 568186 23494
rect 568422 23258 568464 23494
rect 568144 16494 568464 23258
rect 568144 16258 568186 16494
rect 568422 16258 568464 16494
rect 568144 9494 568464 16258
rect 568144 9258 568186 9494
rect 568422 9258 568464 9494
rect 568144 2494 568464 9258
rect 568144 2258 568186 2494
rect 568422 2258 568464 2494
rect 568144 -746 568464 2258
rect 568144 -982 568186 -746
rect 568422 -982 568464 -746
rect 568144 -1066 568464 -982
rect 568144 -1302 568186 -1066
rect 568422 -1302 568464 -1066
rect 568144 -2294 568464 -1302
rect 569876 706198 570196 706230
rect 569876 705962 569918 706198
rect 570154 705962 570196 706198
rect 569876 705878 570196 705962
rect 569876 705642 569918 705878
rect 570154 705642 570196 705878
rect 569876 696434 570196 705642
rect 569876 696198 569918 696434
rect 570154 696198 570196 696434
rect 569876 689434 570196 696198
rect 569876 689198 569918 689434
rect 570154 689198 570196 689434
rect 569876 682434 570196 689198
rect 569876 682198 569918 682434
rect 570154 682198 570196 682434
rect 569876 675434 570196 682198
rect 569876 675198 569918 675434
rect 570154 675198 570196 675434
rect 569876 668434 570196 675198
rect 569876 668198 569918 668434
rect 570154 668198 570196 668434
rect 569876 661434 570196 668198
rect 569876 661198 569918 661434
rect 570154 661198 570196 661434
rect 569876 654434 570196 661198
rect 569876 654198 569918 654434
rect 570154 654198 570196 654434
rect 569876 647434 570196 654198
rect 569876 647198 569918 647434
rect 570154 647198 570196 647434
rect 569876 640434 570196 647198
rect 569876 640198 569918 640434
rect 570154 640198 570196 640434
rect 569876 633434 570196 640198
rect 569876 633198 569918 633434
rect 570154 633198 570196 633434
rect 569876 626434 570196 633198
rect 569876 626198 569918 626434
rect 570154 626198 570196 626434
rect 569876 619434 570196 626198
rect 569876 619198 569918 619434
rect 570154 619198 570196 619434
rect 569876 612434 570196 619198
rect 569876 612198 569918 612434
rect 570154 612198 570196 612434
rect 569876 605434 570196 612198
rect 569876 605198 569918 605434
rect 570154 605198 570196 605434
rect 569876 598434 570196 605198
rect 569876 598198 569918 598434
rect 570154 598198 570196 598434
rect 569876 591434 570196 598198
rect 569876 591198 569918 591434
rect 570154 591198 570196 591434
rect 569876 584434 570196 591198
rect 569876 584198 569918 584434
rect 570154 584198 570196 584434
rect 569876 577434 570196 584198
rect 569876 577198 569918 577434
rect 570154 577198 570196 577434
rect 569876 570434 570196 577198
rect 569876 570198 569918 570434
rect 570154 570198 570196 570434
rect 569876 563434 570196 570198
rect 569876 563198 569918 563434
rect 570154 563198 570196 563434
rect 569876 556434 570196 563198
rect 569876 556198 569918 556434
rect 570154 556198 570196 556434
rect 569876 549434 570196 556198
rect 569876 549198 569918 549434
rect 570154 549198 570196 549434
rect 569876 542434 570196 549198
rect 569876 542198 569918 542434
rect 570154 542198 570196 542434
rect 569876 535434 570196 542198
rect 569876 535198 569918 535434
rect 570154 535198 570196 535434
rect 569876 528434 570196 535198
rect 569876 528198 569918 528434
rect 570154 528198 570196 528434
rect 569876 521434 570196 528198
rect 569876 521198 569918 521434
rect 570154 521198 570196 521434
rect 569876 514434 570196 521198
rect 569876 514198 569918 514434
rect 570154 514198 570196 514434
rect 569876 507434 570196 514198
rect 569876 507198 569918 507434
rect 570154 507198 570196 507434
rect 569876 500434 570196 507198
rect 569876 500198 569918 500434
rect 570154 500198 570196 500434
rect 569876 493434 570196 500198
rect 569876 493198 569918 493434
rect 570154 493198 570196 493434
rect 569876 486434 570196 493198
rect 569876 486198 569918 486434
rect 570154 486198 570196 486434
rect 569876 479434 570196 486198
rect 569876 479198 569918 479434
rect 570154 479198 570196 479434
rect 569876 472434 570196 479198
rect 569876 472198 569918 472434
rect 570154 472198 570196 472434
rect 569876 465434 570196 472198
rect 569876 465198 569918 465434
rect 570154 465198 570196 465434
rect 569876 458434 570196 465198
rect 569876 458198 569918 458434
rect 570154 458198 570196 458434
rect 569876 451434 570196 458198
rect 569876 451198 569918 451434
rect 570154 451198 570196 451434
rect 569876 444434 570196 451198
rect 569876 444198 569918 444434
rect 570154 444198 570196 444434
rect 569876 437434 570196 444198
rect 569876 437198 569918 437434
rect 570154 437198 570196 437434
rect 569876 430434 570196 437198
rect 569876 430198 569918 430434
rect 570154 430198 570196 430434
rect 569876 423434 570196 430198
rect 569876 423198 569918 423434
rect 570154 423198 570196 423434
rect 569876 416434 570196 423198
rect 569876 416198 569918 416434
rect 570154 416198 570196 416434
rect 569876 409434 570196 416198
rect 569876 409198 569918 409434
rect 570154 409198 570196 409434
rect 569876 402434 570196 409198
rect 569876 402198 569918 402434
rect 570154 402198 570196 402434
rect 569876 395434 570196 402198
rect 569876 395198 569918 395434
rect 570154 395198 570196 395434
rect 569876 388434 570196 395198
rect 569876 388198 569918 388434
rect 570154 388198 570196 388434
rect 569876 381434 570196 388198
rect 569876 381198 569918 381434
rect 570154 381198 570196 381434
rect 569876 374434 570196 381198
rect 569876 374198 569918 374434
rect 570154 374198 570196 374434
rect 569876 367434 570196 374198
rect 569876 367198 569918 367434
rect 570154 367198 570196 367434
rect 569876 360434 570196 367198
rect 569876 360198 569918 360434
rect 570154 360198 570196 360434
rect 569876 353434 570196 360198
rect 569876 353198 569918 353434
rect 570154 353198 570196 353434
rect 569876 346434 570196 353198
rect 569876 346198 569918 346434
rect 570154 346198 570196 346434
rect 569876 339434 570196 346198
rect 569876 339198 569918 339434
rect 570154 339198 570196 339434
rect 569876 332434 570196 339198
rect 569876 332198 569918 332434
rect 570154 332198 570196 332434
rect 569876 325434 570196 332198
rect 569876 325198 569918 325434
rect 570154 325198 570196 325434
rect 569876 318434 570196 325198
rect 569876 318198 569918 318434
rect 570154 318198 570196 318434
rect 569876 311434 570196 318198
rect 569876 311198 569918 311434
rect 570154 311198 570196 311434
rect 569876 304434 570196 311198
rect 569876 304198 569918 304434
rect 570154 304198 570196 304434
rect 569876 297434 570196 304198
rect 569876 297198 569918 297434
rect 570154 297198 570196 297434
rect 569876 290434 570196 297198
rect 569876 290198 569918 290434
rect 570154 290198 570196 290434
rect 569876 283434 570196 290198
rect 569876 283198 569918 283434
rect 570154 283198 570196 283434
rect 569876 276434 570196 283198
rect 569876 276198 569918 276434
rect 570154 276198 570196 276434
rect 569876 269434 570196 276198
rect 569876 269198 569918 269434
rect 570154 269198 570196 269434
rect 569876 262434 570196 269198
rect 569876 262198 569918 262434
rect 570154 262198 570196 262434
rect 569876 255434 570196 262198
rect 569876 255198 569918 255434
rect 570154 255198 570196 255434
rect 569876 248434 570196 255198
rect 569876 248198 569918 248434
rect 570154 248198 570196 248434
rect 569876 241434 570196 248198
rect 569876 241198 569918 241434
rect 570154 241198 570196 241434
rect 569876 234434 570196 241198
rect 569876 234198 569918 234434
rect 570154 234198 570196 234434
rect 569876 227434 570196 234198
rect 569876 227198 569918 227434
rect 570154 227198 570196 227434
rect 569876 220434 570196 227198
rect 569876 220198 569918 220434
rect 570154 220198 570196 220434
rect 569876 213434 570196 220198
rect 569876 213198 569918 213434
rect 570154 213198 570196 213434
rect 569876 206434 570196 213198
rect 569876 206198 569918 206434
rect 570154 206198 570196 206434
rect 569876 199434 570196 206198
rect 569876 199198 569918 199434
rect 570154 199198 570196 199434
rect 569876 192434 570196 199198
rect 569876 192198 569918 192434
rect 570154 192198 570196 192434
rect 569876 185434 570196 192198
rect 569876 185198 569918 185434
rect 570154 185198 570196 185434
rect 569876 178434 570196 185198
rect 569876 178198 569918 178434
rect 570154 178198 570196 178434
rect 569876 171434 570196 178198
rect 569876 171198 569918 171434
rect 570154 171198 570196 171434
rect 569876 164434 570196 171198
rect 569876 164198 569918 164434
rect 570154 164198 570196 164434
rect 569876 157434 570196 164198
rect 569876 157198 569918 157434
rect 570154 157198 570196 157434
rect 569876 150434 570196 157198
rect 569876 150198 569918 150434
rect 570154 150198 570196 150434
rect 569876 143434 570196 150198
rect 569876 143198 569918 143434
rect 570154 143198 570196 143434
rect 569876 136434 570196 143198
rect 569876 136198 569918 136434
rect 570154 136198 570196 136434
rect 569876 129434 570196 136198
rect 569876 129198 569918 129434
rect 570154 129198 570196 129434
rect 569876 122434 570196 129198
rect 569876 122198 569918 122434
rect 570154 122198 570196 122434
rect 569876 115434 570196 122198
rect 569876 115198 569918 115434
rect 570154 115198 570196 115434
rect 569876 108434 570196 115198
rect 569876 108198 569918 108434
rect 570154 108198 570196 108434
rect 569876 101434 570196 108198
rect 569876 101198 569918 101434
rect 570154 101198 570196 101434
rect 569876 94434 570196 101198
rect 569876 94198 569918 94434
rect 570154 94198 570196 94434
rect 569876 87434 570196 94198
rect 569876 87198 569918 87434
rect 570154 87198 570196 87434
rect 569876 80434 570196 87198
rect 569876 80198 569918 80434
rect 570154 80198 570196 80434
rect 569876 73434 570196 80198
rect 569876 73198 569918 73434
rect 570154 73198 570196 73434
rect 569876 66434 570196 73198
rect 569876 66198 569918 66434
rect 570154 66198 570196 66434
rect 569876 59434 570196 66198
rect 569876 59198 569918 59434
rect 570154 59198 570196 59434
rect 569876 52434 570196 59198
rect 569876 52198 569918 52434
rect 570154 52198 570196 52434
rect 569876 45434 570196 52198
rect 569876 45198 569918 45434
rect 570154 45198 570196 45434
rect 569876 38434 570196 45198
rect 569876 38198 569918 38434
rect 570154 38198 570196 38434
rect 569876 31434 570196 38198
rect 569876 31198 569918 31434
rect 570154 31198 570196 31434
rect 569876 24434 570196 31198
rect 569876 24198 569918 24434
rect 570154 24198 570196 24434
rect 569876 17434 570196 24198
rect 569876 17198 569918 17434
rect 570154 17198 570196 17434
rect 569876 10434 570196 17198
rect 569876 10198 569918 10434
rect 570154 10198 570196 10434
rect 569876 3434 570196 10198
rect 569876 3198 569918 3434
rect 570154 3198 570196 3434
rect 569876 -1706 570196 3198
rect 569876 -1942 569918 -1706
rect 570154 -1942 570196 -1706
rect 569876 -2026 570196 -1942
rect 569876 -2262 569918 -2026
rect 570154 -2262 570196 -2026
rect 569876 -2294 570196 -2262
rect 575144 705238 575464 706230
rect 575144 705002 575186 705238
rect 575422 705002 575464 705238
rect 575144 704918 575464 705002
rect 575144 704682 575186 704918
rect 575422 704682 575464 704918
rect 575144 695494 575464 704682
rect 575144 695258 575186 695494
rect 575422 695258 575464 695494
rect 575144 688494 575464 695258
rect 575144 688258 575186 688494
rect 575422 688258 575464 688494
rect 575144 681494 575464 688258
rect 575144 681258 575186 681494
rect 575422 681258 575464 681494
rect 575144 674494 575464 681258
rect 575144 674258 575186 674494
rect 575422 674258 575464 674494
rect 575144 667494 575464 674258
rect 575144 667258 575186 667494
rect 575422 667258 575464 667494
rect 575144 660494 575464 667258
rect 575144 660258 575186 660494
rect 575422 660258 575464 660494
rect 575144 653494 575464 660258
rect 575144 653258 575186 653494
rect 575422 653258 575464 653494
rect 575144 646494 575464 653258
rect 575144 646258 575186 646494
rect 575422 646258 575464 646494
rect 575144 639494 575464 646258
rect 575144 639258 575186 639494
rect 575422 639258 575464 639494
rect 575144 632494 575464 639258
rect 575144 632258 575186 632494
rect 575422 632258 575464 632494
rect 575144 625494 575464 632258
rect 575144 625258 575186 625494
rect 575422 625258 575464 625494
rect 575144 618494 575464 625258
rect 575144 618258 575186 618494
rect 575422 618258 575464 618494
rect 575144 611494 575464 618258
rect 575144 611258 575186 611494
rect 575422 611258 575464 611494
rect 575144 604494 575464 611258
rect 575144 604258 575186 604494
rect 575422 604258 575464 604494
rect 575144 597494 575464 604258
rect 575144 597258 575186 597494
rect 575422 597258 575464 597494
rect 575144 590494 575464 597258
rect 575144 590258 575186 590494
rect 575422 590258 575464 590494
rect 575144 583494 575464 590258
rect 575144 583258 575186 583494
rect 575422 583258 575464 583494
rect 575144 576494 575464 583258
rect 575144 576258 575186 576494
rect 575422 576258 575464 576494
rect 575144 569494 575464 576258
rect 575144 569258 575186 569494
rect 575422 569258 575464 569494
rect 575144 562494 575464 569258
rect 575144 562258 575186 562494
rect 575422 562258 575464 562494
rect 575144 555494 575464 562258
rect 575144 555258 575186 555494
rect 575422 555258 575464 555494
rect 575144 548494 575464 555258
rect 575144 548258 575186 548494
rect 575422 548258 575464 548494
rect 575144 541494 575464 548258
rect 575144 541258 575186 541494
rect 575422 541258 575464 541494
rect 575144 534494 575464 541258
rect 575144 534258 575186 534494
rect 575422 534258 575464 534494
rect 575144 527494 575464 534258
rect 575144 527258 575186 527494
rect 575422 527258 575464 527494
rect 575144 520494 575464 527258
rect 575144 520258 575186 520494
rect 575422 520258 575464 520494
rect 575144 513494 575464 520258
rect 575144 513258 575186 513494
rect 575422 513258 575464 513494
rect 575144 506494 575464 513258
rect 575144 506258 575186 506494
rect 575422 506258 575464 506494
rect 575144 499494 575464 506258
rect 575144 499258 575186 499494
rect 575422 499258 575464 499494
rect 575144 492494 575464 499258
rect 575144 492258 575186 492494
rect 575422 492258 575464 492494
rect 575144 485494 575464 492258
rect 575144 485258 575186 485494
rect 575422 485258 575464 485494
rect 575144 478494 575464 485258
rect 575144 478258 575186 478494
rect 575422 478258 575464 478494
rect 575144 471494 575464 478258
rect 575144 471258 575186 471494
rect 575422 471258 575464 471494
rect 575144 464494 575464 471258
rect 575144 464258 575186 464494
rect 575422 464258 575464 464494
rect 575144 457494 575464 464258
rect 575144 457258 575186 457494
rect 575422 457258 575464 457494
rect 575144 450494 575464 457258
rect 575144 450258 575186 450494
rect 575422 450258 575464 450494
rect 575144 443494 575464 450258
rect 575144 443258 575186 443494
rect 575422 443258 575464 443494
rect 575144 436494 575464 443258
rect 575144 436258 575186 436494
rect 575422 436258 575464 436494
rect 575144 429494 575464 436258
rect 575144 429258 575186 429494
rect 575422 429258 575464 429494
rect 575144 422494 575464 429258
rect 575144 422258 575186 422494
rect 575422 422258 575464 422494
rect 575144 415494 575464 422258
rect 575144 415258 575186 415494
rect 575422 415258 575464 415494
rect 575144 408494 575464 415258
rect 575144 408258 575186 408494
rect 575422 408258 575464 408494
rect 575144 401494 575464 408258
rect 575144 401258 575186 401494
rect 575422 401258 575464 401494
rect 575144 394494 575464 401258
rect 575144 394258 575186 394494
rect 575422 394258 575464 394494
rect 575144 387494 575464 394258
rect 575144 387258 575186 387494
rect 575422 387258 575464 387494
rect 575144 380494 575464 387258
rect 575144 380258 575186 380494
rect 575422 380258 575464 380494
rect 575144 373494 575464 380258
rect 575144 373258 575186 373494
rect 575422 373258 575464 373494
rect 575144 366494 575464 373258
rect 575144 366258 575186 366494
rect 575422 366258 575464 366494
rect 575144 359494 575464 366258
rect 575144 359258 575186 359494
rect 575422 359258 575464 359494
rect 575144 352494 575464 359258
rect 575144 352258 575186 352494
rect 575422 352258 575464 352494
rect 575144 345494 575464 352258
rect 575144 345258 575186 345494
rect 575422 345258 575464 345494
rect 575144 338494 575464 345258
rect 575144 338258 575186 338494
rect 575422 338258 575464 338494
rect 575144 331494 575464 338258
rect 575144 331258 575186 331494
rect 575422 331258 575464 331494
rect 575144 324494 575464 331258
rect 575144 324258 575186 324494
rect 575422 324258 575464 324494
rect 575144 317494 575464 324258
rect 575144 317258 575186 317494
rect 575422 317258 575464 317494
rect 575144 310494 575464 317258
rect 575144 310258 575186 310494
rect 575422 310258 575464 310494
rect 575144 303494 575464 310258
rect 575144 303258 575186 303494
rect 575422 303258 575464 303494
rect 575144 296494 575464 303258
rect 575144 296258 575186 296494
rect 575422 296258 575464 296494
rect 575144 289494 575464 296258
rect 575144 289258 575186 289494
rect 575422 289258 575464 289494
rect 575144 282494 575464 289258
rect 575144 282258 575186 282494
rect 575422 282258 575464 282494
rect 575144 275494 575464 282258
rect 575144 275258 575186 275494
rect 575422 275258 575464 275494
rect 575144 268494 575464 275258
rect 575144 268258 575186 268494
rect 575422 268258 575464 268494
rect 575144 261494 575464 268258
rect 575144 261258 575186 261494
rect 575422 261258 575464 261494
rect 575144 254494 575464 261258
rect 575144 254258 575186 254494
rect 575422 254258 575464 254494
rect 575144 247494 575464 254258
rect 575144 247258 575186 247494
rect 575422 247258 575464 247494
rect 575144 240494 575464 247258
rect 575144 240258 575186 240494
rect 575422 240258 575464 240494
rect 575144 233494 575464 240258
rect 575144 233258 575186 233494
rect 575422 233258 575464 233494
rect 575144 226494 575464 233258
rect 575144 226258 575186 226494
rect 575422 226258 575464 226494
rect 575144 219494 575464 226258
rect 575144 219258 575186 219494
rect 575422 219258 575464 219494
rect 575144 212494 575464 219258
rect 575144 212258 575186 212494
rect 575422 212258 575464 212494
rect 575144 205494 575464 212258
rect 575144 205258 575186 205494
rect 575422 205258 575464 205494
rect 575144 198494 575464 205258
rect 575144 198258 575186 198494
rect 575422 198258 575464 198494
rect 575144 191494 575464 198258
rect 575144 191258 575186 191494
rect 575422 191258 575464 191494
rect 575144 184494 575464 191258
rect 575144 184258 575186 184494
rect 575422 184258 575464 184494
rect 575144 177494 575464 184258
rect 575144 177258 575186 177494
rect 575422 177258 575464 177494
rect 575144 170494 575464 177258
rect 575144 170258 575186 170494
rect 575422 170258 575464 170494
rect 575144 163494 575464 170258
rect 575144 163258 575186 163494
rect 575422 163258 575464 163494
rect 575144 156494 575464 163258
rect 575144 156258 575186 156494
rect 575422 156258 575464 156494
rect 575144 149494 575464 156258
rect 575144 149258 575186 149494
rect 575422 149258 575464 149494
rect 575144 142494 575464 149258
rect 575144 142258 575186 142494
rect 575422 142258 575464 142494
rect 575144 135494 575464 142258
rect 575144 135258 575186 135494
rect 575422 135258 575464 135494
rect 575144 128494 575464 135258
rect 575144 128258 575186 128494
rect 575422 128258 575464 128494
rect 575144 121494 575464 128258
rect 575144 121258 575186 121494
rect 575422 121258 575464 121494
rect 575144 114494 575464 121258
rect 575144 114258 575186 114494
rect 575422 114258 575464 114494
rect 575144 107494 575464 114258
rect 575144 107258 575186 107494
rect 575422 107258 575464 107494
rect 575144 100494 575464 107258
rect 575144 100258 575186 100494
rect 575422 100258 575464 100494
rect 575144 93494 575464 100258
rect 575144 93258 575186 93494
rect 575422 93258 575464 93494
rect 575144 86494 575464 93258
rect 575144 86258 575186 86494
rect 575422 86258 575464 86494
rect 575144 79494 575464 86258
rect 575144 79258 575186 79494
rect 575422 79258 575464 79494
rect 575144 72494 575464 79258
rect 575144 72258 575186 72494
rect 575422 72258 575464 72494
rect 575144 65494 575464 72258
rect 575144 65258 575186 65494
rect 575422 65258 575464 65494
rect 575144 58494 575464 65258
rect 575144 58258 575186 58494
rect 575422 58258 575464 58494
rect 575144 51494 575464 58258
rect 575144 51258 575186 51494
rect 575422 51258 575464 51494
rect 575144 44494 575464 51258
rect 575144 44258 575186 44494
rect 575422 44258 575464 44494
rect 575144 37494 575464 44258
rect 575144 37258 575186 37494
rect 575422 37258 575464 37494
rect 575144 30494 575464 37258
rect 575144 30258 575186 30494
rect 575422 30258 575464 30494
rect 575144 23494 575464 30258
rect 575144 23258 575186 23494
rect 575422 23258 575464 23494
rect 575144 16494 575464 23258
rect 575144 16258 575186 16494
rect 575422 16258 575464 16494
rect 575144 9494 575464 16258
rect 575144 9258 575186 9494
rect 575422 9258 575464 9494
rect 575144 2494 575464 9258
rect 575144 2258 575186 2494
rect 575422 2258 575464 2494
rect 575144 -746 575464 2258
rect 575144 -982 575186 -746
rect 575422 -982 575464 -746
rect 575144 -1066 575464 -982
rect 575144 -1302 575186 -1066
rect 575422 -1302 575464 -1066
rect 575144 -2294 575464 -1302
rect 576876 706198 577196 706230
rect 576876 705962 576918 706198
rect 577154 705962 577196 706198
rect 576876 705878 577196 705962
rect 576876 705642 576918 705878
rect 577154 705642 577196 705878
rect 576876 696434 577196 705642
rect 576876 696198 576918 696434
rect 577154 696198 577196 696434
rect 576876 689434 577196 696198
rect 576876 689198 576918 689434
rect 577154 689198 577196 689434
rect 576876 682434 577196 689198
rect 576876 682198 576918 682434
rect 577154 682198 577196 682434
rect 576876 675434 577196 682198
rect 576876 675198 576918 675434
rect 577154 675198 577196 675434
rect 576876 668434 577196 675198
rect 576876 668198 576918 668434
rect 577154 668198 577196 668434
rect 576876 661434 577196 668198
rect 576876 661198 576918 661434
rect 577154 661198 577196 661434
rect 576876 654434 577196 661198
rect 576876 654198 576918 654434
rect 577154 654198 577196 654434
rect 576876 647434 577196 654198
rect 576876 647198 576918 647434
rect 577154 647198 577196 647434
rect 576876 640434 577196 647198
rect 576876 640198 576918 640434
rect 577154 640198 577196 640434
rect 576876 633434 577196 640198
rect 576876 633198 576918 633434
rect 577154 633198 577196 633434
rect 576876 626434 577196 633198
rect 576876 626198 576918 626434
rect 577154 626198 577196 626434
rect 576876 619434 577196 626198
rect 576876 619198 576918 619434
rect 577154 619198 577196 619434
rect 576876 612434 577196 619198
rect 576876 612198 576918 612434
rect 577154 612198 577196 612434
rect 576876 605434 577196 612198
rect 576876 605198 576918 605434
rect 577154 605198 577196 605434
rect 576876 598434 577196 605198
rect 576876 598198 576918 598434
rect 577154 598198 577196 598434
rect 576876 591434 577196 598198
rect 576876 591198 576918 591434
rect 577154 591198 577196 591434
rect 576876 584434 577196 591198
rect 576876 584198 576918 584434
rect 577154 584198 577196 584434
rect 576876 577434 577196 584198
rect 576876 577198 576918 577434
rect 577154 577198 577196 577434
rect 576876 570434 577196 577198
rect 576876 570198 576918 570434
rect 577154 570198 577196 570434
rect 576876 563434 577196 570198
rect 576876 563198 576918 563434
rect 577154 563198 577196 563434
rect 576876 556434 577196 563198
rect 576876 556198 576918 556434
rect 577154 556198 577196 556434
rect 576876 549434 577196 556198
rect 576876 549198 576918 549434
rect 577154 549198 577196 549434
rect 576876 542434 577196 549198
rect 576876 542198 576918 542434
rect 577154 542198 577196 542434
rect 576876 535434 577196 542198
rect 576876 535198 576918 535434
rect 577154 535198 577196 535434
rect 576876 528434 577196 535198
rect 576876 528198 576918 528434
rect 577154 528198 577196 528434
rect 576876 521434 577196 528198
rect 576876 521198 576918 521434
rect 577154 521198 577196 521434
rect 576876 514434 577196 521198
rect 576876 514198 576918 514434
rect 577154 514198 577196 514434
rect 576876 507434 577196 514198
rect 576876 507198 576918 507434
rect 577154 507198 577196 507434
rect 576876 500434 577196 507198
rect 576876 500198 576918 500434
rect 577154 500198 577196 500434
rect 576876 493434 577196 500198
rect 576876 493198 576918 493434
rect 577154 493198 577196 493434
rect 576876 486434 577196 493198
rect 576876 486198 576918 486434
rect 577154 486198 577196 486434
rect 576876 479434 577196 486198
rect 576876 479198 576918 479434
rect 577154 479198 577196 479434
rect 576876 472434 577196 479198
rect 576876 472198 576918 472434
rect 577154 472198 577196 472434
rect 576876 465434 577196 472198
rect 576876 465198 576918 465434
rect 577154 465198 577196 465434
rect 576876 458434 577196 465198
rect 576876 458198 576918 458434
rect 577154 458198 577196 458434
rect 576876 451434 577196 458198
rect 576876 451198 576918 451434
rect 577154 451198 577196 451434
rect 576876 444434 577196 451198
rect 576876 444198 576918 444434
rect 577154 444198 577196 444434
rect 576876 437434 577196 444198
rect 576876 437198 576918 437434
rect 577154 437198 577196 437434
rect 576876 430434 577196 437198
rect 576876 430198 576918 430434
rect 577154 430198 577196 430434
rect 576876 423434 577196 430198
rect 576876 423198 576918 423434
rect 577154 423198 577196 423434
rect 576876 416434 577196 423198
rect 576876 416198 576918 416434
rect 577154 416198 577196 416434
rect 576876 409434 577196 416198
rect 576876 409198 576918 409434
rect 577154 409198 577196 409434
rect 576876 402434 577196 409198
rect 576876 402198 576918 402434
rect 577154 402198 577196 402434
rect 576876 395434 577196 402198
rect 576876 395198 576918 395434
rect 577154 395198 577196 395434
rect 576876 388434 577196 395198
rect 576876 388198 576918 388434
rect 577154 388198 577196 388434
rect 576876 381434 577196 388198
rect 576876 381198 576918 381434
rect 577154 381198 577196 381434
rect 576876 374434 577196 381198
rect 576876 374198 576918 374434
rect 577154 374198 577196 374434
rect 576876 367434 577196 374198
rect 576876 367198 576918 367434
rect 577154 367198 577196 367434
rect 576876 360434 577196 367198
rect 576876 360198 576918 360434
rect 577154 360198 577196 360434
rect 576876 353434 577196 360198
rect 576876 353198 576918 353434
rect 577154 353198 577196 353434
rect 576876 346434 577196 353198
rect 576876 346198 576918 346434
rect 577154 346198 577196 346434
rect 576876 339434 577196 346198
rect 576876 339198 576918 339434
rect 577154 339198 577196 339434
rect 576876 332434 577196 339198
rect 576876 332198 576918 332434
rect 577154 332198 577196 332434
rect 576876 325434 577196 332198
rect 576876 325198 576918 325434
rect 577154 325198 577196 325434
rect 576876 318434 577196 325198
rect 576876 318198 576918 318434
rect 577154 318198 577196 318434
rect 576876 311434 577196 318198
rect 576876 311198 576918 311434
rect 577154 311198 577196 311434
rect 576876 304434 577196 311198
rect 576876 304198 576918 304434
rect 577154 304198 577196 304434
rect 576876 297434 577196 304198
rect 576876 297198 576918 297434
rect 577154 297198 577196 297434
rect 576876 290434 577196 297198
rect 576876 290198 576918 290434
rect 577154 290198 577196 290434
rect 576876 283434 577196 290198
rect 576876 283198 576918 283434
rect 577154 283198 577196 283434
rect 576876 276434 577196 283198
rect 576876 276198 576918 276434
rect 577154 276198 577196 276434
rect 576876 269434 577196 276198
rect 576876 269198 576918 269434
rect 577154 269198 577196 269434
rect 576876 262434 577196 269198
rect 576876 262198 576918 262434
rect 577154 262198 577196 262434
rect 576876 255434 577196 262198
rect 576876 255198 576918 255434
rect 577154 255198 577196 255434
rect 576876 248434 577196 255198
rect 576876 248198 576918 248434
rect 577154 248198 577196 248434
rect 576876 241434 577196 248198
rect 576876 241198 576918 241434
rect 577154 241198 577196 241434
rect 576876 234434 577196 241198
rect 576876 234198 576918 234434
rect 577154 234198 577196 234434
rect 576876 227434 577196 234198
rect 576876 227198 576918 227434
rect 577154 227198 577196 227434
rect 576876 220434 577196 227198
rect 576876 220198 576918 220434
rect 577154 220198 577196 220434
rect 576876 213434 577196 220198
rect 576876 213198 576918 213434
rect 577154 213198 577196 213434
rect 576876 206434 577196 213198
rect 576876 206198 576918 206434
rect 577154 206198 577196 206434
rect 576876 199434 577196 206198
rect 576876 199198 576918 199434
rect 577154 199198 577196 199434
rect 576876 192434 577196 199198
rect 576876 192198 576918 192434
rect 577154 192198 577196 192434
rect 576876 185434 577196 192198
rect 576876 185198 576918 185434
rect 577154 185198 577196 185434
rect 576876 178434 577196 185198
rect 576876 178198 576918 178434
rect 577154 178198 577196 178434
rect 576876 171434 577196 178198
rect 576876 171198 576918 171434
rect 577154 171198 577196 171434
rect 576876 164434 577196 171198
rect 576876 164198 576918 164434
rect 577154 164198 577196 164434
rect 576876 157434 577196 164198
rect 576876 157198 576918 157434
rect 577154 157198 577196 157434
rect 576876 150434 577196 157198
rect 576876 150198 576918 150434
rect 577154 150198 577196 150434
rect 576876 143434 577196 150198
rect 576876 143198 576918 143434
rect 577154 143198 577196 143434
rect 576876 136434 577196 143198
rect 576876 136198 576918 136434
rect 577154 136198 577196 136434
rect 576876 129434 577196 136198
rect 576876 129198 576918 129434
rect 577154 129198 577196 129434
rect 576876 122434 577196 129198
rect 576876 122198 576918 122434
rect 577154 122198 577196 122434
rect 576876 115434 577196 122198
rect 576876 115198 576918 115434
rect 577154 115198 577196 115434
rect 576876 108434 577196 115198
rect 576876 108198 576918 108434
rect 577154 108198 577196 108434
rect 576876 101434 577196 108198
rect 576876 101198 576918 101434
rect 577154 101198 577196 101434
rect 576876 94434 577196 101198
rect 576876 94198 576918 94434
rect 577154 94198 577196 94434
rect 576876 87434 577196 94198
rect 576876 87198 576918 87434
rect 577154 87198 577196 87434
rect 576876 80434 577196 87198
rect 576876 80198 576918 80434
rect 577154 80198 577196 80434
rect 576876 73434 577196 80198
rect 576876 73198 576918 73434
rect 577154 73198 577196 73434
rect 576876 66434 577196 73198
rect 576876 66198 576918 66434
rect 577154 66198 577196 66434
rect 576876 59434 577196 66198
rect 576876 59198 576918 59434
rect 577154 59198 577196 59434
rect 576876 52434 577196 59198
rect 576876 52198 576918 52434
rect 577154 52198 577196 52434
rect 576876 45434 577196 52198
rect 576876 45198 576918 45434
rect 577154 45198 577196 45434
rect 576876 38434 577196 45198
rect 576876 38198 576918 38434
rect 577154 38198 577196 38434
rect 576876 31434 577196 38198
rect 576876 31198 576918 31434
rect 577154 31198 577196 31434
rect 576876 24434 577196 31198
rect 576876 24198 576918 24434
rect 577154 24198 577196 24434
rect 576876 17434 577196 24198
rect 576876 17198 576918 17434
rect 577154 17198 577196 17434
rect 576876 10434 577196 17198
rect 576876 10198 576918 10434
rect 577154 10198 577196 10434
rect 576876 3434 577196 10198
rect 576876 3198 576918 3434
rect 577154 3198 577196 3434
rect 576876 -1706 577196 3198
rect 576876 -1942 576918 -1706
rect 577154 -1942 577196 -1706
rect 576876 -2026 577196 -1942
rect 576876 -2262 576918 -2026
rect 577154 -2262 577196 -2026
rect 576876 -2294 577196 -2262
rect 582144 705238 582464 706230
rect 582144 705002 582186 705238
rect 582422 705002 582464 705238
rect 582144 704918 582464 705002
rect 582144 704682 582186 704918
rect 582422 704682 582464 704918
rect 582144 695494 582464 704682
rect 582144 695258 582186 695494
rect 582422 695258 582464 695494
rect 582144 688494 582464 695258
rect 582144 688258 582186 688494
rect 582422 688258 582464 688494
rect 582144 681494 582464 688258
rect 582144 681258 582186 681494
rect 582422 681258 582464 681494
rect 582144 674494 582464 681258
rect 582144 674258 582186 674494
rect 582422 674258 582464 674494
rect 582144 667494 582464 674258
rect 582144 667258 582186 667494
rect 582422 667258 582464 667494
rect 582144 660494 582464 667258
rect 582144 660258 582186 660494
rect 582422 660258 582464 660494
rect 582144 653494 582464 660258
rect 582144 653258 582186 653494
rect 582422 653258 582464 653494
rect 582144 646494 582464 653258
rect 582144 646258 582186 646494
rect 582422 646258 582464 646494
rect 582144 639494 582464 646258
rect 582144 639258 582186 639494
rect 582422 639258 582464 639494
rect 582144 632494 582464 639258
rect 582144 632258 582186 632494
rect 582422 632258 582464 632494
rect 582144 625494 582464 632258
rect 582144 625258 582186 625494
rect 582422 625258 582464 625494
rect 582144 618494 582464 625258
rect 582144 618258 582186 618494
rect 582422 618258 582464 618494
rect 582144 611494 582464 618258
rect 582144 611258 582186 611494
rect 582422 611258 582464 611494
rect 582144 604494 582464 611258
rect 582144 604258 582186 604494
rect 582422 604258 582464 604494
rect 582144 597494 582464 604258
rect 582144 597258 582186 597494
rect 582422 597258 582464 597494
rect 582144 590494 582464 597258
rect 582144 590258 582186 590494
rect 582422 590258 582464 590494
rect 582144 583494 582464 590258
rect 582144 583258 582186 583494
rect 582422 583258 582464 583494
rect 582144 576494 582464 583258
rect 582144 576258 582186 576494
rect 582422 576258 582464 576494
rect 582144 569494 582464 576258
rect 582144 569258 582186 569494
rect 582422 569258 582464 569494
rect 582144 562494 582464 569258
rect 582144 562258 582186 562494
rect 582422 562258 582464 562494
rect 582144 555494 582464 562258
rect 582144 555258 582186 555494
rect 582422 555258 582464 555494
rect 582144 548494 582464 555258
rect 582144 548258 582186 548494
rect 582422 548258 582464 548494
rect 582144 541494 582464 548258
rect 582144 541258 582186 541494
rect 582422 541258 582464 541494
rect 582144 534494 582464 541258
rect 582144 534258 582186 534494
rect 582422 534258 582464 534494
rect 582144 527494 582464 534258
rect 582144 527258 582186 527494
rect 582422 527258 582464 527494
rect 582144 520494 582464 527258
rect 582144 520258 582186 520494
rect 582422 520258 582464 520494
rect 582144 513494 582464 520258
rect 582144 513258 582186 513494
rect 582422 513258 582464 513494
rect 582144 506494 582464 513258
rect 582144 506258 582186 506494
rect 582422 506258 582464 506494
rect 582144 499494 582464 506258
rect 582144 499258 582186 499494
rect 582422 499258 582464 499494
rect 582144 492494 582464 499258
rect 582144 492258 582186 492494
rect 582422 492258 582464 492494
rect 582144 485494 582464 492258
rect 582144 485258 582186 485494
rect 582422 485258 582464 485494
rect 582144 478494 582464 485258
rect 582144 478258 582186 478494
rect 582422 478258 582464 478494
rect 582144 471494 582464 478258
rect 582144 471258 582186 471494
rect 582422 471258 582464 471494
rect 582144 464494 582464 471258
rect 582144 464258 582186 464494
rect 582422 464258 582464 464494
rect 582144 457494 582464 464258
rect 582144 457258 582186 457494
rect 582422 457258 582464 457494
rect 582144 450494 582464 457258
rect 582144 450258 582186 450494
rect 582422 450258 582464 450494
rect 582144 443494 582464 450258
rect 582144 443258 582186 443494
rect 582422 443258 582464 443494
rect 582144 436494 582464 443258
rect 582144 436258 582186 436494
rect 582422 436258 582464 436494
rect 582144 429494 582464 436258
rect 582144 429258 582186 429494
rect 582422 429258 582464 429494
rect 582144 422494 582464 429258
rect 582144 422258 582186 422494
rect 582422 422258 582464 422494
rect 582144 415494 582464 422258
rect 582144 415258 582186 415494
rect 582422 415258 582464 415494
rect 582144 408494 582464 415258
rect 582144 408258 582186 408494
rect 582422 408258 582464 408494
rect 582144 401494 582464 408258
rect 582144 401258 582186 401494
rect 582422 401258 582464 401494
rect 582144 394494 582464 401258
rect 582144 394258 582186 394494
rect 582422 394258 582464 394494
rect 582144 387494 582464 394258
rect 582144 387258 582186 387494
rect 582422 387258 582464 387494
rect 582144 380494 582464 387258
rect 582144 380258 582186 380494
rect 582422 380258 582464 380494
rect 582144 373494 582464 380258
rect 582144 373258 582186 373494
rect 582422 373258 582464 373494
rect 582144 366494 582464 373258
rect 582144 366258 582186 366494
rect 582422 366258 582464 366494
rect 582144 359494 582464 366258
rect 582144 359258 582186 359494
rect 582422 359258 582464 359494
rect 582144 352494 582464 359258
rect 582144 352258 582186 352494
rect 582422 352258 582464 352494
rect 582144 345494 582464 352258
rect 582144 345258 582186 345494
rect 582422 345258 582464 345494
rect 582144 338494 582464 345258
rect 582144 338258 582186 338494
rect 582422 338258 582464 338494
rect 582144 331494 582464 338258
rect 582144 331258 582186 331494
rect 582422 331258 582464 331494
rect 582144 324494 582464 331258
rect 582144 324258 582186 324494
rect 582422 324258 582464 324494
rect 582144 317494 582464 324258
rect 582144 317258 582186 317494
rect 582422 317258 582464 317494
rect 582144 310494 582464 317258
rect 582144 310258 582186 310494
rect 582422 310258 582464 310494
rect 582144 303494 582464 310258
rect 582144 303258 582186 303494
rect 582422 303258 582464 303494
rect 582144 296494 582464 303258
rect 582144 296258 582186 296494
rect 582422 296258 582464 296494
rect 582144 289494 582464 296258
rect 582144 289258 582186 289494
rect 582422 289258 582464 289494
rect 582144 282494 582464 289258
rect 582144 282258 582186 282494
rect 582422 282258 582464 282494
rect 582144 275494 582464 282258
rect 582144 275258 582186 275494
rect 582422 275258 582464 275494
rect 582144 268494 582464 275258
rect 582144 268258 582186 268494
rect 582422 268258 582464 268494
rect 582144 261494 582464 268258
rect 582144 261258 582186 261494
rect 582422 261258 582464 261494
rect 582144 254494 582464 261258
rect 582144 254258 582186 254494
rect 582422 254258 582464 254494
rect 582144 247494 582464 254258
rect 582144 247258 582186 247494
rect 582422 247258 582464 247494
rect 582144 240494 582464 247258
rect 582144 240258 582186 240494
rect 582422 240258 582464 240494
rect 582144 233494 582464 240258
rect 582144 233258 582186 233494
rect 582422 233258 582464 233494
rect 582144 226494 582464 233258
rect 582144 226258 582186 226494
rect 582422 226258 582464 226494
rect 582144 219494 582464 226258
rect 582144 219258 582186 219494
rect 582422 219258 582464 219494
rect 582144 212494 582464 219258
rect 582144 212258 582186 212494
rect 582422 212258 582464 212494
rect 582144 205494 582464 212258
rect 582144 205258 582186 205494
rect 582422 205258 582464 205494
rect 582144 198494 582464 205258
rect 582144 198258 582186 198494
rect 582422 198258 582464 198494
rect 582144 191494 582464 198258
rect 582144 191258 582186 191494
rect 582422 191258 582464 191494
rect 582144 184494 582464 191258
rect 582144 184258 582186 184494
rect 582422 184258 582464 184494
rect 582144 177494 582464 184258
rect 582144 177258 582186 177494
rect 582422 177258 582464 177494
rect 582144 170494 582464 177258
rect 582144 170258 582186 170494
rect 582422 170258 582464 170494
rect 582144 163494 582464 170258
rect 582144 163258 582186 163494
rect 582422 163258 582464 163494
rect 582144 156494 582464 163258
rect 582144 156258 582186 156494
rect 582422 156258 582464 156494
rect 582144 149494 582464 156258
rect 582144 149258 582186 149494
rect 582422 149258 582464 149494
rect 582144 142494 582464 149258
rect 582144 142258 582186 142494
rect 582422 142258 582464 142494
rect 582144 135494 582464 142258
rect 582144 135258 582186 135494
rect 582422 135258 582464 135494
rect 582144 128494 582464 135258
rect 582144 128258 582186 128494
rect 582422 128258 582464 128494
rect 582144 121494 582464 128258
rect 582144 121258 582186 121494
rect 582422 121258 582464 121494
rect 582144 114494 582464 121258
rect 582144 114258 582186 114494
rect 582422 114258 582464 114494
rect 582144 107494 582464 114258
rect 582144 107258 582186 107494
rect 582422 107258 582464 107494
rect 582144 100494 582464 107258
rect 582144 100258 582186 100494
rect 582422 100258 582464 100494
rect 582144 93494 582464 100258
rect 582144 93258 582186 93494
rect 582422 93258 582464 93494
rect 582144 86494 582464 93258
rect 582144 86258 582186 86494
rect 582422 86258 582464 86494
rect 582144 79494 582464 86258
rect 582144 79258 582186 79494
rect 582422 79258 582464 79494
rect 582144 72494 582464 79258
rect 582144 72258 582186 72494
rect 582422 72258 582464 72494
rect 582144 65494 582464 72258
rect 582144 65258 582186 65494
rect 582422 65258 582464 65494
rect 582144 58494 582464 65258
rect 582144 58258 582186 58494
rect 582422 58258 582464 58494
rect 582144 51494 582464 58258
rect 582144 51258 582186 51494
rect 582422 51258 582464 51494
rect 582144 44494 582464 51258
rect 582144 44258 582186 44494
rect 582422 44258 582464 44494
rect 582144 37494 582464 44258
rect 582144 37258 582186 37494
rect 582422 37258 582464 37494
rect 582144 30494 582464 37258
rect 582144 30258 582186 30494
rect 582422 30258 582464 30494
rect 582144 23494 582464 30258
rect 582144 23258 582186 23494
rect 582422 23258 582464 23494
rect 582144 16494 582464 23258
rect 582144 16258 582186 16494
rect 582422 16258 582464 16494
rect 582144 9494 582464 16258
rect 582144 9258 582186 9494
rect 582422 9258 582464 9494
rect 582144 2494 582464 9258
rect 582144 2258 582186 2494
rect 582422 2258 582464 2494
rect 582144 -746 582464 2258
rect 582144 -982 582186 -746
rect 582422 -982 582464 -746
rect 582144 -1066 582464 -982
rect 582144 -1302 582186 -1066
rect 582422 -1302 582464 -1066
rect 582144 -2294 582464 -1302
rect 585710 705238 587122 706062
rect 585710 705002 585818 705238
rect 586054 705002 586138 705238
rect 586374 705002 586458 705238
rect 586694 705002 586778 705238
rect 587014 705002 587122 705238
rect 585710 704918 587122 705002
rect 585710 704682 585818 704918
rect 586054 704682 586138 704918
rect 586374 704682 586458 704918
rect 586694 704682 586778 704918
rect 587014 704682 587122 704918
rect 585710 695494 587122 704682
rect 585710 695258 585818 695494
rect 586054 695258 586138 695494
rect 586374 695258 586458 695494
rect 586694 695258 586778 695494
rect 587014 695258 587122 695494
rect 585710 688494 587122 695258
rect 585710 688258 585818 688494
rect 586054 688258 586138 688494
rect 586374 688258 586458 688494
rect 586694 688258 586778 688494
rect 587014 688258 587122 688494
rect 585710 681494 587122 688258
rect 585710 681258 585818 681494
rect 586054 681258 586138 681494
rect 586374 681258 586458 681494
rect 586694 681258 586778 681494
rect 587014 681258 587122 681494
rect 585710 674494 587122 681258
rect 585710 674258 585818 674494
rect 586054 674258 586138 674494
rect 586374 674258 586458 674494
rect 586694 674258 586778 674494
rect 587014 674258 587122 674494
rect 585710 667494 587122 674258
rect 585710 667258 585818 667494
rect 586054 667258 586138 667494
rect 586374 667258 586458 667494
rect 586694 667258 586778 667494
rect 587014 667258 587122 667494
rect 585710 660494 587122 667258
rect 585710 660258 585818 660494
rect 586054 660258 586138 660494
rect 586374 660258 586458 660494
rect 586694 660258 586778 660494
rect 587014 660258 587122 660494
rect 585710 653494 587122 660258
rect 585710 653258 585818 653494
rect 586054 653258 586138 653494
rect 586374 653258 586458 653494
rect 586694 653258 586778 653494
rect 587014 653258 587122 653494
rect 585710 646494 587122 653258
rect 585710 646258 585818 646494
rect 586054 646258 586138 646494
rect 586374 646258 586458 646494
rect 586694 646258 586778 646494
rect 587014 646258 587122 646494
rect 585710 639494 587122 646258
rect 585710 639258 585818 639494
rect 586054 639258 586138 639494
rect 586374 639258 586458 639494
rect 586694 639258 586778 639494
rect 587014 639258 587122 639494
rect 585710 632494 587122 639258
rect 585710 632258 585818 632494
rect 586054 632258 586138 632494
rect 586374 632258 586458 632494
rect 586694 632258 586778 632494
rect 587014 632258 587122 632494
rect 585710 625494 587122 632258
rect 585710 625258 585818 625494
rect 586054 625258 586138 625494
rect 586374 625258 586458 625494
rect 586694 625258 586778 625494
rect 587014 625258 587122 625494
rect 585710 618494 587122 625258
rect 585710 618258 585818 618494
rect 586054 618258 586138 618494
rect 586374 618258 586458 618494
rect 586694 618258 586778 618494
rect 587014 618258 587122 618494
rect 585710 611494 587122 618258
rect 585710 611258 585818 611494
rect 586054 611258 586138 611494
rect 586374 611258 586458 611494
rect 586694 611258 586778 611494
rect 587014 611258 587122 611494
rect 585710 604494 587122 611258
rect 585710 604258 585818 604494
rect 586054 604258 586138 604494
rect 586374 604258 586458 604494
rect 586694 604258 586778 604494
rect 587014 604258 587122 604494
rect 585710 597494 587122 604258
rect 585710 597258 585818 597494
rect 586054 597258 586138 597494
rect 586374 597258 586458 597494
rect 586694 597258 586778 597494
rect 587014 597258 587122 597494
rect 585710 590494 587122 597258
rect 585710 590258 585818 590494
rect 586054 590258 586138 590494
rect 586374 590258 586458 590494
rect 586694 590258 586778 590494
rect 587014 590258 587122 590494
rect 585710 583494 587122 590258
rect 585710 583258 585818 583494
rect 586054 583258 586138 583494
rect 586374 583258 586458 583494
rect 586694 583258 586778 583494
rect 587014 583258 587122 583494
rect 585710 576494 587122 583258
rect 585710 576258 585818 576494
rect 586054 576258 586138 576494
rect 586374 576258 586458 576494
rect 586694 576258 586778 576494
rect 587014 576258 587122 576494
rect 585710 569494 587122 576258
rect 585710 569258 585818 569494
rect 586054 569258 586138 569494
rect 586374 569258 586458 569494
rect 586694 569258 586778 569494
rect 587014 569258 587122 569494
rect 585710 562494 587122 569258
rect 585710 562258 585818 562494
rect 586054 562258 586138 562494
rect 586374 562258 586458 562494
rect 586694 562258 586778 562494
rect 587014 562258 587122 562494
rect 585710 555494 587122 562258
rect 585710 555258 585818 555494
rect 586054 555258 586138 555494
rect 586374 555258 586458 555494
rect 586694 555258 586778 555494
rect 587014 555258 587122 555494
rect 585710 548494 587122 555258
rect 585710 548258 585818 548494
rect 586054 548258 586138 548494
rect 586374 548258 586458 548494
rect 586694 548258 586778 548494
rect 587014 548258 587122 548494
rect 585710 541494 587122 548258
rect 585710 541258 585818 541494
rect 586054 541258 586138 541494
rect 586374 541258 586458 541494
rect 586694 541258 586778 541494
rect 587014 541258 587122 541494
rect 585710 534494 587122 541258
rect 585710 534258 585818 534494
rect 586054 534258 586138 534494
rect 586374 534258 586458 534494
rect 586694 534258 586778 534494
rect 587014 534258 587122 534494
rect 585710 527494 587122 534258
rect 585710 527258 585818 527494
rect 586054 527258 586138 527494
rect 586374 527258 586458 527494
rect 586694 527258 586778 527494
rect 587014 527258 587122 527494
rect 585710 520494 587122 527258
rect 585710 520258 585818 520494
rect 586054 520258 586138 520494
rect 586374 520258 586458 520494
rect 586694 520258 586778 520494
rect 587014 520258 587122 520494
rect 585710 513494 587122 520258
rect 585710 513258 585818 513494
rect 586054 513258 586138 513494
rect 586374 513258 586458 513494
rect 586694 513258 586778 513494
rect 587014 513258 587122 513494
rect 585710 506494 587122 513258
rect 585710 506258 585818 506494
rect 586054 506258 586138 506494
rect 586374 506258 586458 506494
rect 586694 506258 586778 506494
rect 587014 506258 587122 506494
rect 585710 499494 587122 506258
rect 585710 499258 585818 499494
rect 586054 499258 586138 499494
rect 586374 499258 586458 499494
rect 586694 499258 586778 499494
rect 587014 499258 587122 499494
rect 585710 492494 587122 499258
rect 585710 492258 585818 492494
rect 586054 492258 586138 492494
rect 586374 492258 586458 492494
rect 586694 492258 586778 492494
rect 587014 492258 587122 492494
rect 585710 485494 587122 492258
rect 585710 485258 585818 485494
rect 586054 485258 586138 485494
rect 586374 485258 586458 485494
rect 586694 485258 586778 485494
rect 587014 485258 587122 485494
rect 585710 478494 587122 485258
rect 585710 478258 585818 478494
rect 586054 478258 586138 478494
rect 586374 478258 586458 478494
rect 586694 478258 586778 478494
rect 587014 478258 587122 478494
rect 585710 471494 587122 478258
rect 585710 471258 585818 471494
rect 586054 471258 586138 471494
rect 586374 471258 586458 471494
rect 586694 471258 586778 471494
rect 587014 471258 587122 471494
rect 585710 464494 587122 471258
rect 585710 464258 585818 464494
rect 586054 464258 586138 464494
rect 586374 464258 586458 464494
rect 586694 464258 586778 464494
rect 587014 464258 587122 464494
rect 585710 457494 587122 464258
rect 585710 457258 585818 457494
rect 586054 457258 586138 457494
rect 586374 457258 586458 457494
rect 586694 457258 586778 457494
rect 587014 457258 587122 457494
rect 585710 450494 587122 457258
rect 585710 450258 585818 450494
rect 586054 450258 586138 450494
rect 586374 450258 586458 450494
rect 586694 450258 586778 450494
rect 587014 450258 587122 450494
rect 585710 443494 587122 450258
rect 585710 443258 585818 443494
rect 586054 443258 586138 443494
rect 586374 443258 586458 443494
rect 586694 443258 586778 443494
rect 587014 443258 587122 443494
rect 585710 436494 587122 443258
rect 585710 436258 585818 436494
rect 586054 436258 586138 436494
rect 586374 436258 586458 436494
rect 586694 436258 586778 436494
rect 587014 436258 587122 436494
rect 585710 429494 587122 436258
rect 585710 429258 585818 429494
rect 586054 429258 586138 429494
rect 586374 429258 586458 429494
rect 586694 429258 586778 429494
rect 587014 429258 587122 429494
rect 585710 422494 587122 429258
rect 585710 422258 585818 422494
rect 586054 422258 586138 422494
rect 586374 422258 586458 422494
rect 586694 422258 586778 422494
rect 587014 422258 587122 422494
rect 585710 415494 587122 422258
rect 585710 415258 585818 415494
rect 586054 415258 586138 415494
rect 586374 415258 586458 415494
rect 586694 415258 586778 415494
rect 587014 415258 587122 415494
rect 585710 408494 587122 415258
rect 585710 408258 585818 408494
rect 586054 408258 586138 408494
rect 586374 408258 586458 408494
rect 586694 408258 586778 408494
rect 587014 408258 587122 408494
rect 585710 401494 587122 408258
rect 585710 401258 585818 401494
rect 586054 401258 586138 401494
rect 586374 401258 586458 401494
rect 586694 401258 586778 401494
rect 587014 401258 587122 401494
rect 585710 394494 587122 401258
rect 585710 394258 585818 394494
rect 586054 394258 586138 394494
rect 586374 394258 586458 394494
rect 586694 394258 586778 394494
rect 587014 394258 587122 394494
rect 585710 387494 587122 394258
rect 585710 387258 585818 387494
rect 586054 387258 586138 387494
rect 586374 387258 586458 387494
rect 586694 387258 586778 387494
rect 587014 387258 587122 387494
rect 585710 380494 587122 387258
rect 585710 380258 585818 380494
rect 586054 380258 586138 380494
rect 586374 380258 586458 380494
rect 586694 380258 586778 380494
rect 587014 380258 587122 380494
rect 585710 373494 587122 380258
rect 585710 373258 585818 373494
rect 586054 373258 586138 373494
rect 586374 373258 586458 373494
rect 586694 373258 586778 373494
rect 587014 373258 587122 373494
rect 585710 366494 587122 373258
rect 585710 366258 585818 366494
rect 586054 366258 586138 366494
rect 586374 366258 586458 366494
rect 586694 366258 586778 366494
rect 587014 366258 587122 366494
rect 585710 359494 587122 366258
rect 585710 359258 585818 359494
rect 586054 359258 586138 359494
rect 586374 359258 586458 359494
rect 586694 359258 586778 359494
rect 587014 359258 587122 359494
rect 585710 352494 587122 359258
rect 585710 352258 585818 352494
rect 586054 352258 586138 352494
rect 586374 352258 586458 352494
rect 586694 352258 586778 352494
rect 587014 352258 587122 352494
rect 585710 345494 587122 352258
rect 585710 345258 585818 345494
rect 586054 345258 586138 345494
rect 586374 345258 586458 345494
rect 586694 345258 586778 345494
rect 587014 345258 587122 345494
rect 585710 338494 587122 345258
rect 585710 338258 585818 338494
rect 586054 338258 586138 338494
rect 586374 338258 586458 338494
rect 586694 338258 586778 338494
rect 587014 338258 587122 338494
rect 585710 331494 587122 338258
rect 585710 331258 585818 331494
rect 586054 331258 586138 331494
rect 586374 331258 586458 331494
rect 586694 331258 586778 331494
rect 587014 331258 587122 331494
rect 585710 324494 587122 331258
rect 585710 324258 585818 324494
rect 586054 324258 586138 324494
rect 586374 324258 586458 324494
rect 586694 324258 586778 324494
rect 587014 324258 587122 324494
rect 585710 317494 587122 324258
rect 585710 317258 585818 317494
rect 586054 317258 586138 317494
rect 586374 317258 586458 317494
rect 586694 317258 586778 317494
rect 587014 317258 587122 317494
rect 585710 310494 587122 317258
rect 585710 310258 585818 310494
rect 586054 310258 586138 310494
rect 586374 310258 586458 310494
rect 586694 310258 586778 310494
rect 587014 310258 587122 310494
rect 585710 303494 587122 310258
rect 585710 303258 585818 303494
rect 586054 303258 586138 303494
rect 586374 303258 586458 303494
rect 586694 303258 586778 303494
rect 587014 303258 587122 303494
rect 585710 296494 587122 303258
rect 585710 296258 585818 296494
rect 586054 296258 586138 296494
rect 586374 296258 586458 296494
rect 586694 296258 586778 296494
rect 587014 296258 587122 296494
rect 585710 289494 587122 296258
rect 585710 289258 585818 289494
rect 586054 289258 586138 289494
rect 586374 289258 586458 289494
rect 586694 289258 586778 289494
rect 587014 289258 587122 289494
rect 585710 282494 587122 289258
rect 585710 282258 585818 282494
rect 586054 282258 586138 282494
rect 586374 282258 586458 282494
rect 586694 282258 586778 282494
rect 587014 282258 587122 282494
rect 585710 275494 587122 282258
rect 585710 275258 585818 275494
rect 586054 275258 586138 275494
rect 586374 275258 586458 275494
rect 586694 275258 586778 275494
rect 587014 275258 587122 275494
rect 585710 268494 587122 275258
rect 585710 268258 585818 268494
rect 586054 268258 586138 268494
rect 586374 268258 586458 268494
rect 586694 268258 586778 268494
rect 587014 268258 587122 268494
rect 585710 261494 587122 268258
rect 585710 261258 585818 261494
rect 586054 261258 586138 261494
rect 586374 261258 586458 261494
rect 586694 261258 586778 261494
rect 587014 261258 587122 261494
rect 585710 254494 587122 261258
rect 585710 254258 585818 254494
rect 586054 254258 586138 254494
rect 586374 254258 586458 254494
rect 586694 254258 586778 254494
rect 587014 254258 587122 254494
rect 585710 247494 587122 254258
rect 585710 247258 585818 247494
rect 586054 247258 586138 247494
rect 586374 247258 586458 247494
rect 586694 247258 586778 247494
rect 587014 247258 587122 247494
rect 585710 240494 587122 247258
rect 585710 240258 585818 240494
rect 586054 240258 586138 240494
rect 586374 240258 586458 240494
rect 586694 240258 586778 240494
rect 587014 240258 587122 240494
rect 585710 233494 587122 240258
rect 585710 233258 585818 233494
rect 586054 233258 586138 233494
rect 586374 233258 586458 233494
rect 586694 233258 586778 233494
rect 587014 233258 587122 233494
rect 585710 226494 587122 233258
rect 585710 226258 585818 226494
rect 586054 226258 586138 226494
rect 586374 226258 586458 226494
rect 586694 226258 586778 226494
rect 587014 226258 587122 226494
rect 585710 219494 587122 226258
rect 585710 219258 585818 219494
rect 586054 219258 586138 219494
rect 586374 219258 586458 219494
rect 586694 219258 586778 219494
rect 587014 219258 587122 219494
rect 585710 212494 587122 219258
rect 585710 212258 585818 212494
rect 586054 212258 586138 212494
rect 586374 212258 586458 212494
rect 586694 212258 586778 212494
rect 587014 212258 587122 212494
rect 585710 205494 587122 212258
rect 585710 205258 585818 205494
rect 586054 205258 586138 205494
rect 586374 205258 586458 205494
rect 586694 205258 586778 205494
rect 587014 205258 587122 205494
rect 585710 198494 587122 205258
rect 585710 198258 585818 198494
rect 586054 198258 586138 198494
rect 586374 198258 586458 198494
rect 586694 198258 586778 198494
rect 587014 198258 587122 198494
rect 585710 191494 587122 198258
rect 585710 191258 585818 191494
rect 586054 191258 586138 191494
rect 586374 191258 586458 191494
rect 586694 191258 586778 191494
rect 587014 191258 587122 191494
rect 585710 184494 587122 191258
rect 585710 184258 585818 184494
rect 586054 184258 586138 184494
rect 586374 184258 586458 184494
rect 586694 184258 586778 184494
rect 587014 184258 587122 184494
rect 585710 177494 587122 184258
rect 585710 177258 585818 177494
rect 586054 177258 586138 177494
rect 586374 177258 586458 177494
rect 586694 177258 586778 177494
rect 587014 177258 587122 177494
rect 585710 170494 587122 177258
rect 585710 170258 585818 170494
rect 586054 170258 586138 170494
rect 586374 170258 586458 170494
rect 586694 170258 586778 170494
rect 587014 170258 587122 170494
rect 585710 163494 587122 170258
rect 585710 163258 585818 163494
rect 586054 163258 586138 163494
rect 586374 163258 586458 163494
rect 586694 163258 586778 163494
rect 587014 163258 587122 163494
rect 585710 156494 587122 163258
rect 585710 156258 585818 156494
rect 586054 156258 586138 156494
rect 586374 156258 586458 156494
rect 586694 156258 586778 156494
rect 587014 156258 587122 156494
rect 585710 149494 587122 156258
rect 585710 149258 585818 149494
rect 586054 149258 586138 149494
rect 586374 149258 586458 149494
rect 586694 149258 586778 149494
rect 587014 149258 587122 149494
rect 585710 142494 587122 149258
rect 585710 142258 585818 142494
rect 586054 142258 586138 142494
rect 586374 142258 586458 142494
rect 586694 142258 586778 142494
rect 587014 142258 587122 142494
rect 585710 135494 587122 142258
rect 585710 135258 585818 135494
rect 586054 135258 586138 135494
rect 586374 135258 586458 135494
rect 586694 135258 586778 135494
rect 587014 135258 587122 135494
rect 585710 128494 587122 135258
rect 585710 128258 585818 128494
rect 586054 128258 586138 128494
rect 586374 128258 586458 128494
rect 586694 128258 586778 128494
rect 587014 128258 587122 128494
rect 585710 121494 587122 128258
rect 585710 121258 585818 121494
rect 586054 121258 586138 121494
rect 586374 121258 586458 121494
rect 586694 121258 586778 121494
rect 587014 121258 587122 121494
rect 585710 114494 587122 121258
rect 585710 114258 585818 114494
rect 586054 114258 586138 114494
rect 586374 114258 586458 114494
rect 586694 114258 586778 114494
rect 587014 114258 587122 114494
rect 585710 107494 587122 114258
rect 585710 107258 585818 107494
rect 586054 107258 586138 107494
rect 586374 107258 586458 107494
rect 586694 107258 586778 107494
rect 587014 107258 587122 107494
rect 585710 100494 587122 107258
rect 585710 100258 585818 100494
rect 586054 100258 586138 100494
rect 586374 100258 586458 100494
rect 586694 100258 586778 100494
rect 587014 100258 587122 100494
rect 585710 93494 587122 100258
rect 585710 93258 585818 93494
rect 586054 93258 586138 93494
rect 586374 93258 586458 93494
rect 586694 93258 586778 93494
rect 587014 93258 587122 93494
rect 585710 86494 587122 93258
rect 585710 86258 585818 86494
rect 586054 86258 586138 86494
rect 586374 86258 586458 86494
rect 586694 86258 586778 86494
rect 587014 86258 587122 86494
rect 585710 79494 587122 86258
rect 585710 79258 585818 79494
rect 586054 79258 586138 79494
rect 586374 79258 586458 79494
rect 586694 79258 586778 79494
rect 587014 79258 587122 79494
rect 585710 72494 587122 79258
rect 585710 72258 585818 72494
rect 586054 72258 586138 72494
rect 586374 72258 586458 72494
rect 586694 72258 586778 72494
rect 587014 72258 587122 72494
rect 585710 65494 587122 72258
rect 585710 65258 585818 65494
rect 586054 65258 586138 65494
rect 586374 65258 586458 65494
rect 586694 65258 586778 65494
rect 587014 65258 587122 65494
rect 585710 58494 587122 65258
rect 585710 58258 585818 58494
rect 586054 58258 586138 58494
rect 586374 58258 586458 58494
rect 586694 58258 586778 58494
rect 587014 58258 587122 58494
rect 585710 51494 587122 58258
rect 585710 51258 585818 51494
rect 586054 51258 586138 51494
rect 586374 51258 586458 51494
rect 586694 51258 586778 51494
rect 587014 51258 587122 51494
rect 585710 44494 587122 51258
rect 585710 44258 585818 44494
rect 586054 44258 586138 44494
rect 586374 44258 586458 44494
rect 586694 44258 586778 44494
rect 587014 44258 587122 44494
rect 585710 37494 587122 44258
rect 585710 37258 585818 37494
rect 586054 37258 586138 37494
rect 586374 37258 586458 37494
rect 586694 37258 586778 37494
rect 587014 37258 587122 37494
rect 585710 30494 587122 37258
rect 585710 30258 585818 30494
rect 586054 30258 586138 30494
rect 586374 30258 586458 30494
rect 586694 30258 586778 30494
rect 587014 30258 587122 30494
rect 585710 23494 587122 30258
rect 585710 23258 585818 23494
rect 586054 23258 586138 23494
rect 586374 23258 586458 23494
rect 586694 23258 586778 23494
rect 587014 23258 587122 23494
rect 585710 16494 587122 23258
rect 585710 16258 585818 16494
rect 586054 16258 586138 16494
rect 586374 16258 586458 16494
rect 586694 16258 586778 16494
rect 587014 16258 587122 16494
rect 585710 9494 587122 16258
rect 585710 9258 585818 9494
rect 586054 9258 586138 9494
rect 586374 9258 586458 9494
rect 586694 9258 586778 9494
rect 587014 9258 587122 9494
rect 585710 2494 587122 9258
rect 585710 2258 585818 2494
rect 586054 2258 586138 2494
rect 586374 2258 586458 2494
rect 586694 2258 586778 2494
rect 587014 2258 587122 2494
rect 585710 -746 587122 2258
rect 585710 -982 585818 -746
rect 586054 -982 586138 -746
rect 586374 -982 586458 -746
rect 586694 -982 586778 -746
rect 587014 -982 587122 -746
rect 585710 -1066 587122 -982
rect 585710 -1302 585818 -1066
rect 586054 -1302 586138 -1066
rect 586374 -1302 586458 -1066
rect 586694 -1302 586778 -1066
rect 587014 -1302 587122 -1066
rect 585710 -2126 587122 -1302
rect 587462 696434 588874 707814
rect 587462 696198 587570 696434
rect 587806 696198 587890 696434
rect 588126 696198 588210 696434
rect 588446 696198 588530 696434
rect 588766 696198 588874 696434
rect 587462 689434 588874 696198
rect 587462 689198 587570 689434
rect 587806 689198 587890 689434
rect 588126 689198 588210 689434
rect 588446 689198 588530 689434
rect 588766 689198 588874 689434
rect 587462 682434 588874 689198
rect 587462 682198 587570 682434
rect 587806 682198 587890 682434
rect 588126 682198 588210 682434
rect 588446 682198 588530 682434
rect 588766 682198 588874 682434
rect 587462 675434 588874 682198
rect 587462 675198 587570 675434
rect 587806 675198 587890 675434
rect 588126 675198 588210 675434
rect 588446 675198 588530 675434
rect 588766 675198 588874 675434
rect 587462 668434 588874 675198
rect 587462 668198 587570 668434
rect 587806 668198 587890 668434
rect 588126 668198 588210 668434
rect 588446 668198 588530 668434
rect 588766 668198 588874 668434
rect 587462 661434 588874 668198
rect 587462 661198 587570 661434
rect 587806 661198 587890 661434
rect 588126 661198 588210 661434
rect 588446 661198 588530 661434
rect 588766 661198 588874 661434
rect 587462 654434 588874 661198
rect 587462 654198 587570 654434
rect 587806 654198 587890 654434
rect 588126 654198 588210 654434
rect 588446 654198 588530 654434
rect 588766 654198 588874 654434
rect 587462 647434 588874 654198
rect 587462 647198 587570 647434
rect 587806 647198 587890 647434
rect 588126 647198 588210 647434
rect 588446 647198 588530 647434
rect 588766 647198 588874 647434
rect 587462 640434 588874 647198
rect 587462 640198 587570 640434
rect 587806 640198 587890 640434
rect 588126 640198 588210 640434
rect 588446 640198 588530 640434
rect 588766 640198 588874 640434
rect 587462 633434 588874 640198
rect 587462 633198 587570 633434
rect 587806 633198 587890 633434
rect 588126 633198 588210 633434
rect 588446 633198 588530 633434
rect 588766 633198 588874 633434
rect 587462 626434 588874 633198
rect 587462 626198 587570 626434
rect 587806 626198 587890 626434
rect 588126 626198 588210 626434
rect 588446 626198 588530 626434
rect 588766 626198 588874 626434
rect 587462 619434 588874 626198
rect 587462 619198 587570 619434
rect 587806 619198 587890 619434
rect 588126 619198 588210 619434
rect 588446 619198 588530 619434
rect 588766 619198 588874 619434
rect 587462 612434 588874 619198
rect 587462 612198 587570 612434
rect 587806 612198 587890 612434
rect 588126 612198 588210 612434
rect 588446 612198 588530 612434
rect 588766 612198 588874 612434
rect 587462 605434 588874 612198
rect 587462 605198 587570 605434
rect 587806 605198 587890 605434
rect 588126 605198 588210 605434
rect 588446 605198 588530 605434
rect 588766 605198 588874 605434
rect 587462 598434 588874 605198
rect 587462 598198 587570 598434
rect 587806 598198 587890 598434
rect 588126 598198 588210 598434
rect 588446 598198 588530 598434
rect 588766 598198 588874 598434
rect 587462 591434 588874 598198
rect 587462 591198 587570 591434
rect 587806 591198 587890 591434
rect 588126 591198 588210 591434
rect 588446 591198 588530 591434
rect 588766 591198 588874 591434
rect 587462 584434 588874 591198
rect 587462 584198 587570 584434
rect 587806 584198 587890 584434
rect 588126 584198 588210 584434
rect 588446 584198 588530 584434
rect 588766 584198 588874 584434
rect 587462 577434 588874 584198
rect 587462 577198 587570 577434
rect 587806 577198 587890 577434
rect 588126 577198 588210 577434
rect 588446 577198 588530 577434
rect 588766 577198 588874 577434
rect 587462 570434 588874 577198
rect 587462 570198 587570 570434
rect 587806 570198 587890 570434
rect 588126 570198 588210 570434
rect 588446 570198 588530 570434
rect 588766 570198 588874 570434
rect 587462 563434 588874 570198
rect 587462 563198 587570 563434
rect 587806 563198 587890 563434
rect 588126 563198 588210 563434
rect 588446 563198 588530 563434
rect 588766 563198 588874 563434
rect 587462 556434 588874 563198
rect 587462 556198 587570 556434
rect 587806 556198 587890 556434
rect 588126 556198 588210 556434
rect 588446 556198 588530 556434
rect 588766 556198 588874 556434
rect 587462 549434 588874 556198
rect 587462 549198 587570 549434
rect 587806 549198 587890 549434
rect 588126 549198 588210 549434
rect 588446 549198 588530 549434
rect 588766 549198 588874 549434
rect 587462 542434 588874 549198
rect 587462 542198 587570 542434
rect 587806 542198 587890 542434
rect 588126 542198 588210 542434
rect 588446 542198 588530 542434
rect 588766 542198 588874 542434
rect 587462 535434 588874 542198
rect 587462 535198 587570 535434
rect 587806 535198 587890 535434
rect 588126 535198 588210 535434
rect 588446 535198 588530 535434
rect 588766 535198 588874 535434
rect 587462 528434 588874 535198
rect 587462 528198 587570 528434
rect 587806 528198 587890 528434
rect 588126 528198 588210 528434
rect 588446 528198 588530 528434
rect 588766 528198 588874 528434
rect 587462 521434 588874 528198
rect 587462 521198 587570 521434
rect 587806 521198 587890 521434
rect 588126 521198 588210 521434
rect 588446 521198 588530 521434
rect 588766 521198 588874 521434
rect 587462 514434 588874 521198
rect 587462 514198 587570 514434
rect 587806 514198 587890 514434
rect 588126 514198 588210 514434
rect 588446 514198 588530 514434
rect 588766 514198 588874 514434
rect 587462 507434 588874 514198
rect 587462 507198 587570 507434
rect 587806 507198 587890 507434
rect 588126 507198 588210 507434
rect 588446 507198 588530 507434
rect 588766 507198 588874 507434
rect 587462 500434 588874 507198
rect 587462 500198 587570 500434
rect 587806 500198 587890 500434
rect 588126 500198 588210 500434
rect 588446 500198 588530 500434
rect 588766 500198 588874 500434
rect 587462 493434 588874 500198
rect 587462 493198 587570 493434
rect 587806 493198 587890 493434
rect 588126 493198 588210 493434
rect 588446 493198 588530 493434
rect 588766 493198 588874 493434
rect 587462 486434 588874 493198
rect 587462 486198 587570 486434
rect 587806 486198 587890 486434
rect 588126 486198 588210 486434
rect 588446 486198 588530 486434
rect 588766 486198 588874 486434
rect 587462 479434 588874 486198
rect 587462 479198 587570 479434
rect 587806 479198 587890 479434
rect 588126 479198 588210 479434
rect 588446 479198 588530 479434
rect 588766 479198 588874 479434
rect 587462 472434 588874 479198
rect 587462 472198 587570 472434
rect 587806 472198 587890 472434
rect 588126 472198 588210 472434
rect 588446 472198 588530 472434
rect 588766 472198 588874 472434
rect 587462 465434 588874 472198
rect 587462 465198 587570 465434
rect 587806 465198 587890 465434
rect 588126 465198 588210 465434
rect 588446 465198 588530 465434
rect 588766 465198 588874 465434
rect 587462 458434 588874 465198
rect 587462 458198 587570 458434
rect 587806 458198 587890 458434
rect 588126 458198 588210 458434
rect 588446 458198 588530 458434
rect 588766 458198 588874 458434
rect 587462 451434 588874 458198
rect 587462 451198 587570 451434
rect 587806 451198 587890 451434
rect 588126 451198 588210 451434
rect 588446 451198 588530 451434
rect 588766 451198 588874 451434
rect 587462 444434 588874 451198
rect 587462 444198 587570 444434
rect 587806 444198 587890 444434
rect 588126 444198 588210 444434
rect 588446 444198 588530 444434
rect 588766 444198 588874 444434
rect 587462 437434 588874 444198
rect 587462 437198 587570 437434
rect 587806 437198 587890 437434
rect 588126 437198 588210 437434
rect 588446 437198 588530 437434
rect 588766 437198 588874 437434
rect 587462 430434 588874 437198
rect 587462 430198 587570 430434
rect 587806 430198 587890 430434
rect 588126 430198 588210 430434
rect 588446 430198 588530 430434
rect 588766 430198 588874 430434
rect 587462 423434 588874 430198
rect 587462 423198 587570 423434
rect 587806 423198 587890 423434
rect 588126 423198 588210 423434
rect 588446 423198 588530 423434
rect 588766 423198 588874 423434
rect 587462 416434 588874 423198
rect 587462 416198 587570 416434
rect 587806 416198 587890 416434
rect 588126 416198 588210 416434
rect 588446 416198 588530 416434
rect 588766 416198 588874 416434
rect 587462 409434 588874 416198
rect 587462 409198 587570 409434
rect 587806 409198 587890 409434
rect 588126 409198 588210 409434
rect 588446 409198 588530 409434
rect 588766 409198 588874 409434
rect 587462 402434 588874 409198
rect 587462 402198 587570 402434
rect 587806 402198 587890 402434
rect 588126 402198 588210 402434
rect 588446 402198 588530 402434
rect 588766 402198 588874 402434
rect 587462 395434 588874 402198
rect 587462 395198 587570 395434
rect 587806 395198 587890 395434
rect 588126 395198 588210 395434
rect 588446 395198 588530 395434
rect 588766 395198 588874 395434
rect 587462 388434 588874 395198
rect 587462 388198 587570 388434
rect 587806 388198 587890 388434
rect 588126 388198 588210 388434
rect 588446 388198 588530 388434
rect 588766 388198 588874 388434
rect 587462 381434 588874 388198
rect 587462 381198 587570 381434
rect 587806 381198 587890 381434
rect 588126 381198 588210 381434
rect 588446 381198 588530 381434
rect 588766 381198 588874 381434
rect 587462 374434 588874 381198
rect 587462 374198 587570 374434
rect 587806 374198 587890 374434
rect 588126 374198 588210 374434
rect 588446 374198 588530 374434
rect 588766 374198 588874 374434
rect 587462 367434 588874 374198
rect 587462 367198 587570 367434
rect 587806 367198 587890 367434
rect 588126 367198 588210 367434
rect 588446 367198 588530 367434
rect 588766 367198 588874 367434
rect 587462 360434 588874 367198
rect 587462 360198 587570 360434
rect 587806 360198 587890 360434
rect 588126 360198 588210 360434
rect 588446 360198 588530 360434
rect 588766 360198 588874 360434
rect 587462 353434 588874 360198
rect 587462 353198 587570 353434
rect 587806 353198 587890 353434
rect 588126 353198 588210 353434
rect 588446 353198 588530 353434
rect 588766 353198 588874 353434
rect 587462 346434 588874 353198
rect 587462 346198 587570 346434
rect 587806 346198 587890 346434
rect 588126 346198 588210 346434
rect 588446 346198 588530 346434
rect 588766 346198 588874 346434
rect 587462 339434 588874 346198
rect 587462 339198 587570 339434
rect 587806 339198 587890 339434
rect 588126 339198 588210 339434
rect 588446 339198 588530 339434
rect 588766 339198 588874 339434
rect 587462 332434 588874 339198
rect 587462 332198 587570 332434
rect 587806 332198 587890 332434
rect 588126 332198 588210 332434
rect 588446 332198 588530 332434
rect 588766 332198 588874 332434
rect 587462 325434 588874 332198
rect 587462 325198 587570 325434
rect 587806 325198 587890 325434
rect 588126 325198 588210 325434
rect 588446 325198 588530 325434
rect 588766 325198 588874 325434
rect 587462 318434 588874 325198
rect 587462 318198 587570 318434
rect 587806 318198 587890 318434
rect 588126 318198 588210 318434
rect 588446 318198 588530 318434
rect 588766 318198 588874 318434
rect 587462 311434 588874 318198
rect 587462 311198 587570 311434
rect 587806 311198 587890 311434
rect 588126 311198 588210 311434
rect 588446 311198 588530 311434
rect 588766 311198 588874 311434
rect 587462 304434 588874 311198
rect 587462 304198 587570 304434
rect 587806 304198 587890 304434
rect 588126 304198 588210 304434
rect 588446 304198 588530 304434
rect 588766 304198 588874 304434
rect 587462 297434 588874 304198
rect 587462 297198 587570 297434
rect 587806 297198 587890 297434
rect 588126 297198 588210 297434
rect 588446 297198 588530 297434
rect 588766 297198 588874 297434
rect 587462 290434 588874 297198
rect 587462 290198 587570 290434
rect 587806 290198 587890 290434
rect 588126 290198 588210 290434
rect 588446 290198 588530 290434
rect 588766 290198 588874 290434
rect 587462 283434 588874 290198
rect 587462 283198 587570 283434
rect 587806 283198 587890 283434
rect 588126 283198 588210 283434
rect 588446 283198 588530 283434
rect 588766 283198 588874 283434
rect 587462 276434 588874 283198
rect 587462 276198 587570 276434
rect 587806 276198 587890 276434
rect 588126 276198 588210 276434
rect 588446 276198 588530 276434
rect 588766 276198 588874 276434
rect 587462 269434 588874 276198
rect 587462 269198 587570 269434
rect 587806 269198 587890 269434
rect 588126 269198 588210 269434
rect 588446 269198 588530 269434
rect 588766 269198 588874 269434
rect 587462 262434 588874 269198
rect 587462 262198 587570 262434
rect 587806 262198 587890 262434
rect 588126 262198 588210 262434
rect 588446 262198 588530 262434
rect 588766 262198 588874 262434
rect 587462 255434 588874 262198
rect 587462 255198 587570 255434
rect 587806 255198 587890 255434
rect 588126 255198 588210 255434
rect 588446 255198 588530 255434
rect 588766 255198 588874 255434
rect 587462 248434 588874 255198
rect 587462 248198 587570 248434
rect 587806 248198 587890 248434
rect 588126 248198 588210 248434
rect 588446 248198 588530 248434
rect 588766 248198 588874 248434
rect 587462 241434 588874 248198
rect 587462 241198 587570 241434
rect 587806 241198 587890 241434
rect 588126 241198 588210 241434
rect 588446 241198 588530 241434
rect 588766 241198 588874 241434
rect 587462 234434 588874 241198
rect 587462 234198 587570 234434
rect 587806 234198 587890 234434
rect 588126 234198 588210 234434
rect 588446 234198 588530 234434
rect 588766 234198 588874 234434
rect 587462 227434 588874 234198
rect 587462 227198 587570 227434
rect 587806 227198 587890 227434
rect 588126 227198 588210 227434
rect 588446 227198 588530 227434
rect 588766 227198 588874 227434
rect 587462 220434 588874 227198
rect 587462 220198 587570 220434
rect 587806 220198 587890 220434
rect 588126 220198 588210 220434
rect 588446 220198 588530 220434
rect 588766 220198 588874 220434
rect 587462 213434 588874 220198
rect 587462 213198 587570 213434
rect 587806 213198 587890 213434
rect 588126 213198 588210 213434
rect 588446 213198 588530 213434
rect 588766 213198 588874 213434
rect 587462 206434 588874 213198
rect 587462 206198 587570 206434
rect 587806 206198 587890 206434
rect 588126 206198 588210 206434
rect 588446 206198 588530 206434
rect 588766 206198 588874 206434
rect 587462 199434 588874 206198
rect 587462 199198 587570 199434
rect 587806 199198 587890 199434
rect 588126 199198 588210 199434
rect 588446 199198 588530 199434
rect 588766 199198 588874 199434
rect 587462 192434 588874 199198
rect 587462 192198 587570 192434
rect 587806 192198 587890 192434
rect 588126 192198 588210 192434
rect 588446 192198 588530 192434
rect 588766 192198 588874 192434
rect 587462 185434 588874 192198
rect 587462 185198 587570 185434
rect 587806 185198 587890 185434
rect 588126 185198 588210 185434
rect 588446 185198 588530 185434
rect 588766 185198 588874 185434
rect 587462 178434 588874 185198
rect 587462 178198 587570 178434
rect 587806 178198 587890 178434
rect 588126 178198 588210 178434
rect 588446 178198 588530 178434
rect 588766 178198 588874 178434
rect 587462 171434 588874 178198
rect 587462 171198 587570 171434
rect 587806 171198 587890 171434
rect 588126 171198 588210 171434
rect 588446 171198 588530 171434
rect 588766 171198 588874 171434
rect 587462 164434 588874 171198
rect 587462 164198 587570 164434
rect 587806 164198 587890 164434
rect 588126 164198 588210 164434
rect 588446 164198 588530 164434
rect 588766 164198 588874 164434
rect 587462 157434 588874 164198
rect 587462 157198 587570 157434
rect 587806 157198 587890 157434
rect 588126 157198 588210 157434
rect 588446 157198 588530 157434
rect 588766 157198 588874 157434
rect 587462 150434 588874 157198
rect 587462 150198 587570 150434
rect 587806 150198 587890 150434
rect 588126 150198 588210 150434
rect 588446 150198 588530 150434
rect 588766 150198 588874 150434
rect 587462 143434 588874 150198
rect 587462 143198 587570 143434
rect 587806 143198 587890 143434
rect 588126 143198 588210 143434
rect 588446 143198 588530 143434
rect 588766 143198 588874 143434
rect 587462 136434 588874 143198
rect 587462 136198 587570 136434
rect 587806 136198 587890 136434
rect 588126 136198 588210 136434
rect 588446 136198 588530 136434
rect 588766 136198 588874 136434
rect 587462 129434 588874 136198
rect 587462 129198 587570 129434
rect 587806 129198 587890 129434
rect 588126 129198 588210 129434
rect 588446 129198 588530 129434
rect 588766 129198 588874 129434
rect 587462 122434 588874 129198
rect 587462 122198 587570 122434
rect 587806 122198 587890 122434
rect 588126 122198 588210 122434
rect 588446 122198 588530 122434
rect 588766 122198 588874 122434
rect 587462 115434 588874 122198
rect 587462 115198 587570 115434
rect 587806 115198 587890 115434
rect 588126 115198 588210 115434
rect 588446 115198 588530 115434
rect 588766 115198 588874 115434
rect 587462 108434 588874 115198
rect 587462 108198 587570 108434
rect 587806 108198 587890 108434
rect 588126 108198 588210 108434
rect 588446 108198 588530 108434
rect 588766 108198 588874 108434
rect 587462 101434 588874 108198
rect 587462 101198 587570 101434
rect 587806 101198 587890 101434
rect 588126 101198 588210 101434
rect 588446 101198 588530 101434
rect 588766 101198 588874 101434
rect 587462 94434 588874 101198
rect 587462 94198 587570 94434
rect 587806 94198 587890 94434
rect 588126 94198 588210 94434
rect 588446 94198 588530 94434
rect 588766 94198 588874 94434
rect 587462 87434 588874 94198
rect 587462 87198 587570 87434
rect 587806 87198 587890 87434
rect 588126 87198 588210 87434
rect 588446 87198 588530 87434
rect 588766 87198 588874 87434
rect 587462 80434 588874 87198
rect 587462 80198 587570 80434
rect 587806 80198 587890 80434
rect 588126 80198 588210 80434
rect 588446 80198 588530 80434
rect 588766 80198 588874 80434
rect 587462 73434 588874 80198
rect 587462 73198 587570 73434
rect 587806 73198 587890 73434
rect 588126 73198 588210 73434
rect 588446 73198 588530 73434
rect 588766 73198 588874 73434
rect 587462 66434 588874 73198
rect 587462 66198 587570 66434
rect 587806 66198 587890 66434
rect 588126 66198 588210 66434
rect 588446 66198 588530 66434
rect 588766 66198 588874 66434
rect 587462 59434 588874 66198
rect 587462 59198 587570 59434
rect 587806 59198 587890 59434
rect 588126 59198 588210 59434
rect 588446 59198 588530 59434
rect 588766 59198 588874 59434
rect 587462 52434 588874 59198
rect 587462 52198 587570 52434
rect 587806 52198 587890 52434
rect 588126 52198 588210 52434
rect 588446 52198 588530 52434
rect 588766 52198 588874 52434
rect 587462 45434 588874 52198
rect 587462 45198 587570 45434
rect 587806 45198 587890 45434
rect 588126 45198 588210 45434
rect 588446 45198 588530 45434
rect 588766 45198 588874 45434
rect 587462 38434 588874 45198
rect 587462 38198 587570 38434
rect 587806 38198 587890 38434
rect 588126 38198 588210 38434
rect 588446 38198 588530 38434
rect 588766 38198 588874 38434
rect 587462 31434 588874 38198
rect 587462 31198 587570 31434
rect 587806 31198 587890 31434
rect 588126 31198 588210 31434
rect 588446 31198 588530 31434
rect 588766 31198 588874 31434
rect 587462 24434 588874 31198
rect 587462 24198 587570 24434
rect 587806 24198 587890 24434
rect 588126 24198 588210 24434
rect 588446 24198 588530 24434
rect 588766 24198 588874 24434
rect 587462 17434 588874 24198
rect 587462 17198 587570 17434
rect 587806 17198 587890 17434
rect 588126 17198 588210 17434
rect 588446 17198 588530 17434
rect 588766 17198 588874 17434
rect 587462 10434 588874 17198
rect 587462 10198 587570 10434
rect 587806 10198 587890 10434
rect 588126 10198 588210 10434
rect 588446 10198 588530 10434
rect 588766 10198 588874 10434
rect 587462 3434 588874 10198
rect 587462 3198 587570 3434
rect 587806 3198 587890 3434
rect 588126 3198 588210 3434
rect 588446 3198 588530 3434
rect 588766 3198 588874 3434
rect 587462 -3878 588874 3198
<< via4 >>
rect -4842 696198 -4606 696434
rect -4522 696198 -4286 696434
rect -4202 696198 -3966 696434
rect -3882 696198 -3646 696434
rect -4842 689198 -4606 689434
rect -4522 689198 -4286 689434
rect -4202 689198 -3966 689434
rect -3882 689198 -3646 689434
rect -4842 682198 -4606 682434
rect -4522 682198 -4286 682434
rect -4202 682198 -3966 682434
rect -3882 682198 -3646 682434
rect -4842 675198 -4606 675434
rect -4522 675198 -4286 675434
rect -4202 675198 -3966 675434
rect -3882 675198 -3646 675434
rect -4842 668198 -4606 668434
rect -4522 668198 -4286 668434
rect -4202 668198 -3966 668434
rect -3882 668198 -3646 668434
rect -4842 661198 -4606 661434
rect -4522 661198 -4286 661434
rect -4202 661198 -3966 661434
rect -3882 661198 -3646 661434
rect -4842 654198 -4606 654434
rect -4522 654198 -4286 654434
rect -4202 654198 -3966 654434
rect -3882 654198 -3646 654434
rect -4842 647198 -4606 647434
rect -4522 647198 -4286 647434
rect -4202 647198 -3966 647434
rect -3882 647198 -3646 647434
rect -4842 640198 -4606 640434
rect -4522 640198 -4286 640434
rect -4202 640198 -3966 640434
rect -3882 640198 -3646 640434
rect -4842 633198 -4606 633434
rect -4522 633198 -4286 633434
rect -4202 633198 -3966 633434
rect -3882 633198 -3646 633434
rect -4842 626198 -4606 626434
rect -4522 626198 -4286 626434
rect -4202 626198 -3966 626434
rect -3882 626198 -3646 626434
rect -4842 619198 -4606 619434
rect -4522 619198 -4286 619434
rect -4202 619198 -3966 619434
rect -3882 619198 -3646 619434
rect -4842 612198 -4606 612434
rect -4522 612198 -4286 612434
rect -4202 612198 -3966 612434
rect -3882 612198 -3646 612434
rect -4842 605198 -4606 605434
rect -4522 605198 -4286 605434
rect -4202 605198 -3966 605434
rect -3882 605198 -3646 605434
rect -4842 598198 -4606 598434
rect -4522 598198 -4286 598434
rect -4202 598198 -3966 598434
rect -3882 598198 -3646 598434
rect -4842 591198 -4606 591434
rect -4522 591198 -4286 591434
rect -4202 591198 -3966 591434
rect -3882 591198 -3646 591434
rect -4842 584198 -4606 584434
rect -4522 584198 -4286 584434
rect -4202 584198 -3966 584434
rect -3882 584198 -3646 584434
rect -4842 577198 -4606 577434
rect -4522 577198 -4286 577434
rect -4202 577198 -3966 577434
rect -3882 577198 -3646 577434
rect -4842 570198 -4606 570434
rect -4522 570198 -4286 570434
rect -4202 570198 -3966 570434
rect -3882 570198 -3646 570434
rect -4842 563198 -4606 563434
rect -4522 563198 -4286 563434
rect -4202 563198 -3966 563434
rect -3882 563198 -3646 563434
rect -4842 556198 -4606 556434
rect -4522 556198 -4286 556434
rect -4202 556198 -3966 556434
rect -3882 556198 -3646 556434
rect -4842 549198 -4606 549434
rect -4522 549198 -4286 549434
rect -4202 549198 -3966 549434
rect -3882 549198 -3646 549434
rect -4842 542198 -4606 542434
rect -4522 542198 -4286 542434
rect -4202 542198 -3966 542434
rect -3882 542198 -3646 542434
rect -4842 535198 -4606 535434
rect -4522 535198 -4286 535434
rect -4202 535198 -3966 535434
rect -3882 535198 -3646 535434
rect -4842 528198 -4606 528434
rect -4522 528198 -4286 528434
rect -4202 528198 -3966 528434
rect -3882 528198 -3646 528434
rect -4842 521198 -4606 521434
rect -4522 521198 -4286 521434
rect -4202 521198 -3966 521434
rect -3882 521198 -3646 521434
rect -4842 514198 -4606 514434
rect -4522 514198 -4286 514434
rect -4202 514198 -3966 514434
rect -3882 514198 -3646 514434
rect -4842 507198 -4606 507434
rect -4522 507198 -4286 507434
rect -4202 507198 -3966 507434
rect -3882 507198 -3646 507434
rect -4842 500198 -4606 500434
rect -4522 500198 -4286 500434
rect -4202 500198 -3966 500434
rect -3882 500198 -3646 500434
rect -4842 493198 -4606 493434
rect -4522 493198 -4286 493434
rect -4202 493198 -3966 493434
rect -3882 493198 -3646 493434
rect -4842 486198 -4606 486434
rect -4522 486198 -4286 486434
rect -4202 486198 -3966 486434
rect -3882 486198 -3646 486434
rect -4842 479198 -4606 479434
rect -4522 479198 -4286 479434
rect -4202 479198 -3966 479434
rect -3882 479198 -3646 479434
rect -4842 472198 -4606 472434
rect -4522 472198 -4286 472434
rect -4202 472198 -3966 472434
rect -3882 472198 -3646 472434
rect -4842 465198 -4606 465434
rect -4522 465198 -4286 465434
rect -4202 465198 -3966 465434
rect -3882 465198 -3646 465434
rect -4842 458198 -4606 458434
rect -4522 458198 -4286 458434
rect -4202 458198 -3966 458434
rect -3882 458198 -3646 458434
rect -4842 451198 -4606 451434
rect -4522 451198 -4286 451434
rect -4202 451198 -3966 451434
rect -3882 451198 -3646 451434
rect -4842 444198 -4606 444434
rect -4522 444198 -4286 444434
rect -4202 444198 -3966 444434
rect -3882 444198 -3646 444434
rect -4842 437198 -4606 437434
rect -4522 437198 -4286 437434
rect -4202 437198 -3966 437434
rect -3882 437198 -3646 437434
rect -4842 430198 -4606 430434
rect -4522 430198 -4286 430434
rect -4202 430198 -3966 430434
rect -3882 430198 -3646 430434
rect -4842 423198 -4606 423434
rect -4522 423198 -4286 423434
rect -4202 423198 -3966 423434
rect -3882 423198 -3646 423434
rect -4842 416198 -4606 416434
rect -4522 416198 -4286 416434
rect -4202 416198 -3966 416434
rect -3882 416198 -3646 416434
rect -4842 409198 -4606 409434
rect -4522 409198 -4286 409434
rect -4202 409198 -3966 409434
rect -3882 409198 -3646 409434
rect -4842 402198 -4606 402434
rect -4522 402198 -4286 402434
rect -4202 402198 -3966 402434
rect -3882 402198 -3646 402434
rect -4842 395198 -4606 395434
rect -4522 395198 -4286 395434
rect -4202 395198 -3966 395434
rect -3882 395198 -3646 395434
rect -4842 388198 -4606 388434
rect -4522 388198 -4286 388434
rect -4202 388198 -3966 388434
rect -3882 388198 -3646 388434
rect -4842 381198 -4606 381434
rect -4522 381198 -4286 381434
rect -4202 381198 -3966 381434
rect -3882 381198 -3646 381434
rect -4842 374198 -4606 374434
rect -4522 374198 -4286 374434
rect -4202 374198 -3966 374434
rect -3882 374198 -3646 374434
rect -4842 367198 -4606 367434
rect -4522 367198 -4286 367434
rect -4202 367198 -3966 367434
rect -3882 367198 -3646 367434
rect -4842 360198 -4606 360434
rect -4522 360198 -4286 360434
rect -4202 360198 -3966 360434
rect -3882 360198 -3646 360434
rect -4842 353198 -4606 353434
rect -4522 353198 -4286 353434
rect -4202 353198 -3966 353434
rect -3882 353198 -3646 353434
rect -4842 346198 -4606 346434
rect -4522 346198 -4286 346434
rect -4202 346198 -3966 346434
rect -3882 346198 -3646 346434
rect -4842 339198 -4606 339434
rect -4522 339198 -4286 339434
rect -4202 339198 -3966 339434
rect -3882 339198 -3646 339434
rect -4842 332198 -4606 332434
rect -4522 332198 -4286 332434
rect -4202 332198 -3966 332434
rect -3882 332198 -3646 332434
rect -4842 325198 -4606 325434
rect -4522 325198 -4286 325434
rect -4202 325198 -3966 325434
rect -3882 325198 -3646 325434
rect -4842 318198 -4606 318434
rect -4522 318198 -4286 318434
rect -4202 318198 -3966 318434
rect -3882 318198 -3646 318434
rect -4842 311198 -4606 311434
rect -4522 311198 -4286 311434
rect -4202 311198 -3966 311434
rect -3882 311198 -3646 311434
rect -4842 304198 -4606 304434
rect -4522 304198 -4286 304434
rect -4202 304198 -3966 304434
rect -3882 304198 -3646 304434
rect -4842 297198 -4606 297434
rect -4522 297198 -4286 297434
rect -4202 297198 -3966 297434
rect -3882 297198 -3646 297434
rect -4842 290198 -4606 290434
rect -4522 290198 -4286 290434
rect -4202 290198 -3966 290434
rect -3882 290198 -3646 290434
rect -4842 283198 -4606 283434
rect -4522 283198 -4286 283434
rect -4202 283198 -3966 283434
rect -3882 283198 -3646 283434
rect -4842 276198 -4606 276434
rect -4522 276198 -4286 276434
rect -4202 276198 -3966 276434
rect -3882 276198 -3646 276434
rect -4842 269198 -4606 269434
rect -4522 269198 -4286 269434
rect -4202 269198 -3966 269434
rect -3882 269198 -3646 269434
rect -4842 262198 -4606 262434
rect -4522 262198 -4286 262434
rect -4202 262198 -3966 262434
rect -3882 262198 -3646 262434
rect -4842 255198 -4606 255434
rect -4522 255198 -4286 255434
rect -4202 255198 -3966 255434
rect -3882 255198 -3646 255434
rect -4842 248198 -4606 248434
rect -4522 248198 -4286 248434
rect -4202 248198 -3966 248434
rect -3882 248198 -3646 248434
rect -4842 241198 -4606 241434
rect -4522 241198 -4286 241434
rect -4202 241198 -3966 241434
rect -3882 241198 -3646 241434
rect -4842 234198 -4606 234434
rect -4522 234198 -4286 234434
rect -4202 234198 -3966 234434
rect -3882 234198 -3646 234434
rect -4842 227198 -4606 227434
rect -4522 227198 -4286 227434
rect -4202 227198 -3966 227434
rect -3882 227198 -3646 227434
rect -4842 220198 -4606 220434
rect -4522 220198 -4286 220434
rect -4202 220198 -3966 220434
rect -3882 220198 -3646 220434
rect -4842 213198 -4606 213434
rect -4522 213198 -4286 213434
rect -4202 213198 -3966 213434
rect -3882 213198 -3646 213434
rect -4842 206198 -4606 206434
rect -4522 206198 -4286 206434
rect -4202 206198 -3966 206434
rect -3882 206198 -3646 206434
rect -4842 199198 -4606 199434
rect -4522 199198 -4286 199434
rect -4202 199198 -3966 199434
rect -3882 199198 -3646 199434
rect -4842 192198 -4606 192434
rect -4522 192198 -4286 192434
rect -4202 192198 -3966 192434
rect -3882 192198 -3646 192434
rect -4842 185198 -4606 185434
rect -4522 185198 -4286 185434
rect -4202 185198 -3966 185434
rect -3882 185198 -3646 185434
rect -4842 178198 -4606 178434
rect -4522 178198 -4286 178434
rect -4202 178198 -3966 178434
rect -3882 178198 -3646 178434
rect -4842 171198 -4606 171434
rect -4522 171198 -4286 171434
rect -4202 171198 -3966 171434
rect -3882 171198 -3646 171434
rect -4842 164198 -4606 164434
rect -4522 164198 -4286 164434
rect -4202 164198 -3966 164434
rect -3882 164198 -3646 164434
rect -4842 157198 -4606 157434
rect -4522 157198 -4286 157434
rect -4202 157198 -3966 157434
rect -3882 157198 -3646 157434
rect -4842 150198 -4606 150434
rect -4522 150198 -4286 150434
rect -4202 150198 -3966 150434
rect -3882 150198 -3646 150434
rect -4842 143198 -4606 143434
rect -4522 143198 -4286 143434
rect -4202 143198 -3966 143434
rect -3882 143198 -3646 143434
rect -4842 136198 -4606 136434
rect -4522 136198 -4286 136434
rect -4202 136198 -3966 136434
rect -3882 136198 -3646 136434
rect -4842 129198 -4606 129434
rect -4522 129198 -4286 129434
rect -4202 129198 -3966 129434
rect -3882 129198 -3646 129434
rect -4842 122198 -4606 122434
rect -4522 122198 -4286 122434
rect -4202 122198 -3966 122434
rect -3882 122198 -3646 122434
rect -4842 115198 -4606 115434
rect -4522 115198 -4286 115434
rect -4202 115198 -3966 115434
rect -3882 115198 -3646 115434
rect -4842 108198 -4606 108434
rect -4522 108198 -4286 108434
rect -4202 108198 -3966 108434
rect -3882 108198 -3646 108434
rect -4842 101198 -4606 101434
rect -4522 101198 -4286 101434
rect -4202 101198 -3966 101434
rect -3882 101198 -3646 101434
rect -4842 94198 -4606 94434
rect -4522 94198 -4286 94434
rect -4202 94198 -3966 94434
rect -3882 94198 -3646 94434
rect -4842 87198 -4606 87434
rect -4522 87198 -4286 87434
rect -4202 87198 -3966 87434
rect -3882 87198 -3646 87434
rect -4842 80198 -4606 80434
rect -4522 80198 -4286 80434
rect -4202 80198 -3966 80434
rect -3882 80198 -3646 80434
rect -4842 73198 -4606 73434
rect -4522 73198 -4286 73434
rect -4202 73198 -3966 73434
rect -3882 73198 -3646 73434
rect -4842 66198 -4606 66434
rect -4522 66198 -4286 66434
rect -4202 66198 -3966 66434
rect -3882 66198 -3646 66434
rect -4842 59198 -4606 59434
rect -4522 59198 -4286 59434
rect -4202 59198 -3966 59434
rect -3882 59198 -3646 59434
rect -4842 52198 -4606 52434
rect -4522 52198 -4286 52434
rect -4202 52198 -3966 52434
rect -3882 52198 -3646 52434
rect -4842 45198 -4606 45434
rect -4522 45198 -4286 45434
rect -4202 45198 -3966 45434
rect -3882 45198 -3646 45434
rect -4842 38198 -4606 38434
rect -4522 38198 -4286 38434
rect -4202 38198 -3966 38434
rect -3882 38198 -3646 38434
rect -4842 31198 -4606 31434
rect -4522 31198 -4286 31434
rect -4202 31198 -3966 31434
rect -3882 31198 -3646 31434
rect -4842 24198 -4606 24434
rect -4522 24198 -4286 24434
rect -4202 24198 -3966 24434
rect -3882 24198 -3646 24434
rect -4842 17198 -4606 17434
rect -4522 17198 -4286 17434
rect -4202 17198 -3966 17434
rect -3882 17198 -3646 17434
rect -4842 10198 -4606 10434
rect -4522 10198 -4286 10434
rect -4202 10198 -3966 10434
rect -3882 10198 -3646 10434
rect -4842 3198 -4606 3434
rect -4522 3198 -4286 3434
rect -4202 3198 -3966 3434
rect -3882 3198 -3646 3434
rect -2374 705002 -2138 705238
rect -2054 705002 -1818 705238
rect -2374 704682 -2138 704918
rect -2054 704682 -1818 704918
rect -3090 695258 -2854 695494
rect -2770 695258 -2534 695494
rect -2450 695258 -2214 695494
rect -2130 695258 -1894 695494
rect -3090 688258 -2854 688494
rect -2770 688258 -2534 688494
rect -2450 688258 -2214 688494
rect -2130 688258 -1894 688494
rect -3090 681258 -2854 681494
rect -2770 681258 -2534 681494
rect -2450 681258 -2214 681494
rect -2130 681258 -1894 681494
rect -3090 674258 -2854 674494
rect -2770 674258 -2534 674494
rect -2450 674258 -2214 674494
rect -2130 674258 -1894 674494
rect -3090 667258 -2854 667494
rect -2770 667258 -2534 667494
rect -2450 667258 -2214 667494
rect -2130 667258 -1894 667494
rect -3090 660258 -2854 660494
rect -2770 660258 -2534 660494
rect -2450 660258 -2214 660494
rect -2130 660258 -1894 660494
rect -3090 653258 -2854 653494
rect -2770 653258 -2534 653494
rect -2450 653258 -2214 653494
rect -2130 653258 -1894 653494
rect -3090 646258 -2854 646494
rect -2770 646258 -2534 646494
rect -2450 646258 -2214 646494
rect -2130 646258 -1894 646494
rect -3090 639258 -2854 639494
rect -2770 639258 -2534 639494
rect -2450 639258 -2214 639494
rect -2130 639258 -1894 639494
rect -3090 632258 -2854 632494
rect -2770 632258 -2534 632494
rect -2450 632258 -2214 632494
rect -2130 632258 -1894 632494
rect -3090 625258 -2854 625494
rect -2770 625258 -2534 625494
rect -2450 625258 -2214 625494
rect -2130 625258 -1894 625494
rect -3090 618258 -2854 618494
rect -2770 618258 -2534 618494
rect -2450 618258 -2214 618494
rect -2130 618258 -1894 618494
rect -3090 611258 -2854 611494
rect -2770 611258 -2534 611494
rect -2450 611258 -2214 611494
rect -2130 611258 -1894 611494
rect -3090 604258 -2854 604494
rect -2770 604258 -2534 604494
rect -2450 604258 -2214 604494
rect -2130 604258 -1894 604494
rect -3090 597258 -2854 597494
rect -2770 597258 -2534 597494
rect -2450 597258 -2214 597494
rect -2130 597258 -1894 597494
rect -3090 590258 -2854 590494
rect -2770 590258 -2534 590494
rect -2450 590258 -2214 590494
rect -2130 590258 -1894 590494
rect -3090 583258 -2854 583494
rect -2770 583258 -2534 583494
rect -2450 583258 -2214 583494
rect -2130 583258 -1894 583494
rect -3090 576258 -2854 576494
rect -2770 576258 -2534 576494
rect -2450 576258 -2214 576494
rect -2130 576258 -1894 576494
rect -3090 569258 -2854 569494
rect -2770 569258 -2534 569494
rect -2450 569258 -2214 569494
rect -2130 569258 -1894 569494
rect -3090 562258 -2854 562494
rect -2770 562258 -2534 562494
rect -2450 562258 -2214 562494
rect -2130 562258 -1894 562494
rect -3090 555258 -2854 555494
rect -2770 555258 -2534 555494
rect -2450 555258 -2214 555494
rect -2130 555258 -1894 555494
rect -3090 548258 -2854 548494
rect -2770 548258 -2534 548494
rect -2450 548258 -2214 548494
rect -2130 548258 -1894 548494
rect -3090 541258 -2854 541494
rect -2770 541258 -2534 541494
rect -2450 541258 -2214 541494
rect -2130 541258 -1894 541494
rect -3090 534258 -2854 534494
rect -2770 534258 -2534 534494
rect -2450 534258 -2214 534494
rect -2130 534258 -1894 534494
rect -3090 527258 -2854 527494
rect -2770 527258 -2534 527494
rect -2450 527258 -2214 527494
rect -2130 527258 -1894 527494
rect -3090 520258 -2854 520494
rect -2770 520258 -2534 520494
rect -2450 520258 -2214 520494
rect -2130 520258 -1894 520494
rect -3090 513258 -2854 513494
rect -2770 513258 -2534 513494
rect -2450 513258 -2214 513494
rect -2130 513258 -1894 513494
rect -3090 506258 -2854 506494
rect -2770 506258 -2534 506494
rect -2450 506258 -2214 506494
rect -2130 506258 -1894 506494
rect -3090 499258 -2854 499494
rect -2770 499258 -2534 499494
rect -2450 499258 -2214 499494
rect -2130 499258 -1894 499494
rect -3090 492258 -2854 492494
rect -2770 492258 -2534 492494
rect -2450 492258 -2214 492494
rect -2130 492258 -1894 492494
rect -3090 485258 -2854 485494
rect -2770 485258 -2534 485494
rect -2450 485258 -2214 485494
rect -2130 485258 -1894 485494
rect -3090 478258 -2854 478494
rect -2770 478258 -2534 478494
rect -2450 478258 -2214 478494
rect -2130 478258 -1894 478494
rect -3090 471258 -2854 471494
rect -2770 471258 -2534 471494
rect -2450 471258 -2214 471494
rect -2130 471258 -1894 471494
rect -3090 464258 -2854 464494
rect -2770 464258 -2534 464494
rect -2450 464258 -2214 464494
rect -2130 464258 -1894 464494
rect -3090 457258 -2854 457494
rect -2770 457258 -2534 457494
rect -2450 457258 -2214 457494
rect -2130 457258 -1894 457494
rect -3090 450258 -2854 450494
rect -2770 450258 -2534 450494
rect -2450 450258 -2214 450494
rect -2130 450258 -1894 450494
rect -3090 443258 -2854 443494
rect -2770 443258 -2534 443494
rect -2450 443258 -2214 443494
rect -2130 443258 -1894 443494
rect -3090 436258 -2854 436494
rect -2770 436258 -2534 436494
rect -2450 436258 -2214 436494
rect -2130 436258 -1894 436494
rect -3090 429258 -2854 429494
rect -2770 429258 -2534 429494
rect -2450 429258 -2214 429494
rect -2130 429258 -1894 429494
rect -3090 422258 -2854 422494
rect -2770 422258 -2534 422494
rect -2450 422258 -2214 422494
rect -2130 422258 -1894 422494
rect -3090 415258 -2854 415494
rect -2770 415258 -2534 415494
rect -2450 415258 -2214 415494
rect -2130 415258 -1894 415494
rect -3090 408258 -2854 408494
rect -2770 408258 -2534 408494
rect -2450 408258 -2214 408494
rect -2130 408258 -1894 408494
rect -3090 401258 -2854 401494
rect -2770 401258 -2534 401494
rect -2450 401258 -2214 401494
rect -2130 401258 -1894 401494
rect -3090 394258 -2854 394494
rect -2770 394258 -2534 394494
rect -2450 394258 -2214 394494
rect -2130 394258 -1894 394494
rect -3090 387258 -2854 387494
rect -2770 387258 -2534 387494
rect -2450 387258 -2214 387494
rect -2130 387258 -1894 387494
rect -3090 380258 -2854 380494
rect -2770 380258 -2534 380494
rect -2450 380258 -2214 380494
rect -2130 380258 -1894 380494
rect -3090 373258 -2854 373494
rect -2770 373258 -2534 373494
rect -2450 373258 -2214 373494
rect -2130 373258 -1894 373494
rect -3090 366258 -2854 366494
rect -2770 366258 -2534 366494
rect -2450 366258 -2214 366494
rect -2130 366258 -1894 366494
rect -3090 359258 -2854 359494
rect -2770 359258 -2534 359494
rect -2450 359258 -2214 359494
rect -2130 359258 -1894 359494
rect -3090 352258 -2854 352494
rect -2770 352258 -2534 352494
rect -2450 352258 -2214 352494
rect -2130 352258 -1894 352494
rect -3090 345258 -2854 345494
rect -2770 345258 -2534 345494
rect -2450 345258 -2214 345494
rect -2130 345258 -1894 345494
rect -3090 338258 -2854 338494
rect -2770 338258 -2534 338494
rect -2450 338258 -2214 338494
rect -2130 338258 -1894 338494
rect -3090 331258 -2854 331494
rect -2770 331258 -2534 331494
rect -2450 331258 -2214 331494
rect -2130 331258 -1894 331494
rect -3090 324258 -2854 324494
rect -2770 324258 -2534 324494
rect -2450 324258 -2214 324494
rect -2130 324258 -1894 324494
rect -3090 317258 -2854 317494
rect -2770 317258 -2534 317494
rect -2450 317258 -2214 317494
rect -2130 317258 -1894 317494
rect -3090 310258 -2854 310494
rect -2770 310258 -2534 310494
rect -2450 310258 -2214 310494
rect -2130 310258 -1894 310494
rect -3090 303258 -2854 303494
rect -2770 303258 -2534 303494
rect -2450 303258 -2214 303494
rect -2130 303258 -1894 303494
rect -3090 296258 -2854 296494
rect -2770 296258 -2534 296494
rect -2450 296258 -2214 296494
rect -2130 296258 -1894 296494
rect -3090 289258 -2854 289494
rect -2770 289258 -2534 289494
rect -2450 289258 -2214 289494
rect -2130 289258 -1894 289494
rect -3090 282258 -2854 282494
rect -2770 282258 -2534 282494
rect -2450 282258 -2214 282494
rect -2130 282258 -1894 282494
rect -3090 275258 -2854 275494
rect -2770 275258 -2534 275494
rect -2450 275258 -2214 275494
rect -2130 275258 -1894 275494
rect -3090 268258 -2854 268494
rect -2770 268258 -2534 268494
rect -2450 268258 -2214 268494
rect -2130 268258 -1894 268494
rect -3090 261258 -2854 261494
rect -2770 261258 -2534 261494
rect -2450 261258 -2214 261494
rect -2130 261258 -1894 261494
rect -3090 254258 -2854 254494
rect -2770 254258 -2534 254494
rect -2450 254258 -2214 254494
rect -2130 254258 -1894 254494
rect -3090 247258 -2854 247494
rect -2770 247258 -2534 247494
rect -2450 247258 -2214 247494
rect -2130 247258 -1894 247494
rect -3090 240258 -2854 240494
rect -2770 240258 -2534 240494
rect -2450 240258 -2214 240494
rect -2130 240258 -1894 240494
rect -3090 233258 -2854 233494
rect -2770 233258 -2534 233494
rect -2450 233258 -2214 233494
rect -2130 233258 -1894 233494
rect -3090 226258 -2854 226494
rect -2770 226258 -2534 226494
rect -2450 226258 -2214 226494
rect -2130 226258 -1894 226494
rect -3090 219258 -2854 219494
rect -2770 219258 -2534 219494
rect -2450 219258 -2214 219494
rect -2130 219258 -1894 219494
rect -3090 212258 -2854 212494
rect -2770 212258 -2534 212494
rect -2450 212258 -2214 212494
rect -2130 212258 -1894 212494
rect -3090 205258 -2854 205494
rect -2770 205258 -2534 205494
rect -2450 205258 -2214 205494
rect -2130 205258 -1894 205494
rect -3090 198258 -2854 198494
rect -2770 198258 -2534 198494
rect -2450 198258 -2214 198494
rect -2130 198258 -1894 198494
rect -3090 191258 -2854 191494
rect -2770 191258 -2534 191494
rect -2450 191258 -2214 191494
rect -2130 191258 -1894 191494
rect -3090 184258 -2854 184494
rect -2770 184258 -2534 184494
rect -2450 184258 -2214 184494
rect -2130 184258 -1894 184494
rect -3090 177258 -2854 177494
rect -2770 177258 -2534 177494
rect -2450 177258 -2214 177494
rect -2130 177258 -1894 177494
rect -3090 170258 -2854 170494
rect -2770 170258 -2534 170494
rect -2450 170258 -2214 170494
rect -2130 170258 -1894 170494
rect -3090 163258 -2854 163494
rect -2770 163258 -2534 163494
rect -2450 163258 -2214 163494
rect -2130 163258 -1894 163494
rect -3090 156258 -2854 156494
rect -2770 156258 -2534 156494
rect -2450 156258 -2214 156494
rect -2130 156258 -1894 156494
rect -3090 149258 -2854 149494
rect -2770 149258 -2534 149494
rect -2450 149258 -2214 149494
rect -2130 149258 -1894 149494
rect -3090 142258 -2854 142494
rect -2770 142258 -2534 142494
rect -2450 142258 -2214 142494
rect -2130 142258 -1894 142494
rect -3090 135258 -2854 135494
rect -2770 135258 -2534 135494
rect -2450 135258 -2214 135494
rect -2130 135258 -1894 135494
rect -3090 128258 -2854 128494
rect -2770 128258 -2534 128494
rect -2450 128258 -2214 128494
rect -2130 128258 -1894 128494
rect -3090 121258 -2854 121494
rect -2770 121258 -2534 121494
rect -2450 121258 -2214 121494
rect -2130 121258 -1894 121494
rect -3090 114258 -2854 114494
rect -2770 114258 -2534 114494
rect -2450 114258 -2214 114494
rect -2130 114258 -1894 114494
rect -3090 107258 -2854 107494
rect -2770 107258 -2534 107494
rect -2450 107258 -2214 107494
rect -2130 107258 -1894 107494
rect -3090 100258 -2854 100494
rect -2770 100258 -2534 100494
rect -2450 100258 -2214 100494
rect -2130 100258 -1894 100494
rect -3090 93258 -2854 93494
rect -2770 93258 -2534 93494
rect -2450 93258 -2214 93494
rect -2130 93258 -1894 93494
rect -3090 86258 -2854 86494
rect -2770 86258 -2534 86494
rect -2450 86258 -2214 86494
rect -2130 86258 -1894 86494
rect -3090 79258 -2854 79494
rect -2770 79258 -2534 79494
rect -2450 79258 -2214 79494
rect -2130 79258 -1894 79494
rect -3090 72258 -2854 72494
rect -2770 72258 -2534 72494
rect -2450 72258 -2214 72494
rect -2130 72258 -1894 72494
rect -3090 65258 -2854 65494
rect -2770 65258 -2534 65494
rect -2450 65258 -2214 65494
rect -2130 65258 -1894 65494
rect -3090 58258 -2854 58494
rect -2770 58258 -2534 58494
rect -2450 58258 -2214 58494
rect -2130 58258 -1894 58494
rect -3090 51258 -2854 51494
rect -2770 51258 -2534 51494
rect -2450 51258 -2214 51494
rect -2130 51258 -1894 51494
rect -3090 44258 -2854 44494
rect -2770 44258 -2534 44494
rect -2450 44258 -2214 44494
rect -2130 44258 -1894 44494
rect -3090 37258 -2854 37494
rect -2770 37258 -2534 37494
rect -2450 37258 -2214 37494
rect -2130 37258 -1894 37494
rect -3090 30258 -2854 30494
rect -2770 30258 -2534 30494
rect -2450 30258 -2214 30494
rect -2130 30258 -1894 30494
rect -3090 23258 -2854 23494
rect -2770 23258 -2534 23494
rect -2450 23258 -2214 23494
rect -2130 23258 -1894 23494
rect -3090 16258 -2854 16494
rect -2770 16258 -2534 16494
rect -2450 16258 -2214 16494
rect -2130 16258 -1894 16494
rect -3090 9258 -2854 9494
rect -2770 9258 -2534 9494
rect -2450 9258 -2214 9494
rect -2130 9258 -1894 9494
rect -3090 2258 -2854 2494
rect -2770 2258 -2534 2494
rect -2450 2258 -2214 2494
rect -2130 2258 -1894 2494
rect -2374 -982 -2138 -746
rect -2054 -982 -1818 -746
rect -2374 -1302 -2138 -1066
rect -2054 -1302 -1818 -1066
rect 1186 705002 1422 705238
rect 1186 704682 1422 704918
rect 1186 695258 1422 695494
rect 1186 688258 1422 688494
rect 1186 681258 1422 681494
rect 1186 674258 1422 674494
rect 1186 667258 1422 667494
rect 1186 660258 1422 660494
rect 1186 653258 1422 653494
rect 1186 646258 1422 646494
rect 1186 639258 1422 639494
rect 1186 632258 1422 632494
rect 1186 625258 1422 625494
rect 1186 618258 1422 618494
rect 1186 611258 1422 611494
rect 1186 604258 1422 604494
rect 1186 597258 1422 597494
rect 1186 590258 1422 590494
rect 1186 583258 1422 583494
rect 1186 576258 1422 576494
rect 1186 569258 1422 569494
rect 1186 562258 1422 562494
rect 1186 555258 1422 555494
rect 1186 548258 1422 548494
rect 1186 541258 1422 541494
rect 1186 534258 1422 534494
rect 1186 527258 1422 527494
rect 1186 520258 1422 520494
rect 1186 513258 1422 513494
rect 1186 506258 1422 506494
rect 1186 499258 1422 499494
rect 1186 492258 1422 492494
rect 1186 485258 1422 485494
rect 1186 478258 1422 478494
rect 1186 471258 1422 471494
rect 1186 464258 1422 464494
rect 1186 457258 1422 457494
rect 1186 450258 1422 450494
rect 1186 443258 1422 443494
rect 1186 436258 1422 436494
rect 1186 429258 1422 429494
rect 1186 422258 1422 422494
rect 1186 415258 1422 415494
rect 1186 408258 1422 408494
rect 1186 401258 1422 401494
rect 1186 394258 1422 394494
rect 1186 387258 1422 387494
rect 1186 380258 1422 380494
rect 1186 373258 1422 373494
rect 1186 366258 1422 366494
rect 1186 359258 1422 359494
rect 1186 352258 1422 352494
rect 1186 345258 1422 345494
rect 1186 338258 1422 338494
rect 1186 331258 1422 331494
rect 1186 324258 1422 324494
rect 1186 317258 1422 317494
rect 1186 310258 1422 310494
rect 1186 303258 1422 303494
rect 1186 296258 1422 296494
rect 1186 289258 1422 289494
rect 1186 282258 1422 282494
rect 1186 275258 1422 275494
rect 1186 268258 1422 268494
rect 1186 261258 1422 261494
rect 1186 254258 1422 254494
rect 1186 247258 1422 247494
rect 1186 240258 1422 240494
rect 1186 233258 1422 233494
rect 1186 226258 1422 226494
rect 1186 219258 1422 219494
rect 1186 212258 1422 212494
rect 1186 205258 1422 205494
rect 1186 198258 1422 198494
rect 1186 191258 1422 191494
rect 1186 184258 1422 184494
rect 1186 177258 1422 177494
rect 1186 170258 1422 170494
rect 1186 163258 1422 163494
rect 1186 156258 1422 156494
rect 1186 149258 1422 149494
rect 1186 142258 1422 142494
rect 1186 135258 1422 135494
rect 1186 128258 1422 128494
rect 1186 121258 1422 121494
rect 1186 114258 1422 114494
rect 1186 107258 1422 107494
rect 1186 100258 1422 100494
rect 1186 93258 1422 93494
rect 1186 86258 1422 86494
rect 1186 79258 1422 79494
rect 1186 72258 1422 72494
rect 1186 65258 1422 65494
rect 1186 58258 1422 58494
rect 1186 51258 1422 51494
rect 1186 44258 1422 44494
rect 1186 37258 1422 37494
rect 1186 30258 1422 30494
rect 1186 23258 1422 23494
rect 1186 16258 1422 16494
rect 1186 9258 1422 9494
rect 1186 2258 1422 2494
rect 1186 -982 1422 -746
rect 1186 -1302 1422 -1066
rect 2918 705962 3154 706198
rect 2918 705642 3154 705878
rect 2918 696198 3154 696434
rect 2918 689198 3154 689434
rect 2918 682198 3154 682434
rect 2918 675198 3154 675434
rect 2918 668198 3154 668434
rect 2918 661198 3154 661434
rect 2918 654198 3154 654434
rect 2918 647198 3154 647434
rect 2918 640198 3154 640434
rect 2918 633198 3154 633434
rect 2918 626198 3154 626434
rect 2918 619198 3154 619434
rect 2918 612198 3154 612434
rect 2918 605198 3154 605434
rect 2918 598198 3154 598434
rect 2918 591198 3154 591434
rect 2918 584198 3154 584434
rect 2918 577198 3154 577434
rect 2918 570198 3154 570434
rect 2918 563198 3154 563434
rect 2918 556198 3154 556434
rect 2918 549198 3154 549434
rect 2918 542198 3154 542434
rect 2918 535198 3154 535434
rect 2918 528198 3154 528434
rect 2918 521198 3154 521434
rect 2918 514198 3154 514434
rect 2918 507198 3154 507434
rect 2918 500198 3154 500434
rect 2918 493198 3154 493434
rect 2918 486198 3154 486434
rect 2918 479198 3154 479434
rect 2918 472198 3154 472434
rect 2918 465198 3154 465434
rect 2918 458198 3154 458434
rect 2918 451198 3154 451434
rect 2918 444198 3154 444434
rect 2918 437198 3154 437434
rect 2918 430198 3154 430434
rect 2918 423198 3154 423434
rect 2918 416198 3154 416434
rect 2918 409198 3154 409434
rect 2918 402198 3154 402434
rect 2918 395198 3154 395434
rect 2918 388198 3154 388434
rect 2918 381198 3154 381434
rect 2918 374198 3154 374434
rect 2918 367198 3154 367434
rect 2918 360198 3154 360434
rect 2918 353198 3154 353434
rect 2918 346198 3154 346434
rect 2918 339198 3154 339434
rect 2918 332198 3154 332434
rect 2918 325198 3154 325434
rect 2918 318198 3154 318434
rect 2918 311198 3154 311434
rect 2918 304198 3154 304434
rect 2918 297198 3154 297434
rect 2918 290198 3154 290434
rect 2918 283198 3154 283434
rect 2918 276198 3154 276434
rect 2918 269198 3154 269434
rect 2918 262198 3154 262434
rect 2918 255198 3154 255434
rect 2918 248198 3154 248434
rect 2918 241198 3154 241434
rect 2918 234198 3154 234434
rect 2918 227198 3154 227434
rect 2918 220198 3154 220434
rect 2918 213198 3154 213434
rect 2918 206198 3154 206434
rect 2918 199198 3154 199434
rect 2918 192198 3154 192434
rect 2918 185198 3154 185434
rect 2918 178198 3154 178434
rect 2918 171198 3154 171434
rect 2918 164198 3154 164434
rect 2918 157198 3154 157434
rect 2918 150198 3154 150434
rect 2918 143198 3154 143434
rect 2918 136198 3154 136434
rect 2918 129198 3154 129434
rect 2918 122198 3154 122434
rect 2918 115198 3154 115434
rect 2918 108198 3154 108434
rect 2918 101198 3154 101434
rect 2918 94198 3154 94434
rect 2918 87198 3154 87434
rect 2918 80198 3154 80434
rect 2918 73198 3154 73434
rect 2918 66198 3154 66434
rect 2918 59198 3154 59434
rect 2918 52198 3154 52434
rect 2918 45198 3154 45434
rect 2918 38198 3154 38434
rect 2918 31198 3154 31434
rect 2918 24198 3154 24434
rect 2918 17198 3154 17434
rect 2918 10198 3154 10434
rect 2918 3198 3154 3434
rect 2918 -1942 3154 -1706
rect 2918 -2262 3154 -2026
rect 8186 705002 8422 705238
rect 8186 704682 8422 704918
rect 8186 695258 8422 695494
rect 8186 688258 8422 688494
rect 8186 681258 8422 681494
rect 8186 674258 8422 674494
rect 8186 667258 8422 667494
rect 8186 660258 8422 660494
rect 8186 653258 8422 653494
rect 8186 646258 8422 646494
rect 8186 639258 8422 639494
rect 8186 632258 8422 632494
rect 8186 625258 8422 625494
rect 8186 618258 8422 618494
rect 8186 611258 8422 611494
rect 8186 604258 8422 604494
rect 8186 597258 8422 597494
rect 8186 590258 8422 590494
rect 8186 583258 8422 583494
rect 8186 576258 8422 576494
rect 8186 569258 8422 569494
rect 8186 562258 8422 562494
rect 8186 555258 8422 555494
rect 8186 548258 8422 548494
rect 8186 541258 8422 541494
rect 8186 534258 8422 534494
rect 8186 527258 8422 527494
rect 8186 520258 8422 520494
rect 8186 513258 8422 513494
rect 8186 506258 8422 506494
rect 8186 499258 8422 499494
rect 8186 492258 8422 492494
rect 8186 485258 8422 485494
rect 8186 478258 8422 478494
rect 8186 471258 8422 471494
rect 8186 464258 8422 464494
rect 8186 457258 8422 457494
rect 8186 450258 8422 450494
rect 8186 443258 8422 443494
rect 8186 436258 8422 436494
rect 8186 429258 8422 429494
rect 8186 422258 8422 422494
rect 8186 415258 8422 415494
rect 8186 408258 8422 408494
rect 8186 401258 8422 401494
rect 8186 394258 8422 394494
rect 8186 387258 8422 387494
rect 8186 380258 8422 380494
rect 8186 373258 8422 373494
rect 8186 366258 8422 366494
rect 8186 359258 8422 359494
rect 8186 352258 8422 352494
rect 8186 345258 8422 345494
rect 8186 338258 8422 338494
rect 8186 331258 8422 331494
rect 8186 324258 8422 324494
rect 8186 317258 8422 317494
rect 8186 310258 8422 310494
rect 8186 303258 8422 303494
rect 8186 296258 8422 296494
rect 8186 289258 8422 289494
rect 8186 282258 8422 282494
rect 8186 275258 8422 275494
rect 8186 268258 8422 268494
rect 8186 261258 8422 261494
rect 8186 254258 8422 254494
rect 8186 247258 8422 247494
rect 8186 240258 8422 240494
rect 8186 233258 8422 233494
rect 8186 226258 8422 226494
rect 8186 219258 8422 219494
rect 8186 212258 8422 212494
rect 8186 205258 8422 205494
rect 8186 198258 8422 198494
rect 8186 191258 8422 191494
rect 8186 184258 8422 184494
rect 8186 177258 8422 177494
rect 8186 170258 8422 170494
rect 8186 163258 8422 163494
rect 8186 156258 8422 156494
rect 8186 149258 8422 149494
rect 8186 142258 8422 142494
rect 8186 135258 8422 135494
rect 8186 128258 8422 128494
rect 8186 121258 8422 121494
rect 8186 114258 8422 114494
rect 8186 107258 8422 107494
rect 8186 100258 8422 100494
rect 8186 93258 8422 93494
rect 8186 86258 8422 86494
rect 8186 79258 8422 79494
rect 8186 72258 8422 72494
rect 8186 65258 8422 65494
rect 8186 58258 8422 58494
rect 8186 51258 8422 51494
rect 8186 44258 8422 44494
rect 8186 37258 8422 37494
rect 8186 30258 8422 30494
rect 8186 23258 8422 23494
rect 8186 16258 8422 16494
rect 8186 9258 8422 9494
rect 8186 2258 8422 2494
rect 8186 -982 8422 -746
rect 8186 -1302 8422 -1066
rect 9918 705962 10154 706198
rect 9918 705642 10154 705878
rect 9918 696198 10154 696434
rect 9918 689198 10154 689434
rect 9918 682198 10154 682434
rect 9918 675198 10154 675434
rect 9918 668198 10154 668434
rect 9918 661198 10154 661434
rect 9918 654198 10154 654434
rect 9918 647198 10154 647434
rect 9918 640198 10154 640434
rect 9918 633198 10154 633434
rect 9918 626198 10154 626434
rect 9918 619198 10154 619434
rect 9918 612198 10154 612434
rect 9918 605198 10154 605434
rect 9918 598198 10154 598434
rect 9918 591198 10154 591434
rect 9918 584198 10154 584434
rect 9918 577198 10154 577434
rect 9918 570198 10154 570434
rect 9918 563198 10154 563434
rect 9918 556198 10154 556434
rect 9918 549198 10154 549434
rect 9918 542198 10154 542434
rect 9918 535198 10154 535434
rect 9918 528198 10154 528434
rect 9918 521198 10154 521434
rect 9918 514198 10154 514434
rect 9918 507198 10154 507434
rect 9918 500198 10154 500434
rect 9918 493198 10154 493434
rect 9918 486198 10154 486434
rect 9918 479198 10154 479434
rect 9918 472198 10154 472434
rect 9918 465198 10154 465434
rect 9918 458198 10154 458434
rect 9918 451198 10154 451434
rect 9918 444198 10154 444434
rect 9918 437198 10154 437434
rect 9918 430198 10154 430434
rect 9918 423198 10154 423434
rect 9918 416198 10154 416434
rect 9918 409198 10154 409434
rect 9918 402198 10154 402434
rect 9918 395198 10154 395434
rect 9918 388198 10154 388434
rect 9918 381198 10154 381434
rect 9918 374198 10154 374434
rect 9918 367198 10154 367434
rect 9918 360198 10154 360434
rect 9918 353198 10154 353434
rect 9918 346198 10154 346434
rect 9918 339198 10154 339434
rect 9918 332198 10154 332434
rect 9918 325198 10154 325434
rect 9918 318198 10154 318434
rect 9918 311198 10154 311434
rect 9918 304198 10154 304434
rect 9918 297198 10154 297434
rect 9918 290198 10154 290434
rect 9918 283198 10154 283434
rect 9918 276198 10154 276434
rect 9918 269198 10154 269434
rect 9918 262198 10154 262434
rect 9918 255198 10154 255434
rect 9918 248198 10154 248434
rect 9918 241198 10154 241434
rect 9918 234198 10154 234434
rect 9918 227198 10154 227434
rect 9918 220198 10154 220434
rect 9918 213198 10154 213434
rect 9918 206198 10154 206434
rect 9918 199198 10154 199434
rect 9918 192198 10154 192434
rect 9918 185198 10154 185434
rect 9918 178198 10154 178434
rect 9918 171198 10154 171434
rect 9918 164198 10154 164434
rect 9918 157198 10154 157434
rect 9918 150198 10154 150434
rect 9918 143198 10154 143434
rect 9918 136198 10154 136434
rect 9918 129198 10154 129434
rect 9918 122198 10154 122434
rect 9918 115198 10154 115434
rect 9918 108198 10154 108434
rect 9918 101198 10154 101434
rect 9918 94198 10154 94434
rect 9918 87198 10154 87434
rect 9918 80198 10154 80434
rect 9918 73198 10154 73434
rect 9918 66198 10154 66434
rect 9918 59198 10154 59434
rect 9918 52198 10154 52434
rect 9918 45198 10154 45434
rect 9918 38198 10154 38434
rect 9918 31198 10154 31434
rect 9918 24198 10154 24434
rect 9918 17198 10154 17434
rect 9918 10198 10154 10434
rect 9918 3198 10154 3434
rect 9918 -1942 10154 -1706
rect 9918 -2262 10154 -2026
rect 15186 705002 15422 705238
rect 15186 704682 15422 704918
rect 15186 695258 15422 695494
rect 15186 688258 15422 688494
rect 15186 681258 15422 681494
rect 15186 674258 15422 674494
rect 15186 667258 15422 667494
rect 15186 660258 15422 660494
rect 15186 653258 15422 653494
rect 15186 646258 15422 646494
rect 15186 639258 15422 639494
rect 15186 632258 15422 632494
rect 15186 625258 15422 625494
rect 15186 618258 15422 618494
rect 15186 611258 15422 611494
rect 15186 604258 15422 604494
rect 15186 597258 15422 597494
rect 15186 590258 15422 590494
rect 15186 583258 15422 583494
rect 15186 576258 15422 576494
rect 15186 569258 15422 569494
rect 15186 562258 15422 562494
rect 15186 555258 15422 555494
rect 15186 548258 15422 548494
rect 15186 541258 15422 541494
rect 15186 534258 15422 534494
rect 15186 527258 15422 527494
rect 15186 520258 15422 520494
rect 15186 513258 15422 513494
rect 15186 506258 15422 506494
rect 15186 499258 15422 499494
rect 15186 492258 15422 492494
rect 15186 485258 15422 485494
rect 15186 478258 15422 478494
rect 15186 471258 15422 471494
rect 15186 464258 15422 464494
rect 15186 457258 15422 457494
rect 15186 450258 15422 450494
rect 15186 443258 15422 443494
rect 15186 436258 15422 436494
rect 15186 429258 15422 429494
rect 15186 422258 15422 422494
rect 15186 415258 15422 415494
rect 15186 408258 15422 408494
rect 15186 401258 15422 401494
rect 15186 394258 15422 394494
rect 15186 387258 15422 387494
rect 15186 380258 15422 380494
rect 15186 373258 15422 373494
rect 15186 366258 15422 366494
rect 15186 359258 15422 359494
rect 15186 352258 15422 352494
rect 15186 345258 15422 345494
rect 15186 338258 15422 338494
rect 15186 331258 15422 331494
rect 15186 324258 15422 324494
rect 15186 317258 15422 317494
rect 15186 310258 15422 310494
rect 15186 303258 15422 303494
rect 15186 296258 15422 296494
rect 15186 289258 15422 289494
rect 15186 282258 15422 282494
rect 15186 275258 15422 275494
rect 15186 268258 15422 268494
rect 15186 261258 15422 261494
rect 15186 254258 15422 254494
rect 15186 247258 15422 247494
rect 15186 240258 15422 240494
rect 15186 233258 15422 233494
rect 15186 226258 15422 226494
rect 15186 219258 15422 219494
rect 15186 212258 15422 212494
rect 15186 205258 15422 205494
rect 15186 198258 15422 198494
rect 15186 191258 15422 191494
rect 15186 184258 15422 184494
rect 15186 177258 15422 177494
rect 15186 170258 15422 170494
rect 15186 163258 15422 163494
rect 15186 156258 15422 156494
rect 15186 149258 15422 149494
rect 15186 142258 15422 142494
rect 15186 135258 15422 135494
rect 15186 128258 15422 128494
rect 15186 121258 15422 121494
rect 15186 114258 15422 114494
rect 15186 107258 15422 107494
rect 15186 100258 15422 100494
rect 15186 93258 15422 93494
rect 15186 86258 15422 86494
rect 15186 79258 15422 79494
rect 15186 72258 15422 72494
rect 15186 65258 15422 65494
rect 15186 58258 15422 58494
rect 15186 51258 15422 51494
rect 15186 44258 15422 44494
rect 15186 37258 15422 37494
rect 15186 30258 15422 30494
rect 15186 23258 15422 23494
rect 15186 16258 15422 16494
rect 15186 9258 15422 9494
rect 15186 2258 15422 2494
rect 15186 -982 15422 -746
rect 15186 -1302 15422 -1066
rect 16918 705962 17154 706198
rect 16918 705642 17154 705878
rect 16918 696198 17154 696434
rect 16918 689198 17154 689434
rect 16918 682198 17154 682434
rect 16918 675198 17154 675434
rect 16918 668198 17154 668434
rect 16918 661198 17154 661434
rect 16918 654198 17154 654434
rect 16918 647198 17154 647434
rect 16918 640198 17154 640434
rect 16918 633198 17154 633434
rect 16918 626198 17154 626434
rect 16918 619198 17154 619434
rect 16918 612198 17154 612434
rect 16918 605198 17154 605434
rect 16918 598198 17154 598434
rect 16918 591198 17154 591434
rect 16918 584198 17154 584434
rect 16918 577198 17154 577434
rect 16918 570198 17154 570434
rect 16918 563198 17154 563434
rect 16918 556198 17154 556434
rect 16918 549198 17154 549434
rect 16918 542198 17154 542434
rect 16918 535198 17154 535434
rect 16918 528198 17154 528434
rect 16918 521198 17154 521434
rect 16918 514198 17154 514434
rect 16918 507198 17154 507434
rect 16918 500198 17154 500434
rect 16918 493198 17154 493434
rect 16918 486198 17154 486434
rect 16918 479198 17154 479434
rect 16918 472198 17154 472434
rect 16918 465198 17154 465434
rect 16918 458198 17154 458434
rect 16918 451198 17154 451434
rect 16918 444198 17154 444434
rect 16918 437198 17154 437434
rect 16918 430198 17154 430434
rect 16918 423198 17154 423434
rect 16918 416198 17154 416434
rect 16918 409198 17154 409434
rect 16918 402198 17154 402434
rect 16918 395198 17154 395434
rect 16918 388198 17154 388434
rect 16918 381198 17154 381434
rect 16918 374198 17154 374434
rect 16918 367198 17154 367434
rect 16918 360198 17154 360434
rect 16918 353198 17154 353434
rect 16918 346198 17154 346434
rect 16918 339198 17154 339434
rect 16918 332198 17154 332434
rect 16918 325198 17154 325434
rect 16918 318198 17154 318434
rect 16918 311198 17154 311434
rect 16918 304198 17154 304434
rect 16918 297198 17154 297434
rect 16918 290198 17154 290434
rect 16918 283198 17154 283434
rect 16918 276198 17154 276434
rect 16918 269198 17154 269434
rect 16918 262198 17154 262434
rect 16918 255198 17154 255434
rect 16918 248198 17154 248434
rect 16918 241198 17154 241434
rect 16918 234198 17154 234434
rect 16918 227198 17154 227434
rect 16918 220198 17154 220434
rect 16918 213198 17154 213434
rect 16918 206198 17154 206434
rect 16918 199198 17154 199434
rect 16918 192198 17154 192434
rect 16918 185198 17154 185434
rect 16918 178198 17154 178434
rect 16918 171198 17154 171434
rect 16918 164198 17154 164434
rect 16918 157198 17154 157434
rect 16918 150198 17154 150434
rect 16918 143198 17154 143434
rect 16918 136198 17154 136434
rect 16918 129198 17154 129434
rect 16918 122198 17154 122434
rect 16918 115198 17154 115434
rect 16918 108198 17154 108434
rect 16918 101198 17154 101434
rect 16918 94198 17154 94434
rect 16918 87198 17154 87434
rect 16918 80198 17154 80434
rect 16918 73198 17154 73434
rect 16918 66198 17154 66434
rect 16918 59198 17154 59434
rect 16918 52198 17154 52434
rect 16918 45198 17154 45434
rect 16918 38198 17154 38434
rect 16918 31198 17154 31434
rect 16918 24198 17154 24434
rect 16918 17198 17154 17434
rect 16918 10198 17154 10434
rect 16918 3198 17154 3434
rect 16918 -1942 17154 -1706
rect 16918 -2262 17154 -2026
rect 22186 705002 22422 705238
rect 22186 704682 22422 704918
rect 22186 695258 22422 695494
rect 22186 688258 22422 688494
rect 22186 681258 22422 681494
rect 22186 674258 22422 674494
rect 22186 667258 22422 667494
rect 22186 660258 22422 660494
rect 22186 653258 22422 653494
rect 22186 646258 22422 646494
rect 22186 639258 22422 639494
rect 22186 632258 22422 632494
rect 22186 625258 22422 625494
rect 22186 618258 22422 618494
rect 22186 611258 22422 611494
rect 22186 604258 22422 604494
rect 22186 597258 22422 597494
rect 22186 590258 22422 590494
rect 22186 583258 22422 583494
rect 22186 576258 22422 576494
rect 22186 569258 22422 569494
rect 22186 562258 22422 562494
rect 22186 555258 22422 555494
rect 22186 548258 22422 548494
rect 22186 541258 22422 541494
rect 22186 534258 22422 534494
rect 22186 527258 22422 527494
rect 22186 520258 22422 520494
rect 22186 513258 22422 513494
rect 22186 506258 22422 506494
rect 22186 499258 22422 499494
rect 22186 492258 22422 492494
rect 22186 485258 22422 485494
rect 22186 478258 22422 478494
rect 22186 471258 22422 471494
rect 22186 464258 22422 464494
rect 22186 457258 22422 457494
rect 22186 450258 22422 450494
rect 22186 443258 22422 443494
rect 22186 436258 22422 436494
rect 22186 429258 22422 429494
rect 22186 422258 22422 422494
rect 22186 415258 22422 415494
rect 22186 408258 22422 408494
rect 22186 401258 22422 401494
rect 22186 394258 22422 394494
rect 22186 387258 22422 387494
rect 22186 380258 22422 380494
rect 22186 373258 22422 373494
rect 22186 366258 22422 366494
rect 22186 359258 22422 359494
rect 22186 352258 22422 352494
rect 22186 345258 22422 345494
rect 22186 338258 22422 338494
rect 22186 331258 22422 331494
rect 22186 324258 22422 324494
rect 22186 317258 22422 317494
rect 22186 310258 22422 310494
rect 22186 303258 22422 303494
rect 22186 296258 22422 296494
rect 22186 289258 22422 289494
rect 22186 282258 22422 282494
rect 22186 275258 22422 275494
rect 22186 268258 22422 268494
rect 22186 261258 22422 261494
rect 22186 254258 22422 254494
rect 22186 247258 22422 247494
rect 22186 240258 22422 240494
rect 22186 233258 22422 233494
rect 22186 226258 22422 226494
rect 22186 219258 22422 219494
rect 22186 212258 22422 212494
rect 22186 205258 22422 205494
rect 22186 198258 22422 198494
rect 22186 191258 22422 191494
rect 22186 184258 22422 184494
rect 22186 177258 22422 177494
rect 22186 170258 22422 170494
rect 22186 163258 22422 163494
rect 22186 156258 22422 156494
rect 22186 149258 22422 149494
rect 22186 142258 22422 142494
rect 22186 135258 22422 135494
rect 22186 128258 22422 128494
rect 22186 121258 22422 121494
rect 22186 114258 22422 114494
rect 22186 107258 22422 107494
rect 22186 100258 22422 100494
rect 22186 93258 22422 93494
rect 22186 86258 22422 86494
rect 22186 79258 22422 79494
rect 22186 72258 22422 72494
rect 22186 65258 22422 65494
rect 22186 58258 22422 58494
rect 22186 51258 22422 51494
rect 22186 44258 22422 44494
rect 22186 37258 22422 37494
rect 22186 30258 22422 30494
rect 22186 23258 22422 23494
rect 22186 16258 22422 16494
rect 22186 9258 22422 9494
rect 22186 2258 22422 2494
rect 22186 -982 22422 -746
rect 22186 -1302 22422 -1066
rect 23918 705962 24154 706198
rect 23918 705642 24154 705878
rect 23918 696198 24154 696434
rect 23918 689198 24154 689434
rect 23918 682198 24154 682434
rect 23918 675198 24154 675434
rect 23918 668198 24154 668434
rect 23918 661198 24154 661434
rect 23918 654198 24154 654434
rect 23918 647198 24154 647434
rect 23918 640198 24154 640434
rect 23918 633198 24154 633434
rect 23918 626198 24154 626434
rect 23918 619198 24154 619434
rect 23918 612198 24154 612434
rect 23918 605198 24154 605434
rect 23918 598198 24154 598434
rect 23918 591198 24154 591434
rect 23918 584198 24154 584434
rect 23918 577198 24154 577434
rect 23918 570198 24154 570434
rect 23918 563198 24154 563434
rect 23918 556198 24154 556434
rect 23918 549198 24154 549434
rect 23918 542198 24154 542434
rect 23918 535198 24154 535434
rect 23918 528198 24154 528434
rect 23918 521198 24154 521434
rect 23918 514198 24154 514434
rect 23918 507198 24154 507434
rect 23918 500198 24154 500434
rect 23918 493198 24154 493434
rect 23918 486198 24154 486434
rect 23918 479198 24154 479434
rect 23918 472198 24154 472434
rect 23918 465198 24154 465434
rect 23918 458198 24154 458434
rect 23918 451198 24154 451434
rect 23918 444198 24154 444434
rect 23918 437198 24154 437434
rect 23918 430198 24154 430434
rect 23918 423198 24154 423434
rect 23918 416198 24154 416434
rect 23918 409198 24154 409434
rect 23918 402198 24154 402434
rect 23918 395198 24154 395434
rect 23918 388198 24154 388434
rect 23918 381198 24154 381434
rect 23918 374198 24154 374434
rect 23918 367198 24154 367434
rect 23918 360198 24154 360434
rect 23918 353198 24154 353434
rect 23918 346198 24154 346434
rect 23918 339198 24154 339434
rect 23918 332198 24154 332434
rect 23918 325198 24154 325434
rect 23918 318198 24154 318434
rect 23918 311198 24154 311434
rect 23918 304198 24154 304434
rect 23918 297198 24154 297434
rect 23918 290198 24154 290434
rect 23918 283198 24154 283434
rect 23918 276198 24154 276434
rect 23918 269198 24154 269434
rect 23918 262198 24154 262434
rect 23918 255198 24154 255434
rect 23918 248198 24154 248434
rect 23918 241198 24154 241434
rect 23918 234198 24154 234434
rect 23918 227198 24154 227434
rect 23918 220198 24154 220434
rect 23918 213198 24154 213434
rect 23918 206198 24154 206434
rect 23918 199198 24154 199434
rect 23918 192198 24154 192434
rect 23918 185198 24154 185434
rect 23918 178198 24154 178434
rect 23918 171198 24154 171434
rect 23918 164198 24154 164434
rect 23918 157198 24154 157434
rect 23918 150198 24154 150434
rect 23918 143198 24154 143434
rect 23918 136198 24154 136434
rect 23918 129198 24154 129434
rect 23918 122198 24154 122434
rect 23918 115198 24154 115434
rect 23918 108198 24154 108434
rect 23918 101198 24154 101434
rect 23918 94198 24154 94434
rect 23918 87198 24154 87434
rect 23918 80198 24154 80434
rect 23918 73198 24154 73434
rect 23918 66198 24154 66434
rect 23918 59198 24154 59434
rect 23918 52198 24154 52434
rect 23918 45198 24154 45434
rect 23918 38198 24154 38434
rect 23918 31198 24154 31434
rect 23918 24198 24154 24434
rect 23918 17198 24154 17434
rect 23918 10198 24154 10434
rect 23918 3198 24154 3434
rect 23918 -1942 24154 -1706
rect 23918 -2262 24154 -2026
rect 29186 705002 29422 705238
rect 29186 704682 29422 704918
rect 29186 695258 29422 695494
rect 29186 688258 29422 688494
rect 29186 681258 29422 681494
rect 29186 674258 29422 674494
rect 29186 667258 29422 667494
rect 29186 660258 29422 660494
rect 29186 653258 29422 653494
rect 29186 646258 29422 646494
rect 29186 639258 29422 639494
rect 29186 632258 29422 632494
rect 29186 625258 29422 625494
rect 29186 618258 29422 618494
rect 29186 611258 29422 611494
rect 29186 604258 29422 604494
rect 29186 597258 29422 597494
rect 29186 590258 29422 590494
rect 29186 583258 29422 583494
rect 29186 576258 29422 576494
rect 29186 569258 29422 569494
rect 29186 562258 29422 562494
rect 29186 555258 29422 555494
rect 29186 548258 29422 548494
rect 29186 541258 29422 541494
rect 29186 534258 29422 534494
rect 29186 527258 29422 527494
rect 29186 520258 29422 520494
rect 29186 513258 29422 513494
rect 29186 506258 29422 506494
rect 29186 499258 29422 499494
rect 29186 492258 29422 492494
rect 29186 485258 29422 485494
rect 29186 478258 29422 478494
rect 29186 471258 29422 471494
rect 29186 464258 29422 464494
rect 29186 457258 29422 457494
rect 29186 450258 29422 450494
rect 29186 443258 29422 443494
rect 29186 436258 29422 436494
rect 29186 429258 29422 429494
rect 29186 422258 29422 422494
rect 29186 415258 29422 415494
rect 29186 408258 29422 408494
rect 29186 401258 29422 401494
rect 29186 394258 29422 394494
rect 29186 387258 29422 387494
rect 29186 380258 29422 380494
rect 29186 373258 29422 373494
rect 29186 366258 29422 366494
rect 29186 359258 29422 359494
rect 29186 352258 29422 352494
rect 29186 345258 29422 345494
rect 29186 338258 29422 338494
rect 29186 331258 29422 331494
rect 29186 324258 29422 324494
rect 29186 317258 29422 317494
rect 29186 310258 29422 310494
rect 29186 303258 29422 303494
rect 29186 296258 29422 296494
rect 29186 289258 29422 289494
rect 29186 282258 29422 282494
rect 29186 275258 29422 275494
rect 29186 268258 29422 268494
rect 29186 261258 29422 261494
rect 29186 254258 29422 254494
rect 29186 247258 29422 247494
rect 29186 240258 29422 240494
rect 29186 233258 29422 233494
rect 29186 226258 29422 226494
rect 29186 219258 29422 219494
rect 29186 212258 29422 212494
rect 29186 205258 29422 205494
rect 29186 198258 29422 198494
rect 29186 191258 29422 191494
rect 29186 184258 29422 184494
rect 29186 177258 29422 177494
rect 29186 170258 29422 170494
rect 29186 163258 29422 163494
rect 29186 156258 29422 156494
rect 29186 149258 29422 149494
rect 29186 142258 29422 142494
rect 29186 135258 29422 135494
rect 29186 128258 29422 128494
rect 29186 121258 29422 121494
rect 29186 114258 29422 114494
rect 29186 107258 29422 107494
rect 29186 100258 29422 100494
rect 29186 93258 29422 93494
rect 29186 86258 29422 86494
rect 29186 79258 29422 79494
rect 29186 72258 29422 72494
rect 29186 65258 29422 65494
rect 29186 58258 29422 58494
rect 29186 51258 29422 51494
rect 29186 44258 29422 44494
rect 29186 37258 29422 37494
rect 29186 30258 29422 30494
rect 29186 23258 29422 23494
rect 29186 16258 29422 16494
rect 29186 9258 29422 9494
rect 29186 2258 29422 2494
rect 29186 -982 29422 -746
rect 29186 -1302 29422 -1066
rect 30918 705962 31154 706198
rect 30918 705642 31154 705878
rect 30918 696198 31154 696434
rect 30918 689198 31154 689434
rect 30918 682198 31154 682434
rect 30918 675198 31154 675434
rect 30918 668198 31154 668434
rect 30918 661198 31154 661434
rect 30918 654198 31154 654434
rect 30918 647198 31154 647434
rect 30918 640198 31154 640434
rect 30918 633198 31154 633434
rect 30918 626198 31154 626434
rect 30918 619198 31154 619434
rect 30918 612198 31154 612434
rect 30918 605198 31154 605434
rect 30918 598198 31154 598434
rect 30918 591198 31154 591434
rect 30918 584198 31154 584434
rect 30918 577198 31154 577434
rect 30918 570198 31154 570434
rect 30918 563198 31154 563434
rect 30918 556198 31154 556434
rect 30918 549198 31154 549434
rect 30918 542198 31154 542434
rect 30918 535198 31154 535434
rect 30918 528198 31154 528434
rect 30918 521198 31154 521434
rect 30918 514198 31154 514434
rect 30918 507198 31154 507434
rect 30918 500198 31154 500434
rect 30918 493198 31154 493434
rect 30918 486198 31154 486434
rect 30918 479198 31154 479434
rect 30918 472198 31154 472434
rect 30918 465198 31154 465434
rect 30918 458198 31154 458434
rect 30918 451198 31154 451434
rect 30918 444198 31154 444434
rect 30918 437198 31154 437434
rect 30918 430198 31154 430434
rect 30918 423198 31154 423434
rect 30918 416198 31154 416434
rect 30918 409198 31154 409434
rect 30918 402198 31154 402434
rect 30918 395198 31154 395434
rect 30918 388198 31154 388434
rect 30918 381198 31154 381434
rect 30918 374198 31154 374434
rect 30918 367198 31154 367434
rect 30918 360198 31154 360434
rect 30918 353198 31154 353434
rect 30918 346198 31154 346434
rect 30918 339198 31154 339434
rect 30918 332198 31154 332434
rect 30918 325198 31154 325434
rect 30918 318198 31154 318434
rect 30918 311198 31154 311434
rect 30918 304198 31154 304434
rect 30918 297198 31154 297434
rect 30918 290198 31154 290434
rect 30918 283198 31154 283434
rect 30918 276198 31154 276434
rect 30918 269198 31154 269434
rect 30918 262198 31154 262434
rect 30918 255198 31154 255434
rect 30918 248198 31154 248434
rect 30918 241198 31154 241434
rect 30918 234198 31154 234434
rect 30918 227198 31154 227434
rect 30918 220198 31154 220434
rect 30918 213198 31154 213434
rect 30918 206198 31154 206434
rect 30918 199198 31154 199434
rect 30918 192198 31154 192434
rect 30918 185198 31154 185434
rect 30918 178198 31154 178434
rect 30918 171198 31154 171434
rect 30918 164198 31154 164434
rect 30918 157198 31154 157434
rect 30918 150198 31154 150434
rect 30918 143198 31154 143434
rect 30918 136198 31154 136434
rect 30918 129198 31154 129434
rect 30918 122198 31154 122434
rect 30918 115198 31154 115434
rect 30918 108198 31154 108434
rect 30918 101198 31154 101434
rect 30918 94198 31154 94434
rect 30918 87198 31154 87434
rect 30918 80198 31154 80434
rect 30918 73198 31154 73434
rect 30918 66198 31154 66434
rect 30918 59198 31154 59434
rect 30918 52198 31154 52434
rect 30918 45198 31154 45434
rect 30918 38198 31154 38434
rect 30918 31198 31154 31434
rect 30918 24198 31154 24434
rect 30918 17198 31154 17434
rect 30918 10198 31154 10434
rect 30918 3198 31154 3434
rect 30918 -1942 31154 -1706
rect 30918 -2262 31154 -2026
rect 36186 705002 36422 705238
rect 36186 704682 36422 704918
rect 36186 695258 36422 695494
rect 36186 688258 36422 688494
rect 36186 681258 36422 681494
rect 36186 674258 36422 674494
rect 36186 667258 36422 667494
rect 36186 660258 36422 660494
rect 36186 653258 36422 653494
rect 36186 646258 36422 646494
rect 36186 639258 36422 639494
rect 36186 632258 36422 632494
rect 36186 625258 36422 625494
rect 36186 618258 36422 618494
rect 36186 611258 36422 611494
rect 36186 604258 36422 604494
rect 36186 597258 36422 597494
rect 36186 590258 36422 590494
rect 36186 583258 36422 583494
rect 36186 576258 36422 576494
rect 36186 569258 36422 569494
rect 36186 562258 36422 562494
rect 36186 555258 36422 555494
rect 36186 548258 36422 548494
rect 36186 541258 36422 541494
rect 36186 534258 36422 534494
rect 36186 527258 36422 527494
rect 36186 520258 36422 520494
rect 36186 513258 36422 513494
rect 36186 506258 36422 506494
rect 36186 499258 36422 499494
rect 36186 492258 36422 492494
rect 36186 485258 36422 485494
rect 36186 478258 36422 478494
rect 36186 471258 36422 471494
rect 36186 464258 36422 464494
rect 36186 457258 36422 457494
rect 36186 450258 36422 450494
rect 36186 443258 36422 443494
rect 36186 436258 36422 436494
rect 36186 429258 36422 429494
rect 36186 422258 36422 422494
rect 36186 415258 36422 415494
rect 36186 408258 36422 408494
rect 36186 401258 36422 401494
rect 36186 394258 36422 394494
rect 36186 387258 36422 387494
rect 36186 380258 36422 380494
rect 36186 373258 36422 373494
rect 36186 366258 36422 366494
rect 36186 359258 36422 359494
rect 36186 352258 36422 352494
rect 36186 345258 36422 345494
rect 36186 338258 36422 338494
rect 36186 331258 36422 331494
rect 36186 324258 36422 324494
rect 36186 317258 36422 317494
rect 36186 310258 36422 310494
rect 36186 303258 36422 303494
rect 36186 296258 36422 296494
rect 36186 289258 36422 289494
rect 36186 282258 36422 282494
rect 36186 275258 36422 275494
rect 36186 268258 36422 268494
rect 36186 261258 36422 261494
rect 36186 254258 36422 254494
rect 36186 247258 36422 247494
rect 36186 240258 36422 240494
rect 36186 233258 36422 233494
rect 36186 226258 36422 226494
rect 36186 219258 36422 219494
rect 36186 212258 36422 212494
rect 36186 205258 36422 205494
rect 36186 198258 36422 198494
rect 36186 191258 36422 191494
rect 36186 184258 36422 184494
rect 36186 177258 36422 177494
rect 36186 170258 36422 170494
rect 36186 163258 36422 163494
rect 36186 156258 36422 156494
rect 36186 149258 36422 149494
rect 36186 142258 36422 142494
rect 36186 135258 36422 135494
rect 36186 128258 36422 128494
rect 36186 121258 36422 121494
rect 36186 114258 36422 114494
rect 36186 107258 36422 107494
rect 36186 100258 36422 100494
rect 36186 93258 36422 93494
rect 36186 86258 36422 86494
rect 36186 79258 36422 79494
rect 36186 72258 36422 72494
rect 36186 65258 36422 65494
rect 36186 58258 36422 58494
rect 36186 51258 36422 51494
rect 36186 44258 36422 44494
rect 36186 37258 36422 37494
rect 36186 30258 36422 30494
rect 36186 23258 36422 23494
rect 36186 16258 36422 16494
rect 36186 9258 36422 9494
rect 36186 2258 36422 2494
rect 36186 -982 36422 -746
rect 36186 -1302 36422 -1066
rect 37918 705962 38154 706198
rect 37918 705642 38154 705878
rect 37918 696198 38154 696434
rect 37918 689198 38154 689434
rect 37918 682198 38154 682434
rect 37918 675198 38154 675434
rect 37918 668198 38154 668434
rect 37918 661198 38154 661434
rect 37918 654198 38154 654434
rect 37918 647198 38154 647434
rect 37918 640198 38154 640434
rect 37918 633198 38154 633434
rect 37918 626198 38154 626434
rect 37918 619198 38154 619434
rect 37918 612198 38154 612434
rect 37918 605198 38154 605434
rect 37918 598198 38154 598434
rect 37918 591198 38154 591434
rect 37918 584198 38154 584434
rect 37918 577198 38154 577434
rect 37918 570198 38154 570434
rect 37918 563198 38154 563434
rect 37918 556198 38154 556434
rect 37918 549198 38154 549434
rect 37918 542198 38154 542434
rect 37918 535198 38154 535434
rect 37918 528198 38154 528434
rect 37918 521198 38154 521434
rect 37918 514198 38154 514434
rect 37918 507198 38154 507434
rect 37918 500198 38154 500434
rect 37918 493198 38154 493434
rect 37918 486198 38154 486434
rect 37918 479198 38154 479434
rect 37918 472198 38154 472434
rect 37918 465198 38154 465434
rect 37918 458198 38154 458434
rect 37918 451198 38154 451434
rect 37918 444198 38154 444434
rect 37918 437198 38154 437434
rect 37918 430198 38154 430434
rect 37918 423198 38154 423434
rect 37918 416198 38154 416434
rect 37918 409198 38154 409434
rect 37918 402198 38154 402434
rect 37918 395198 38154 395434
rect 37918 388198 38154 388434
rect 37918 381198 38154 381434
rect 37918 374198 38154 374434
rect 37918 367198 38154 367434
rect 37918 360198 38154 360434
rect 37918 353198 38154 353434
rect 37918 346198 38154 346434
rect 37918 339198 38154 339434
rect 37918 332198 38154 332434
rect 37918 325198 38154 325434
rect 37918 318198 38154 318434
rect 37918 311198 38154 311434
rect 37918 304198 38154 304434
rect 37918 297198 38154 297434
rect 37918 290198 38154 290434
rect 37918 283198 38154 283434
rect 37918 276198 38154 276434
rect 37918 269198 38154 269434
rect 37918 262198 38154 262434
rect 37918 255198 38154 255434
rect 37918 248198 38154 248434
rect 37918 241198 38154 241434
rect 37918 234198 38154 234434
rect 37918 227198 38154 227434
rect 37918 220198 38154 220434
rect 37918 213198 38154 213434
rect 37918 206198 38154 206434
rect 37918 199198 38154 199434
rect 37918 192198 38154 192434
rect 37918 185198 38154 185434
rect 37918 178198 38154 178434
rect 37918 171198 38154 171434
rect 37918 164198 38154 164434
rect 37918 157198 38154 157434
rect 37918 150198 38154 150434
rect 37918 143198 38154 143434
rect 37918 136198 38154 136434
rect 37918 129198 38154 129434
rect 37918 122198 38154 122434
rect 37918 115198 38154 115434
rect 37918 108198 38154 108434
rect 37918 101198 38154 101434
rect 37918 94198 38154 94434
rect 37918 87198 38154 87434
rect 37918 80198 38154 80434
rect 37918 73198 38154 73434
rect 37918 66198 38154 66434
rect 37918 59198 38154 59434
rect 37918 52198 38154 52434
rect 37918 45198 38154 45434
rect 37918 38198 38154 38434
rect 37918 31198 38154 31434
rect 37918 24198 38154 24434
rect 37918 17198 38154 17434
rect 37918 10198 38154 10434
rect 37918 3198 38154 3434
rect 37918 -1942 38154 -1706
rect 37918 -2262 38154 -2026
rect 43186 705002 43422 705238
rect 43186 704682 43422 704918
rect 43186 695258 43422 695494
rect 43186 688258 43422 688494
rect 43186 681258 43422 681494
rect 43186 674258 43422 674494
rect 43186 667258 43422 667494
rect 43186 660258 43422 660494
rect 43186 653258 43422 653494
rect 43186 646258 43422 646494
rect 43186 639258 43422 639494
rect 43186 632258 43422 632494
rect 43186 625258 43422 625494
rect 43186 618258 43422 618494
rect 43186 611258 43422 611494
rect 43186 604258 43422 604494
rect 43186 597258 43422 597494
rect 43186 590258 43422 590494
rect 43186 583258 43422 583494
rect 43186 576258 43422 576494
rect 43186 569258 43422 569494
rect 43186 562258 43422 562494
rect 43186 555258 43422 555494
rect 43186 548258 43422 548494
rect 43186 541258 43422 541494
rect 43186 534258 43422 534494
rect 43186 527258 43422 527494
rect 43186 520258 43422 520494
rect 43186 513258 43422 513494
rect 43186 506258 43422 506494
rect 43186 499258 43422 499494
rect 43186 492258 43422 492494
rect 43186 485258 43422 485494
rect 43186 478258 43422 478494
rect 43186 471258 43422 471494
rect 43186 464258 43422 464494
rect 43186 457258 43422 457494
rect 43186 450258 43422 450494
rect 43186 443258 43422 443494
rect 43186 436258 43422 436494
rect 43186 429258 43422 429494
rect 43186 422258 43422 422494
rect 43186 415258 43422 415494
rect 43186 408258 43422 408494
rect 43186 401258 43422 401494
rect 43186 394258 43422 394494
rect 43186 387258 43422 387494
rect 43186 380258 43422 380494
rect 43186 373258 43422 373494
rect 43186 366258 43422 366494
rect 43186 359258 43422 359494
rect 43186 352258 43422 352494
rect 43186 345258 43422 345494
rect 43186 338258 43422 338494
rect 43186 331258 43422 331494
rect 43186 324258 43422 324494
rect 43186 317258 43422 317494
rect 43186 310258 43422 310494
rect 43186 303258 43422 303494
rect 43186 296258 43422 296494
rect 43186 289258 43422 289494
rect 43186 282258 43422 282494
rect 43186 275258 43422 275494
rect 43186 268258 43422 268494
rect 43186 261258 43422 261494
rect 43186 254258 43422 254494
rect 43186 247258 43422 247494
rect 43186 240258 43422 240494
rect 43186 233258 43422 233494
rect 43186 226258 43422 226494
rect 43186 219258 43422 219494
rect 43186 212258 43422 212494
rect 43186 205258 43422 205494
rect 43186 198258 43422 198494
rect 43186 191258 43422 191494
rect 43186 184258 43422 184494
rect 43186 177258 43422 177494
rect 43186 170258 43422 170494
rect 43186 163258 43422 163494
rect 43186 156258 43422 156494
rect 43186 149258 43422 149494
rect 43186 142258 43422 142494
rect 43186 135258 43422 135494
rect 43186 128258 43422 128494
rect 43186 121258 43422 121494
rect 43186 114258 43422 114494
rect 43186 107258 43422 107494
rect 43186 100258 43422 100494
rect 43186 93258 43422 93494
rect 43186 86258 43422 86494
rect 43186 79258 43422 79494
rect 43186 72258 43422 72494
rect 43186 65258 43422 65494
rect 43186 58258 43422 58494
rect 43186 51258 43422 51494
rect 43186 44258 43422 44494
rect 43186 37258 43422 37494
rect 43186 30258 43422 30494
rect 43186 23258 43422 23494
rect 43186 16258 43422 16494
rect 43186 9258 43422 9494
rect 43186 2258 43422 2494
rect 43186 -982 43422 -746
rect 43186 -1302 43422 -1066
rect 44918 705962 45154 706198
rect 44918 705642 45154 705878
rect 44918 696198 45154 696434
rect 44918 689198 45154 689434
rect 44918 682198 45154 682434
rect 44918 675198 45154 675434
rect 44918 668198 45154 668434
rect 44918 661198 45154 661434
rect 44918 654198 45154 654434
rect 44918 647198 45154 647434
rect 44918 640198 45154 640434
rect 44918 633198 45154 633434
rect 44918 626198 45154 626434
rect 44918 619198 45154 619434
rect 44918 612198 45154 612434
rect 44918 605198 45154 605434
rect 44918 598198 45154 598434
rect 44918 591198 45154 591434
rect 44918 584198 45154 584434
rect 44918 577198 45154 577434
rect 44918 570198 45154 570434
rect 44918 563198 45154 563434
rect 44918 556198 45154 556434
rect 44918 549198 45154 549434
rect 44918 542198 45154 542434
rect 44918 535198 45154 535434
rect 44918 528198 45154 528434
rect 44918 521198 45154 521434
rect 44918 514198 45154 514434
rect 44918 507198 45154 507434
rect 44918 500198 45154 500434
rect 44918 493198 45154 493434
rect 44918 486198 45154 486434
rect 44918 479198 45154 479434
rect 44918 472198 45154 472434
rect 44918 465198 45154 465434
rect 44918 458198 45154 458434
rect 44918 451198 45154 451434
rect 44918 444198 45154 444434
rect 44918 437198 45154 437434
rect 44918 430198 45154 430434
rect 44918 423198 45154 423434
rect 44918 416198 45154 416434
rect 44918 409198 45154 409434
rect 44918 402198 45154 402434
rect 44918 395198 45154 395434
rect 44918 388198 45154 388434
rect 44918 381198 45154 381434
rect 44918 374198 45154 374434
rect 44918 367198 45154 367434
rect 44918 360198 45154 360434
rect 44918 353198 45154 353434
rect 44918 346198 45154 346434
rect 44918 339198 45154 339434
rect 44918 332198 45154 332434
rect 44918 325198 45154 325434
rect 44918 318198 45154 318434
rect 44918 311198 45154 311434
rect 44918 304198 45154 304434
rect 44918 297198 45154 297434
rect 44918 290198 45154 290434
rect 44918 283198 45154 283434
rect 44918 276198 45154 276434
rect 44918 269198 45154 269434
rect 44918 262198 45154 262434
rect 44918 255198 45154 255434
rect 44918 248198 45154 248434
rect 44918 241198 45154 241434
rect 44918 234198 45154 234434
rect 44918 227198 45154 227434
rect 44918 220198 45154 220434
rect 44918 213198 45154 213434
rect 44918 206198 45154 206434
rect 44918 199198 45154 199434
rect 44918 192198 45154 192434
rect 44918 185198 45154 185434
rect 44918 178198 45154 178434
rect 44918 171198 45154 171434
rect 44918 164198 45154 164434
rect 44918 157198 45154 157434
rect 44918 150198 45154 150434
rect 44918 143198 45154 143434
rect 44918 136198 45154 136434
rect 44918 129198 45154 129434
rect 44918 122198 45154 122434
rect 44918 115198 45154 115434
rect 44918 108198 45154 108434
rect 44918 101198 45154 101434
rect 44918 94198 45154 94434
rect 44918 87198 45154 87434
rect 44918 80198 45154 80434
rect 44918 73198 45154 73434
rect 44918 66198 45154 66434
rect 44918 59198 45154 59434
rect 44918 52198 45154 52434
rect 44918 45198 45154 45434
rect 44918 38198 45154 38434
rect 44918 31198 45154 31434
rect 44918 24198 45154 24434
rect 44918 17198 45154 17434
rect 44918 10198 45154 10434
rect 44918 3198 45154 3434
rect 44918 -1942 45154 -1706
rect 44918 -2262 45154 -2026
rect 50186 705002 50422 705238
rect 50186 704682 50422 704918
rect 50186 695258 50422 695494
rect 50186 688258 50422 688494
rect 50186 681258 50422 681494
rect 50186 674258 50422 674494
rect 50186 667258 50422 667494
rect 50186 660258 50422 660494
rect 50186 653258 50422 653494
rect 50186 646258 50422 646494
rect 50186 639258 50422 639494
rect 50186 632258 50422 632494
rect 50186 625258 50422 625494
rect 50186 618258 50422 618494
rect 50186 611258 50422 611494
rect 50186 604258 50422 604494
rect 50186 597258 50422 597494
rect 50186 590258 50422 590494
rect 50186 583258 50422 583494
rect 50186 576258 50422 576494
rect 50186 569258 50422 569494
rect 50186 562258 50422 562494
rect 50186 555258 50422 555494
rect 50186 548258 50422 548494
rect 50186 541258 50422 541494
rect 50186 534258 50422 534494
rect 50186 527258 50422 527494
rect 50186 520258 50422 520494
rect 50186 513258 50422 513494
rect 50186 506258 50422 506494
rect 50186 499258 50422 499494
rect 50186 492258 50422 492494
rect 50186 485258 50422 485494
rect 50186 478258 50422 478494
rect 50186 471258 50422 471494
rect 50186 464258 50422 464494
rect 50186 457258 50422 457494
rect 50186 450258 50422 450494
rect 50186 443258 50422 443494
rect 50186 436258 50422 436494
rect 50186 429258 50422 429494
rect 50186 422258 50422 422494
rect 50186 415258 50422 415494
rect 50186 408258 50422 408494
rect 50186 401258 50422 401494
rect 50186 394258 50422 394494
rect 50186 387258 50422 387494
rect 50186 380258 50422 380494
rect 50186 373258 50422 373494
rect 50186 366258 50422 366494
rect 50186 359258 50422 359494
rect 50186 352258 50422 352494
rect 50186 345258 50422 345494
rect 50186 338258 50422 338494
rect 50186 331258 50422 331494
rect 50186 324258 50422 324494
rect 50186 317258 50422 317494
rect 50186 310258 50422 310494
rect 50186 303258 50422 303494
rect 50186 296258 50422 296494
rect 50186 289258 50422 289494
rect 50186 282258 50422 282494
rect 50186 275258 50422 275494
rect 50186 268258 50422 268494
rect 50186 261258 50422 261494
rect 50186 254258 50422 254494
rect 50186 247258 50422 247494
rect 50186 240258 50422 240494
rect 50186 233258 50422 233494
rect 50186 226258 50422 226494
rect 50186 219258 50422 219494
rect 50186 212258 50422 212494
rect 50186 205258 50422 205494
rect 50186 198258 50422 198494
rect 50186 191258 50422 191494
rect 50186 184258 50422 184494
rect 50186 177258 50422 177494
rect 50186 170258 50422 170494
rect 50186 163258 50422 163494
rect 50186 156258 50422 156494
rect 50186 149258 50422 149494
rect 50186 142258 50422 142494
rect 50186 135258 50422 135494
rect 50186 128258 50422 128494
rect 50186 121258 50422 121494
rect 50186 114258 50422 114494
rect 50186 107258 50422 107494
rect 50186 100258 50422 100494
rect 50186 93258 50422 93494
rect 50186 86258 50422 86494
rect 50186 79258 50422 79494
rect 50186 72258 50422 72494
rect 50186 65258 50422 65494
rect 50186 58258 50422 58494
rect 50186 51258 50422 51494
rect 50186 44258 50422 44494
rect 50186 37258 50422 37494
rect 50186 30258 50422 30494
rect 50186 23258 50422 23494
rect 50186 16258 50422 16494
rect 50186 9258 50422 9494
rect 50186 2258 50422 2494
rect 50186 -982 50422 -746
rect 50186 -1302 50422 -1066
rect 51918 705962 52154 706198
rect 51918 705642 52154 705878
rect 51918 696198 52154 696434
rect 51918 689198 52154 689434
rect 51918 682198 52154 682434
rect 51918 675198 52154 675434
rect 51918 668198 52154 668434
rect 51918 661198 52154 661434
rect 51918 654198 52154 654434
rect 51918 647198 52154 647434
rect 51918 640198 52154 640434
rect 51918 633198 52154 633434
rect 51918 626198 52154 626434
rect 51918 619198 52154 619434
rect 51918 612198 52154 612434
rect 51918 605198 52154 605434
rect 51918 598198 52154 598434
rect 51918 591198 52154 591434
rect 51918 584198 52154 584434
rect 51918 577198 52154 577434
rect 51918 570198 52154 570434
rect 51918 563198 52154 563434
rect 51918 556198 52154 556434
rect 51918 549198 52154 549434
rect 51918 542198 52154 542434
rect 51918 535198 52154 535434
rect 51918 528198 52154 528434
rect 51918 521198 52154 521434
rect 51918 514198 52154 514434
rect 51918 507198 52154 507434
rect 51918 500198 52154 500434
rect 51918 493198 52154 493434
rect 51918 486198 52154 486434
rect 51918 479198 52154 479434
rect 51918 472198 52154 472434
rect 51918 465198 52154 465434
rect 51918 458198 52154 458434
rect 51918 451198 52154 451434
rect 51918 444198 52154 444434
rect 51918 437198 52154 437434
rect 51918 430198 52154 430434
rect 51918 423198 52154 423434
rect 51918 416198 52154 416434
rect 51918 409198 52154 409434
rect 51918 402198 52154 402434
rect 51918 395198 52154 395434
rect 51918 388198 52154 388434
rect 51918 381198 52154 381434
rect 51918 374198 52154 374434
rect 51918 367198 52154 367434
rect 51918 360198 52154 360434
rect 51918 353198 52154 353434
rect 51918 346198 52154 346434
rect 51918 339198 52154 339434
rect 51918 332198 52154 332434
rect 51918 325198 52154 325434
rect 51918 318198 52154 318434
rect 51918 311198 52154 311434
rect 51918 304198 52154 304434
rect 51918 297198 52154 297434
rect 51918 290198 52154 290434
rect 51918 283198 52154 283434
rect 51918 276198 52154 276434
rect 51918 269198 52154 269434
rect 51918 262198 52154 262434
rect 51918 255198 52154 255434
rect 51918 248198 52154 248434
rect 51918 241198 52154 241434
rect 51918 234198 52154 234434
rect 51918 227198 52154 227434
rect 51918 220198 52154 220434
rect 51918 213198 52154 213434
rect 51918 206198 52154 206434
rect 51918 199198 52154 199434
rect 51918 192198 52154 192434
rect 51918 185198 52154 185434
rect 51918 178198 52154 178434
rect 51918 171198 52154 171434
rect 51918 164198 52154 164434
rect 51918 157198 52154 157434
rect 51918 150198 52154 150434
rect 51918 143198 52154 143434
rect 51918 136198 52154 136434
rect 51918 129198 52154 129434
rect 51918 122198 52154 122434
rect 51918 115198 52154 115434
rect 51918 108198 52154 108434
rect 51918 101198 52154 101434
rect 51918 94198 52154 94434
rect 51918 87198 52154 87434
rect 51918 80198 52154 80434
rect 51918 73198 52154 73434
rect 51918 66198 52154 66434
rect 51918 59198 52154 59434
rect 51918 52198 52154 52434
rect 51918 45198 52154 45434
rect 51918 38198 52154 38434
rect 51918 31198 52154 31434
rect 51918 24198 52154 24434
rect 51918 17198 52154 17434
rect 51918 10198 52154 10434
rect 51918 3198 52154 3434
rect 51918 -1942 52154 -1706
rect 51918 -2262 52154 -2026
rect 57186 705002 57422 705238
rect 57186 704682 57422 704918
rect 57186 695258 57422 695494
rect 57186 688258 57422 688494
rect 57186 681258 57422 681494
rect 57186 674258 57422 674494
rect 57186 667258 57422 667494
rect 57186 660258 57422 660494
rect 57186 653258 57422 653494
rect 57186 646258 57422 646494
rect 57186 639258 57422 639494
rect 57186 632258 57422 632494
rect 57186 625258 57422 625494
rect 57186 618258 57422 618494
rect 57186 611258 57422 611494
rect 57186 604258 57422 604494
rect 57186 597258 57422 597494
rect 57186 590258 57422 590494
rect 57186 583258 57422 583494
rect 57186 576258 57422 576494
rect 57186 569258 57422 569494
rect 57186 562258 57422 562494
rect 57186 555258 57422 555494
rect 57186 548258 57422 548494
rect 57186 541258 57422 541494
rect 57186 534258 57422 534494
rect 57186 527258 57422 527494
rect 57186 520258 57422 520494
rect 57186 513258 57422 513494
rect 57186 506258 57422 506494
rect 57186 499258 57422 499494
rect 57186 492258 57422 492494
rect 57186 485258 57422 485494
rect 57186 478258 57422 478494
rect 57186 471258 57422 471494
rect 57186 464258 57422 464494
rect 57186 457258 57422 457494
rect 57186 450258 57422 450494
rect 57186 443258 57422 443494
rect 57186 436258 57422 436494
rect 57186 429258 57422 429494
rect 57186 422258 57422 422494
rect 57186 415258 57422 415494
rect 57186 408258 57422 408494
rect 57186 401258 57422 401494
rect 57186 394258 57422 394494
rect 57186 387258 57422 387494
rect 57186 380258 57422 380494
rect 57186 373258 57422 373494
rect 57186 366258 57422 366494
rect 57186 359258 57422 359494
rect 57186 352258 57422 352494
rect 57186 345258 57422 345494
rect 57186 338258 57422 338494
rect 57186 331258 57422 331494
rect 57186 324258 57422 324494
rect 57186 317258 57422 317494
rect 57186 310258 57422 310494
rect 57186 303258 57422 303494
rect 57186 296258 57422 296494
rect 57186 289258 57422 289494
rect 57186 282258 57422 282494
rect 57186 275258 57422 275494
rect 57186 268258 57422 268494
rect 57186 261258 57422 261494
rect 57186 254258 57422 254494
rect 57186 247258 57422 247494
rect 57186 240258 57422 240494
rect 57186 233258 57422 233494
rect 57186 226258 57422 226494
rect 57186 219258 57422 219494
rect 57186 212258 57422 212494
rect 57186 205258 57422 205494
rect 57186 198258 57422 198494
rect 57186 191258 57422 191494
rect 57186 184258 57422 184494
rect 57186 177258 57422 177494
rect 57186 170258 57422 170494
rect 57186 163258 57422 163494
rect 57186 156258 57422 156494
rect 57186 149258 57422 149494
rect 57186 142258 57422 142494
rect 57186 135258 57422 135494
rect 57186 128258 57422 128494
rect 57186 121258 57422 121494
rect 57186 114258 57422 114494
rect 57186 107258 57422 107494
rect 57186 100258 57422 100494
rect 57186 93258 57422 93494
rect 57186 86258 57422 86494
rect 57186 79258 57422 79494
rect 57186 72258 57422 72494
rect 57186 65258 57422 65494
rect 57186 58258 57422 58494
rect 57186 51258 57422 51494
rect 57186 44258 57422 44494
rect 57186 37258 57422 37494
rect 57186 30258 57422 30494
rect 57186 23258 57422 23494
rect 57186 16258 57422 16494
rect 57186 9258 57422 9494
rect 57186 2258 57422 2494
rect 57186 -982 57422 -746
rect 57186 -1302 57422 -1066
rect 58918 705962 59154 706198
rect 58918 705642 59154 705878
rect 58918 696198 59154 696434
rect 58918 689198 59154 689434
rect 58918 682198 59154 682434
rect 58918 675198 59154 675434
rect 58918 668198 59154 668434
rect 58918 661198 59154 661434
rect 58918 654198 59154 654434
rect 58918 647198 59154 647434
rect 58918 640198 59154 640434
rect 58918 633198 59154 633434
rect 58918 626198 59154 626434
rect 58918 619198 59154 619434
rect 58918 612198 59154 612434
rect 58918 605198 59154 605434
rect 58918 598198 59154 598434
rect 58918 591198 59154 591434
rect 58918 584198 59154 584434
rect 58918 577198 59154 577434
rect 58918 570198 59154 570434
rect 58918 563198 59154 563434
rect 58918 556198 59154 556434
rect 58918 549198 59154 549434
rect 58918 542198 59154 542434
rect 58918 535198 59154 535434
rect 58918 528198 59154 528434
rect 58918 521198 59154 521434
rect 58918 514198 59154 514434
rect 58918 507198 59154 507434
rect 58918 500198 59154 500434
rect 58918 493198 59154 493434
rect 58918 486198 59154 486434
rect 58918 479198 59154 479434
rect 58918 472198 59154 472434
rect 58918 465198 59154 465434
rect 58918 458198 59154 458434
rect 58918 451198 59154 451434
rect 58918 444198 59154 444434
rect 58918 437198 59154 437434
rect 58918 430198 59154 430434
rect 58918 423198 59154 423434
rect 58918 416198 59154 416434
rect 58918 409198 59154 409434
rect 58918 402198 59154 402434
rect 58918 395198 59154 395434
rect 58918 388198 59154 388434
rect 58918 381198 59154 381434
rect 58918 374198 59154 374434
rect 58918 367198 59154 367434
rect 58918 360198 59154 360434
rect 58918 353198 59154 353434
rect 58918 346198 59154 346434
rect 58918 339198 59154 339434
rect 58918 332198 59154 332434
rect 58918 325198 59154 325434
rect 58918 318198 59154 318434
rect 58918 311198 59154 311434
rect 58918 304198 59154 304434
rect 58918 297198 59154 297434
rect 58918 290198 59154 290434
rect 58918 283198 59154 283434
rect 58918 276198 59154 276434
rect 58918 269198 59154 269434
rect 58918 262198 59154 262434
rect 58918 255198 59154 255434
rect 58918 248198 59154 248434
rect 58918 241198 59154 241434
rect 58918 234198 59154 234434
rect 58918 227198 59154 227434
rect 58918 220198 59154 220434
rect 58918 213198 59154 213434
rect 58918 206198 59154 206434
rect 58918 199198 59154 199434
rect 58918 192198 59154 192434
rect 58918 185198 59154 185434
rect 58918 178198 59154 178434
rect 58918 171198 59154 171434
rect 58918 164198 59154 164434
rect 58918 157198 59154 157434
rect 58918 150198 59154 150434
rect 58918 143198 59154 143434
rect 58918 136198 59154 136434
rect 58918 129198 59154 129434
rect 58918 122198 59154 122434
rect 58918 115198 59154 115434
rect 58918 108198 59154 108434
rect 58918 101198 59154 101434
rect 58918 94198 59154 94434
rect 58918 87198 59154 87434
rect 58918 80198 59154 80434
rect 58918 73198 59154 73434
rect 58918 66198 59154 66434
rect 58918 59198 59154 59434
rect 58918 52198 59154 52434
rect 58918 45198 59154 45434
rect 58918 38198 59154 38434
rect 58918 31198 59154 31434
rect 58918 24198 59154 24434
rect 58918 17198 59154 17434
rect 58918 10198 59154 10434
rect 58918 3198 59154 3434
rect 58918 -1942 59154 -1706
rect 58918 -2262 59154 -2026
rect 64186 705002 64422 705238
rect 64186 704682 64422 704918
rect 64186 695258 64422 695494
rect 64186 688258 64422 688494
rect 64186 681258 64422 681494
rect 64186 674258 64422 674494
rect 64186 667258 64422 667494
rect 64186 660258 64422 660494
rect 64186 653258 64422 653494
rect 64186 646258 64422 646494
rect 64186 639258 64422 639494
rect 64186 632258 64422 632494
rect 64186 625258 64422 625494
rect 64186 618258 64422 618494
rect 64186 611258 64422 611494
rect 64186 604258 64422 604494
rect 64186 597258 64422 597494
rect 64186 590258 64422 590494
rect 64186 583258 64422 583494
rect 64186 576258 64422 576494
rect 64186 569258 64422 569494
rect 64186 562258 64422 562494
rect 64186 555258 64422 555494
rect 64186 548258 64422 548494
rect 64186 541258 64422 541494
rect 64186 534258 64422 534494
rect 64186 527258 64422 527494
rect 64186 520258 64422 520494
rect 64186 513258 64422 513494
rect 64186 506258 64422 506494
rect 64186 499258 64422 499494
rect 64186 492258 64422 492494
rect 64186 485258 64422 485494
rect 64186 478258 64422 478494
rect 64186 471258 64422 471494
rect 64186 464258 64422 464494
rect 64186 457258 64422 457494
rect 64186 450258 64422 450494
rect 64186 443258 64422 443494
rect 64186 436258 64422 436494
rect 64186 429258 64422 429494
rect 64186 422258 64422 422494
rect 64186 415258 64422 415494
rect 64186 408258 64422 408494
rect 64186 401258 64422 401494
rect 64186 394258 64422 394494
rect 64186 387258 64422 387494
rect 64186 380258 64422 380494
rect 64186 373258 64422 373494
rect 64186 366258 64422 366494
rect 64186 359258 64422 359494
rect 64186 352258 64422 352494
rect 64186 345258 64422 345494
rect 64186 338258 64422 338494
rect 64186 331258 64422 331494
rect 64186 324258 64422 324494
rect 64186 317258 64422 317494
rect 64186 310258 64422 310494
rect 64186 303258 64422 303494
rect 64186 296258 64422 296494
rect 64186 289258 64422 289494
rect 64186 282258 64422 282494
rect 64186 275258 64422 275494
rect 64186 268258 64422 268494
rect 64186 261258 64422 261494
rect 64186 254258 64422 254494
rect 64186 247258 64422 247494
rect 64186 240258 64422 240494
rect 64186 233258 64422 233494
rect 64186 226258 64422 226494
rect 64186 219258 64422 219494
rect 64186 212258 64422 212494
rect 64186 205258 64422 205494
rect 64186 198258 64422 198494
rect 64186 191258 64422 191494
rect 64186 184258 64422 184494
rect 64186 177258 64422 177494
rect 64186 170258 64422 170494
rect 64186 163258 64422 163494
rect 64186 156258 64422 156494
rect 64186 149258 64422 149494
rect 64186 142258 64422 142494
rect 64186 135258 64422 135494
rect 64186 128258 64422 128494
rect 64186 121258 64422 121494
rect 64186 114258 64422 114494
rect 64186 107258 64422 107494
rect 64186 100258 64422 100494
rect 64186 93258 64422 93494
rect 64186 86258 64422 86494
rect 64186 79258 64422 79494
rect 64186 72258 64422 72494
rect 64186 65258 64422 65494
rect 64186 58258 64422 58494
rect 64186 51258 64422 51494
rect 64186 44258 64422 44494
rect 64186 37258 64422 37494
rect 64186 30258 64422 30494
rect 64186 23258 64422 23494
rect 64186 16258 64422 16494
rect 64186 9258 64422 9494
rect 64186 2258 64422 2494
rect 64186 -982 64422 -746
rect 64186 -1302 64422 -1066
rect 65918 705962 66154 706198
rect 65918 705642 66154 705878
rect 65918 696198 66154 696434
rect 65918 689198 66154 689434
rect 65918 682198 66154 682434
rect 65918 675198 66154 675434
rect 65918 668198 66154 668434
rect 65918 661198 66154 661434
rect 65918 654198 66154 654434
rect 65918 647198 66154 647434
rect 65918 640198 66154 640434
rect 65918 633198 66154 633434
rect 65918 626198 66154 626434
rect 65918 619198 66154 619434
rect 65918 612198 66154 612434
rect 65918 605198 66154 605434
rect 65918 598198 66154 598434
rect 65918 591198 66154 591434
rect 65918 584198 66154 584434
rect 65918 577198 66154 577434
rect 65918 570198 66154 570434
rect 65918 563198 66154 563434
rect 65918 556198 66154 556434
rect 65918 549198 66154 549434
rect 65918 542198 66154 542434
rect 65918 535198 66154 535434
rect 65918 528198 66154 528434
rect 65918 521198 66154 521434
rect 65918 514198 66154 514434
rect 65918 507198 66154 507434
rect 65918 500198 66154 500434
rect 65918 493198 66154 493434
rect 65918 486198 66154 486434
rect 65918 479198 66154 479434
rect 65918 472198 66154 472434
rect 65918 465198 66154 465434
rect 65918 458198 66154 458434
rect 65918 451198 66154 451434
rect 65918 444198 66154 444434
rect 65918 437198 66154 437434
rect 65918 430198 66154 430434
rect 65918 423198 66154 423434
rect 65918 416198 66154 416434
rect 65918 409198 66154 409434
rect 65918 402198 66154 402434
rect 65918 395198 66154 395434
rect 65918 388198 66154 388434
rect 65918 381198 66154 381434
rect 65918 374198 66154 374434
rect 65918 367198 66154 367434
rect 65918 360198 66154 360434
rect 65918 353198 66154 353434
rect 65918 346198 66154 346434
rect 65918 339198 66154 339434
rect 65918 332198 66154 332434
rect 65918 325198 66154 325434
rect 65918 318198 66154 318434
rect 65918 311198 66154 311434
rect 65918 304198 66154 304434
rect 65918 297198 66154 297434
rect 65918 290198 66154 290434
rect 65918 283198 66154 283434
rect 65918 276198 66154 276434
rect 65918 269198 66154 269434
rect 65918 262198 66154 262434
rect 65918 255198 66154 255434
rect 65918 248198 66154 248434
rect 65918 241198 66154 241434
rect 65918 234198 66154 234434
rect 65918 227198 66154 227434
rect 65918 220198 66154 220434
rect 65918 213198 66154 213434
rect 65918 206198 66154 206434
rect 65918 199198 66154 199434
rect 65918 192198 66154 192434
rect 65918 185198 66154 185434
rect 65918 178198 66154 178434
rect 65918 171198 66154 171434
rect 65918 164198 66154 164434
rect 65918 157198 66154 157434
rect 65918 150198 66154 150434
rect 65918 143198 66154 143434
rect 65918 136198 66154 136434
rect 65918 129198 66154 129434
rect 65918 122198 66154 122434
rect 65918 115198 66154 115434
rect 65918 108198 66154 108434
rect 65918 101198 66154 101434
rect 65918 94198 66154 94434
rect 65918 87198 66154 87434
rect 65918 80198 66154 80434
rect 65918 73198 66154 73434
rect 65918 66198 66154 66434
rect 65918 59198 66154 59434
rect 65918 52198 66154 52434
rect 65918 45198 66154 45434
rect 65918 38198 66154 38434
rect 65918 31198 66154 31434
rect 65918 24198 66154 24434
rect 65918 17198 66154 17434
rect 65918 10198 66154 10434
rect 65918 3198 66154 3434
rect 65918 -1942 66154 -1706
rect 65918 -2262 66154 -2026
rect 71186 705002 71422 705238
rect 71186 704682 71422 704918
rect 71186 695258 71422 695494
rect 71186 688258 71422 688494
rect 71186 681258 71422 681494
rect 71186 674258 71422 674494
rect 71186 667258 71422 667494
rect 71186 660258 71422 660494
rect 71186 653258 71422 653494
rect 71186 646258 71422 646494
rect 71186 639258 71422 639494
rect 71186 632258 71422 632494
rect 71186 625258 71422 625494
rect 71186 618258 71422 618494
rect 71186 611258 71422 611494
rect 71186 604258 71422 604494
rect 71186 597258 71422 597494
rect 71186 590258 71422 590494
rect 71186 583258 71422 583494
rect 71186 576258 71422 576494
rect 71186 569258 71422 569494
rect 71186 562258 71422 562494
rect 71186 555258 71422 555494
rect 71186 548258 71422 548494
rect 71186 541258 71422 541494
rect 71186 534258 71422 534494
rect 71186 527258 71422 527494
rect 71186 520258 71422 520494
rect 71186 513258 71422 513494
rect 71186 506258 71422 506494
rect 71186 499258 71422 499494
rect 71186 492258 71422 492494
rect 71186 485258 71422 485494
rect 71186 478258 71422 478494
rect 71186 471258 71422 471494
rect 71186 464258 71422 464494
rect 71186 457258 71422 457494
rect 71186 450258 71422 450494
rect 71186 443258 71422 443494
rect 71186 436258 71422 436494
rect 71186 429258 71422 429494
rect 71186 422258 71422 422494
rect 71186 415258 71422 415494
rect 71186 408258 71422 408494
rect 71186 401258 71422 401494
rect 71186 394258 71422 394494
rect 71186 387258 71422 387494
rect 71186 380258 71422 380494
rect 71186 373258 71422 373494
rect 71186 366258 71422 366494
rect 71186 359258 71422 359494
rect 71186 352258 71422 352494
rect 71186 345258 71422 345494
rect 71186 338258 71422 338494
rect 71186 331258 71422 331494
rect 71186 324258 71422 324494
rect 71186 317258 71422 317494
rect 71186 310258 71422 310494
rect 71186 303258 71422 303494
rect 71186 296258 71422 296494
rect 71186 289258 71422 289494
rect 71186 282258 71422 282494
rect 71186 275258 71422 275494
rect 71186 268258 71422 268494
rect 71186 261258 71422 261494
rect 71186 254258 71422 254494
rect 71186 247258 71422 247494
rect 71186 240258 71422 240494
rect 71186 233258 71422 233494
rect 71186 226258 71422 226494
rect 71186 219258 71422 219494
rect 71186 212258 71422 212494
rect 71186 205258 71422 205494
rect 71186 198258 71422 198494
rect 71186 191258 71422 191494
rect 71186 184258 71422 184494
rect 71186 177258 71422 177494
rect 71186 170258 71422 170494
rect 71186 163258 71422 163494
rect 71186 156258 71422 156494
rect 71186 149258 71422 149494
rect 71186 142258 71422 142494
rect 71186 135258 71422 135494
rect 71186 128258 71422 128494
rect 71186 121258 71422 121494
rect 71186 114258 71422 114494
rect 71186 107258 71422 107494
rect 71186 100258 71422 100494
rect 71186 93258 71422 93494
rect 71186 86258 71422 86494
rect 71186 79258 71422 79494
rect 71186 72258 71422 72494
rect 71186 65258 71422 65494
rect 71186 58258 71422 58494
rect 71186 51258 71422 51494
rect 71186 44258 71422 44494
rect 71186 37258 71422 37494
rect 71186 30258 71422 30494
rect 71186 23258 71422 23494
rect 71186 16258 71422 16494
rect 71186 9258 71422 9494
rect 71186 2258 71422 2494
rect 71186 -982 71422 -746
rect 71186 -1302 71422 -1066
rect 72918 705962 73154 706198
rect 72918 705642 73154 705878
rect 72918 696198 73154 696434
rect 72918 689198 73154 689434
rect 72918 682198 73154 682434
rect 72918 675198 73154 675434
rect 72918 668198 73154 668434
rect 72918 661198 73154 661434
rect 72918 654198 73154 654434
rect 72918 647198 73154 647434
rect 72918 640198 73154 640434
rect 72918 633198 73154 633434
rect 72918 626198 73154 626434
rect 72918 619198 73154 619434
rect 72918 612198 73154 612434
rect 72918 605198 73154 605434
rect 72918 598198 73154 598434
rect 72918 591198 73154 591434
rect 72918 584198 73154 584434
rect 72918 577198 73154 577434
rect 72918 570198 73154 570434
rect 72918 563198 73154 563434
rect 72918 556198 73154 556434
rect 72918 549198 73154 549434
rect 72918 542198 73154 542434
rect 72918 535198 73154 535434
rect 72918 528198 73154 528434
rect 72918 521198 73154 521434
rect 72918 514198 73154 514434
rect 72918 507198 73154 507434
rect 72918 500198 73154 500434
rect 72918 493198 73154 493434
rect 72918 486198 73154 486434
rect 72918 479198 73154 479434
rect 72918 472198 73154 472434
rect 72918 465198 73154 465434
rect 72918 458198 73154 458434
rect 72918 451198 73154 451434
rect 72918 444198 73154 444434
rect 72918 437198 73154 437434
rect 72918 430198 73154 430434
rect 72918 423198 73154 423434
rect 72918 416198 73154 416434
rect 72918 409198 73154 409434
rect 72918 402198 73154 402434
rect 72918 395198 73154 395434
rect 72918 388198 73154 388434
rect 72918 381198 73154 381434
rect 72918 374198 73154 374434
rect 72918 367198 73154 367434
rect 72918 360198 73154 360434
rect 72918 353198 73154 353434
rect 72918 346198 73154 346434
rect 72918 339198 73154 339434
rect 72918 332198 73154 332434
rect 72918 325198 73154 325434
rect 72918 318198 73154 318434
rect 72918 311198 73154 311434
rect 72918 304198 73154 304434
rect 72918 297198 73154 297434
rect 72918 290198 73154 290434
rect 72918 283198 73154 283434
rect 72918 276198 73154 276434
rect 72918 269198 73154 269434
rect 72918 262198 73154 262434
rect 72918 255198 73154 255434
rect 72918 248198 73154 248434
rect 72918 241198 73154 241434
rect 72918 234198 73154 234434
rect 72918 227198 73154 227434
rect 72918 220198 73154 220434
rect 72918 213198 73154 213434
rect 72918 206198 73154 206434
rect 72918 199198 73154 199434
rect 72918 192198 73154 192434
rect 72918 185198 73154 185434
rect 72918 178198 73154 178434
rect 72918 171198 73154 171434
rect 72918 164198 73154 164434
rect 72918 157198 73154 157434
rect 72918 150198 73154 150434
rect 72918 143198 73154 143434
rect 72918 136198 73154 136434
rect 72918 129198 73154 129434
rect 72918 122198 73154 122434
rect 72918 115198 73154 115434
rect 72918 108198 73154 108434
rect 72918 101198 73154 101434
rect 72918 94198 73154 94434
rect 72918 87198 73154 87434
rect 72918 80198 73154 80434
rect 72918 73198 73154 73434
rect 72918 66198 73154 66434
rect 72918 59198 73154 59434
rect 72918 52198 73154 52434
rect 72918 45198 73154 45434
rect 72918 38198 73154 38434
rect 72918 31198 73154 31434
rect 72918 24198 73154 24434
rect 72918 17198 73154 17434
rect 72918 10198 73154 10434
rect 72918 3198 73154 3434
rect 72918 -1942 73154 -1706
rect 72918 -2262 73154 -2026
rect 78186 705002 78422 705238
rect 78186 704682 78422 704918
rect 78186 695258 78422 695494
rect 78186 688258 78422 688494
rect 78186 681258 78422 681494
rect 78186 674258 78422 674494
rect 78186 667258 78422 667494
rect 78186 660258 78422 660494
rect 78186 653258 78422 653494
rect 78186 646258 78422 646494
rect 78186 639258 78422 639494
rect 78186 632258 78422 632494
rect 78186 625258 78422 625494
rect 78186 618258 78422 618494
rect 78186 611258 78422 611494
rect 78186 604258 78422 604494
rect 78186 597258 78422 597494
rect 78186 590258 78422 590494
rect 78186 583258 78422 583494
rect 78186 576258 78422 576494
rect 78186 569258 78422 569494
rect 78186 562258 78422 562494
rect 78186 555258 78422 555494
rect 78186 548258 78422 548494
rect 78186 541258 78422 541494
rect 78186 534258 78422 534494
rect 78186 527258 78422 527494
rect 78186 520258 78422 520494
rect 78186 513258 78422 513494
rect 78186 506258 78422 506494
rect 78186 499258 78422 499494
rect 78186 492258 78422 492494
rect 78186 485258 78422 485494
rect 78186 478258 78422 478494
rect 78186 471258 78422 471494
rect 78186 464258 78422 464494
rect 78186 457258 78422 457494
rect 78186 450258 78422 450494
rect 78186 443258 78422 443494
rect 78186 436258 78422 436494
rect 78186 429258 78422 429494
rect 78186 422258 78422 422494
rect 78186 415258 78422 415494
rect 78186 408258 78422 408494
rect 78186 401258 78422 401494
rect 78186 394258 78422 394494
rect 78186 387258 78422 387494
rect 78186 380258 78422 380494
rect 78186 373258 78422 373494
rect 78186 366258 78422 366494
rect 78186 359258 78422 359494
rect 78186 352258 78422 352494
rect 78186 345258 78422 345494
rect 78186 338258 78422 338494
rect 78186 331258 78422 331494
rect 78186 324258 78422 324494
rect 78186 317258 78422 317494
rect 78186 310258 78422 310494
rect 78186 303258 78422 303494
rect 78186 296258 78422 296494
rect 78186 289258 78422 289494
rect 78186 282258 78422 282494
rect 78186 275258 78422 275494
rect 78186 268258 78422 268494
rect 78186 261258 78422 261494
rect 78186 254258 78422 254494
rect 78186 247258 78422 247494
rect 78186 240258 78422 240494
rect 78186 233258 78422 233494
rect 78186 226258 78422 226494
rect 78186 219258 78422 219494
rect 78186 212258 78422 212494
rect 78186 205258 78422 205494
rect 78186 198258 78422 198494
rect 78186 191258 78422 191494
rect 78186 184258 78422 184494
rect 78186 177258 78422 177494
rect 78186 170258 78422 170494
rect 78186 163258 78422 163494
rect 78186 156258 78422 156494
rect 78186 149258 78422 149494
rect 78186 142258 78422 142494
rect 78186 135258 78422 135494
rect 78186 128258 78422 128494
rect 78186 121258 78422 121494
rect 78186 114258 78422 114494
rect 78186 107258 78422 107494
rect 78186 100258 78422 100494
rect 78186 93258 78422 93494
rect 78186 86258 78422 86494
rect 78186 79258 78422 79494
rect 78186 72258 78422 72494
rect 78186 65258 78422 65494
rect 78186 58258 78422 58494
rect 78186 51258 78422 51494
rect 78186 44258 78422 44494
rect 78186 37258 78422 37494
rect 78186 30258 78422 30494
rect 78186 23258 78422 23494
rect 78186 16258 78422 16494
rect 78186 9258 78422 9494
rect 78186 2258 78422 2494
rect 78186 -982 78422 -746
rect 78186 -1302 78422 -1066
rect 79918 705962 80154 706198
rect 79918 705642 80154 705878
rect 79918 696198 80154 696434
rect 79918 689198 80154 689434
rect 79918 682198 80154 682434
rect 79918 675198 80154 675434
rect 79918 668198 80154 668434
rect 79918 661198 80154 661434
rect 79918 654198 80154 654434
rect 79918 647198 80154 647434
rect 79918 640198 80154 640434
rect 79918 633198 80154 633434
rect 79918 626198 80154 626434
rect 79918 619198 80154 619434
rect 79918 612198 80154 612434
rect 79918 605198 80154 605434
rect 79918 598198 80154 598434
rect 79918 591198 80154 591434
rect 79918 584198 80154 584434
rect 79918 577198 80154 577434
rect 79918 570198 80154 570434
rect 79918 563198 80154 563434
rect 79918 556198 80154 556434
rect 79918 549198 80154 549434
rect 79918 542198 80154 542434
rect 79918 535198 80154 535434
rect 79918 528198 80154 528434
rect 79918 521198 80154 521434
rect 79918 514198 80154 514434
rect 79918 507198 80154 507434
rect 79918 500198 80154 500434
rect 79918 493198 80154 493434
rect 79918 486198 80154 486434
rect 79918 479198 80154 479434
rect 79918 472198 80154 472434
rect 79918 465198 80154 465434
rect 79918 458198 80154 458434
rect 79918 451198 80154 451434
rect 79918 444198 80154 444434
rect 79918 437198 80154 437434
rect 79918 430198 80154 430434
rect 79918 423198 80154 423434
rect 79918 416198 80154 416434
rect 79918 409198 80154 409434
rect 79918 402198 80154 402434
rect 79918 395198 80154 395434
rect 79918 388198 80154 388434
rect 79918 381198 80154 381434
rect 79918 374198 80154 374434
rect 79918 367198 80154 367434
rect 79918 360198 80154 360434
rect 79918 353198 80154 353434
rect 79918 346198 80154 346434
rect 79918 339198 80154 339434
rect 79918 332198 80154 332434
rect 79918 325198 80154 325434
rect 79918 318198 80154 318434
rect 79918 311198 80154 311434
rect 79918 304198 80154 304434
rect 79918 297198 80154 297434
rect 79918 290198 80154 290434
rect 79918 283198 80154 283434
rect 79918 276198 80154 276434
rect 79918 269198 80154 269434
rect 79918 262198 80154 262434
rect 79918 255198 80154 255434
rect 79918 248198 80154 248434
rect 79918 241198 80154 241434
rect 79918 234198 80154 234434
rect 79918 227198 80154 227434
rect 79918 220198 80154 220434
rect 79918 213198 80154 213434
rect 79918 206198 80154 206434
rect 79918 199198 80154 199434
rect 79918 192198 80154 192434
rect 79918 185198 80154 185434
rect 79918 178198 80154 178434
rect 79918 171198 80154 171434
rect 79918 164198 80154 164434
rect 79918 157198 80154 157434
rect 79918 150198 80154 150434
rect 79918 143198 80154 143434
rect 79918 136198 80154 136434
rect 79918 129198 80154 129434
rect 79918 122198 80154 122434
rect 79918 115198 80154 115434
rect 79918 108198 80154 108434
rect 79918 101198 80154 101434
rect 79918 94198 80154 94434
rect 79918 87198 80154 87434
rect 79918 80198 80154 80434
rect 79918 73198 80154 73434
rect 79918 66198 80154 66434
rect 79918 59198 80154 59434
rect 79918 52198 80154 52434
rect 79918 45198 80154 45434
rect 79918 38198 80154 38434
rect 79918 31198 80154 31434
rect 79918 24198 80154 24434
rect 79918 17198 80154 17434
rect 79918 10198 80154 10434
rect 79918 3198 80154 3434
rect 79918 -1942 80154 -1706
rect 79918 -2262 80154 -2026
rect 85186 705002 85422 705238
rect 85186 704682 85422 704918
rect 85186 695258 85422 695494
rect 85186 688258 85422 688494
rect 85186 681258 85422 681494
rect 85186 674258 85422 674494
rect 85186 667258 85422 667494
rect 85186 660258 85422 660494
rect 85186 653258 85422 653494
rect 85186 646258 85422 646494
rect 85186 639258 85422 639494
rect 85186 632258 85422 632494
rect 85186 625258 85422 625494
rect 85186 618258 85422 618494
rect 85186 611258 85422 611494
rect 85186 604258 85422 604494
rect 85186 597258 85422 597494
rect 85186 590258 85422 590494
rect 85186 583258 85422 583494
rect 85186 576258 85422 576494
rect 85186 569258 85422 569494
rect 85186 562258 85422 562494
rect 85186 555258 85422 555494
rect 85186 548258 85422 548494
rect 85186 541258 85422 541494
rect 85186 534258 85422 534494
rect 85186 527258 85422 527494
rect 85186 520258 85422 520494
rect 85186 513258 85422 513494
rect 85186 506258 85422 506494
rect 85186 499258 85422 499494
rect 85186 492258 85422 492494
rect 85186 485258 85422 485494
rect 85186 478258 85422 478494
rect 85186 471258 85422 471494
rect 85186 464258 85422 464494
rect 85186 457258 85422 457494
rect 85186 450258 85422 450494
rect 85186 443258 85422 443494
rect 85186 436258 85422 436494
rect 85186 429258 85422 429494
rect 85186 422258 85422 422494
rect 85186 415258 85422 415494
rect 85186 408258 85422 408494
rect 85186 401258 85422 401494
rect 85186 394258 85422 394494
rect 85186 387258 85422 387494
rect 85186 380258 85422 380494
rect 85186 373258 85422 373494
rect 85186 366258 85422 366494
rect 85186 359258 85422 359494
rect 85186 352258 85422 352494
rect 85186 345258 85422 345494
rect 85186 338258 85422 338494
rect 85186 331258 85422 331494
rect 85186 324258 85422 324494
rect 85186 317258 85422 317494
rect 85186 310258 85422 310494
rect 85186 303258 85422 303494
rect 85186 296258 85422 296494
rect 85186 289258 85422 289494
rect 85186 282258 85422 282494
rect 85186 275258 85422 275494
rect 85186 268258 85422 268494
rect 85186 261258 85422 261494
rect 85186 254258 85422 254494
rect 85186 247258 85422 247494
rect 85186 240258 85422 240494
rect 85186 233258 85422 233494
rect 85186 226258 85422 226494
rect 85186 219258 85422 219494
rect 85186 212258 85422 212494
rect 85186 205258 85422 205494
rect 85186 198258 85422 198494
rect 85186 191258 85422 191494
rect 85186 184258 85422 184494
rect 85186 177258 85422 177494
rect 85186 170258 85422 170494
rect 85186 163258 85422 163494
rect 85186 156258 85422 156494
rect 85186 149258 85422 149494
rect 85186 142258 85422 142494
rect 85186 135258 85422 135494
rect 85186 128258 85422 128494
rect 85186 121258 85422 121494
rect 85186 114258 85422 114494
rect 85186 107258 85422 107494
rect 85186 100258 85422 100494
rect 85186 93258 85422 93494
rect 85186 86258 85422 86494
rect 85186 79258 85422 79494
rect 85186 72258 85422 72494
rect 85186 65258 85422 65494
rect 85186 58258 85422 58494
rect 85186 51258 85422 51494
rect 85186 44258 85422 44494
rect 85186 37258 85422 37494
rect 85186 30258 85422 30494
rect 85186 23258 85422 23494
rect 85186 16258 85422 16494
rect 85186 9258 85422 9494
rect 85186 2258 85422 2494
rect 85186 -982 85422 -746
rect 85186 -1302 85422 -1066
rect 86918 705962 87154 706198
rect 86918 705642 87154 705878
rect 86918 696198 87154 696434
rect 86918 689198 87154 689434
rect 86918 682198 87154 682434
rect 86918 675198 87154 675434
rect 86918 668198 87154 668434
rect 86918 661198 87154 661434
rect 86918 654198 87154 654434
rect 86918 647198 87154 647434
rect 86918 640198 87154 640434
rect 86918 633198 87154 633434
rect 86918 626198 87154 626434
rect 86918 619198 87154 619434
rect 86918 612198 87154 612434
rect 86918 605198 87154 605434
rect 86918 598198 87154 598434
rect 86918 591198 87154 591434
rect 86918 584198 87154 584434
rect 86918 577198 87154 577434
rect 86918 570198 87154 570434
rect 86918 563198 87154 563434
rect 86918 556198 87154 556434
rect 86918 549198 87154 549434
rect 86918 542198 87154 542434
rect 86918 535198 87154 535434
rect 86918 528198 87154 528434
rect 86918 521198 87154 521434
rect 86918 514198 87154 514434
rect 86918 507198 87154 507434
rect 86918 500198 87154 500434
rect 86918 493198 87154 493434
rect 86918 486198 87154 486434
rect 86918 479198 87154 479434
rect 86918 472198 87154 472434
rect 86918 465198 87154 465434
rect 86918 458198 87154 458434
rect 86918 451198 87154 451434
rect 86918 444198 87154 444434
rect 86918 437198 87154 437434
rect 86918 430198 87154 430434
rect 86918 423198 87154 423434
rect 86918 416198 87154 416434
rect 86918 409198 87154 409434
rect 86918 402198 87154 402434
rect 86918 395198 87154 395434
rect 86918 388198 87154 388434
rect 86918 381198 87154 381434
rect 86918 374198 87154 374434
rect 86918 367198 87154 367434
rect 86918 360198 87154 360434
rect 86918 353198 87154 353434
rect 86918 346198 87154 346434
rect 86918 339198 87154 339434
rect 86918 332198 87154 332434
rect 86918 325198 87154 325434
rect 86918 318198 87154 318434
rect 86918 311198 87154 311434
rect 86918 304198 87154 304434
rect 86918 297198 87154 297434
rect 86918 290198 87154 290434
rect 86918 283198 87154 283434
rect 86918 276198 87154 276434
rect 86918 269198 87154 269434
rect 86918 262198 87154 262434
rect 86918 255198 87154 255434
rect 86918 248198 87154 248434
rect 86918 241198 87154 241434
rect 86918 234198 87154 234434
rect 86918 227198 87154 227434
rect 86918 220198 87154 220434
rect 86918 213198 87154 213434
rect 86918 206198 87154 206434
rect 86918 199198 87154 199434
rect 86918 192198 87154 192434
rect 86918 185198 87154 185434
rect 86918 178198 87154 178434
rect 86918 171198 87154 171434
rect 86918 164198 87154 164434
rect 86918 157198 87154 157434
rect 86918 150198 87154 150434
rect 86918 143198 87154 143434
rect 86918 136198 87154 136434
rect 86918 129198 87154 129434
rect 86918 122198 87154 122434
rect 86918 115198 87154 115434
rect 86918 108198 87154 108434
rect 86918 101198 87154 101434
rect 86918 94198 87154 94434
rect 86918 87198 87154 87434
rect 86918 80198 87154 80434
rect 86918 73198 87154 73434
rect 86918 66198 87154 66434
rect 86918 59198 87154 59434
rect 86918 52198 87154 52434
rect 86918 45198 87154 45434
rect 86918 38198 87154 38434
rect 86918 31198 87154 31434
rect 86918 24198 87154 24434
rect 86918 17198 87154 17434
rect 86918 10198 87154 10434
rect 86918 3198 87154 3434
rect 86918 -1942 87154 -1706
rect 86918 -2262 87154 -2026
rect 92186 705002 92422 705238
rect 92186 704682 92422 704918
rect 92186 695258 92422 695494
rect 92186 688258 92422 688494
rect 92186 681258 92422 681494
rect 92186 674258 92422 674494
rect 92186 667258 92422 667494
rect 92186 660258 92422 660494
rect 92186 653258 92422 653494
rect 92186 646258 92422 646494
rect 92186 639258 92422 639494
rect 92186 632258 92422 632494
rect 92186 625258 92422 625494
rect 92186 618258 92422 618494
rect 92186 611258 92422 611494
rect 92186 604258 92422 604494
rect 92186 597258 92422 597494
rect 92186 590258 92422 590494
rect 92186 583258 92422 583494
rect 92186 576258 92422 576494
rect 92186 569258 92422 569494
rect 92186 562258 92422 562494
rect 92186 555258 92422 555494
rect 92186 548258 92422 548494
rect 92186 541258 92422 541494
rect 92186 534258 92422 534494
rect 92186 527258 92422 527494
rect 92186 520258 92422 520494
rect 92186 513258 92422 513494
rect 92186 506258 92422 506494
rect 92186 499258 92422 499494
rect 92186 492258 92422 492494
rect 92186 485258 92422 485494
rect 92186 478258 92422 478494
rect 92186 471258 92422 471494
rect 92186 464258 92422 464494
rect 92186 457258 92422 457494
rect 92186 450258 92422 450494
rect 92186 443258 92422 443494
rect 92186 436258 92422 436494
rect 92186 429258 92422 429494
rect 92186 422258 92422 422494
rect 92186 415258 92422 415494
rect 92186 408258 92422 408494
rect 92186 401258 92422 401494
rect 92186 394258 92422 394494
rect 92186 387258 92422 387494
rect 92186 380258 92422 380494
rect 92186 373258 92422 373494
rect 92186 366258 92422 366494
rect 92186 359258 92422 359494
rect 92186 352258 92422 352494
rect 92186 345258 92422 345494
rect 92186 338258 92422 338494
rect 92186 331258 92422 331494
rect 92186 324258 92422 324494
rect 92186 317258 92422 317494
rect 92186 310258 92422 310494
rect 92186 303258 92422 303494
rect 92186 296258 92422 296494
rect 92186 289258 92422 289494
rect 92186 282258 92422 282494
rect 92186 275258 92422 275494
rect 92186 268258 92422 268494
rect 92186 261258 92422 261494
rect 92186 254258 92422 254494
rect 92186 247258 92422 247494
rect 92186 240258 92422 240494
rect 92186 233258 92422 233494
rect 92186 226258 92422 226494
rect 92186 219258 92422 219494
rect 92186 212258 92422 212494
rect 92186 205258 92422 205494
rect 92186 198258 92422 198494
rect 92186 191258 92422 191494
rect 92186 184258 92422 184494
rect 92186 177258 92422 177494
rect 92186 170258 92422 170494
rect 92186 163258 92422 163494
rect 92186 156258 92422 156494
rect 92186 149258 92422 149494
rect 92186 142258 92422 142494
rect 92186 135258 92422 135494
rect 92186 128258 92422 128494
rect 92186 121258 92422 121494
rect 92186 114258 92422 114494
rect 92186 107258 92422 107494
rect 92186 100258 92422 100494
rect 92186 93258 92422 93494
rect 92186 86258 92422 86494
rect 92186 79258 92422 79494
rect 92186 72258 92422 72494
rect 92186 65258 92422 65494
rect 92186 58258 92422 58494
rect 92186 51258 92422 51494
rect 92186 44258 92422 44494
rect 92186 37258 92422 37494
rect 92186 30258 92422 30494
rect 92186 23258 92422 23494
rect 92186 16258 92422 16494
rect 92186 9258 92422 9494
rect 92186 2258 92422 2494
rect 92186 -982 92422 -746
rect 92186 -1302 92422 -1066
rect 93918 705962 94154 706198
rect 93918 705642 94154 705878
rect 93918 696198 94154 696434
rect 93918 689198 94154 689434
rect 93918 682198 94154 682434
rect 93918 675198 94154 675434
rect 93918 668198 94154 668434
rect 93918 661198 94154 661434
rect 93918 654198 94154 654434
rect 93918 647198 94154 647434
rect 93918 640198 94154 640434
rect 93918 633198 94154 633434
rect 93918 626198 94154 626434
rect 93918 619198 94154 619434
rect 93918 612198 94154 612434
rect 93918 605198 94154 605434
rect 93918 598198 94154 598434
rect 93918 591198 94154 591434
rect 93918 584198 94154 584434
rect 93918 577198 94154 577434
rect 93918 570198 94154 570434
rect 93918 563198 94154 563434
rect 93918 556198 94154 556434
rect 93918 549198 94154 549434
rect 93918 542198 94154 542434
rect 93918 535198 94154 535434
rect 93918 528198 94154 528434
rect 93918 521198 94154 521434
rect 93918 514198 94154 514434
rect 93918 507198 94154 507434
rect 93918 500198 94154 500434
rect 93918 493198 94154 493434
rect 93918 486198 94154 486434
rect 93918 479198 94154 479434
rect 93918 472198 94154 472434
rect 93918 465198 94154 465434
rect 93918 458198 94154 458434
rect 93918 451198 94154 451434
rect 93918 444198 94154 444434
rect 93918 437198 94154 437434
rect 93918 430198 94154 430434
rect 93918 423198 94154 423434
rect 93918 416198 94154 416434
rect 93918 409198 94154 409434
rect 93918 402198 94154 402434
rect 93918 395198 94154 395434
rect 93918 388198 94154 388434
rect 93918 381198 94154 381434
rect 93918 374198 94154 374434
rect 93918 367198 94154 367434
rect 93918 360198 94154 360434
rect 93918 353198 94154 353434
rect 93918 346198 94154 346434
rect 93918 339198 94154 339434
rect 93918 332198 94154 332434
rect 93918 325198 94154 325434
rect 93918 318198 94154 318434
rect 93918 311198 94154 311434
rect 93918 304198 94154 304434
rect 93918 297198 94154 297434
rect 93918 290198 94154 290434
rect 93918 283198 94154 283434
rect 93918 276198 94154 276434
rect 93918 269198 94154 269434
rect 93918 262198 94154 262434
rect 93918 255198 94154 255434
rect 93918 248198 94154 248434
rect 93918 241198 94154 241434
rect 93918 234198 94154 234434
rect 93918 227198 94154 227434
rect 93918 220198 94154 220434
rect 93918 213198 94154 213434
rect 93918 206198 94154 206434
rect 93918 199198 94154 199434
rect 93918 192198 94154 192434
rect 93918 185198 94154 185434
rect 93918 178198 94154 178434
rect 93918 171198 94154 171434
rect 93918 164198 94154 164434
rect 93918 157198 94154 157434
rect 93918 150198 94154 150434
rect 93918 143198 94154 143434
rect 93918 136198 94154 136434
rect 93918 129198 94154 129434
rect 93918 122198 94154 122434
rect 93918 115198 94154 115434
rect 93918 108198 94154 108434
rect 93918 101198 94154 101434
rect 93918 94198 94154 94434
rect 93918 87198 94154 87434
rect 93918 80198 94154 80434
rect 93918 73198 94154 73434
rect 93918 66198 94154 66434
rect 93918 59198 94154 59434
rect 93918 52198 94154 52434
rect 93918 45198 94154 45434
rect 93918 38198 94154 38434
rect 93918 31198 94154 31434
rect 93918 24198 94154 24434
rect 93918 17198 94154 17434
rect 93918 10198 94154 10434
rect 93918 3198 94154 3434
rect 93918 -1942 94154 -1706
rect 93918 -2262 94154 -2026
rect 99186 705002 99422 705238
rect 99186 704682 99422 704918
rect 99186 695258 99422 695494
rect 99186 688258 99422 688494
rect 99186 681258 99422 681494
rect 99186 674258 99422 674494
rect 99186 667258 99422 667494
rect 99186 660258 99422 660494
rect 99186 653258 99422 653494
rect 99186 646258 99422 646494
rect 99186 639258 99422 639494
rect 99186 632258 99422 632494
rect 99186 625258 99422 625494
rect 99186 618258 99422 618494
rect 99186 611258 99422 611494
rect 99186 604258 99422 604494
rect 99186 597258 99422 597494
rect 99186 590258 99422 590494
rect 99186 583258 99422 583494
rect 99186 576258 99422 576494
rect 99186 569258 99422 569494
rect 99186 562258 99422 562494
rect 99186 555258 99422 555494
rect 99186 548258 99422 548494
rect 99186 541258 99422 541494
rect 99186 534258 99422 534494
rect 99186 527258 99422 527494
rect 99186 520258 99422 520494
rect 99186 513258 99422 513494
rect 99186 506258 99422 506494
rect 99186 499258 99422 499494
rect 99186 492258 99422 492494
rect 99186 485258 99422 485494
rect 99186 478258 99422 478494
rect 99186 471258 99422 471494
rect 99186 464258 99422 464494
rect 99186 457258 99422 457494
rect 99186 450258 99422 450494
rect 99186 443258 99422 443494
rect 99186 436258 99422 436494
rect 99186 429258 99422 429494
rect 99186 422258 99422 422494
rect 99186 415258 99422 415494
rect 99186 408258 99422 408494
rect 99186 401258 99422 401494
rect 99186 394258 99422 394494
rect 99186 387258 99422 387494
rect 99186 380258 99422 380494
rect 99186 373258 99422 373494
rect 99186 366258 99422 366494
rect 99186 359258 99422 359494
rect 99186 352258 99422 352494
rect 99186 345258 99422 345494
rect 99186 338258 99422 338494
rect 99186 331258 99422 331494
rect 99186 324258 99422 324494
rect 99186 317258 99422 317494
rect 99186 310258 99422 310494
rect 99186 303258 99422 303494
rect 99186 296258 99422 296494
rect 99186 289258 99422 289494
rect 99186 282258 99422 282494
rect 99186 275258 99422 275494
rect 99186 268258 99422 268494
rect 99186 261258 99422 261494
rect 99186 254258 99422 254494
rect 99186 247258 99422 247494
rect 99186 240258 99422 240494
rect 99186 233258 99422 233494
rect 99186 226258 99422 226494
rect 99186 219258 99422 219494
rect 99186 212258 99422 212494
rect 99186 205258 99422 205494
rect 99186 198258 99422 198494
rect 99186 191258 99422 191494
rect 99186 184258 99422 184494
rect 99186 177258 99422 177494
rect 99186 170258 99422 170494
rect 99186 163258 99422 163494
rect 99186 156258 99422 156494
rect 99186 149258 99422 149494
rect 99186 142258 99422 142494
rect 99186 135258 99422 135494
rect 99186 128258 99422 128494
rect 99186 121258 99422 121494
rect 99186 114258 99422 114494
rect 99186 107258 99422 107494
rect 99186 100258 99422 100494
rect 99186 93258 99422 93494
rect 99186 86258 99422 86494
rect 99186 79258 99422 79494
rect 99186 72258 99422 72494
rect 99186 65258 99422 65494
rect 99186 58258 99422 58494
rect 99186 51258 99422 51494
rect 99186 44258 99422 44494
rect 99186 37258 99422 37494
rect 99186 30258 99422 30494
rect 99186 23258 99422 23494
rect 99186 16258 99422 16494
rect 99186 9258 99422 9494
rect 99186 2258 99422 2494
rect 99186 -982 99422 -746
rect 99186 -1302 99422 -1066
rect 100918 705962 101154 706198
rect 100918 705642 101154 705878
rect 100918 696198 101154 696434
rect 100918 689198 101154 689434
rect 100918 682198 101154 682434
rect 100918 675198 101154 675434
rect 100918 668198 101154 668434
rect 100918 661198 101154 661434
rect 100918 654198 101154 654434
rect 100918 647198 101154 647434
rect 100918 640198 101154 640434
rect 100918 633198 101154 633434
rect 100918 626198 101154 626434
rect 100918 619198 101154 619434
rect 100918 612198 101154 612434
rect 100918 605198 101154 605434
rect 100918 598198 101154 598434
rect 100918 591198 101154 591434
rect 100918 584198 101154 584434
rect 100918 577198 101154 577434
rect 100918 570198 101154 570434
rect 100918 563198 101154 563434
rect 100918 556198 101154 556434
rect 100918 549198 101154 549434
rect 100918 542198 101154 542434
rect 100918 535198 101154 535434
rect 100918 528198 101154 528434
rect 100918 521198 101154 521434
rect 100918 514198 101154 514434
rect 100918 507198 101154 507434
rect 100918 500198 101154 500434
rect 100918 493198 101154 493434
rect 100918 486198 101154 486434
rect 100918 479198 101154 479434
rect 100918 472198 101154 472434
rect 100918 465198 101154 465434
rect 100918 458198 101154 458434
rect 100918 451198 101154 451434
rect 100918 444198 101154 444434
rect 100918 437198 101154 437434
rect 100918 430198 101154 430434
rect 100918 423198 101154 423434
rect 100918 416198 101154 416434
rect 100918 409198 101154 409434
rect 100918 402198 101154 402434
rect 100918 395198 101154 395434
rect 100918 388198 101154 388434
rect 100918 381198 101154 381434
rect 100918 374198 101154 374434
rect 100918 367198 101154 367434
rect 100918 360198 101154 360434
rect 100918 353198 101154 353434
rect 100918 346198 101154 346434
rect 100918 339198 101154 339434
rect 100918 332198 101154 332434
rect 100918 325198 101154 325434
rect 100918 318198 101154 318434
rect 100918 311198 101154 311434
rect 100918 304198 101154 304434
rect 100918 297198 101154 297434
rect 100918 290198 101154 290434
rect 100918 283198 101154 283434
rect 100918 276198 101154 276434
rect 100918 269198 101154 269434
rect 100918 262198 101154 262434
rect 100918 255198 101154 255434
rect 100918 248198 101154 248434
rect 100918 241198 101154 241434
rect 100918 234198 101154 234434
rect 100918 227198 101154 227434
rect 100918 220198 101154 220434
rect 100918 213198 101154 213434
rect 100918 206198 101154 206434
rect 100918 199198 101154 199434
rect 100918 192198 101154 192434
rect 100918 185198 101154 185434
rect 100918 178198 101154 178434
rect 100918 171198 101154 171434
rect 100918 164198 101154 164434
rect 100918 157198 101154 157434
rect 100918 150198 101154 150434
rect 100918 143198 101154 143434
rect 100918 136198 101154 136434
rect 100918 129198 101154 129434
rect 100918 122198 101154 122434
rect 100918 115198 101154 115434
rect 100918 108198 101154 108434
rect 100918 101198 101154 101434
rect 100918 94198 101154 94434
rect 100918 87198 101154 87434
rect 100918 80198 101154 80434
rect 100918 73198 101154 73434
rect 100918 66198 101154 66434
rect 100918 59198 101154 59434
rect 100918 52198 101154 52434
rect 100918 45198 101154 45434
rect 100918 38198 101154 38434
rect 100918 31198 101154 31434
rect 100918 24198 101154 24434
rect 100918 17198 101154 17434
rect 100918 10198 101154 10434
rect 100918 3198 101154 3434
rect 100918 -1942 101154 -1706
rect 100918 -2262 101154 -2026
rect 106186 705002 106422 705238
rect 106186 704682 106422 704918
rect 106186 695258 106422 695494
rect 106186 688258 106422 688494
rect 106186 681258 106422 681494
rect 106186 674258 106422 674494
rect 106186 667258 106422 667494
rect 106186 660258 106422 660494
rect 106186 653258 106422 653494
rect 106186 646258 106422 646494
rect 106186 639258 106422 639494
rect 106186 632258 106422 632494
rect 106186 625258 106422 625494
rect 106186 618258 106422 618494
rect 106186 611258 106422 611494
rect 106186 604258 106422 604494
rect 106186 597258 106422 597494
rect 106186 590258 106422 590494
rect 106186 583258 106422 583494
rect 106186 576258 106422 576494
rect 106186 569258 106422 569494
rect 106186 562258 106422 562494
rect 106186 555258 106422 555494
rect 106186 548258 106422 548494
rect 106186 541258 106422 541494
rect 106186 534258 106422 534494
rect 106186 527258 106422 527494
rect 106186 520258 106422 520494
rect 106186 513258 106422 513494
rect 106186 506258 106422 506494
rect 106186 499258 106422 499494
rect 106186 492258 106422 492494
rect 106186 485258 106422 485494
rect 106186 478258 106422 478494
rect 106186 471258 106422 471494
rect 106186 464258 106422 464494
rect 106186 457258 106422 457494
rect 106186 450258 106422 450494
rect 106186 443258 106422 443494
rect 106186 436258 106422 436494
rect 106186 429258 106422 429494
rect 106186 422258 106422 422494
rect 106186 415258 106422 415494
rect 106186 408258 106422 408494
rect 106186 401258 106422 401494
rect 106186 394258 106422 394494
rect 106186 387258 106422 387494
rect 106186 380258 106422 380494
rect 106186 373258 106422 373494
rect 106186 366258 106422 366494
rect 106186 359258 106422 359494
rect 106186 352258 106422 352494
rect 106186 345258 106422 345494
rect 106186 338258 106422 338494
rect 106186 331258 106422 331494
rect 106186 324258 106422 324494
rect 106186 317258 106422 317494
rect 106186 310258 106422 310494
rect 106186 303258 106422 303494
rect 106186 296258 106422 296494
rect 106186 289258 106422 289494
rect 106186 282258 106422 282494
rect 106186 275258 106422 275494
rect 106186 268258 106422 268494
rect 106186 261258 106422 261494
rect 106186 254258 106422 254494
rect 106186 247258 106422 247494
rect 106186 240258 106422 240494
rect 106186 233258 106422 233494
rect 106186 226258 106422 226494
rect 106186 219258 106422 219494
rect 106186 212258 106422 212494
rect 106186 205258 106422 205494
rect 106186 198258 106422 198494
rect 106186 191258 106422 191494
rect 106186 184258 106422 184494
rect 106186 177258 106422 177494
rect 106186 170258 106422 170494
rect 106186 163258 106422 163494
rect 106186 156258 106422 156494
rect 106186 149258 106422 149494
rect 106186 142258 106422 142494
rect 106186 135258 106422 135494
rect 106186 128258 106422 128494
rect 106186 121258 106422 121494
rect 106186 114258 106422 114494
rect 106186 107258 106422 107494
rect 106186 100258 106422 100494
rect 106186 93258 106422 93494
rect 106186 86258 106422 86494
rect 106186 79258 106422 79494
rect 106186 72258 106422 72494
rect 106186 65258 106422 65494
rect 106186 58258 106422 58494
rect 106186 51258 106422 51494
rect 106186 44258 106422 44494
rect 106186 37258 106422 37494
rect 106186 30258 106422 30494
rect 106186 23258 106422 23494
rect 106186 16258 106422 16494
rect 106186 9258 106422 9494
rect 106186 2258 106422 2494
rect 106186 -982 106422 -746
rect 106186 -1302 106422 -1066
rect 107918 705962 108154 706198
rect 107918 705642 108154 705878
rect 107918 696198 108154 696434
rect 107918 689198 108154 689434
rect 107918 682198 108154 682434
rect 107918 675198 108154 675434
rect 107918 668198 108154 668434
rect 107918 661198 108154 661434
rect 107918 654198 108154 654434
rect 107918 647198 108154 647434
rect 107918 640198 108154 640434
rect 107918 633198 108154 633434
rect 107918 626198 108154 626434
rect 107918 619198 108154 619434
rect 107918 612198 108154 612434
rect 107918 605198 108154 605434
rect 107918 598198 108154 598434
rect 107918 591198 108154 591434
rect 107918 584198 108154 584434
rect 107918 577198 108154 577434
rect 107918 570198 108154 570434
rect 107918 563198 108154 563434
rect 107918 556198 108154 556434
rect 107918 549198 108154 549434
rect 107918 542198 108154 542434
rect 107918 535198 108154 535434
rect 107918 528198 108154 528434
rect 107918 521198 108154 521434
rect 107918 514198 108154 514434
rect 107918 507198 108154 507434
rect 107918 500198 108154 500434
rect 107918 493198 108154 493434
rect 107918 486198 108154 486434
rect 107918 479198 108154 479434
rect 107918 472198 108154 472434
rect 107918 465198 108154 465434
rect 107918 458198 108154 458434
rect 107918 451198 108154 451434
rect 107918 444198 108154 444434
rect 107918 437198 108154 437434
rect 107918 430198 108154 430434
rect 107918 423198 108154 423434
rect 107918 416198 108154 416434
rect 107918 409198 108154 409434
rect 107918 402198 108154 402434
rect 107918 395198 108154 395434
rect 107918 388198 108154 388434
rect 107918 381198 108154 381434
rect 107918 374198 108154 374434
rect 107918 367198 108154 367434
rect 107918 360198 108154 360434
rect 107918 353198 108154 353434
rect 107918 346198 108154 346434
rect 107918 339198 108154 339434
rect 107918 332198 108154 332434
rect 107918 325198 108154 325434
rect 107918 318198 108154 318434
rect 107918 311198 108154 311434
rect 107918 304198 108154 304434
rect 107918 297198 108154 297434
rect 107918 290198 108154 290434
rect 107918 283198 108154 283434
rect 107918 276198 108154 276434
rect 107918 269198 108154 269434
rect 107918 262198 108154 262434
rect 107918 255198 108154 255434
rect 107918 248198 108154 248434
rect 107918 241198 108154 241434
rect 107918 234198 108154 234434
rect 107918 227198 108154 227434
rect 107918 220198 108154 220434
rect 107918 213198 108154 213434
rect 107918 206198 108154 206434
rect 107918 199198 108154 199434
rect 107918 192198 108154 192434
rect 107918 185198 108154 185434
rect 107918 178198 108154 178434
rect 107918 171198 108154 171434
rect 107918 164198 108154 164434
rect 107918 157198 108154 157434
rect 107918 150198 108154 150434
rect 107918 143198 108154 143434
rect 107918 136198 108154 136434
rect 107918 129198 108154 129434
rect 107918 122198 108154 122434
rect 107918 115198 108154 115434
rect 107918 108198 108154 108434
rect 107918 101198 108154 101434
rect 107918 94198 108154 94434
rect 107918 87198 108154 87434
rect 107918 80198 108154 80434
rect 107918 73198 108154 73434
rect 107918 66198 108154 66434
rect 107918 59198 108154 59434
rect 107918 52198 108154 52434
rect 107918 45198 108154 45434
rect 107918 38198 108154 38434
rect 107918 31198 108154 31434
rect 107918 24198 108154 24434
rect 107918 17198 108154 17434
rect 107918 10198 108154 10434
rect 107918 3198 108154 3434
rect 107918 -1942 108154 -1706
rect 107918 -2262 108154 -2026
rect 113186 705002 113422 705238
rect 113186 704682 113422 704918
rect 113186 695258 113422 695494
rect 113186 688258 113422 688494
rect 113186 681258 113422 681494
rect 113186 674258 113422 674494
rect 113186 667258 113422 667494
rect 113186 660258 113422 660494
rect 113186 653258 113422 653494
rect 113186 646258 113422 646494
rect 113186 639258 113422 639494
rect 113186 632258 113422 632494
rect 113186 625258 113422 625494
rect 113186 618258 113422 618494
rect 113186 611258 113422 611494
rect 113186 604258 113422 604494
rect 113186 597258 113422 597494
rect 113186 590258 113422 590494
rect 113186 583258 113422 583494
rect 113186 576258 113422 576494
rect 113186 569258 113422 569494
rect 113186 562258 113422 562494
rect 113186 555258 113422 555494
rect 113186 548258 113422 548494
rect 113186 541258 113422 541494
rect 113186 534258 113422 534494
rect 113186 527258 113422 527494
rect 113186 520258 113422 520494
rect 113186 513258 113422 513494
rect 113186 506258 113422 506494
rect 113186 499258 113422 499494
rect 113186 492258 113422 492494
rect 113186 485258 113422 485494
rect 113186 478258 113422 478494
rect 113186 471258 113422 471494
rect 113186 464258 113422 464494
rect 113186 457258 113422 457494
rect 113186 450258 113422 450494
rect 113186 443258 113422 443494
rect 113186 436258 113422 436494
rect 113186 429258 113422 429494
rect 113186 422258 113422 422494
rect 113186 415258 113422 415494
rect 113186 408258 113422 408494
rect 113186 401258 113422 401494
rect 113186 394258 113422 394494
rect 113186 387258 113422 387494
rect 113186 380258 113422 380494
rect 113186 373258 113422 373494
rect 113186 366258 113422 366494
rect 113186 359258 113422 359494
rect 113186 352258 113422 352494
rect 113186 345258 113422 345494
rect 113186 338258 113422 338494
rect 113186 331258 113422 331494
rect 113186 324258 113422 324494
rect 113186 317258 113422 317494
rect 113186 310258 113422 310494
rect 113186 303258 113422 303494
rect 113186 296258 113422 296494
rect 113186 289258 113422 289494
rect 113186 282258 113422 282494
rect 113186 275258 113422 275494
rect 113186 268258 113422 268494
rect 113186 261258 113422 261494
rect 113186 254258 113422 254494
rect 113186 247258 113422 247494
rect 113186 240258 113422 240494
rect 113186 233258 113422 233494
rect 113186 226258 113422 226494
rect 113186 219258 113422 219494
rect 113186 212258 113422 212494
rect 113186 205258 113422 205494
rect 113186 198258 113422 198494
rect 113186 191258 113422 191494
rect 113186 184258 113422 184494
rect 113186 177258 113422 177494
rect 113186 170258 113422 170494
rect 113186 163258 113422 163494
rect 113186 156258 113422 156494
rect 113186 149258 113422 149494
rect 113186 142258 113422 142494
rect 113186 135258 113422 135494
rect 113186 128258 113422 128494
rect 113186 121258 113422 121494
rect 113186 114258 113422 114494
rect 113186 107258 113422 107494
rect 113186 100258 113422 100494
rect 113186 93258 113422 93494
rect 113186 86258 113422 86494
rect 113186 79258 113422 79494
rect 113186 72258 113422 72494
rect 113186 65258 113422 65494
rect 113186 58258 113422 58494
rect 113186 51258 113422 51494
rect 113186 44258 113422 44494
rect 113186 37258 113422 37494
rect 113186 30258 113422 30494
rect 113186 23258 113422 23494
rect 113186 16258 113422 16494
rect 113186 9258 113422 9494
rect 113186 2258 113422 2494
rect 113186 -982 113422 -746
rect 113186 -1302 113422 -1066
rect 114918 705962 115154 706198
rect 114918 705642 115154 705878
rect 114918 696198 115154 696434
rect 114918 689198 115154 689434
rect 114918 682198 115154 682434
rect 114918 675198 115154 675434
rect 114918 668198 115154 668434
rect 114918 661198 115154 661434
rect 114918 654198 115154 654434
rect 114918 647198 115154 647434
rect 114918 640198 115154 640434
rect 114918 633198 115154 633434
rect 114918 626198 115154 626434
rect 114918 619198 115154 619434
rect 114918 612198 115154 612434
rect 114918 605198 115154 605434
rect 114918 598198 115154 598434
rect 114918 591198 115154 591434
rect 114918 584198 115154 584434
rect 114918 577198 115154 577434
rect 114918 570198 115154 570434
rect 114918 563198 115154 563434
rect 114918 556198 115154 556434
rect 114918 549198 115154 549434
rect 114918 542198 115154 542434
rect 114918 535198 115154 535434
rect 114918 528198 115154 528434
rect 114918 521198 115154 521434
rect 114918 514198 115154 514434
rect 114918 507198 115154 507434
rect 114918 500198 115154 500434
rect 114918 493198 115154 493434
rect 114918 486198 115154 486434
rect 114918 479198 115154 479434
rect 114918 472198 115154 472434
rect 114918 465198 115154 465434
rect 114918 458198 115154 458434
rect 114918 451198 115154 451434
rect 114918 444198 115154 444434
rect 114918 437198 115154 437434
rect 114918 430198 115154 430434
rect 114918 423198 115154 423434
rect 114918 416198 115154 416434
rect 114918 409198 115154 409434
rect 114918 402198 115154 402434
rect 114918 395198 115154 395434
rect 114918 388198 115154 388434
rect 114918 381198 115154 381434
rect 114918 374198 115154 374434
rect 114918 367198 115154 367434
rect 114918 360198 115154 360434
rect 114918 353198 115154 353434
rect 114918 346198 115154 346434
rect 114918 339198 115154 339434
rect 114918 332198 115154 332434
rect 114918 325198 115154 325434
rect 114918 318198 115154 318434
rect 114918 311198 115154 311434
rect 114918 304198 115154 304434
rect 114918 297198 115154 297434
rect 114918 290198 115154 290434
rect 114918 283198 115154 283434
rect 114918 276198 115154 276434
rect 114918 269198 115154 269434
rect 114918 262198 115154 262434
rect 114918 255198 115154 255434
rect 114918 248198 115154 248434
rect 114918 241198 115154 241434
rect 114918 234198 115154 234434
rect 114918 227198 115154 227434
rect 114918 220198 115154 220434
rect 114918 213198 115154 213434
rect 114918 206198 115154 206434
rect 114918 199198 115154 199434
rect 114918 192198 115154 192434
rect 114918 185198 115154 185434
rect 114918 178198 115154 178434
rect 114918 171198 115154 171434
rect 114918 164198 115154 164434
rect 114918 157198 115154 157434
rect 114918 150198 115154 150434
rect 114918 143198 115154 143434
rect 114918 136198 115154 136434
rect 114918 129198 115154 129434
rect 114918 122198 115154 122434
rect 114918 115198 115154 115434
rect 114918 108198 115154 108434
rect 114918 101198 115154 101434
rect 114918 94198 115154 94434
rect 114918 87198 115154 87434
rect 114918 80198 115154 80434
rect 114918 73198 115154 73434
rect 114918 66198 115154 66434
rect 114918 59198 115154 59434
rect 114918 52198 115154 52434
rect 114918 45198 115154 45434
rect 114918 38198 115154 38434
rect 114918 31198 115154 31434
rect 114918 24198 115154 24434
rect 114918 17198 115154 17434
rect 114918 10198 115154 10434
rect 114918 3198 115154 3434
rect 114918 -1942 115154 -1706
rect 114918 -2262 115154 -2026
rect 120186 705002 120422 705238
rect 120186 704682 120422 704918
rect 120186 695258 120422 695494
rect 120186 688258 120422 688494
rect 120186 681258 120422 681494
rect 120186 674258 120422 674494
rect 120186 667258 120422 667494
rect 120186 660258 120422 660494
rect 120186 653258 120422 653494
rect 120186 646258 120422 646494
rect 120186 639258 120422 639494
rect 120186 632258 120422 632494
rect 120186 625258 120422 625494
rect 120186 618258 120422 618494
rect 120186 611258 120422 611494
rect 120186 604258 120422 604494
rect 120186 597258 120422 597494
rect 120186 590258 120422 590494
rect 120186 583258 120422 583494
rect 120186 576258 120422 576494
rect 120186 569258 120422 569494
rect 120186 562258 120422 562494
rect 120186 555258 120422 555494
rect 120186 548258 120422 548494
rect 120186 541258 120422 541494
rect 120186 534258 120422 534494
rect 120186 527258 120422 527494
rect 120186 520258 120422 520494
rect 120186 513258 120422 513494
rect 120186 506258 120422 506494
rect 120186 499258 120422 499494
rect 120186 492258 120422 492494
rect 120186 485258 120422 485494
rect 120186 478258 120422 478494
rect 120186 471258 120422 471494
rect 120186 464258 120422 464494
rect 120186 457258 120422 457494
rect 120186 450258 120422 450494
rect 120186 443258 120422 443494
rect 120186 436258 120422 436494
rect 120186 429258 120422 429494
rect 120186 422258 120422 422494
rect 120186 415258 120422 415494
rect 120186 408258 120422 408494
rect 120186 401258 120422 401494
rect 120186 394258 120422 394494
rect 120186 387258 120422 387494
rect 120186 380258 120422 380494
rect 120186 373258 120422 373494
rect 120186 366258 120422 366494
rect 120186 359258 120422 359494
rect 120186 352258 120422 352494
rect 120186 345258 120422 345494
rect 120186 338258 120422 338494
rect 120186 331258 120422 331494
rect 120186 324258 120422 324494
rect 120186 317258 120422 317494
rect 120186 310258 120422 310494
rect 120186 303258 120422 303494
rect 120186 296258 120422 296494
rect 120186 289258 120422 289494
rect 120186 282258 120422 282494
rect 120186 275258 120422 275494
rect 120186 268258 120422 268494
rect 120186 261258 120422 261494
rect 120186 254258 120422 254494
rect 120186 247258 120422 247494
rect 120186 240258 120422 240494
rect 120186 233258 120422 233494
rect 120186 226258 120422 226494
rect 120186 219258 120422 219494
rect 120186 212258 120422 212494
rect 120186 205258 120422 205494
rect 120186 198258 120422 198494
rect 120186 191258 120422 191494
rect 120186 184258 120422 184494
rect 120186 177258 120422 177494
rect 120186 170258 120422 170494
rect 120186 163258 120422 163494
rect 120186 156258 120422 156494
rect 120186 149258 120422 149494
rect 120186 142258 120422 142494
rect 120186 135258 120422 135494
rect 120186 128258 120422 128494
rect 120186 121258 120422 121494
rect 120186 114258 120422 114494
rect 120186 107258 120422 107494
rect 120186 100258 120422 100494
rect 120186 93258 120422 93494
rect 120186 86258 120422 86494
rect 120186 79258 120422 79494
rect 120186 72258 120422 72494
rect 120186 65258 120422 65494
rect 120186 58258 120422 58494
rect 120186 51258 120422 51494
rect 120186 44258 120422 44494
rect 120186 37258 120422 37494
rect 120186 30258 120422 30494
rect 120186 23258 120422 23494
rect 120186 16258 120422 16494
rect 120186 9258 120422 9494
rect 120186 2258 120422 2494
rect 120186 -982 120422 -746
rect 120186 -1302 120422 -1066
rect 121918 705962 122154 706198
rect 121918 705642 122154 705878
rect 121918 696198 122154 696434
rect 121918 689198 122154 689434
rect 121918 682198 122154 682434
rect 121918 675198 122154 675434
rect 121918 668198 122154 668434
rect 121918 661198 122154 661434
rect 121918 654198 122154 654434
rect 121918 647198 122154 647434
rect 121918 640198 122154 640434
rect 121918 633198 122154 633434
rect 121918 626198 122154 626434
rect 121918 619198 122154 619434
rect 121918 612198 122154 612434
rect 121918 605198 122154 605434
rect 121918 598198 122154 598434
rect 121918 591198 122154 591434
rect 121918 584198 122154 584434
rect 121918 577198 122154 577434
rect 121918 570198 122154 570434
rect 121918 563198 122154 563434
rect 121918 556198 122154 556434
rect 121918 549198 122154 549434
rect 121918 542198 122154 542434
rect 121918 535198 122154 535434
rect 121918 528198 122154 528434
rect 121918 521198 122154 521434
rect 121918 514198 122154 514434
rect 121918 507198 122154 507434
rect 121918 500198 122154 500434
rect 121918 493198 122154 493434
rect 121918 486198 122154 486434
rect 121918 479198 122154 479434
rect 121918 472198 122154 472434
rect 121918 465198 122154 465434
rect 121918 458198 122154 458434
rect 121918 451198 122154 451434
rect 121918 444198 122154 444434
rect 121918 437198 122154 437434
rect 121918 430198 122154 430434
rect 121918 423198 122154 423434
rect 121918 416198 122154 416434
rect 121918 409198 122154 409434
rect 121918 402198 122154 402434
rect 121918 395198 122154 395434
rect 121918 388198 122154 388434
rect 121918 381198 122154 381434
rect 121918 374198 122154 374434
rect 121918 367198 122154 367434
rect 121918 360198 122154 360434
rect 121918 353198 122154 353434
rect 121918 346198 122154 346434
rect 121918 339198 122154 339434
rect 121918 332198 122154 332434
rect 121918 325198 122154 325434
rect 121918 318198 122154 318434
rect 121918 311198 122154 311434
rect 121918 304198 122154 304434
rect 121918 297198 122154 297434
rect 121918 290198 122154 290434
rect 121918 283198 122154 283434
rect 121918 276198 122154 276434
rect 121918 269198 122154 269434
rect 121918 262198 122154 262434
rect 121918 255198 122154 255434
rect 121918 248198 122154 248434
rect 121918 241198 122154 241434
rect 121918 234198 122154 234434
rect 121918 227198 122154 227434
rect 121918 220198 122154 220434
rect 121918 213198 122154 213434
rect 121918 206198 122154 206434
rect 121918 199198 122154 199434
rect 121918 192198 122154 192434
rect 121918 185198 122154 185434
rect 121918 178198 122154 178434
rect 121918 171198 122154 171434
rect 121918 164198 122154 164434
rect 121918 157198 122154 157434
rect 121918 150198 122154 150434
rect 121918 143198 122154 143434
rect 121918 136198 122154 136434
rect 121918 129198 122154 129434
rect 121918 122198 122154 122434
rect 121918 115198 122154 115434
rect 121918 108198 122154 108434
rect 121918 101198 122154 101434
rect 121918 94198 122154 94434
rect 121918 87198 122154 87434
rect 121918 80198 122154 80434
rect 121918 73198 122154 73434
rect 121918 66198 122154 66434
rect 121918 59198 122154 59434
rect 121918 52198 122154 52434
rect 121918 45198 122154 45434
rect 121918 38198 122154 38434
rect 121918 31198 122154 31434
rect 121918 24198 122154 24434
rect 121918 17198 122154 17434
rect 121918 10198 122154 10434
rect 121918 3198 122154 3434
rect 121918 -1942 122154 -1706
rect 121918 -2262 122154 -2026
rect 127186 705002 127422 705238
rect 127186 704682 127422 704918
rect 127186 695258 127422 695494
rect 127186 688258 127422 688494
rect 127186 681258 127422 681494
rect 127186 674258 127422 674494
rect 127186 667258 127422 667494
rect 127186 660258 127422 660494
rect 127186 653258 127422 653494
rect 127186 646258 127422 646494
rect 127186 639258 127422 639494
rect 127186 632258 127422 632494
rect 127186 625258 127422 625494
rect 127186 618258 127422 618494
rect 127186 611258 127422 611494
rect 127186 604258 127422 604494
rect 127186 597258 127422 597494
rect 127186 590258 127422 590494
rect 127186 583258 127422 583494
rect 127186 576258 127422 576494
rect 127186 569258 127422 569494
rect 127186 562258 127422 562494
rect 127186 555258 127422 555494
rect 127186 548258 127422 548494
rect 127186 541258 127422 541494
rect 127186 534258 127422 534494
rect 127186 527258 127422 527494
rect 127186 520258 127422 520494
rect 127186 513258 127422 513494
rect 127186 506258 127422 506494
rect 127186 499258 127422 499494
rect 127186 492258 127422 492494
rect 127186 485258 127422 485494
rect 127186 478258 127422 478494
rect 127186 471258 127422 471494
rect 127186 464258 127422 464494
rect 127186 457258 127422 457494
rect 127186 450258 127422 450494
rect 127186 443258 127422 443494
rect 127186 436258 127422 436494
rect 127186 429258 127422 429494
rect 127186 422258 127422 422494
rect 127186 415258 127422 415494
rect 127186 408258 127422 408494
rect 127186 401258 127422 401494
rect 127186 394258 127422 394494
rect 127186 387258 127422 387494
rect 127186 380258 127422 380494
rect 127186 373258 127422 373494
rect 127186 366258 127422 366494
rect 127186 359258 127422 359494
rect 127186 352258 127422 352494
rect 127186 345258 127422 345494
rect 127186 338258 127422 338494
rect 127186 331258 127422 331494
rect 127186 324258 127422 324494
rect 127186 317258 127422 317494
rect 127186 310258 127422 310494
rect 127186 303258 127422 303494
rect 127186 296258 127422 296494
rect 127186 289258 127422 289494
rect 127186 282258 127422 282494
rect 127186 275258 127422 275494
rect 127186 268258 127422 268494
rect 127186 261258 127422 261494
rect 127186 254258 127422 254494
rect 127186 247258 127422 247494
rect 127186 240258 127422 240494
rect 127186 233258 127422 233494
rect 127186 226258 127422 226494
rect 127186 219258 127422 219494
rect 127186 212258 127422 212494
rect 127186 205258 127422 205494
rect 127186 198258 127422 198494
rect 127186 191258 127422 191494
rect 127186 184258 127422 184494
rect 127186 177258 127422 177494
rect 127186 170258 127422 170494
rect 127186 163258 127422 163494
rect 127186 156258 127422 156494
rect 127186 149258 127422 149494
rect 127186 142258 127422 142494
rect 127186 135258 127422 135494
rect 127186 128258 127422 128494
rect 127186 121258 127422 121494
rect 127186 114258 127422 114494
rect 127186 107258 127422 107494
rect 127186 100258 127422 100494
rect 127186 93258 127422 93494
rect 127186 86258 127422 86494
rect 127186 79258 127422 79494
rect 127186 72258 127422 72494
rect 127186 65258 127422 65494
rect 127186 58258 127422 58494
rect 127186 51258 127422 51494
rect 127186 44258 127422 44494
rect 127186 37258 127422 37494
rect 127186 30258 127422 30494
rect 127186 23258 127422 23494
rect 127186 16258 127422 16494
rect 127186 9258 127422 9494
rect 127186 2258 127422 2494
rect 127186 -982 127422 -746
rect 127186 -1302 127422 -1066
rect 128918 705962 129154 706198
rect 128918 705642 129154 705878
rect 128918 696198 129154 696434
rect 128918 689198 129154 689434
rect 128918 682198 129154 682434
rect 128918 675198 129154 675434
rect 128918 668198 129154 668434
rect 128918 661198 129154 661434
rect 128918 654198 129154 654434
rect 128918 647198 129154 647434
rect 128918 640198 129154 640434
rect 128918 633198 129154 633434
rect 128918 626198 129154 626434
rect 128918 619198 129154 619434
rect 128918 612198 129154 612434
rect 128918 605198 129154 605434
rect 128918 598198 129154 598434
rect 128918 591198 129154 591434
rect 128918 584198 129154 584434
rect 128918 577198 129154 577434
rect 128918 570198 129154 570434
rect 128918 563198 129154 563434
rect 128918 556198 129154 556434
rect 128918 549198 129154 549434
rect 128918 542198 129154 542434
rect 128918 535198 129154 535434
rect 128918 528198 129154 528434
rect 128918 521198 129154 521434
rect 128918 514198 129154 514434
rect 128918 507198 129154 507434
rect 128918 500198 129154 500434
rect 128918 493198 129154 493434
rect 128918 486198 129154 486434
rect 128918 479198 129154 479434
rect 128918 472198 129154 472434
rect 128918 465198 129154 465434
rect 128918 458198 129154 458434
rect 128918 451198 129154 451434
rect 128918 444198 129154 444434
rect 128918 437198 129154 437434
rect 128918 430198 129154 430434
rect 128918 423198 129154 423434
rect 128918 416198 129154 416434
rect 128918 409198 129154 409434
rect 128918 402198 129154 402434
rect 128918 395198 129154 395434
rect 128918 388198 129154 388434
rect 128918 381198 129154 381434
rect 128918 374198 129154 374434
rect 128918 367198 129154 367434
rect 128918 360198 129154 360434
rect 128918 353198 129154 353434
rect 128918 346198 129154 346434
rect 128918 339198 129154 339434
rect 128918 332198 129154 332434
rect 128918 325198 129154 325434
rect 128918 318198 129154 318434
rect 128918 311198 129154 311434
rect 128918 304198 129154 304434
rect 128918 297198 129154 297434
rect 128918 290198 129154 290434
rect 128918 283198 129154 283434
rect 128918 276198 129154 276434
rect 128918 269198 129154 269434
rect 128918 262198 129154 262434
rect 128918 255198 129154 255434
rect 128918 248198 129154 248434
rect 128918 241198 129154 241434
rect 128918 234198 129154 234434
rect 128918 227198 129154 227434
rect 128918 220198 129154 220434
rect 128918 213198 129154 213434
rect 128918 206198 129154 206434
rect 128918 199198 129154 199434
rect 128918 192198 129154 192434
rect 128918 185198 129154 185434
rect 128918 178198 129154 178434
rect 128918 171198 129154 171434
rect 128918 164198 129154 164434
rect 128918 157198 129154 157434
rect 128918 150198 129154 150434
rect 128918 143198 129154 143434
rect 128918 136198 129154 136434
rect 128918 129198 129154 129434
rect 128918 122198 129154 122434
rect 128918 115198 129154 115434
rect 128918 108198 129154 108434
rect 128918 101198 129154 101434
rect 128918 94198 129154 94434
rect 128918 87198 129154 87434
rect 128918 80198 129154 80434
rect 128918 73198 129154 73434
rect 128918 66198 129154 66434
rect 128918 59198 129154 59434
rect 128918 52198 129154 52434
rect 128918 45198 129154 45434
rect 128918 38198 129154 38434
rect 128918 31198 129154 31434
rect 128918 24198 129154 24434
rect 128918 17198 129154 17434
rect 128918 10198 129154 10434
rect 128918 3198 129154 3434
rect 128918 -1942 129154 -1706
rect 128918 -2262 129154 -2026
rect 134186 705002 134422 705238
rect 134186 704682 134422 704918
rect 134186 695258 134422 695494
rect 134186 688258 134422 688494
rect 134186 681258 134422 681494
rect 134186 674258 134422 674494
rect 134186 667258 134422 667494
rect 134186 660258 134422 660494
rect 134186 653258 134422 653494
rect 134186 646258 134422 646494
rect 134186 639258 134422 639494
rect 134186 632258 134422 632494
rect 134186 625258 134422 625494
rect 134186 618258 134422 618494
rect 134186 611258 134422 611494
rect 134186 604258 134422 604494
rect 134186 597258 134422 597494
rect 134186 590258 134422 590494
rect 134186 583258 134422 583494
rect 134186 576258 134422 576494
rect 134186 569258 134422 569494
rect 134186 562258 134422 562494
rect 134186 555258 134422 555494
rect 134186 548258 134422 548494
rect 134186 541258 134422 541494
rect 134186 534258 134422 534494
rect 134186 527258 134422 527494
rect 134186 520258 134422 520494
rect 134186 513258 134422 513494
rect 134186 506258 134422 506494
rect 134186 499258 134422 499494
rect 134186 492258 134422 492494
rect 134186 485258 134422 485494
rect 134186 478258 134422 478494
rect 134186 471258 134422 471494
rect 134186 464258 134422 464494
rect 134186 457258 134422 457494
rect 134186 450258 134422 450494
rect 134186 443258 134422 443494
rect 134186 436258 134422 436494
rect 134186 429258 134422 429494
rect 134186 422258 134422 422494
rect 134186 415258 134422 415494
rect 134186 408258 134422 408494
rect 134186 401258 134422 401494
rect 134186 394258 134422 394494
rect 134186 387258 134422 387494
rect 134186 380258 134422 380494
rect 134186 373258 134422 373494
rect 134186 366258 134422 366494
rect 134186 359258 134422 359494
rect 134186 352258 134422 352494
rect 134186 345258 134422 345494
rect 134186 338258 134422 338494
rect 134186 331258 134422 331494
rect 134186 324258 134422 324494
rect 134186 317258 134422 317494
rect 134186 310258 134422 310494
rect 134186 303258 134422 303494
rect 134186 296258 134422 296494
rect 134186 289258 134422 289494
rect 134186 282258 134422 282494
rect 134186 275258 134422 275494
rect 134186 268258 134422 268494
rect 134186 261258 134422 261494
rect 134186 254258 134422 254494
rect 134186 247258 134422 247494
rect 134186 240258 134422 240494
rect 134186 233258 134422 233494
rect 134186 226258 134422 226494
rect 134186 219258 134422 219494
rect 134186 212258 134422 212494
rect 134186 205258 134422 205494
rect 134186 198258 134422 198494
rect 134186 191258 134422 191494
rect 134186 184258 134422 184494
rect 134186 177258 134422 177494
rect 134186 170258 134422 170494
rect 134186 163258 134422 163494
rect 134186 156258 134422 156494
rect 134186 149258 134422 149494
rect 134186 142258 134422 142494
rect 134186 135258 134422 135494
rect 134186 128258 134422 128494
rect 134186 121258 134422 121494
rect 134186 114258 134422 114494
rect 134186 107258 134422 107494
rect 134186 100258 134422 100494
rect 134186 93258 134422 93494
rect 134186 86258 134422 86494
rect 134186 79258 134422 79494
rect 134186 72258 134422 72494
rect 134186 65258 134422 65494
rect 134186 58258 134422 58494
rect 134186 51258 134422 51494
rect 134186 44258 134422 44494
rect 134186 37258 134422 37494
rect 134186 30258 134422 30494
rect 134186 23258 134422 23494
rect 134186 16258 134422 16494
rect 134186 9258 134422 9494
rect 134186 2258 134422 2494
rect 134186 -982 134422 -746
rect 134186 -1302 134422 -1066
rect 135918 705962 136154 706198
rect 135918 705642 136154 705878
rect 135918 696198 136154 696434
rect 135918 689198 136154 689434
rect 135918 682198 136154 682434
rect 135918 675198 136154 675434
rect 135918 668198 136154 668434
rect 135918 661198 136154 661434
rect 135918 654198 136154 654434
rect 135918 647198 136154 647434
rect 135918 640198 136154 640434
rect 135918 633198 136154 633434
rect 135918 626198 136154 626434
rect 135918 619198 136154 619434
rect 135918 612198 136154 612434
rect 135918 605198 136154 605434
rect 135918 598198 136154 598434
rect 135918 591198 136154 591434
rect 135918 584198 136154 584434
rect 135918 577198 136154 577434
rect 135918 570198 136154 570434
rect 135918 563198 136154 563434
rect 135918 556198 136154 556434
rect 135918 549198 136154 549434
rect 135918 542198 136154 542434
rect 135918 535198 136154 535434
rect 135918 528198 136154 528434
rect 135918 521198 136154 521434
rect 135918 514198 136154 514434
rect 135918 507198 136154 507434
rect 135918 500198 136154 500434
rect 135918 493198 136154 493434
rect 135918 486198 136154 486434
rect 135918 479198 136154 479434
rect 135918 472198 136154 472434
rect 135918 465198 136154 465434
rect 135918 458198 136154 458434
rect 135918 451198 136154 451434
rect 135918 444198 136154 444434
rect 135918 437198 136154 437434
rect 135918 430198 136154 430434
rect 135918 423198 136154 423434
rect 135918 416198 136154 416434
rect 135918 409198 136154 409434
rect 135918 402198 136154 402434
rect 135918 395198 136154 395434
rect 135918 388198 136154 388434
rect 135918 381198 136154 381434
rect 135918 374198 136154 374434
rect 135918 367198 136154 367434
rect 135918 360198 136154 360434
rect 135918 353198 136154 353434
rect 135918 346198 136154 346434
rect 135918 339198 136154 339434
rect 135918 332198 136154 332434
rect 135918 325198 136154 325434
rect 135918 318198 136154 318434
rect 135918 311198 136154 311434
rect 135918 304198 136154 304434
rect 135918 297198 136154 297434
rect 135918 290198 136154 290434
rect 135918 283198 136154 283434
rect 135918 276198 136154 276434
rect 135918 269198 136154 269434
rect 135918 262198 136154 262434
rect 135918 255198 136154 255434
rect 135918 248198 136154 248434
rect 135918 241198 136154 241434
rect 135918 234198 136154 234434
rect 135918 227198 136154 227434
rect 135918 220198 136154 220434
rect 135918 213198 136154 213434
rect 135918 206198 136154 206434
rect 135918 199198 136154 199434
rect 135918 192198 136154 192434
rect 135918 185198 136154 185434
rect 135918 178198 136154 178434
rect 135918 171198 136154 171434
rect 135918 164198 136154 164434
rect 135918 157198 136154 157434
rect 135918 150198 136154 150434
rect 135918 143198 136154 143434
rect 135918 136198 136154 136434
rect 135918 129198 136154 129434
rect 135918 122198 136154 122434
rect 135918 115198 136154 115434
rect 135918 108198 136154 108434
rect 135918 101198 136154 101434
rect 135918 94198 136154 94434
rect 135918 87198 136154 87434
rect 135918 80198 136154 80434
rect 135918 73198 136154 73434
rect 135918 66198 136154 66434
rect 135918 59198 136154 59434
rect 135918 52198 136154 52434
rect 135918 45198 136154 45434
rect 135918 38198 136154 38434
rect 135918 31198 136154 31434
rect 135918 24198 136154 24434
rect 135918 17198 136154 17434
rect 135918 10198 136154 10434
rect 135918 3198 136154 3434
rect 135918 -1942 136154 -1706
rect 135918 -2262 136154 -2026
rect 141186 705002 141422 705238
rect 141186 704682 141422 704918
rect 141186 695258 141422 695494
rect 141186 688258 141422 688494
rect 141186 681258 141422 681494
rect 141186 674258 141422 674494
rect 141186 667258 141422 667494
rect 141186 660258 141422 660494
rect 141186 653258 141422 653494
rect 141186 646258 141422 646494
rect 141186 639258 141422 639494
rect 141186 632258 141422 632494
rect 141186 625258 141422 625494
rect 141186 618258 141422 618494
rect 141186 611258 141422 611494
rect 141186 604258 141422 604494
rect 141186 597258 141422 597494
rect 141186 590258 141422 590494
rect 141186 583258 141422 583494
rect 141186 576258 141422 576494
rect 141186 569258 141422 569494
rect 141186 562258 141422 562494
rect 141186 555258 141422 555494
rect 141186 548258 141422 548494
rect 141186 541258 141422 541494
rect 141186 534258 141422 534494
rect 141186 527258 141422 527494
rect 141186 520258 141422 520494
rect 141186 513258 141422 513494
rect 141186 506258 141422 506494
rect 141186 499258 141422 499494
rect 141186 492258 141422 492494
rect 141186 485258 141422 485494
rect 141186 478258 141422 478494
rect 141186 471258 141422 471494
rect 141186 464258 141422 464494
rect 141186 457258 141422 457494
rect 141186 450258 141422 450494
rect 141186 443258 141422 443494
rect 141186 436258 141422 436494
rect 141186 429258 141422 429494
rect 141186 422258 141422 422494
rect 141186 415258 141422 415494
rect 141186 408258 141422 408494
rect 141186 401258 141422 401494
rect 141186 394258 141422 394494
rect 141186 387258 141422 387494
rect 141186 380258 141422 380494
rect 141186 373258 141422 373494
rect 141186 366258 141422 366494
rect 141186 359258 141422 359494
rect 141186 352258 141422 352494
rect 141186 345258 141422 345494
rect 141186 338258 141422 338494
rect 141186 331258 141422 331494
rect 141186 324258 141422 324494
rect 141186 317258 141422 317494
rect 141186 310258 141422 310494
rect 141186 303258 141422 303494
rect 141186 296258 141422 296494
rect 141186 289258 141422 289494
rect 141186 282258 141422 282494
rect 141186 275258 141422 275494
rect 141186 268258 141422 268494
rect 141186 261258 141422 261494
rect 141186 254258 141422 254494
rect 141186 247258 141422 247494
rect 141186 240258 141422 240494
rect 141186 233258 141422 233494
rect 141186 226258 141422 226494
rect 141186 219258 141422 219494
rect 141186 212258 141422 212494
rect 141186 205258 141422 205494
rect 141186 198258 141422 198494
rect 141186 191258 141422 191494
rect 141186 184258 141422 184494
rect 141186 177258 141422 177494
rect 141186 170258 141422 170494
rect 141186 163258 141422 163494
rect 141186 156258 141422 156494
rect 141186 149258 141422 149494
rect 141186 142258 141422 142494
rect 141186 135258 141422 135494
rect 141186 128258 141422 128494
rect 141186 121258 141422 121494
rect 141186 114258 141422 114494
rect 141186 107258 141422 107494
rect 141186 100258 141422 100494
rect 141186 93258 141422 93494
rect 141186 86258 141422 86494
rect 141186 79258 141422 79494
rect 141186 72258 141422 72494
rect 141186 65258 141422 65494
rect 141186 58258 141422 58494
rect 141186 51258 141422 51494
rect 141186 44258 141422 44494
rect 141186 37258 141422 37494
rect 141186 30258 141422 30494
rect 141186 23258 141422 23494
rect 141186 16258 141422 16494
rect 141186 9258 141422 9494
rect 141186 2258 141422 2494
rect 141186 -982 141422 -746
rect 141186 -1302 141422 -1066
rect 142918 705962 143154 706198
rect 142918 705642 143154 705878
rect 142918 696198 143154 696434
rect 142918 689198 143154 689434
rect 142918 682198 143154 682434
rect 142918 675198 143154 675434
rect 142918 668198 143154 668434
rect 142918 661198 143154 661434
rect 142918 654198 143154 654434
rect 142918 647198 143154 647434
rect 142918 640198 143154 640434
rect 142918 633198 143154 633434
rect 142918 626198 143154 626434
rect 142918 619198 143154 619434
rect 142918 612198 143154 612434
rect 142918 605198 143154 605434
rect 142918 598198 143154 598434
rect 142918 591198 143154 591434
rect 142918 584198 143154 584434
rect 142918 577198 143154 577434
rect 142918 570198 143154 570434
rect 142918 563198 143154 563434
rect 142918 556198 143154 556434
rect 142918 549198 143154 549434
rect 142918 542198 143154 542434
rect 142918 535198 143154 535434
rect 142918 528198 143154 528434
rect 142918 521198 143154 521434
rect 142918 514198 143154 514434
rect 142918 507198 143154 507434
rect 142918 500198 143154 500434
rect 142918 493198 143154 493434
rect 142918 486198 143154 486434
rect 142918 479198 143154 479434
rect 142918 472198 143154 472434
rect 142918 465198 143154 465434
rect 142918 458198 143154 458434
rect 142918 451198 143154 451434
rect 142918 444198 143154 444434
rect 142918 437198 143154 437434
rect 142918 430198 143154 430434
rect 142918 423198 143154 423434
rect 142918 416198 143154 416434
rect 142918 409198 143154 409434
rect 142918 402198 143154 402434
rect 142918 395198 143154 395434
rect 142918 388198 143154 388434
rect 142918 381198 143154 381434
rect 142918 374198 143154 374434
rect 142918 367198 143154 367434
rect 142918 360198 143154 360434
rect 142918 353198 143154 353434
rect 142918 346198 143154 346434
rect 142918 339198 143154 339434
rect 142918 332198 143154 332434
rect 142918 325198 143154 325434
rect 142918 318198 143154 318434
rect 142918 311198 143154 311434
rect 142918 304198 143154 304434
rect 142918 297198 143154 297434
rect 142918 290198 143154 290434
rect 142918 283198 143154 283434
rect 142918 276198 143154 276434
rect 142918 269198 143154 269434
rect 142918 262198 143154 262434
rect 142918 255198 143154 255434
rect 142918 248198 143154 248434
rect 142918 241198 143154 241434
rect 142918 234198 143154 234434
rect 142918 227198 143154 227434
rect 142918 220198 143154 220434
rect 142918 213198 143154 213434
rect 142918 206198 143154 206434
rect 142918 199198 143154 199434
rect 142918 192198 143154 192434
rect 142918 185198 143154 185434
rect 142918 178198 143154 178434
rect 142918 171198 143154 171434
rect 142918 164198 143154 164434
rect 142918 157198 143154 157434
rect 142918 150198 143154 150434
rect 142918 143198 143154 143434
rect 142918 136198 143154 136434
rect 142918 129198 143154 129434
rect 142918 122198 143154 122434
rect 142918 115198 143154 115434
rect 142918 108198 143154 108434
rect 142918 101198 143154 101434
rect 142918 94198 143154 94434
rect 142918 87198 143154 87434
rect 142918 80198 143154 80434
rect 142918 73198 143154 73434
rect 142918 66198 143154 66434
rect 142918 59198 143154 59434
rect 142918 52198 143154 52434
rect 142918 45198 143154 45434
rect 142918 38198 143154 38434
rect 142918 31198 143154 31434
rect 142918 24198 143154 24434
rect 142918 17198 143154 17434
rect 142918 10198 143154 10434
rect 142918 3198 143154 3434
rect 142918 -1942 143154 -1706
rect 142918 -2262 143154 -2026
rect 148186 705002 148422 705238
rect 148186 704682 148422 704918
rect 148186 695258 148422 695494
rect 148186 688258 148422 688494
rect 148186 681258 148422 681494
rect 148186 674258 148422 674494
rect 148186 667258 148422 667494
rect 148186 660258 148422 660494
rect 148186 653258 148422 653494
rect 148186 646258 148422 646494
rect 148186 639258 148422 639494
rect 148186 632258 148422 632494
rect 148186 625258 148422 625494
rect 148186 618258 148422 618494
rect 148186 611258 148422 611494
rect 148186 604258 148422 604494
rect 148186 597258 148422 597494
rect 148186 590258 148422 590494
rect 148186 583258 148422 583494
rect 148186 576258 148422 576494
rect 148186 569258 148422 569494
rect 148186 562258 148422 562494
rect 148186 555258 148422 555494
rect 148186 548258 148422 548494
rect 148186 541258 148422 541494
rect 148186 534258 148422 534494
rect 148186 527258 148422 527494
rect 148186 520258 148422 520494
rect 148186 513258 148422 513494
rect 148186 506258 148422 506494
rect 148186 499258 148422 499494
rect 148186 492258 148422 492494
rect 148186 485258 148422 485494
rect 148186 478258 148422 478494
rect 148186 471258 148422 471494
rect 148186 464258 148422 464494
rect 148186 457258 148422 457494
rect 148186 450258 148422 450494
rect 148186 443258 148422 443494
rect 148186 436258 148422 436494
rect 148186 429258 148422 429494
rect 148186 422258 148422 422494
rect 148186 415258 148422 415494
rect 148186 408258 148422 408494
rect 148186 401258 148422 401494
rect 148186 394258 148422 394494
rect 148186 387258 148422 387494
rect 148186 380258 148422 380494
rect 148186 373258 148422 373494
rect 148186 366258 148422 366494
rect 148186 359258 148422 359494
rect 148186 352258 148422 352494
rect 148186 345258 148422 345494
rect 148186 338258 148422 338494
rect 148186 331258 148422 331494
rect 148186 324258 148422 324494
rect 148186 317258 148422 317494
rect 148186 310258 148422 310494
rect 148186 303258 148422 303494
rect 148186 296258 148422 296494
rect 148186 289258 148422 289494
rect 148186 282258 148422 282494
rect 148186 275258 148422 275494
rect 148186 268258 148422 268494
rect 148186 261258 148422 261494
rect 148186 254258 148422 254494
rect 148186 247258 148422 247494
rect 148186 240258 148422 240494
rect 148186 233258 148422 233494
rect 148186 226258 148422 226494
rect 148186 219258 148422 219494
rect 148186 212258 148422 212494
rect 148186 205258 148422 205494
rect 148186 198258 148422 198494
rect 148186 191258 148422 191494
rect 148186 184258 148422 184494
rect 148186 177258 148422 177494
rect 148186 170258 148422 170494
rect 148186 163258 148422 163494
rect 148186 156258 148422 156494
rect 148186 149258 148422 149494
rect 148186 142258 148422 142494
rect 148186 135258 148422 135494
rect 148186 128258 148422 128494
rect 148186 121258 148422 121494
rect 148186 114258 148422 114494
rect 148186 107258 148422 107494
rect 148186 100258 148422 100494
rect 148186 93258 148422 93494
rect 148186 86258 148422 86494
rect 148186 79258 148422 79494
rect 148186 72258 148422 72494
rect 148186 65258 148422 65494
rect 148186 58258 148422 58494
rect 148186 51258 148422 51494
rect 148186 44258 148422 44494
rect 148186 37258 148422 37494
rect 148186 30258 148422 30494
rect 148186 23258 148422 23494
rect 148186 16258 148422 16494
rect 148186 9258 148422 9494
rect 148186 2258 148422 2494
rect 148186 -982 148422 -746
rect 148186 -1302 148422 -1066
rect 149918 705962 150154 706198
rect 149918 705642 150154 705878
rect 149918 696198 150154 696434
rect 149918 689198 150154 689434
rect 149918 682198 150154 682434
rect 149918 675198 150154 675434
rect 149918 668198 150154 668434
rect 149918 661198 150154 661434
rect 149918 654198 150154 654434
rect 149918 647198 150154 647434
rect 149918 640198 150154 640434
rect 149918 633198 150154 633434
rect 149918 626198 150154 626434
rect 149918 619198 150154 619434
rect 149918 612198 150154 612434
rect 149918 605198 150154 605434
rect 149918 598198 150154 598434
rect 149918 591198 150154 591434
rect 149918 584198 150154 584434
rect 149918 577198 150154 577434
rect 149918 570198 150154 570434
rect 149918 563198 150154 563434
rect 149918 556198 150154 556434
rect 149918 549198 150154 549434
rect 149918 542198 150154 542434
rect 149918 535198 150154 535434
rect 149918 528198 150154 528434
rect 149918 521198 150154 521434
rect 149918 514198 150154 514434
rect 149918 507198 150154 507434
rect 149918 500198 150154 500434
rect 149918 493198 150154 493434
rect 149918 486198 150154 486434
rect 149918 479198 150154 479434
rect 149918 472198 150154 472434
rect 149918 465198 150154 465434
rect 149918 458198 150154 458434
rect 149918 451198 150154 451434
rect 149918 444198 150154 444434
rect 149918 437198 150154 437434
rect 149918 430198 150154 430434
rect 149918 423198 150154 423434
rect 149918 416198 150154 416434
rect 149918 409198 150154 409434
rect 149918 402198 150154 402434
rect 149918 395198 150154 395434
rect 149918 388198 150154 388434
rect 149918 381198 150154 381434
rect 149918 374198 150154 374434
rect 149918 367198 150154 367434
rect 149918 360198 150154 360434
rect 149918 353198 150154 353434
rect 149918 346198 150154 346434
rect 149918 339198 150154 339434
rect 149918 332198 150154 332434
rect 149918 325198 150154 325434
rect 149918 318198 150154 318434
rect 149918 311198 150154 311434
rect 149918 304198 150154 304434
rect 149918 297198 150154 297434
rect 149918 290198 150154 290434
rect 149918 283198 150154 283434
rect 149918 276198 150154 276434
rect 149918 269198 150154 269434
rect 149918 262198 150154 262434
rect 149918 255198 150154 255434
rect 149918 248198 150154 248434
rect 149918 241198 150154 241434
rect 149918 234198 150154 234434
rect 149918 227198 150154 227434
rect 149918 220198 150154 220434
rect 149918 213198 150154 213434
rect 149918 206198 150154 206434
rect 149918 199198 150154 199434
rect 149918 192198 150154 192434
rect 149918 185198 150154 185434
rect 149918 178198 150154 178434
rect 149918 171198 150154 171434
rect 149918 164198 150154 164434
rect 149918 157198 150154 157434
rect 149918 150198 150154 150434
rect 149918 143198 150154 143434
rect 149918 136198 150154 136434
rect 149918 129198 150154 129434
rect 149918 122198 150154 122434
rect 149918 115198 150154 115434
rect 149918 108198 150154 108434
rect 149918 101198 150154 101434
rect 149918 94198 150154 94434
rect 149918 87198 150154 87434
rect 149918 80198 150154 80434
rect 149918 73198 150154 73434
rect 149918 66198 150154 66434
rect 149918 59198 150154 59434
rect 149918 52198 150154 52434
rect 149918 45198 150154 45434
rect 149918 38198 150154 38434
rect 149918 31198 150154 31434
rect 149918 24198 150154 24434
rect 149918 17198 150154 17434
rect 149918 10198 150154 10434
rect 149918 3198 150154 3434
rect 149918 -1942 150154 -1706
rect 149918 -2262 150154 -2026
rect 155186 705002 155422 705238
rect 155186 704682 155422 704918
rect 155186 695258 155422 695494
rect 155186 688258 155422 688494
rect 155186 681258 155422 681494
rect 155186 674258 155422 674494
rect 155186 667258 155422 667494
rect 155186 660258 155422 660494
rect 155186 653258 155422 653494
rect 155186 646258 155422 646494
rect 155186 639258 155422 639494
rect 155186 632258 155422 632494
rect 155186 625258 155422 625494
rect 155186 618258 155422 618494
rect 155186 611258 155422 611494
rect 155186 604258 155422 604494
rect 155186 597258 155422 597494
rect 155186 590258 155422 590494
rect 155186 583258 155422 583494
rect 155186 576258 155422 576494
rect 155186 569258 155422 569494
rect 155186 562258 155422 562494
rect 155186 555258 155422 555494
rect 155186 548258 155422 548494
rect 155186 541258 155422 541494
rect 155186 534258 155422 534494
rect 155186 527258 155422 527494
rect 155186 520258 155422 520494
rect 155186 513258 155422 513494
rect 155186 506258 155422 506494
rect 155186 499258 155422 499494
rect 155186 492258 155422 492494
rect 155186 485258 155422 485494
rect 155186 478258 155422 478494
rect 155186 471258 155422 471494
rect 155186 464258 155422 464494
rect 155186 457258 155422 457494
rect 155186 450258 155422 450494
rect 155186 443258 155422 443494
rect 155186 436258 155422 436494
rect 155186 429258 155422 429494
rect 155186 422258 155422 422494
rect 155186 415258 155422 415494
rect 155186 408258 155422 408494
rect 155186 401258 155422 401494
rect 155186 394258 155422 394494
rect 155186 387258 155422 387494
rect 155186 380258 155422 380494
rect 155186 373258 155422 373494
rect 155186 366258 155422 366494
rect 155186 359258 155422 359494
rect 155186 352258 155422 352494
rect 155186 345258 155422 345494
rect 155186 338258 155422 338494
rect 155186 331258 155422 331494
rect 155186 324258 155422 324494
rect 155186 317258 155422 317494
rect 155186 310258 155422 310494
rect 155186 303258 155422 303494
rect 155186 296258 155422 296494
rect 155186 289258 155422 289494
rect 155186 282258 155422 282494
rect 155186 275258 155422 275494
rect 155186 268258 155422 268494
rect 155186 261258 155422 261494
rect 155186 254258 155422 254494
rect 155186 247258 155422 247494
rect 155186 240258 155422 240494
rect 155186 233258 155422 233494
rect 155186 226258 155422 226494
rect 155186 219258 155422 219494
rect 155186 212258 155422 212494
rect 155186 205258 155422 205494
rect 155186 198258 155422 198494
rect 155186 191258 155422 191494
rect 155186 184258 155422 184494
rect 155186 177258 155422 177494
rect 155186 170258 155422 170494
rect 155186 163258 155422 163494
rect 155186 156258 155422 156494
rect 155186 149258 155422 149494
rect 155186 142258 155422 142494
rect 155186 135258 155422 135494
rect 155186 128258 155422 128494
rect 155186 121258 155422 121494
rect 155186 114258 155422 114494
rect 155186 107258 155422 107494
rect 155186 100258 155422 100494
rect 155186 93258 155422 93494
rect 155186 86258 155422 86494
rect 155186 79258 155422 79494
rect 155186 72258 155422 72494
rect 155186 65258 155422 65494
rect 155186 58258 155422 58494
rect 155186 51258 155422 51494
rect 155186 44258 155422 44494
rect 155186 37258 155422 37494
rect 155186 30258 155422 30494
rect 155186 23258 155422 23494
rect 155186 16258 155422 16494
rect 155186 9258 155422 9494
rect 155186 2258 155422 2494
rect 155186 -982 155422 -746
rect 155186 -1302 155422 -1066
rect 156918 705962 157154 706198
rect 156918 705642 157154 705878
rect 156918 696198 157154 696434
rect 156918 689198 157154 689434
rect 156918 682198 157154 682434
rect 156918 675198 157154 675434
rect 156918 668198 157154 668434
rect 156918 661198 157154 661434
rect 156918 654198 157154 654434
rect 156918 647198 157154 647434
rect 156918 640198 157154 640434
rect 156918 633198 157154 633434
rect 156918 626198 157154 626434
rect 156918 619198 157154 619434
rect 156918 612198 157154 612434
rect 156918 605198 157154 605434
rect 156918 598198 157154 598434
rect 156918 591198 157154 591434
rect 156918 584198 157154 584434
rect 156918 577198 157154 577434
rect 156918 570198 157154 570434
rect 156918 563198 157154 563434
rect 156918 556198 157154 556434
rect 156918 549198 157154 549434
rect 156918 542198 157154 542434
rect 156918 535198 157154 535434
rect 156918 528198 157154 528434
rect 156918 521198 157154 521434
rect 156918 514198 157154 514434
rect 156918 507198 157154 507434
rect 156918 500198 157154 500434
rect 156918 493198 157154 493434
rect 156918 486198 157154 486434
rect 156918 479198 157154 479434
rect 156918 472198 157154 472434
rect 156918 465198 157154 465434
rect 156918 458198 157154 458434
rect 156918 451198 157154 451434
rect 156918 444198 157154 444434
rect 156918 437198 157154 437434
rect 156918 430198 157154 430434
rect 156918 423198 157154 423434
rect 156918 416198 157154 416434
rect 156918 409198 157154 409434
rect 156918 402198 157154 402434
rect 156918 395198 157154 395434
rect 156918 388198 157154 388434
rect 156918 381198 157154 381434
rect 156918 374198 157154 374434
rect 156918 367198 157154 367434
rect 156918 360198 157154 360434
rect 156918 353198 157154 353434
rect 156918 346198 157154 346434
rect 156918 339198 157154 339434
rect 156918 332198 157154 332434
rect 156918 325198 157154 325434
rect 156918 318198 157154 318434
rect 156918 311198 157154 311434
rect 156918 304198 157154 304434
rect 156918 297198 157154 297434
rect 156918 290198 157154 290434
rect 156918 283198 157154 283434
rect 156918 276198 157154 276434
rect 156918 269198 157154 269434
rect 156918 262198 157154 262434
rect 156918 255198 157154 255434
rect 156918 248198 157154 248434
rect 156918 241198 157154 241434
rect 156918 234198 157154 234434
rect 156918 227198 157154 227434
rect 156918 220198 157154 220434
rect 156918 213198 157154 213434
rect 156918 206198 157154 206434
rect 156918 199198 157154 199434
rect 156918 192198 157154 192434
rect 156918 185198 157154 185434
rect 156918 178198 157154 178434
rect 156918 171198 157154 171434
rect 156918 164198 157154 164434
rect 156918 157198 157154 157434
rect 156918 150198 157154 150434
rect 156918 143198 157154 143434
rect 156918 136198 157154 136434
rect 156918 129198 157154 129434
rect 156918 122198 157154 122434
rect 156918 115198 157154 115434
rect 156918 108198 157154 108434
rect 156918 101198 157154 101434
rect 156918 94198 157154 94434
rect 156918 87198 157154 87434
rect 156918 80198 157154 80434
rect 156918 73198 157154 73434
rect 156918 66198 157154 66434
rect 156918 59198 157154 59434
rect 156918 52198 157154 52434
rect 156918 45198 157154 45434
rect 156918 38198 157154 38434
rect 156918 31198 157154 31434
rect 156918 24198 157154 24434
rect 156918 17198 157154 17434
rect 156918 10198 157154 10434
rect 156918 3198 157154 3434
rect 156918 -1942 157154 -1706
rect 156918 -2262 157154 -2026
rect 162186 705002 162422 705238
rect 162186 704682 162422 704918
rect 162186 695258 162422 695494
rect 162186 688258 162422 688494
rect 162186 681258 162422 681494
rect 162186 674258 162422 674494
rect 162186 667258 162422 667494
rect 162186 660258 162422 660494
rect 162186 653258 162422 653494
rect 162186 646258 162422 646494
rect 162186 639258 162422 639494
rect 162186 632258 162422 632494
rect 162186 625258 162422 625494
rect 162186 618258 162422 618494
rect 162186 611258 162422 611494
rect 162186 604258 162422 604494
rect 162186 597258 162422 597494
rect 162186 590258 162422 590494
rect 162186 583258 162422 583494
rect 162186 576258 162422 576494
rect 162186 569258 162422 569494
rect 162186 562258 162422 562494
rect 162186 555258 162422 555494
rect 162186 548258 162422 548494
rect 162186 541258 162422 541494
rect 162186 534258 162422 534494
rect 162186 527258 162422 527494
rect 162186 520258 162422 520494
rect 162186 513258 162422 513494
rect 162186 506258 162422 506494
rect 162186 499258 162422 499494
rect 162186 492258 162422 492494
rect 162186 485258 162422 485494
rect 162186 478258 162422 478494
rect 162186 471258 162422 471494
rect 162186 464258 162422 464494
rect 162186 457258 162422 457494
rect 162186 450258 162422 450494
rect 162186 443258 162422 443494
rect 162186 436258 162422 436494
rect 162186 429258 162422 429494
rect 162186 422258 162422 422494
rect 162186 415258 162422 415494
rect 162186 408258 162422 408494
rect 162186 401258 162422 401494
rect 162186 394258 162422 394494
rect 162186 387258 162422 387494
rect 162186 380258 162422 380494
rect 162186 373258 162422 373494
rect 162186 366258 162422 366494
rect 162186 359258 162422 359494
rect 162186 352258 162422 352494
rect 162186 345258 162422 345494
rect 162186 338258 162422 338494
rect 162186 331258 162422 331494
rect 162186 324258 162422 324494
rect 162186 317258 162422 317494
rect 162186 310258 162422 310494
rect 162186 303258 162422 303494
rect 162186 296258 162422 296494
rect 162186 289258 162422 289494
rect 162186 282258 162422 282494
rect 162186 275258 162422 275494
rect 162186 268258 162422 268494
rect 162186 261258 162422 261494
rect 162186 254258 162422 254494
rect 162186 247258 162422 247494
rect 162186 240258 162422 240494
rect 162186 233258 162422 233494
rect 162186 226258 162422 226494
rect 162186 219258 162422 219494
rect 162186 212258 162422 212494
rect 162186 205258 162422 205494
rect 162186 198258 162422 198494
rect 162186 191258 162422 191494
rect 162186 184258 162422 184494
rect 162186 177258 162422 177494
rect 162186 170258 162422 170494
rect 162186 163258 162422 163494
rect 162186 156258 162422 156494
rect 162186 149258 162422 149494
rect 162186 142258 162422 142494
rect 162186 135258 162422 135494
rect 162186 128258 162422 128494
rect 162186 121258 162422 121494
rect 162186 114258 162422 114494
rect 162186 107258 162422 107494
rect 162186 100258 162422 100494
rect 162186 93258 162422 93494
rect 162186 86258 162422 86494
rect 162186 79258 162422 79494
rect 162186 72258 162422 72494
rect 162186 65258 162422 65494
rect 162186 58258 162422 58494
rect 162186 51258 162422 51494
rect 162186 44258 162422 44494
rect 162186 37258 162422 37494
rect 162186 30258 162422 30494
rect 162186 23258 162422 23494
rect 162186 16258 162422 16494
rect 162186 9258 162422 9494
rect 162186 2258 162422 2494
rect 162186 -982 162422 -746
rect 162186 -1302 162422 -1066
rect 163918 705962 164154 706198
rect 163918 705642 164154 705878
rect 163918 696198 164154 696434
rect 163918 689198 164154 689434
rect 163918 682198 164154 682434
rect 163918 675198 164154 675434
rect 163918 668198 164154 668434
rect 163918 661198 164154 661434
rect 163918 654198 164154 654434
rect 163918 647198 164154 647434
rect 163918 640198 164154 640434
rect 163918 633198 164154 633434
rect 163918 626198 164154 626434
rect 163918 619198 164154 619434
rect 163918 612198 164154 612434
rect 163918 605198 164154 605434
rect 163918 598198 164154 598434
rect 163918 591198 164154 591434
rect 163918 584198 164154 584434
rect 163918 577198 164154 577434
rect 163918 570198 164154 570434
rect 163918 563198 164154 563434
rect 163918 556198 164154 556434
rect 163918 549198 164154 549434
rect 163918 542198 164154 542434
rect 163918 535198 164154 535434
rect 163918 528198 164154 528434
rect 163918 521198 164154 521434
rect 163918 514198 164154 514434
rect 163918 507198 164154 507434
rect 163918 500198 164154 500434
rect 163918 493198 164154 493434
rect 163918 486198 164154 486434
rect 163918 479198 164154 479434
rect 163918 472198 164154 472434
rect 163918 465198 164154 465434
rect 163918 458198 164154 458434
rect 163918 451198 164154 451434
rect 163918 444198 164154 444434
rect 163918 437198 164154 437434
rect 163918 430198 164154 430434
rect 163918 423198 164154 423434
rect 163918 416198 164154 416434
rect 163918 409198 164154 409434
rect 163918 402198 164154 402434
rect 163918 395198 164154 395434
rect 163918 388198 164154 388434
rect 163918 381198 164154 381434
rect 163918 374198 164154 374434
rect 163918 367198 164154 367434
rect 163918 360198 164154 360434
rect 163918 353198 164154 353434
rect 163918 346198 164154 346434
rect 163918 339198 164154 339434
rect 163918 332198 164154 332434
rect 163918 325198 164154 325434
rect 163918 318198 164154 318434
rect 163918 311198 164154 311434
rect 163918 304198 164154 304434
rect 163918 297198 164154 297434
rect 163918 290198 164154 290434
rect 163918 283198 164154 283434
rect 163918 276198 164154 276434
rect 163918 269198 164154 269434
rect 163918 262198 164154 262434
rect 163918 255198 164154 255434
rect 163918 248198 164154 248434
rect 163918 241198 164154 241434
rect 163918 234198 164154 234434
rect 163918 227198 164154 227434
rect 163918 220198 164154 220434
rect 163918 213198 164154 213434
rect 163918 206198 164154 206434
rect 163918 199198 164154 199434
rect 163918 192198 164154 192434
rect 163918 185198 164154 185434
rect 163918 178198 164154 178434
rect 163918 171198 164154 171434
rect 163918 164198 164154 164434
rect 163918 157198 164154 157434
rect 163918 150198 164154 150434
rect 163918 143198 164154 143434
rect 163918 136198 164154 136434
rect 163918 129198 164154 129434
rect 163918 122198 164154 122434
rect 163918 115198 164154 115434
rect 163918 108198 164154 108434
rect 163918 101198 164154 101434
rect 163918 94198 164154 94434
rect 163918 87198 164154 87434
rect 163918 80198 164154 80434
rect 163918 73198 164154 73434
rect 163918 66198 164154 66434
rect 163918 59198 164154 59434
rect 163918 52198 164154 52434
rect 163918 45198 164154 45434
rect 163918 38198 164154 38434
rect 163918 31198 164154 31434
rect 163918 24198 164154 24434
rect 163918 17198 164154 17434
rect 163918 10198 164154 10434
rect 163918 3198 164154 3434
rect 163918 -1942 164154 -1706
rect 163918 -2262 164154 -2026
rect 169186 705002 169422 705238
rect 169186 704682 169422 704918
rect 169186 695258 169422 695494
rect 169186 688258 169422 688494
rect 169186 681258 169422 681494
rect 169186 674258 169422 674494
rect 169186 667258 169422 667494
rect 169186 660258 169422 660494
rect 169186 653258 169422 653494
rect 169186 646258 169422 646494
rect 169186 639258 169422 639494
rect 169186 632258 169422 632494
rect 169186 625258 169422 625494
rect 169186 618258 169422 618494
rect 169186 611258 169422 611494
rect 169186 604258 169422 604494
rect 169186 597258 169422 597494
rect 169186 590258 169422 590494
rect 169186 583258 169422 583494
rect 169186 576258 169422 576494
rect 169186 569258 169422 569494
rect 169186 562258 169422 562494
rect 169186 555258 169422 555494
rect 169186 548258 169422 548494
rect 169186 541258 169422 541494
rect 169186 534258 169422 534494
rect 169186 527258 169422 527494
rect 169186 520258 169422 520494
rect 169186 513258 169422 513494
rect 169186 506258 169422 506494
rect 169186 499258 169422 499494
rect 169186 492258 169422 492494
rect 169186 485258 169422 485494
rect 169186 478258 169422 478494
rect 169186 471258 169422 471494
rect 169186 464258 169422 464494
rect 169186 457258 169422 457494
rect 169186 450258 169422 450494
rect 169186 443258 169422 443494
rect 169186 436258 169422 436494
rect 169186 429258 169422 429494
rect 169186 422258 169422 422494
rect 169186 415258 169422 415494
rect 169186 408258 169422 408494
rect 169186 401258 169422 401494
rect 169186 394258 169422 394494
rect 169186 387258 169422 387494
rect 169186 380258 169422 380494
rect 169186 373258 169422 373494
rect 169186 366258 169422 366494
rect 169186 359258 169422 359494
rect 169186 352258 169422 352494
rect 169186 345258 169422 345494
rect 169186 338258 169422 338494
rect 169186 331258 169422 331494
rect 169186 324258 169422 324494
rect 169186 317258 169422 317494
rect 169186 310258 169422 310494
rect 169186 303258 169422 303494
rect 169186 296258 169422 296494
rect 169186 289258 169422 289494
rect 169186 282258 169422 282494
rect 169186 275258 169422 275494
rect 169186 268258 169422 268494
rect 169186 261258 169422 261494
rect 169186 254258 169422 254494
rect 169186 247258 169422 247494
rect 169186 240258 169422 240494
rect 169186 233258 169422 233494
rect 169186 226258 169422 226494
rect 169186 219258 169422 219494
rect 169186 212258 169422 212494
rect 169186 205258 169422 205494
rect 169186 198258 169422 198494
rect 169186 191258 169422 191494
rect 169186 184258 169422 184494
rect 169186 177258 169422 177494
rect 169186 170258 169422 170494
rect 169186 163258 169422 163494
rect 169186 156258 169422 156494
rect 169186 149258 169422 149494
rect 169186 142258 169422 142494
rect 169186 135258 169422 135494
rect 169186 128258 169422 128494
rect 169186 121258 169422 121494
rect 169186 114258 169422 114494
rect 169186 107258 169422 107494
rect 169186 100258 169422 100494
rect 169186 93258 169422 93494
rect 169186 86258 169422 86494
rect 169186 79258 169422 79494
rect 169186 72258 169422 72494
rect 169186 65258 169422 65494
rect 169186 58258 169422 58494
rect 169186 51258 169422 51494
rect 169186 44258 169422 44494
rect 169186 37258 169422 37494
rect 169186 30258 169422 30494
rect 169186 23258 169422 23494
rect 169186 16258 169422 16494
rect 169186 9258 169422 9494
rect 169186 2258 169422 2494
rect 169186 -982 169422 -746
rect 169186 -1302 169422 -1066
rect 170918 705962 171154 706198
rect 170918 705642 171154 705878
rect 170918 696198 171154 696434
rect 170918 689198 171154 689434
rect 170918 682198 171154 682434
rect 170918 675198 171154 675434
rect 170918 668198 171154 668434
rect 170918 661198 171154 661434
rect 170918 654198 171154 654434
rect 170918 647198 171154 647434
rect 170918 640198 171154 640434
rect 170918 633198 171154 633434
rect 170918 626198 171154 626434
rect 170918 619198 171154 619434
rect 170918 612198 171154 612434
rect 170918 605198 171154 605434
rect 170918 598198 171154 598434
rect 170918 591198 171154 591434
rect 170918 584198 171154 584434
rect 170918 577198 171154 577434
rect 170918 570198 171154 570434
rect 170918 563198 171154 563434
rect 170918 556198 171154 556434
rect 170918 549198 171154 549434
rect 170918 542198 171154 542434
rect 170918 535198 171154 535434
rect 170918 528198 171154 528434
rect 170918 521198 171154 521434
rect 170918 514198 171154 514434
rect 170918 507198 171154 507434
rect 170918 500198 171154 500434
rect 170918 493198 171154 493434
rect 170918 486198 171154 486434
rect 170918 479198 171154 479434
rect 170918 472198 171154 472434
rect 170918 465198 171154 465434
rect 170918 458198 171154 458434
rect 170918 451198 171154 451434
rect 170918 444198 171154 444434
rect 170918 437198 171154 437434
rect 170918 430198 171154 430434
rect 170918 423198 171154 423434
rect 170918 416198 171154 416434
rect 170918 409198 171154 409434
rect 170918 402198 171154 402434
rect 170918 395198 171154 395434
rect 170918 388198 171154 388434
rect 170918 381198 171154 381434
rect 170918 374198 171154 374434
rect 170918 367198 171154 367434
rect 170918 360198 171154 360434
rect 170918 353198 171154 353434
rect 170918 346198 171154 346434
rect 170918 339198 171154 339434
rect 170918 332198 171154 332434
rect 170918 325198 171154 325434
rect 170918 318198 171154 318434
rect 170918 311198 171154 311434
rect 170918 304198 171154 304434
rect 170918 297198 171154 297434
rect 170918 290198 171154 290434
rect 170918 283198 171154 283434
rect 170918 276198 171154 276434
rect 170918 269198 171154 269434
rect 170918 262198 171154 262434
rect 170918 255198 171154 255434
rect 170918 248198 171154 248434
rect 170918 241198 171154 241434
rect 170918 234198 171154 234434
rect 170918 227198 171154 227434
rect 170918 220198 171154 220434
rect 170918 213198 171154 213434
rect 170918 206198 171154 206434
rect 170918 199198 171154 199434
rect 170918 192198 171154 192434
rect 170918 185198 171154 185434
rect 170918 178198 171154 178434
rect 170918 171198 171154 171434
rect 170918 164198 171154 164434
rect 170918 157198 171154 157434
rect 170918 150198 171154 150434
rect 170918 143198 171154 143434
rect 170918 136198 171154 136434
rect 170918 129198 171154 129434
rect 170918 122198 171154 122434
rect 170918 115198 171154 115434
rect 170918 108198 171154 108434
rect 170918 101198 171154 101434
rect 170918 94198 171154 94434
rect 170918 87198 171154 87434
rect 170918 80198 171154 80434
rect 170918 73198 171154 73434
rect 170918 66198 171154 66434
rect 170918 59198 171154 59434
rect 170918 52198 171154 52434
rect 170918 45198 171154 45434
rect 170918 38198 171154 38434
rect 170918 31198 171154 31434
rect 170918 24198 171154 24434
rect 170918 17198 171154 17434
rect 170918 10198 171154 10434
rect 170918 3198 171154 3434
rect 170918 -1942 171154 -1706
rect 170918 -2262 171154 -2026
rect 176186 705002 176422 705238
rect 176186 704682 176422 704918
rect 176186 695258 176422 695494
rect 176186 688258 176422 688494
rect 176186 681258 176422 681494
rect 176186 674258 176422 674494
rect 176186 667258 176422 667494
rect 176186 660258 176422 660494
rect 176186 653258 176422 653494
rect 176186 646258 176422 646494
rect 176186 639258 176422 639494
rect 176186 632258 176422 632494
rect 176186 625258 176422 625494
rect 176186 618258 176422 618494
rect 176186 611258 176422 611494
rect 176186 604258 176422 604494
rect 176186 597258 176422 597494
rect 176186 590258 176422 590494
rect 176186 583258 176422 583494
rect 176186 576258 176422 576494
rect 176186 569258 176422 569494
rect 176186 562258 176422 562494
rect 176186 555258 176422 555494
rect 176186 548258 176422 548494
rect 176186 541258 176422 541494
rect 176186 534258 176422 534494
rect 176186 527258 176422 527494
rect 176186 520258 176422 520494
rect 176186 513258 176422 513494
rect 176186 506258 176422 506494
rect 176186 499258 176422 499494
rect 176186 492258 176422 492494
rect 176186 485258 176422 485494
rect 176186 478258 176422 478494
rect 176186 471258 176422 471494
rect 176186 464258 176422 464494
rect 176186 457258 176422 457494
rect 176186 450258 176422 450494
rect 176186 443258 176422 443494
rect 176186 436258 176422 436494
rect 176186 429258 176422 429494
rect 176186 422258 176422 422494
rect 176186 415258 176422 415494
rect 176186 408258 176422 408494
rect 176186 401258 176422 401494
rect 176186 394258 176422 394494
rect 176186 387258 176422 387494
rect 176186 380258 176422 380494
rect 176186 373258 176422 373494
rect 176186 366258 176422 366494
rect 176186 359258 176422 359494
rect 176186 352258 176422 352494
rect 176186 345258 176422 345494
rect 176186 338258 176422 338494
rect 176186 331258 176422 331494
rect 176186 324258 176422 324494
rect 176186 317258 176422 317494
rect 176186 310258 176422 310494
rect 176186 303258 176422 303494
rect 176186 296258 176422 296494
rect 176186 289258 176422 289494
rect 176186 282258 176422 282494
rect 176186 275258 176422 275494
rect 176186 268258 176422 268494
rect 176186 261258 176422 261494
rect 176186 254258 176422 254494
rect 176186 247258 176422 247494
rect 176186 240258 176422 240494
rect 176186 233258 176422 233494
rect 176186 226258 176422 226494
rect 176186 219258 176422 219494
rect 176186 212258 176422 212494
rect 176186 205258 176422 205494
rect 176186 198258 176422 198494
rect 176186 191258 176422 191494
rect 176186 184258 176422 184494
rect 176186 177258 176422 177494
rect 176186 170258 176422 170494
rect 176186 163258 176422 163494
rect 176186 156258 176422 156494
rect 176186 149258 176422 149494
rect 176186 142258 176422 142494
rect 176186 135258 176422 135494
rect 176186 128258 176422 128494
rect 176186 121258 176422 121494
rect 176186 114258 176422 114494
rect 176186 107258 176422 107494
rect 176186 100258 176422 100494
rect 176186 93258 176422 93494
rect 176186 86258 176422 86494
rect 176186 79258 176422 79494
rect 176186 72258 176422 72494
rect 176186 65258 176422 65494
rect 176186 58258 176422 58494
rect 176186 51258 176422 51494
rect 176186 44258 176422 44494
rect 176186 37258 176422 37494
rect 176186 30258 176422 30494
rect 176186 23258 176422 23494
rect 176186 16258 176422 16494
rect 176186 9258 176422 9494
rect 176186 2258 176422 2494
rect 176186 -982 176422 -746
rect 176186 -1302 176422 -1066
rect 177918 705962 178154 706198
rect 177918 705642 178154 705878
rect 177918 696198 178154 696434
rect 177918 689198 178154 689434
rect 177918 682198 178154 682434
rect 177918 675198 178154 675434
rect 177918 668198 178154 668434
rect 177918 661198 178154 661434
rect 177918 654198 178154 654434
rect 177918 647198 178154 647434
rect 177918 640198 178154 640434
rect 177918 633198 178154 633434
rect 177918 626198 178154 626434
rect 177918 619198 178154 619434
rect 177918 612198 178154 612434
rect 177918 605198 178154 605434
rect 177918 598198 178154 598434
rect 177918 591198 178154 591434
rect 177918 584198 178154 584434
rect 177918 577198 178154 577434
rect 177918 570198 178154 570434
rect 177918 563198 178154 563434
rect 177918 556198 178154 556434
rect 177918 549198 178154 549434
rect 177918 542198 178154 542434
rect 177918 535198 178154 535434
rect 177918 528198 178154 528434
rect 177918 521198 178154 521434
rect 177918 514198 178154 514434
rect 177918 507198 178154 507434
rect 177918 500198 178154 500434
rect 177918 493198 178154 493434
rect 177918 486198 178154 486434
rect 177918 479198 178154 479434
rect 177918 472198 178154 472434
rect 177918 465198 178154 465434
rect 177918 458198 178154 458434
rect 177918 451198 178154 451434
rect 177918 444198 178154 444434
rect 177918 437198 178154 437434
rect 177918 430198 178154 430434
rect 177918 423198 178154 423434
rect 177918 416198 178154 416434
rect 177918 409198 178154 409434
rect 177918 402198 178154 402434
rect 177918 395198 178154 395434
rect 177918 388198 178154 388434
rect 177918 381198 178154 381434
rect 177918 374198 178154 374434
rect 177918 367198 178154 367434
rect 177918 360198 178154 360434
rect 177918 353198 178154 353434
rect 177918 346198 178154 346434
rect 177918 339198 178154 339434
rect 177918 332198 178154 332434
rect 177918 325198 178154 325434
rect 177918 318198 178154 318434
rect 177918 311198 178154 311434
rect 177918 304198 178154 304434
rect 177918 297198 178154 297434
rect 177918 290198 178154 290434
rect 177918 283198 178154 283434
rect 177918 276198 178154 276434
rect 177918 269198 178154 269434
rect 177918 262198 178154 262434
rect 177918 255198 178154 255434
rect 177918 248198 178154 248434
rect 177918 241198 178154 241434
rect 177918 234198 178154 234434
rect 177918 227198 178154 227434
rect 177918 220198 178154 220434
rect 177918 213198 178154 213434
rect 177918 206198 178154 206434
rect 177918 199198 178154 199434
rect 177918 192198 178154 192434
rect 177918 185198 178154 185434
rect 177918 178198 178154 178434
rect 177918 171198 178154 171434
rect 177918 164198 178154 164434
rect 177918 157198 178154 157434
rect 177918 150198 178154 150434
rect 177918 143198 178154 143434
rect 177918 136198 178154 136434
rect 177918 129198 178154 129434
rect 177918 122198 178154 122434
rect 177918 115198 178154 115434
rect 177918 108198 178154 108434
rect 177918 101198 178154 101434
rect 177918 94198 178154 94434
rect 177918 87198 178154 87434
rect 177918 80198 178154 80434
rect 177918 73198 178154 73434
rect 177918 66198 178154 66434
rect 177918 59198 178154 59434
rect 177918 52198 178154 52434
rect 177918 45198 178154 45434
rect 177918 38198 178154 38434
rect 177918 31198 178154 31434
rect 177918 24198 178154 24434
rect 177918 17198 178154 17434
rect 177918 10198 178154 10434
rect 177918 3198 178154 3434
rect 177918 -1942 178154 -1706
rect 177918 -2262 178154 -2026
rect 183186 705002 183422 705238
rect 183186 704682 183422 704918
rect 183186 695258 183422 695494
rect 183186 688258 183422 688494
rect 183186 681258 183422 681494
rect 183186 674258 183422 674494
rect 183186 667258 183422 667494
rect 183186 660258 183422 660494
rect 183186 653258 183422 653494
rect 183186 646258 183422 646494
rect 183186 639258 183422 639494
rect 183186 632258 183422 632494
rect 183186 625258 183422 625494
rect 183186 618258 183422 618494
rect 183186 611258 183422 611494
rect 183186 604258 183422 604494
rect 183186 597258 183422 597494
rect 183186 590258 183422 590494
rect 183186 583258 183422 583494
rect 183186 576258 183422 576494
rect 183186 569258 183422 569494
rect 183186 562258 183422 562494
rect 183186 555258 183422 555494
rect 183186 548258 183422 548494
rect 183186 541258 183422 541494
rect 183186 534258 183422 534494
rect 183186 527258 183422 527494
rect 183186 520258 183422 520494
rect 183186 513258 183422 513494
rect 183186 506258 183422 506494
rect 183186 499258 183422 499494
rect 183186 492258 183422 492494
rect 183186 485258 183422 485494
rect 183186 478258 183422 478494
rect 183186 471258 183422 471494
rect 183186 464258 183422 464494
rect 183186 457258 183422 457494
rect 183186 450258 183422 450494
rect 183186 443258 183422 443494
rect 183186 436258 183422 436494
rect 183186 429258 183422 429494
rect 183186 422258 183422 422494
rect 183186 415258 183422 415494
rect 183186 408258 183422 408494
rect 183186 401258 183422 401494
rect 183186 394258 183422 394494
rect 183186 387258 183422 387494
rect 183186 380258 183422 380494
rect 183186 373258 183422 373494
rect 183186 366258 183422 366494
rect 183186 359258 183422 359494
rect 183186 352258 183422 352494
rect 183186 345258 183422 345494
rect 183186 338258 183422 338494
rect 183186 331258 183422 331494
rect 183186 324258 183422 324494
rect 183186 317258 183422 317494
rect 183186 310258 183422 310494
rect 183186 303258 183422 303494
rect 183186 296258 183422 296494
rect 183186 289258 183422 289494
rect 183186 282258 183422 282494
rect 183186 275258 183422 275494
rect 183186 268258 183422 268494
rect 183186 261258 183422 261494
rect 183186 254258 183422 254494
rect 183186 247258 183422 247494
rect 183186 240258 183422 240494
rect 183186 233258 183422 233494
rect 183186 226258 183422 226494
rect 183186 219258 183422 219494
rect 183186 212258 183422 212494
rect 183186 205258 183422 205494
rect 183186 198258 183422 198494
rect 183186 191258 183422 191494
rect 183186 184258 183422 184494
rect 183186 177258 183422 177494
rect 183186 170258 183422 170494
rect 183186 163258 183422 163494
rect 183186 156258 183422 156494
rect 183186 149258 183422 149494
rect 183186 142258 183422 142494
rect 183186 135258 183422 135494
rect 183186 128258 183422 128494
rect 183186 121258 183422 121494
rect 183186 114258 183422 114494
rect 183186 107258 183422 107494
rect 183186 100258 183422 100494
rect 183186 93258 183422 93494
rect 183186 86258 183422 86494
rect 183186 79258 183422 79494
rect 183186 72258 183422 72494
rect 183186 65258 183422 65494
rect 183186 58258 183422 58494
rect 183186 51258 183422 51494
rect 183186 44258 183422 44494
rect 183186 37258 183422 37494
rect 183186 30258 183422 30494
rect 183186 23258 183422 23494
rect 183186 16258 183422 16494
rect 183186 9258 183422 9494
rect 183186 2258 183422 2494
rect 183186 -982 183422 -746
rect 183186 -1302 183422 -1066
rect 184918 705962 185154 706198
rect 184918 705642 185154 705878
rect 184918 696198 185154 696434
rect 184918 689198 185154 689434
rect 184918 682198 185154 682434
rect 184918 675198 185154 675434
rect 184918 668198 185154 668434
rect 184918 661198 185154 661434
rect 184918 654198 185154 654434
rect 184918 647198 185154 647434
rect 184918 640198 185154 640434
rect 184918 633198 185154 633434
rect 184918 626198 185154 626434
rect 184918 619198 185154 619434
rect 184918 612198 185154 612434
rect 184918 605198 185154 605434
rect 184918 598198 185154 598434
rect 184918 591198 185154 591434
rect 184918 584198 185154 584434
rect 184918 577198 185154 577434
rect 184918 570198 185154 570434
rect 184918 563198 185154 563434
rect 184918 556198 185154 556434
rect 184918 549198 185154 549434
rect 184918 542198 185154 542434
rect 184918 535198 185154 535434
rect 184918 528198 185154 528434
rect 184918 521198 185154 521434
rect 184918 514198 185154 514434
rect 184918 507198 185154 507434
rect 184918 500198 185154 500434
rect 184918 493198 185154 493434
rect 184918 486198 185154 486434
rect 184918 479198 185154 479434
rect 184918 472198 185154 472434
rect 184918 465198 185154 465434
rect 184918 458198 185154 458434
rect 184918 451198 185154 451434
rect 184918 444198 185154 444434
rect 184918 437198 185154 437434
rect 184918 430198 185154 430434
rect 184918 423198 185154 423434
rect 184918 416198 185154 416434
rect 184918 409198 185154 409434
rect 184918 402198 185154 402434
rect 184918 395198 185154 395434
rect 184918 388198 185154 388434
rect 184918 381198 185154 381434
rect 184918 374198 185154 374434
rect 184918 367198 185154 367434
rect 184918 360198 185154 360434
rect 184918 353198 185154 353434
rect 184918 346198 185154 346434
rect 184918 339198 185154 339434
rect 184918 332198 185154 332434
rect 184918 325198 185154 325434
rect 184918 318198 185154 318434
rect 184918 311198 185154 311434
rect 184918 304198 185154 304434
rect 184918 297198 185154 297434
rect 184918 290198 185154 290434
rect 184918 283198 185154 283434
rect 184918 276198 185154 276434
rect 184918 269198 185154 269434
rect 184918 262198 185154 262434
rect 184918 255198 185154 255434
rect 184918 248198 185154 248434
rect 184918 241198 185154 241434
rect 184918 234198 185154 234434
rect 184918 227198 185154 227434
rect 184918 220198 185154 220434
rect 184918 213198 185154 213434
rect 184918 206198 185154 206434
rect 184918 199198 185154 199434
rect 184918 192198 185154 192434
rect 184918 185198 185154 185434
rect 184918 178198 185154 178434
rect 184918 171198 185154 171434
rect 184918 164198 185154 164434
rect 184918 157198 185154 157434
rect 184918 150198 185154 150434
rect 184918 143198 185154 143434
rect 184918 136198 185154 136434
rect 184918 129198 185154 129434
rect 184918 122198 185154 122434
rect 184918 115198 185154 115434
rect 184918 108198 185154 108434
rect 184918 101198 185154 101434
rect 184918 94198 185154 94434
rect 184918 87198 185154 87434
rect 184918 80198 185154 80434
rect 184918 73198 185154 73434
rect 184918 66198 185154 66434
rect 184918 59198 185154 59434
rect 184918 52198 185154 52434
rect 184918 45198 185154 45434
rect 184918 38198 185154 38434
rect 184918 31198 185154 31434
rect 184918 24198 185154 24434
rect 184918 17198 185154 17434
rect 184918 10198 185154 10434
rect 184918 3198 185154 3434
rect 184918 -1942 185154 -1706
rect 184918 -2262 185154 -2026
rect 190186 705002 190422 705238
rect 190186 704682 190422 704918
rect 190186 695258 190422 695494
rect 190186 688258 190422 688494
rect 190186 681258 190422 681494
rect 190186 674258 190422 674494
rect 190186 667258 190422 667494
rect 190186 660258 190422 660494
rect 190186 653258 190422 653494
rect 190186 646258 190422 646494
rect 190186 639258 190422 639494
rect 190186 632258 190422 632494
rect 190186 625258 190422 625494
rect 190186 618258 190422 618494
rect 190186 611258 190422 611494
rect 190186 604258 190422 604494
rect 190186 597258 190422 597494
rect 190186 590258 190422 590494
rect 190186 583258 190422 583494
rect 190186 576258 190422 576494
rect 190186 569258 190422 569494
rect 190186 562258 190422 562494
rect 190186 555258 190422 555494
rect 190186 548258 190422 548494
rect 190186 541258 190422 541494
rect 190186 534258 190422 534494
rect 190186 527258 190422 527494
rect 190186 520258 190422 520494
rect 190186 513258 190422 513494
rect 190186 506258 190422 506494
rect 190186 499258 190422 499494
rect 190186 492258 190422 492494
rect 190186 485258 190422 485494
rect 190186 478258 190422 478494
rect 190186 471258 190422 471494
rect 190186 464258 190422 464494
rect 190186 457258 190422 457494
rect 190186 450258 190422 450494
rect 190186 443258 190422 443494
rect 190186 436258 190422 436494
rect 190186 429258 190422 429494
rect 190186 422258 190422 422494
rect 190186 415258 190422 415494
rect 190186 408258 190422 408494
rect 190186 401258 190422 401494
rect 190186 394258 190422 394494
rect 190186 387258 190422 387494
rect 190186 380258 190422 380494
rect 190186 373258 190422 373494
rect 190186 366258 190422 366494
rect 190186 359258 190422 359494
rect 190186 352258 190422 352494
rect 190186 345258 190422 345494
rect 190186 338258 190422 338494
rect 190186 331258 190422 331494
rect 190186 324258 190422 324494
rect 190186 317258 190422 317494
rect 190186 310258 190422 310494
rect 190186 303258 190422 303494
rect 190186 296258 190422 296494
rect 190186 289258 190422 289494
rect 190186 282258 190422 282494
rect 190186 275258 190422 275494
rect 190186 268258 190422 268494
rect 190186 261258 190422 261494
rect 190186 254258 190422 254494
rect 190186 247258 190422 247494
rect 190186 240258 190422 240494
rect 190186 233258 190422 233494
rect 190186 226258 190422 226494
rect 190186 219258 190422 219494
rect 190186 212258 190422 212494
rect 190186 205258 190422 205494
rect 190186 198258 190422 198494
rect 190186 191258 190422 191494
rect 190186 184258 190422 184494
rect 190186 177258 190422 177494
rect 190186 170258 190422 170494
rect 190186 163258 190422 163494
rect 190186 156258 190422 156494
rect 190186 149258 190422 149494
rect 190186 142258 190422 142494
rect 190186 135258 190422 135494
rect 190186 128258 190422 128494
rect 190186 121258 190422 121494
rect 190186 114258 190422 114494
rect 190186 107258 190422 107494
rect 190186 100258 190422 100494
rect 190186 93258 190422 93494
rect 190186 86258 190422 86494
rect 190186 79258 190422 79494
rect 190186 72258 190422 72494
rect 190186 65258 190422 65494
rect 190186 58258 190422 58494
rect 190186 51258 190422 51494
rect 190186 44258 190422 44494
rect 190186 37258 190422 37494
rect 190186 30258 190422 30494
rect 190186 23258 190422 23494
rect 190186 16258 190422 16494
rect 190186 9258 190422 9494
rect 190186 2258 190422 2494
rect 190186 -982 190422 -746
rect 190186 -1302 190422 -1066
rect 191918 705962 192154 706198
rect 191918 705642 192154 705878
rect 191918 696198 192154 696434
rect 191918 689198 192154 689434
rect 191918 682198 192154 682434
rect 191918 675198 192154 675434
rect 191918 668198 192154 668434
rect 191918 661198 192154 661434
rect 191918 654198 192154 654434
rect 191918 647198 192154 647434
rect 191918 640198 192154 640434
rect 191918 633198 192154 633434
rect 191918 626198 192154 626434
rect 191918 619198 192154 619434
rect 191918 612198 192154 612434
rect 191918 605198 192154 605434
rect 191918 598198 192154 598434
rect 191918 591198 192154 591434
rect 191918 584198 192154 584434
rect 191918 577198 192154 577434
rect 191918 570198 192154 570434
rect 191918 563198 192154 563434
rect 191918 556198 192154 556434
rect 191918 549198 192154 549434
rect 191918 542198 192154 542434
rect 191918 535198 192154 535434
rect 191918 528198 192154 528434
rect 191918 521198 192154 521434
rect 191918 514198 192154 514434
rect 191918 507198 192154 507434
rect 191918 500198 192154 500434
rect 191918 493198 192154 493434
rect 191918 486198 192154 486434
rect 191918 479198 192154 479434
rect 191918 472198 192154 472434
rect 191918 465198 192154 465434
rect 191918 458198 192154 458434
rect 191918 451198 192154 451434
rect 191918 444198 192154 444434
rect 191918 437198 192154 437434
rect 191918 430198 192154 430434
rect 191918 423198 192154 423434
rect 191918 416198 192154 416434
rect 191918 409198 192154 409434
rect 191918 402198 192154 402434
rect 191918 395198 192154 395434
rect 191918 388198 192154 388434
rect 191918 381198 192154 381434
rect 191918 374198 192154 374434
rect 191918 367198 192154 367434
rect 191918 360198 192154 360434
rect 191918 353198 192154 353434
rect 191918 346198 192154 346434
rect 191918 339198 192154 339434
rect 191918 332198 192154 332434
rect 191918 325198 192154 325434
rect 191918 318198 192154 318434
rect 191918 311198 192154 311434
rect 191918 304198 192154 304434
rect 191918 297198 192154 297434
rect 191918 290198 192154 290434
rect 191918 283198 192154 283434
rect 191918 276198 192154 276434
rect 191918 269198 192154 269434
rect 191918 262198 192154 262434
rect 191918 255198 192154 255434
rect 191918 248198 192154 248434
rect 191918 241198 192154 241434
rect 191918 234198 192154 234434
rect 191918 227198 192154 227434
rect 191918 220198 192154 220434
rect 191918 213198 192154 213434
rect 191918 206198 192154 206434
rect 191918 199198 192154 199434
rect 191918 192198 192154 192434
rect 191918 185198 192154 185434
rect 191918 178198 192154 178434
rect 191918 171198 192154 171434
rect 191918 164198 192154 164434
rect 191918 157198 192154 157434
rect 191918 150198 192154 150434
rect 191918 143198 192154 143434
rect 191918 136198 192154 136434
rect 191918 129198 192154 129434
rect 191918 122198 192154 122434
rect 191918 115198 192154 115434
rect 191918 108198 192154 108434
rect 191918 101198 192154 101434
rect 191918 94198 192154 94434
rect 191918 87198 192154 87434
rect 191918 80198 192154 80434
rect 191918 73198 192154 73434
rect 191918 66198 192154 66434
rect 191918 59198 192154 59434
rect 191918 52198 192154 52434
rect 191918 45198 192154 45434
rect 191918 38198 192154 38434
rect 191918 31198 192154 31434
rect 191918 24198 192154 24434
rect 191918 17198 192154 17434
rect 191918 10198 192154 10434
rect 191918 3198 192154 3434
rect 191918 -1942 192154 -1706
rect 191918 -2262 192154 -2026
rect 197186 705002 197422 705238
rect 197186 704682 197422 704918
rect 197186 695258 197422 695494
rect 197186 688258 197422 688494
rect 197186 681258 197422 681494
rect 197186 674258 197422 674494
rect 197186 667258 197422 667494
rect 197186 660258 197422 660494
rect 197186 653258 197422 653494
rect 197186 646258 197422 646494
rect 197186 639258 197422 639494
rect 197186 632258 197422 632494
rect 197186 625258 197422 625494
rect 197186 618258 197422 618494
rect 197186 611258 197422 611494
rect 197186 604258 197422 604494
rect 197186 597258 197422 597494
rect 197186 590258 197422 590494
rect 197186 583258 197422 583494
rect 197186 576258 197422 576494
rect 197186 569258 197422 569494
rect 197186 562258 197422 562494
rect 197186 555258 197422 555494
rect 197186 548258 197422 548494
rect 197186 541258 197422 541494
rect 197186 534258 197422 534494
rect 197186 527258 197422 527494
rect 197186 520258 197422 520494
rect 197186 513258 197422 513494
rect 197186 506258 197422 506494
rect 197186 499258 197422 499494
rect 197186 492258 197422 492494
rect 197186 485258 197422 485494
rect 197186 478258 197422 478494
rect 197186 471258 197422 471494
rect 197186 464258 197422 464494
rect 197186 457258 197422 457494
rect 197186 450258 197422 450494
rect 197186 443258 197422 443494
rect 197186 436258 197422 436494
rect 197186 429258 197422 429494
rect 197186 422258 197422 422494
rect 197186 415258 197422 415494
rect 197186 408258 197422 408494
rect 197186 401258 197422 401494
rect 197186 394258 197422 394494
rect 197186 387258 197422 387494
rect 197186 380258 197422 380494
rect 197186 373258 197422 373494
rect 197186 366258 197422 366494
rect 197186 359258 197422 359494
rect 197186 352258 197422 352494
rect 197186 345258 197422 345494
rect 197186 338258 197422 338494
rect 197186 331258 197422 331494
rect 197186 324258 197422 324494
rect 197186 317258 197422 317494
rect 197186 310258 197422 310494
rect 197186 303258 197422 303494
rect 197186 296258 197422 296494
rect 197186 289258 197422 289494
rect 197186 282258 197422 282494
rect 197186 275258 197422 275494
rect 197186 268258 197422 268494
rect 197186 261258 197422 261494
rect 197186 254258 197422 254494
rect 197186 247258 197422 247494
rect 197186 240258 197422 240494
rect 197186 233258 197422 233494
rect 197186 226258 197422 226494
rect 197186 219258 197422 219494
rect 197186 212258 197422 212494
rect 197186 205258 197422 205494
rect 197186 198258 197422 198494
rect 197186 191258 197422 191494
rect 197186 184258 197422 184494
rect 197186 177258 197422 177494
rect 197186 170258 197422 170494
rect 197186 163258 197422 163494
rect 197186 156258 197422 156494
rect 197186 149258 197422 149494
rect 197186 142258 197422 142494
rect 197186 135258 197422 135494
rect 197186 128258 197422 128494
rect 197186 121258 197422 121494
rect 197186 114258 197422 114494
rect 197186 107258 197422 107494
rect 197186 100258 197422 100494
rect 197186 93258 197422 93494
rect 197186 86258 197422 86494
rect 197186 79258 197422 79494
rect 197186 72258 197422 72494
rect 197186 65258 197422 65494
rect 197186 58258 197422 58494
rect 197186 51258 197422 51494
rect 197186 44258 197422 44494
rect 197186 37258 197422 37494
rect 197186 30258 197422 30494
rect 197186 23258 197422 23494
rect 197186 16258 197422 16494
rect 197186 9258 197422 9494
rect 197186 2258 197422 2494
rect 197186 -982 197422 -746
rect 197186 -1302 197422 -1066
rect 198918 705962 199154 706198
rect 198918 705642 199154 705878
rect 198918 696198 199154 696434
rect 198918 689198 199154 689434
rect 198918 682198 199154 682434
rect 198918 675198 199154 675434
rect 198918 668198 199154 668434
rect 198918 661198 199154 661434
rect 198918 654198 199154 654434
rect 198918 647198 199154 647434
rect 198918 640198 199154 640434
rect 198918 633198 199154 633434
rect 198918 626198 199154 626434
rect 198918 619198 199154 619434
rect 198918 612198 199154 612434
rect 198918 605198 199154 605434
rect 198918 598198 199154 598434
rect 198918 591198 199154 591434
rect 198918 584198 199154 584434
rect 198918 577198 199154 577434
rect 198918 570198 199154 570434
rect 198918 563198 199154 563434
rect 198918 556198 199154 556434
rect 198918 549198 199154 549434
rect 198918 542198 199154 542434
rect 198918 535198 199154 535434
rect 198918 528198 199154 528434
rect 198918 521198 199154 521434
rect 198918 514198 199154 514434
rect 198918 507198 199154 507434
rect 198918 500198 199154 500434
rect 198918 493198 199154 493434
rect 198918 486198 199154 486434
rect 198918 479198 199154 479434
rect 198918 472198 199154 472434
rect 198918 465198 199154 465434
rect 198918 458198 199154 458434
rect 198918 451198 199154 451434
rect 198918 444198 199154 444434
rect 198918 437198 199154 437434
rect 198918 430198 199154 430434
rect 198918 423198 199154 423434
rect 198918 416198 199154 416434
rect 198918 409198 199154 409434
rect 198918 402198 199154 402434
rect 198918 395198 199154 395434
rect 198918 388198 199154 388434
rect 198918 381198 199154 381434
rect 198918 374198 199154 374434
rect 198918 367198 199154 367434
rect 198918 360198 199154 360434
rect 198918 353198 199154 353434
rect 198918 346198 199154 346434
rect 198918 339198 199154 339434
rect 198918 332198 199154 332434
rect 198918 325198 199154 325434
rect 198918 318198 199154 318434
rect 198918 311198 199154 311434
rect 198918 304198 199154 304434
rect 198918 297198 199154 297434
rect 198918 290198 199154 290434
rect 198918 283198 199154 283434
rect 198918 276198 199154 276434
rect 198918 269198 199154 269434
rect 198918 262198 199154 262434
rect 198918 255198 199154 255434
rect 198918 248198 199154 248434
rect 198918 241198 199154 241434
rect 198918 234198 199154 234434
rect 198918 227198 199154 227434
rect 198918 220198 199154 220434
rect 198918 213198 199154 213434
rect 198918 206198 199154 206434
rect 198918 199198 199154 199434
rect 198918 192198 199154 192434
rect 198918 185198 199154 185434
rect 198918 178198 199154 178434
rect 198918 171198 199154 171434
rect 198918 164198 199154 164434
rect 198918 157198 199154 157434
rect 198918 150198 199154 150434
rect 198918 143198 199154 143434
rect 198918 136198 199154 136434
rect 198918 129198 199154 129434
rect 198918 122198 199154 122434
rect 198918 115198 199154 115434
rect 198918 108198 199154 108434
rect 198918 101198 199154 101434
rect 198918 94198 199154 94434
rect 198918 87198 199154 87434
rect 198918 80198 199154 80434
rect 198918 73198 199154 73434
rect 198918 66198 199154 66434
rect 198918 59198 199154 59434
rect 198918 52198 199154 52434
rect 198918 45198 199154 45434
rect 198918 38198 199154 38434
rect 198918 31198 199154 31434
rect 198918 24198 199154 24434
rect 198918 17198 199154 17434
rect 198918 10198 199154 10434
rect 198918 3198 199154 3434
rect 198918 -1942 199154 -1706
rect 198918 -2262 199154 -2026
rect 204186 705002 204422 705238
rect 204186 704682 204422 704918
rect 204186 695258 204422 695494
rect 204186 688258 204422 688494
rect 204186 681258 204422 681494
rect 204186 674258 204422 674494
rect 204186 667258 204422 667494
rect 204186 660258 204422 660494
rect 204186 653258 204422 653494
rect 204186 646258 204422 646494
rect 204186 639258 204422 639494
rect 204186 632258 204422 632494
rect 204186 625258 204422 625494
rect 204186 618258 204422 618494
rect 204186 611258 204422 611494
rect 204186 604258 204422 604494
rect 204186 597258 204422 597494
rect 204186 590258 204422 590494
rect 204186 583258 204422 583494
rect 204186 576258 204422 576494
rect 204186 569258 204422 569494
rect 204186 562258 204422 562494
rect 204186 555258 204422 555494
rect 204186 548258 204422 548494
rect 204186 541258 204422 541494
rect 204186 534258 204422 534494
rect 204186 527258 204422 527494
rect 204186 520258 204422 520494
rect 204186 513258 204422 513494
rect 204186 506258 204422 506494
rect 204186 499258 204422 499494
rect 204186 492258 204422 492494
rect 204186 485258 204422 485494
rect 204186 478258 204422 478494
rect 204186 471258 204422 471494
rect 204186 464258 204422 464494
rect 204186 457258 204422 457494
rect 204186 450258 204422 450494
rect 204186 443258 204422 443494
rect 204186 436258 204422 436494
rect 204186 429258 204422 429494
rect 204186 422258 204422 422494
rect 204186 415258 204422 415494
rect 204186 408258 204422 408494
rect 204186 401258 204422 401494
rect 204186 394258 204422 394494
rect 204186 387258 204422 387494
rect 204186 380258 204422 380494
rect 204186 373258 204422 373494
rect 204186 366258 204422 366494
rect 204186 359258 204422 359494
rect 204186 352258 204422 352494
rect 204186 345258 204422 345494
rect 204186 338258 204422 338494
rect 204186 331258 204422 331494
rect 204186 324258 204422 324494
rect 204186 317258 204422 317494
rect 204186 310258 204422 310494
rect 204186 303258 204422 303494
rect 204186 296258 204422 296494
rect 204186 289258 204422 289494
rect 204186 282258 204422 282494
rect 204186 275258 204422 275494
rect 204186 268258 204422 268494
rect 204186 261258 204422 261494
rect 204186 254258 204422 254494
rect 204186 247258 204422 247494
rect 204186 240258 204422 240494
rect 204186 233258 204422 233494
rect 204186 226258 204422 226494
rect 204186 219258 204422 219494
rect 204186 212258 204422 212494
rect 204186 205258 204422 205494
rect 204186 198258 204422 198494
rect 204186 191258 204422 191494
rect 204186 184258 204422 184494
rect 204186 177258 204422 177494
rect 204186 170258 204422 170494
rect 204186 163258 204422 163494
rect 204186 156258 204422 156494
rect 204186 149258 204422 149494
rect 204186 142258 204422 142494
rect 204186 135258 204422 135494
rect 204186 128258 204422 128494
rect 204186 121258 204422 121494
rect 204186 114258 204422 114494
rect 204186 107258 204422 107494
rect 204186 100258 204422 100494
rect 204186 93258 204422 93494
rect 204186 86258 204422 86494
rect 204186 79258 204422 79494
rect 204186 72258 204422 72494
rect 204186 65258 204422 65494
rect 204186 58258 204422 58494
rect 204186 51258 204422 51494
rect 204186 44258 204422 44494
rect 204186 37258 204422 37494
rect 204186 30258 204422 30494
rect 204186 23258 204422 23494
rect 204186 16258 204422 16494
rect 204186 9258 204422 9494
rect 204186 2258 204422 2494
rect 204186 -982 204422 -746
rect 204186 -1302 204422 -1066
rect 205918 705962 206154 706198
rect 205918 705642 206154 705878
rect 205918 696198 206154 696434
rect 205918 689198 206154 689434
rect 205918 682198 206154 682434
rect 205918 675198 206154 675434
rect 205918 668198 206154 668434
rect 205918 661198 206154 661434
rect 205918 654198 206154 654434
rect 205918 647198 206154 647434
rect 205918 640198 206154 640434
rect 205918 633198 206154 633434
rect 205918 626198 206154 626434
rect 205918 619198 206154 619434
rect 205918 612198 206154 612434
rect 205918 605198 206154 605434
rect 205918 598198 206154 598434
rect 205918 591198 206154 591434
rect 205918 584198 206154 584434
rect 205918 577198 206154 577434
rect 205918 570198 206154 570434
rect 205918 563198 206154 563434
rect 205918 556198 206154 556434
rect 205918 549198 206154 549434
rect 205918 542198 206154 542434
rect 205918 535198 206154 535434
rect 205918 528198 206154 528434
rect 205918 521198 206154 521434
rect 205918 514198 206154 514434
rect 205918 507198 206154 507434
rect 205918 500198 206154 500434
rect 205918 493198 206154 493434
rect 205918 486198 206154 486434
rect 205918 479198 206154 479434
rect 205918 472198 206154 472434
rect 205918 465198 206154 465434
rect 205918 458198 206154 458434
rect 205918 451198 206154 451434
rect 205918 444198 206154 444434
rect 205918 437198 206154 437434
rect 205918 430198 206154 430434
rect 205918 423198 206154 423434
rect 205918 416198 206154 416434
rect 205918 409198 206154 409434
rect 205918 402198 206154 402434
rect 205918 395198 206154 395434
rect 205918 388198 206154 388434
rect 205918 381198 206154 381434
rect 205918 374198 206154 374434
rect 205918 367198 206154 367434
rect 205918 360198 206154 360434
rect 205918 353198 206154 353434
rect 205918 346198 206154 346434
rect 205918 339198 206154 339434
rect 205918 332198 206154 332434
rect 205918 325198 206154 325434
rect 205918 318198 206154 318434
rect 205918 311198 206154 311434
rect 205918 304198 206154 304434
rect 205918 297198 206154 297434
rect 205918 290198 206154 290434
rect 205918 283198 206154 283434
rect 205918 276198 206154 276434
rect 205918 269198 206154 269434
rect 205918 262198 206154 262434
rect 205918 255198 206154 255434
rect 205918 248198 206154 248434
rect 205918 241198 206154 241434
rect 205918 234198 206154 234434
rect 205918 227198 206154 227434
rect 205918 220198 206154 220434
rect 205918 213198 206154 213434
rect 205918 206198 206154 206434
rect 205918 199198 206154 199434
rect 205918 192198 206154 192434
rect 205918 185198 206154 185434
rect 205918 178198 206154 178434
rect 205918 171198 206154 171434
rect 205918 164198 206154 164434
rect 205918 157198 206154 157434
rect 205918 150198 206154 150434
rect 205918 143198 206154 143434
rect 205918 136198 206154 136434
rect 205918 129198 206154 129434
rect 205918 122198 206154 122434
rect 205918 115198 206154 115434
rect 205918 108198 206154 108434
rect 205918 101198 206154 101434
rect 205918 94198 206154 94434
rect 205918 87198 206154 87434
rect 205918 80198 206154 80434
rect 205918 73198 206154 73434
rect 205918 66198 206154 66434
rect 205918 59198 206154 59434
rect 205918 52198 206154 52434
rect 205918 45198 206154 45434
rect 205918 38198 206154 38434
rect 205918 31198 206154 31434
rect 205918 24198 206154 24434
rect 205918 17198 206154 17434
rect 205918 10198 206154 10434
rect 205918 3198 206154 3434
rect 205918 -1942 206154 -1706
rect 205918 -2262 206154 -2026
rect 211186 705002 211422 705238
rect 211186 704682 211422 704918
rect 211186 695258 211422 695494
rect 211186 688258 211422 688494
rect 211186 681258 211422 681494
rect 211186 674258 211422 674494
rect 211186 667258 211422 667494
rect 211186 660258 211422 660494
rect 211186 653258 211422 653494
rect 211186 646258 211422 646494
rect 211186 639258 211422 639494
rect 211186 632258 211422 632494
rect 211186 625258 211422 625494
rect 211186 618258 211422 618494
rect 211186 611258 211422 611494
rect 211186 604258 211422 604494
rect 211186 597258 211422 597494
rect 211186 590258 211422 590494
rect 211186 583258 211422 583494
rect 211186 576258 211422 576494
rect 211186 569258 211422 569494
rect 211186 562258 211422 562494
rect 211186 555258 211422 555494
rect 211186 548258 211422 548494
rect 211186 541258 211422 541494
rect 211186 534258 211422 534494
rect 211186 527258 211422 527494
rect 211186 520258 211422 520494
rect 211186 513258 211422 513494
rect 211186 506258 211422 506494
rect 211186 499258 211422 499494
rect 211186 492258 211422 492494
rect 211186 485258 211422 485494
rect 211186 478258 211422 478494
rect 211186 471258 211422 471494
rect 211186 464258 211422 464494
rect 211186 457258 211422 457494
rect 211186 450258 211422 450494
rect 211186 443258 211422 443494
rect 211186 436258 211422 436494
rect 211186 429258 211422 429494
rect 211186 422258 211422 422494
rect 211186 415258 211422 415494
rect 211186 408258 211422 408494
rect 211186 401258 211422 401494
rect 211186 394258 211422 394494
rect 211186 387258 211422 387494
rect 211186 380258 211422 380494
rect 211186 373258 211422 373494
rect 211186 366258 211422 366494
rect 211186 359258 211422 359494
rect 211186 352258 211422 352494
rect 211186 345258 211422 345494
rect 211186 338258 211422 338494
rect 211186 331258 211422 331494
rect 211186 324258 211422 324494
rect 211186 317258 211422 317494
rect 211186 310258 211422 310494
rect 211186 303258 211422 303494
rect 211186 296258 211422 296494
rect 211186 289258 211422 289494
rect 211186 282258 211422 282494
rect 211186 275258 211422 275494
rect 211186 268258 211422 268494
rect 211186 261258 211422 261494
rect 211186 254258 211422 254494
rect 211186 247258 211422 247494
rect 211186 240258 211422 240494
rect 211186 233258 211422 233494
rect 211186 226258 211422 226494
rect 211186 219258 211422 219494
rect 211186 212258 211422 212494
rect 211186 205258 211422 205494
rect 211186 198258 211422 198494
rect 211186 191258 211422 191494
rect 211186 184258 211422 184494
rect 211186 177258 211422 177494
rect 211186 170258 211422 170494
rect 211186 163258 211422 163494
rect 211186 156258 211422 156494
rect 211186 149258 211422 149494
rect 211186 142258 211422 142494
rect 211186 135258 211422 135494
rect 211186 128258 211422 128494
rect 211186 121258 211422 121494
rect 211186 114258 211422 114494
rect 211186 107258 211422 107494
rect 211186 100258 211422 100494
rect 211186 93258 211422 93494
rect 211186 86258 211422 86494
rect 211186 79258 211422 79494
rect 211186 72258 211422 72494
rect 211186 65258 211422 65494
rect 211186 58258 211422 58494
rect 211186 51258 211422 51494
rect 211186 44258 211422 44494
rect 211186 37258 211422 37494
rect 211186 30258 211422 30494
rect 211186 23258 211422 23494
rect 211186 16258 211422 16494
rect 211186 9258 211422 9494
rect 211186 2258 211422 2494
rect 211186 -982 211422 -746
rect 211186 -1302 211422 -1066
rect 212918 705962 213154 706198
rect 212918 705642 213154 705878
rect 212918 696198 213154 696434
rect 212918 689198 213154 689434
rect 212918 682198 213154 682434
rect 212918 675198 213154 675434
rect 212918 668198 213154 668434
rect 212918 661198 213154 661434
rect 212918 654198 213154 654434
rect 212918 647198 213154 647434
rect 212918 640198 213154 640434
rect 212918 633198 213154 633434
rect 212918 626198 213154 626434
rect 212918 619198 213154 619434
rect 212918 612198 213154 612434
rect 212918 605198 213154 605434
rect 212918 598198 213154 598434
rect 212918 591198 213154 591434
rect 212918 584198 213154 584434
rect 212918 577198 213154 577434
rect 212918 570198 213154 570434
rect 212918 563198 213154 563434
rect 212918 556198 213154 556434
rect 212918 549198 213154 549434
rect 212918 542198 213154 542434
rect 212918 535198 213154 535434
rect 212918 528198 213154 528434
rect 212918 521198 213154 521434
rect 212918 514198 213154 514434
rect 212918 507198 213154 507434
rect 212918 500198 213154 500434
rect 212918 493198 213154 493434
rect 212918 486198 213154 486434
rect 212918 479198 213154 479434
rect 212918 472198 213154 472434
rect 212918 465198 213154 465434
rect 212918 458198 213154 458434
rect 212918 451198 213154 451434
rect 212918 444198 213154 444434
rect 212918 437198 213154 437434
rect 212918 430198 213154 430434
rect 212918 423198 213154 423434
rect 212918 416198 213154 416434
rect 212918 409198 213154 409434
rect 212918 402198 213154 402434
rect 212918 395198 213154 395434
rect 212918 388198 213154 388434
rect 212918 381198 213154 381434
rect 212918 374198 213154 374434
rect 212918 367198 213154 367434
rect 212918 360198 213154 360434
rect 212918 353198 213154 353434
rect 212918 346198 213154 346434
rect 212918 339198 213154 339434
rect 212918 332198 213154 332434
rect 212918 325198 213154 325434
rect 212918 318198 213154 318434
rect 212918 311198 213154 311434
rect 212918 304198 213154 304434
rect 212918 297198 213154 297434
rect 212918 290198 213154 290434
rect 212918 283198 213154 283434
rect 212918 276198 213154 276434
rect 212918 269198 213154 269434
rect 212918 262198 213154 262434
rect 212918 255198 213154 255434
rect 212918 248198 213154 248434
rect 212918 241198 213154 241434
rect 212918 234198 213154 234434
rect 212918 227198 213154 227434
rect 212918 220198 213154 220434
rect 212918 213198 213154 213434
rect 212918 206198 213154 206434
rect 212918 199198 213154 199434
rect 212918 192198 213154 192434
rect 212918 185198 213154 185434
rect 212918 178198 213154 178434
rect 212918 171198 213154 171434
rect 212918 164198 213154 164434
rect 212918 157198 213154 157434
rect 212918 150198 213154 150434
rect 212918 143198 213154 143434
rect 212918 136198 213154 136434
rect 212918 129198 213154 129434
rect 212918 122198 213154 122434
rect 212918 115198 213154 115434
rect 212918 108198 213154 108434
rect 212918 101198 213154 101434
rect 212918 94198 213154 94434
rect 212918 87198 213154 87434
rect 212918 80198 213154 80434
rect 212918 73198 213154 73434
rect 212918 66198 213154 66434
rect 212918 59198 213154 59434
rect 212918 52198 213154 52434
rect 212918 45198 213154 45434
rect 212918 38198 213154 38434
rect 212918 31198 213154 31434
rect 212918 24198 213154 24434
rect 212918 17198 213154 17434
rect 212918 10198 213154 10434
rect 212918 3198 213154 3434
rect 212918 -1942 213154 -1706
rect 212918 -2262 213154 -2026
rect 218186 705002 218422 705238
rect 218186 704682 218422 704918
rect 218186 695258 218422 695494
rect 218186 688258 218422 688494
rect 218186 681258 218422 681494
rect 218186 674258 218422 674494
rect 218186 667258 218422 667494
rect 218186 660258 218422 660494
rect 218186 653258 218422 653494
rect 218186 646258 218422 646494
rect 218186 639258 218422 639494
rect 218186 632258 218422 632494
rect 218186 625258 218422 625494
rect 218186 618258 218422 618494
rect 218186 611258 218422 611494
rect 218186 604258 218422 604494
rect 218186 597258 218422 597494
rect 218186 590258 218422 590494
rect 218186 583258 218422 583494
rect 218186 576258 218422 576494
rect 218186 569258 218422 569494
rect 218186 562258 218422 562494
rect 218186 555258 218422 555494
rect 218186 548258 218422 548494
rect 218186 541258 218422 541494
rect 218186 534258 218422 534494
rect 218186 527258 218422 527494
rect 218186 520258 218422 520494
rect 218186 513258 218422 513494
rect 218186 506258 218422 506494
rect 218186 499258 218422 499494
rect 218186 492258 218422 492494
rect 218186 485258 218422 485494
rect 218186 478258 218422 478494
rect 218186 471258 218422 471494
rect 218186 464258 218422 464494
rect 218186 457258 218422 457494
rect 218186 450258 218422 450494
rect 218186 443258 218422 443494
rect 218186 436258 218422 436494
rect 218186 429258 218422 429494
rect 218186 422258 218422 422494
rect 218186 415258 218422 415494
rect 218186 408258 218422 408494
rect 218186 401258 218422 401494
rect 218186 394258 218422 394494
rect 218186 387258 218422 387494
rect 218186 380258 218422 380494
rect 218186 373258 218422 373494
rect 218186 366258 218422 366494
rect 218186 359258 218422 359494
rect 218186 352258 218422 352494
rect 218186 345258 218422 345494
rect 218186 338258 218422 338494
rect 218186 331258 218422 331494
rect 218186 324258 218422 324494
rect 218186 317258 218422 317494
rect 218186 310258 218422 310494
rect 218186 303258 218422 303494
rect 218186 296258 218422 296494
rect 218186 289258 218422 289494
rect 218186 282258 218422 282494
rect 218186 275258 218422 275494
rect 218186 268258 218422 268494
rect 218186 261258 218422 261494
rect 218186 254258 218422 254494
rect 218186 247258 218422 247494
rect 218186 240258 218422 240494
rect 218186 233258 218422 233494
rect 218186 226258 218422 226494
rect 218186 219258 218422 219494
rect 218186 212258 218422 212494
rect 218186 205258 218422 205494
rect 218186 198258 218422 198494
rect 218186 191258 218422 191494
rect 218186 184258 218422 184494
rect 218186 177258 218422 177494
rect 218186 170258 218422 170494
rect 218186 163258 218422 163494
rect 218186 156258 218422 156494
rect 218186 149258 218422 149494
rect 218186 142258 218422 142494
rect 218186 135258 218422 135494
rect 218186 128258 218422 128494
rect 218186 121258 218422 121494
rect 218186 114258 218422 114494
rect 218186 107258 218422 107494
rect 218186 100258 218422 100494
rect 218186 93258 218422 93494
rect 218186 86258 218422 86494
rect 218186 79258 218422 79494
rect 218186 72258 218422 72494
rect 218186 65258 218422 65494
rect 218186 58258 218422 58494
rect 218186 51258 218422 51494
rect 218186 44258 218422 44494
rect 218186 37258 218422 37494
rect 218186 30258 218422 30494
rect 218186 23258 218422 23494
rect 218186 16258 218422 16494
rect 218186 9258 218422 9494
rect 218186 2258 218422 2494
rect 218186 -982 218422 -746
rect 218186 -1302 218422 -1066
rect 219918 705962 220154 706198
rect 219918 705642 220154 705878
rect 219918 696198 220154 696434
rect 219918 689198 220154 689434
rect 219918 682198 220154 682434
rect 219918 675198 220154 675434
rect 219918 668198 220154 668434
rect 219918 661198 220154 661434
rect 219918 654198 220154 654434
rect 219918 647198 220154 647434
rect 219918 640198 220154 640434
rect 219918 633198 220154 633434
rect 219918 626198 220154 626434
rect 219918 619198 220154 619434
rect 219918 612198 220154 612434
rect 219918 605198 220154 605434
rect 219918 598198 220154 598434
rect 219918 591198 220154 591434
rect 219918 584198 220154 584434
rect 219918 577198 220154 577434
rect 219918 570198 220154 570434
rect 219918 563198 220154 563434
rect 219918 556198 220154 556434
rect 219918 549198 220154 549434
rect 219918 542198 220154 542434
rect 219918 535198 220154 535434
rect 219918 528198 220154 528434
rect 219918 521198 220154 521434
rect 219918 514198 220154 514434
rect 219918 507198 220154 507434
rect 219918 500198 220154 500434
rect 219918 493198 220154 493434
rect 219918 486198 220154 486434
rect 219918 479198 220154 479434
rect 219918 472198 220154 472434
rect 219918 465198 220154 465434
rect 219918 458198 220154 458434
rect 219918 451198 220154 451434
rect 219918 444198 220154 444434
rect 219918 437198 220154 437434
rect 219918 430198 220154 430434
rect 219918 423198 220154 423434
rect 219918 416198 220154 416434
rect 219918 409198 220154 409434
rect 219918 402198 220154 402434
rect 219918 395198 220154 395434
rect 219918 388198 220154 388434
rect 219918 381198 220154 381434
rect 219918 374198 220154 374434
rect 219918 367198 220154 367434
rect 219918 360198 220154 360434
rect 219918 353198 220154 353434
rect 219918 346198 220154 346434
rect 219918 339198 220154 339434
rect 219918 332198 220154 332434
rect 219918 325198 220154 325434
rect 219918 318198 220154 318434
rect 219918 311198 220154 311434
rect 219918 304198 220154 304434
rect 219918 297198 220154 297434
rect 219918 290198 220154 290434
rect 219918 283198 220154 283434
rect 219918 276198 220154 276434
rect 219918 269198 220154 269434
rect 219918 262198 220154 262434
rect 219918 255198 220154 255434
rect 219918 248198 220154 248434
rect 219918 241198 220154 241434
rect 219918 234198 220154 234434
rect 219918 227198 220154 227434
rect 219918 220198 220154 220434
rect 219918 213198 220154 213434
rect 219918 206198 220154 206434
rect 219918 199198 220154 199434
rect 219918 192198 220154 192434
rect 219918 185198 220154 185434
rect 219918 178198 220154 178434
rect 219918 171198 220154 171434
rect 219918 164198 220154 164434
rect 219918 157198 220154 157434
rect 219918 150198 220154 150434
rect 219918 143198 220154 143434
rect 219918 136198 220154 136434
rect 219918 129198 220154 129434
rect 219918 122198 220154 122434
rect 219918 115198 220154 115434
rect 219918 108198 220154 108434
rect 219918 101198 220154 101434
rect 219918 94198 220154 94434
rect 219918 87198 220154 87434
rect 219918 80198 220154 80434
rect 219918 73198 220154 73434
rect 219918 66198 220154 66434
rect 219918 59198 220154 59434
rect 219918 52198 220154 52434
rect 219918 45198 220154 45434
rect 219918 38198 220154 38434
rect 219918 31198 220154 31434
rect 219918 24198 220154 24434
rect 219918 17198 220154 17434
rect 219918 10198 220154 10434
rect 219918 3198 220154 3434
rect 219918 -1942 220154 -1706
rect 219918 -2262 220154 -2026
rect 225186 705002 225422 705238
rect 225186 704682 225422 704918
rect 225186 695258 225422 695494
rect 225186 688258 225422 688494
rect 225186 681258 225422 681494
rect 225186 674258 225422 674494
rect 225186 667258 225422 667494
rect 225186 660258 225422 660494
rect 225186 653258 225422 653494
rect 225186 646258 225422 646494
rect 225186 639258 225422 639494
rect 225186 632258 225422 632494
rect 225186 625258 225422 625494
rect 225186 618258 225422 618494
rect 225186 611258 225422 611494
rect 225186 604258 225422 604494
rect 225186 597258 225422 597494
rect 225186 590258 225422 590494
rect 225186 583258 225422 583494
rect 225186 576258 225422 576494
rect 225186 569258 225422 569494
rect 225186 562258 225422 562494
rect 225186 555258 225422 555494
rect 225186 548258 225422 548494
rect 225186 541258 225422 541494
rect 225186 534258 225422 534494
rect 225186 527258 225422 527494
rect 225186 520258 225422 520494
rect 225186 513258 225422 513494
rect 225186 506258 225422 506494
rect 225186 499258 225422 499494
rect 225186 492258 225422 492494
rect 225186 485258 225422 485494
rect 225186 478258 225422 478494
rect 225186 471258 225422 471494
rect 225186 464258 225422 464494
rect 225186 457258 225422 457494
rect 225186 450258 225422 450494
rect 225186 443258 225422 443494
rect 225186 436258 225422 436494
rect 225186 429258 225422 429494
rect 225186 422258 225422 422494
rect 225186 415258 225422 415494
rect 225186 408258 225422 408494
rect 225186 401258 225422 401494
rect 225186 394258 225422 394494
rect 225186 387258 225422 387494
rect 225186 380258 225422 380494
rect 225186 373258 225422 373494
rect 225186 366258 225422 366494
rect 225186 359258 225422 359494
rect 225186 352258 225422 352494
rect 225186 345258 225422 345494
rect 225186 338258 225422 338494
rect 225186 331258 225422 331494
rect 225186 324258 225422 324494
rect 225186 317258 225422 317494
rect 225186 310258 225422 310494
rect 225186 303258 225422 303494
rect 225186 296258 225422 296494
rect 225186 289258 225422 289494
rect 225186 282258 225422 282494
rect 225186 275258 225422 275494
rect 225186 268258 225422 268494
rect 225186 261258 225422 261494
rect 225186 254258 225422 254494
rect 225186 247258 225422 247494
rect 225186 240258 225422 240494
rect 225186 233258 225422 233494
rect 225186 226258 225422 226494
rect 225186 219258 225422 219494
rect 225186 212258 225422 212494
rect 225186 205258 225422 205494
rect 225186 198258 225422 198494
rect 225186 191258 225422 191494
rect 225186 184258 225422 184494
rect 225186 177258 225422 177494
rect 225186 170258 225422 170494
rect 225186 163258 225422 163494
rect 225186 156258 225422 156494
rect 225186 149258 225422 149494
rect 225186 142258 225422 142494
rect 225186 135258 225422 135494
rect 225186 128258 225422 128494
rect 225186 121258 225422 121494
rect 225186 114258 225422 114494
rect 225186 107258 225422 107494
rect 225186 100258 225422 100494
rect 225186 93258 225422 93494
rect 225186 86258 225422 86494
rect 225186 79258 225422 79494
rect 225186 72258 225422 72494
rect 225186 65258 225422 65494
rect 225186 58258 225422 58494
rect 225186 51258 225422 51494
rect 225186 44258 225422 44494
rect 225186 37258 225422 37494
rect 225186 30258 225422 30494
rect 225186 23258 225422 23494
rect 225186 16258 225422 16494
rect 225186 9258 225422 9494
rect 225186 2258 225422 2494
rect 225186 -982 225422 -746
rect 225186 -1302 225422 -1066
rect 226918 705962 227154 706198
rect 226918 705642 227154 705878
rect 226918 696198 227154 696434
rect 226918 689198 227154 689434
rect 226918 682198 227154 682434
rect 226918 675198 227154 675434
rect 226918 668198 227154 668434
rect 226918 661198 227154 661434
rect 226918 654198 227154 654434
rect 226918 647198 227154 647434
rect 226918 640198 227154 640434
rect 226918 633198 227154 633434
rect 226918 626198 227154 626434
rect 226918 619198 227154 619434
rect 226918 612198 227154 612434
rect 226918 605198 227154 605434
rect 226918 598198 227154 598434
rect 226918 591198 227154 591434
rect 226918 584198 227154 584434
rect 226918 577198 227154 577434
rect 226918 570198 227154 570434
rect 226918 563198 227154 563434
rect 226918 556198 227154 556434
rect 226918 549198 227154 549434
rect 226918 542198 227154 542434
rect 226918 535198 227154 535434
rect 226918 528198 227154 528434
rect 226918 521198 227154 521434
rect 226918 514198 227154 514434
rect 226918 507198 227154 507434
rect 226918 500198 227154 500434
rect 226918 493198 227154 493434
rect 226918 486198 227154 486434
rect 226918 479198 227154 479434
rect 226918 472198 227154 472434
rect 226918 465198 227154 465434
rect 226918 458198 227154 458434
rect 226918 451198 227154 451434
rect 226918 444198 227154 444434
rect 226918 437198 227154 437434
rect 226918 430198 227154 430434
rect 226918 423198 227154 423434
rect 226918 416198 227154 416434
rect 226918 409198 227154 409434
rect 226918 402198 227154 402434
rect 226918 395198 227154 395434
rect 226918 388198 227154 388434
rect 226918 381198 227154 381434
rect 226918 374198 227154 374434
rect 226918 367198 227154 367434
rect 226918 360198 227154 360434
rect 226918 353198 227154 353434
rect 226918 346198 227154 346434
rect 226918 339198 227154 339434
rect 226918 332198 227154 332434
rect 226918 325198 227154 325434
rect 226918 318198 227154 318434
rect 226918 311198 227154 311434
rect 226918 304198 227154 304434
rect 226918 297198 227154 297434
rect 226918 290198 227154 290434
rect 226918 283198 227154 283434
rect 226918 276198 227154 276434
rect 226918 269198 227154 269434
rect 226918 262198 227154 262434
rect 226918 255198 227154 255434
rect 226918 248198 227154 248434
rect 226918 241198 227154 241434
rect 226918 234198 227154 234434
rect 226918 227198 227154 227434
rect 226918 220198 227154 220434
rect 226918 213198 227154 213434
rect 226918 206198 227154 206434
rect 226918 199198 227154 199434
rect 226918 192198 227154 192434
rect 226918 185198 227154 185434
rect 226918 178198 227154 178434
rect 226918 171198 227154 171434
rect 226918 164198 227154 164434
rect 226918 157198 227154 157434
rect 226918 150198 227154 150434
rect 226918 143198 227154 143434
rect 226918 136198 227154 136434
rect 226918 129198 227154 129434
rect 226918 122198 227154 122434
rect 226918 115198 227154 115434
rect 226918 108198 227154 108434
rect 226918 101198 227154 101434
rect 226918 94198 227154 94434
rect 226918 87198 227154 87434
rect 226918 80198 227154 80434
rect 226918 73198 227154 73434
rect 226918 66198 227154 66434
rect 226918 59198 227154 59434
rect 226918 52198 227154 52434
rect 226918 45198 227154 45434
rect 226918 38198 227154 38434
rect 226918 31198 227154 31434
rect 226918 24198 227154 24434
rect 226918 17198 227154 17434
rect 226918 10198 227154 10434
rect 226918 3198 227154 3434
rect 226918 -1942 227154 -1706
rect 226918 -2262 227154 -2026
rect 232186 705002 232422 705238
rect 232186 704682 232422 704918
rect 232186 695258 232422 695494
rect 232186 688258 232422 688494
rect 232186 681258 232422 681494
rect 232186 674258 232422 674494
rect 232186 667258 232422 667494
rect 232186 660258 232422 660494
rect 232186 653258 232422 653494
rect 232186 646258 232422 646494
rect 232186 639258 232422 639494
rect 232186 632258 232422 632494
rect 232186 625258 232422 625494
rect 232186 618258 232422 618494
rect 232186 611258 232422 611494
rect 232186 604258 232422 604494
rect 232186 597258 232422 597494
rect 232186 590258 232422 590494
rect 232186 583258 232422 583494
rect 232186 576258 232422 576494
rect 232186 569258 232422 569494
rect 232186 562258 232422 562494
rect 232186 555258 232422 555494
rect 232186 548258 232422 548494
rect 232186 541258 232422 541494
rect 232186 534258 232422 534494
rect 232186 527258 232422 527494
rect 232186 520258 232422 520494
rect 232186 513258 232422 513494
rect 232186 506258 232422 506494
rect 232186 499258 232422 499494
rect 232186 492258 232422 492494
rect 232186 485258 232422 485494
rect 232186 478258 232422 478494
rect 232186 471258 232422 471494
rect 232186 464258 232422 464494
rect 232186 457258 232422 457494
rect 232186 450258 232422 450494
rect 232186 443258 232422 443494
rect 232186 436258 232422 436494
rect 232186 429258 232422 429494
rect 232186 422258 232422 422494
rect 232186 415258 232422 415494
rect 232186 408258 232422 408494
rect 232186 401258 232422 401494
rect 232186 394258 232422 394494
rect 232186 387258 232422 387494
rect 232186 380258 232422 380494
rect 232186 373258 232422 373494
rect 232186 366258 232422 366494
rect 232186 359258 232422 359494
rect 232186 352258 232422 352494
rect 232186 345258 232422 345494
rect 232186 338258 232422 338494
rect 232186 331258 232422 331494
rect 232186 324258 232422 324494
rect 232186 317258 232422 317494
rect 232186 310258 232422 310494
rect 232186 303258 232422 303494
rect 232186 296258 232422 296494
rect 232186 289258 232422 289494
rect 232186 282258 232422 282494
rect 232186 275258 232422 275494
rect 232186 268258 232422 268494
rect 232186 261258 232422 261494
rect 232186 254258 232422 254494
rect 232186 247258 232422 247494
rect 232186 240258 232422 240494
rect 232186 233258 232422 233494
rect 232186 226258 232422 226494
rect 232186 219258 232422 219494
rect 232186 212258 232422 212494
rect 232186 205258 232422 205494
rect 232186 198258 232422 198494
rect 232186 191258 232422 191494
rect 232186 184258 232422 184494
rect 232186 177258 232422 177494
rect 232186 170258 232422 170494
rect 232186 163258 232422 163494
rect 232186 156258 232422 156494
rect 232186 149258 232422 149494
rect 232186 142258 232422 142494
rect 232186 135258 232422 135494
rect 232186 128258 232422 128494
rect 232186 121258 232422 121494
rect 232186 114258 232422 114494
rect 232186 107258 232422 107494
rect 232186 100258 232422 100494
rect 232186 93258 232422 93494
rect 232186 86258 232422 86494
rect 232186 79258 232422 79494
rect 232186 72258 232422 72494
rect 232186 65258 232422 65494
rect 232186 58258 232422 58494
rect 232186 51258 232422 51494
rect 232186 44258 232422 44494
rect 232186 37258 232422 37494
rect 232186 30258 232422 30494
rect 232186 23258 232422 23494
rect 232186 16258 232422 16494
rect 232186 9258 232422 9494
rect 232186 2258 232422 2494
rect 232186 -982 232422 -746
rect 232186 -1302 232422 -1066
rect 233918 705962 234154 706198
rect 233918 705642 234154 705878
rect 233918 696198 234154 696434
rect 233918 689198 234154 689434
rect 233918 682198 234154 682434
rect 233918 675198 234154 675434
rect 233918 668198 234154 668434
rect 233918 661198 234154 661434
rect 233918 654198 234154 654434
rect 233918 647198 234154 647434
rect 233918 640198 234154 640434
rect 233918 633198 234154 633434
rect 233918 626198 234154 626434
rect 233918 619198 234154 619434
rect 233918 612198 234154 612434
rect 233918 605198 234154 605434
rect 233918 598198 234154 598434
rect 233918 591198 234154 591434
rect 233918 584198 234154 584434
rect 233918 577198 234154 577434
rect 233918 570198 234154 570434
rect 233918 563198 234154 563434
rect 233918 556198 234154 556434
rect 233918 549198 234154 549434
rect 233918 542198 234154 542434
rect 233918 535198 234154 535434
rect 233918 528198 234154 528434
rect 233918 521198 234154 521434
rect 233918 514198 234154 514434
rect 233918 507198 234154 507434
rect 233918 500198 234154 500434
rect 233918 493198 234154 493434
rect 233918 486198 234154 486434
rect 233918 479198 234154 479434
rect 233918 472198 234154 472434
rect 233918 465198 234154 465434
rect 233918 458198 234154 458434
rect 233918 451198 234154 451434
rect 233918 444198 234154 444434
rect 233918 437198 234154 437434
rect 233918 430198 234154 430434
rect 233918 423198 234154 423434
rect 233918 416198 234154 416434
rect 233918 409198 234154 409434
rect 233918 402198 234154 402434
rect 233918 395198 234154 395434
rect 233918 388198 234154 388434
rect 233918 381198 234154 381434
rect 233918 374198 234154 374434
rect 233918 367198 234154 367434
rect 233918 360198 234154 360434
rect 233918 353198 234154 353434
rect 233918 346198 234154 346434
rect 233918 339198 234154 339434
rect 233918 332198 234154 332434
rect 233918 325198 234154 325434
rect 233918 318198 234154 318434
rect 233918 311198 234154 311434
rect 233918 304198 234154 304434
rect 233918 297198 234154 297434
rect 233918 290198 234154 290434
rect 233918 283198 234154 283434
rect 233918 276198 234154 276434
rect 233918 269198 234154 269434
rect 233918 262198 234154 262434
rect 233918 255198 234154 255434
rect 233918 248198 234154 248434
rect 233918 241198 234154 241434
rect 233918 234198 234154 234434
rect 233918 227198 234154 227434
rect 233918 220198 234154 220434
rect 233918 213198 234154 213434
rect 233918 206198 234154 206434
rect 233918 199198 234154 199434
rect 233918 192198 234154 192434
rect 233918 185198 234154 185434
rect 233918 178198 234154 178434
rect 233918 171198 234154 171434
rect 233918 164198 234154 164434
rect 233918 157198 234154 157434
rect 233918 150198 234154 150434
rect 233918 143198 234154 143434
rect 233918 136198 234154 136434
rect 233918 129198 234154 129434
rect 233918 122198 234154 122434
rect 233918 115198 234154 115434
rect 233918 108198 234154 108434
rect 233918 101198 234154 101434
rect 233918 94198 234154 94434
rect 233918 87198 234154 87434
rect 233918 80198 234154 80434
rect 233918 73198 234154 73434
rect 233918 66198 234154 66434
rect 233918 59198 234154 59434
rect 233918 52198 234154 52434
rect 233918 45198 234154 45434
rect 233918 38198 234154 38434
rect 233918 31198 234154 31434
rect 233918 24198 234154 24434
rect 233918 17198 234154 17434
rect 233918 10198 234154 10434
rect 233918 3198 234154 3434
rect 233918 -1942 234154 -1706
rect 233918 -2262 234154 -2026
rect 239186 705002 239422 705238
rect 239186 704682 239422 704918
rect 239186 695258 239422 695494
rect 239186 688258 239422 688494
rect 239186 681258 239422 681494
rect 239186 674258 239422 674494
rect 239186 667258 239422 667494
rect 239186 660258 239422 660494
rect 239186 653258 239422 653494
rect 239186 646258 239422 646494
rect 239186 639258 239422 639494
rect 239186 632258 239422 632494
rect 239186 625258 239422 625494
rect 239186 618258 239422 618494
rect 239186 611258 239422 611494
rect 239186 604258 239422 604494
rect 239186 597258 239422 597494
rect 239186 590258 239422 590494
rect 239186 583258 239422 583494
rect 239186 576258 239422 576494
rect 239186 569258 239422 569494
rect 239186 562258 239422 562494
rect 239186 555258 239422 555494
rect 239186 548258 239422 548494
rect 239186 541258 239422 541494
rect 239186 534258 239422 534494
rect 239186 527258 239422 527494
rect 239186 520258 239422 520494
rect 239186 513258 239422 513494
rect 239186 506258 239422 506494
rect 239186 499258 239422 499494
rect 239186 492258 239422 492494
rect 239186 485258 239422 485494
rect 239186 478258 239422 478494
rect 239186 471258 239422 471494
rect 239186 464258 239422 464494
rect 239186 457258 239422 457494
rect 239186 450258 239422 450494
rect 239186 443258 239422 443494
rect 239186 436258 239422 436494
rect 239186 429258 239422 429494
rect 239186 422258 239422 422494
rect 239186 415258 239422 415494
rect 239186 408258 239422 408494
rect 239186 401258 239422 401494
rect 239186 394258 239422 394494
rect 239186 387258 239422 387494
rect 239186 380258 239422 380494
rect 239186 373258 239422 373494
rect 239186 366258 239422 366494
rect 239186 359258 239422 359494
rect 239186 352258 239422 352494
rect 239186 345258 239422 345494
rect 239186 338258 239422 338494
rect 239186 331258 239422 331494
rect 239186 324258 239422 324494
rect 239186 317258 239422 317494
rect 239186 310258 239422 310494
rect 239186 303258 239422 303494
rect 239186 296258 239422 296494
rect 239186 289258 239422 289494
rect 239186 282258 239422 282494
rect 239186 275258 239422 275494
rect 239186 268258 239422 268494
rect 239186 261258 239422 261494
rect 239186 254258 239422 254494
rect 239186 247258 239422 247494
rect 239186 240258 239422 240494
rect 239186 233258 239422 233494
rect 239186 226258 239422 226494
rect 239186 219258 239422 219494
rect 239186 212258 239422 212494
rect 239186 205258 239422 205494
rect 239186 198258 239422 198494
rect 239186 191258 239422 191494
rect 239186 184258 239422 184494
rect 239186 177258 239422 177494
rect 239186 170258 239422 170494
rect 239186 163258 239422 163494
rect 239186 156258 239422 156494
rect 239186 149258 239422 149494
rect 239186 142258 239422 142494
rect 239186 135258 239422 135494
rect 239186 128258 239422 128494
rect 239186 121258 239422 121494
rect 239186 114258 239422 114494
rect 239186 107258 239422 107494
rect 239186 100258 239422 100494
rect 239186 93258 239422 93494
rect 239186 86258 239422 86494
rect 239186 79258 239422 79494
rect 239186 72258 239422 72494
rect 239186 65258 239422 65494
rect 239186 58258 239422 58494
rect 239186 51258 239422 51494
rect 239186 44258 239422 44494
rect 239186 37258 239422 37494
rect 239186 30258 239422 30494
rect 239186 23258 239422 23494
rect 239186 16258 239422 16494
rect 239186 9258 239422 9494
rect 239186 2258 239422 2494
rect 239186 -982 239422 -746
rect 239186 -1302 239422 -1066
rect 240918 705962 241154 706198
rect 240918 705642 241154 705878
rect 240918 696198 241154 696434
rect 240918 689198 241154 689434
rect 240918 682198 241154 682434
rect 240918 675198 241154 675434
rect 240918 668198 241154 668434
rect 240918 661198 241154 661434
rect 240918 654198 241154 654434
rect 240918 647198 241154 647434
rect 240918 640198 241154 640434
rect 240918 633198 241154 633434
rect 240918 626198 241154 626434
rect 240918 619198 241154 619434
rect 240918 612198 241154 612434
rect 240918 605198 241154 605434
rect 240918 598198 241154 598434
rect 240918 591198 241154 591434
rect 240918 584198 241154 584434
rect 240918 577198 241154 577434
rect 240918 570198 241154 570434
rect 240918 563198 241154 563434
rect 240918 556198 241154 556434
rect 240918 549198 241154 549434
rect 240918 542198 241154 542434
rect 240918 535198 241154 535434
rect 240918 528198 241154 528434
rect 240918 521198 241154 521434
rect 240918 514198 241154 514434
rect 240918 507198 241154 507434
rect 240918 500198 241154 500434
rect 240918 493198 241154 493434
rect 240918 486198 241154 486434
rect 240918 479198 241154 479434
rect 240918 472198 241154 472434
rect 240918 465198 241154 465434
rect 240918 458198 241154 458434
rect 240918 451198 241154 451434
rect 240918 444198 241154 444434
rect 240918 437198 241154 437434
rect 240918 430198 241154 430434
rect 240918 423198 241154 423434
rect 240918 416198 241154 416434
rect 240918 409198 241154 409434
rect 240918 402198 241154 402434
rect 240918 395198 241154 395434
rect 240918 388198 241154 388434
rect 240918 381198 241154 381434
rect 240918 374198 241154 374434
rect 240918 367198 241154 367434
rect 240918 360198 241154 360434
rect 240918 353198 241154 353434
rect 240918 346198 241154 346434
rect 240918 339198 241154 339434
rect 240918 332198 241154 332434
rect 240918 325198 241154 325434
rect 240918 318198 241154 318434
rect 240918 311198 241154 311434
rect 240918 304198 241154 304434
rect 240918 297198 241154 297434
rect 240918 290198 241154 290434
rect 240918 283198 241154 283434
rect 240918 276198 241154 276434
rect 240918 269198 241154 269434
rect 240918 262198 241154 262434
rect 240918 255198 241154 255434
rect 240918 248198 241154 248434
rect 240918 241198 241154 241434
rect 240918 234198 241154 234434
rect 240918 227198 241154 227434
rect 240918 220198 241154 220434
rect 240918 213198 241154 213434
rect 240918 206198 241154 206434
rect 240918 199198 241154 199434
rect 240918 192198 241154 192434
rect 240918 185198 241154 185434
rect 240918 178198 241154 178434
rect 240918 171198 241154 171434
rect 240918 164198 241154 164434
rect 240918 157198 241154 157434
rect 240918 150198 241154 150434
rect 240918 143198 241154 143434
rect 240918 136198 241154 136434
rect 240918 129198 241154 129434
rect 240918 122198 241154 122434
rect 240918 115198 241154 115434
rect 240918 108198 241154 108434
rect 240918 101198 241154 101434
rect 240918 94198 241154 94434
rect 240918 87198 241154 87434
rect 240918 80198 241154 80434
rect 240918 73198 241154 73434
rect 240918 66198 241154 66434
rect 240918 59198 241154 59434
rect 240918 52198 241154 52434
rect 240918 45198 241154 45434
rect 240918 38198 241154 38434
rect 240918 31198 241154 31434
rect 240918 24198 241154 24434
rect 240918 17198 241154 17434
rect 240918 10198 241154 10434
rect 240918 3198 241154 3434
rect 240918 -1942 241154 -1706
rect 240918 -2262 241154 -2026
rect 246186 705002 246422 705238
rect 246186 704682 246422 704918
rect 246186 695258 246422 695494
rect 246186 688258 246422 688494
rect 246186 681258 246422 681494
rect 246186 674258 246422 674494
rect 246186 667258 246422 667494
rect 246186 660258 246422 660494
rect 246186 653258 246422 653494
rect 246186 646258 246422 646494
rect 246186 639258 246422 639494
rect 246186 632258 246422 632494
rect 246186 625258 246422 625494
rect 246186 618258 246422 618494
rect 246186 611258 246422 611494
rect 246186 604258 246422 604494
rect 246186 597258 246422 597494
rect 246186 590258 246422 590494
rect 246186 583258 246422 583494
rect 246186 576258 246422 576494
rect 246186 569258 246422 569494
rect 246186 562258 246422 562494
rect 246186 555258 246422 555494
rect 246186 548258 246422 548494
rect 246186 541258 246422 541494
rect 246186 534258 246422 534494
rect 246186 527258 246422 527494
rect 246186 520258 246422 520494
rect 246186 513258 246422 513494
rect 246186 506258 246422 506494
rect 246186 499258 246422 499494
rect 246186 492258 246422 492494
rect 246186 485258 246422 485494
rect 246186 478258 246422 478494
rect 246186 471258 246422 471494
rect 246186 464258 246422 464494
rect 246186 457258 246422 457494
rect 246186 450258 246422 450494
rect 246186 443258 246422 443494
rect 246186 436258 246422 436494
rect 246186 429258 246422 429494
rect 246186 422258 246422 422494
rect 246186 415258 246422 415494
rect 246186 408258 246422 408494
rect 246186 401258 246422 401494
rect 246186 394258 246422 394494
rect 246186 387258 246422 387494
rect 246186 380258 246422 380494
rect 246186 373258 246422 373494
rect 246186 366258 246422 366494
rect 246186 359258 246422 359494
rect 246186 352258 246422 352494
rect 246186 345258 246422 345494
rect 246186 338258 246422 338494
rect 246186 331258 246422 331494
rect 246186 324258 246422 324494
rect 246186 317258 246422 317494
rect 246186 310258 246422 310494
rect 246186 303258 246422 303494
rect 246186 296258 246422 296494
rect 246186 289258 246422 289494
rect 246186 282258 246422 282494
rect 246186 275258 246422 275494
rect 246186 268258 246422 268494
rect 246186 261258 246422 261494
rect 246186 254258 246422 254494
rect 246186 247258 246422 247494
rect 246186 240258 246422 240494
rect 246186 233258 246422 233494
rect 246186 226258 246422 226494
rect 246186 219258 246422 219494
rect 246186 212258 246422 212494
rect 246186 205258 246422 205494
rect 246186 198258 246422 198494
rect 246186 191258 246422 191494
rect 246186 184258 246422 184494
rect 246186 177258 246422 177494
rect 246186 170258 246422 170494
rect 246186 163258 246422 163494
rect 246186 156258 246422 156494
rect 246186 149258 246422 149494
rect 246186 142258 246422 142494
rect 246186 135258 246422 135494
rect 246186 128258 246422 128494
rect 246186 121258 246422 121494
rect 246186 114258 246422 114494
rect 246186 107258 246422 107494
rect 246186 100258 246422 100494
rect 246186 93258 246422 93494
rect 246186 86258 246422 86494
rect 246186 79258 246422 79494
rect 246186 72258 246422 72494
rect 246186 65258 246422 65494
rect 246186 58258 246422 58494
rect 246186 51258 246422 51494
rect 246186 44258 246422 44494
rect 246186 37258 246422 37494
rect 246186 30258 246422 30494
rect 246186 23258 246422 23494
rect 246186 16258 246422 16494
rect 246186 9258 246422 9494
rect 246186 2258 246422 2494
rect 246186 -982 246422 -746
rect 246186 -1302 246422 -1066
rect 247918 705962 248154 706198
rect 247918 705642 248154 705878
rect 247918 696198 248154 696434
rect 247918 689198 248154 689434
rect 247918 682198 248154 682434
rect 247918 675198 248154 675434
rect 247918 668198 248154 668434
rect 247918 661198 248154 661434
rect 247918 654198 248154 654434
rect 247918 647198 248154 647434
rect 247918 640198 248154 640434
rect 247918 633198 248154 633434
rect 247918 626198 248154 626434
rect 247918 619198 248154 619434
rect 247918 612198 248154 612434
rect 247918 605198 248154 605434
rect 247918 598198 248154 598434
rect 247918 591198 248154 591434
rect 247918 584198 248154 584434
rect 247918 577198 248154 577434
rect 247918 570198 248154 570434
rect 247918 563198 248154 563434
rect 247918 556198 248154 556434
rect 247918 549198 248154 549434
rect 247918 542198 248154 542434
rect 247918 535198 248154 535434
rect 247918 528198 248154 528434
rect 247918 521198 248154 521434
rect 247918 514198 248154 514434
rect 247918 507198 248154 507434
rect 247918 500198 248154 500434
rect 247918 493198 248154 493434
rect 247918 486198 248154 486434
rect 247918 479198 248154 479434
rect 247918 472198 248154 472434
rect 247918 465198 248154 465434
rect 247918 458198 248154 458434
rect 247918 451198 248154 451434
rect 247918 444198 248154 444434
rect 247918 437198 248154 437434
rect 247918 430198 248154 430434
rect 247918 423198 248154 423434
rect 247918 416198 248154 416434
rect 247918 409198 248154 409434
rect 247918 402198 248154 402434
rect 247918 395198 248154 395434
rect 247918 388198 248154 388434
rect 247918 381198 248154 381434
rect 247918 374198 248154 374434
rect 247918 367198 248154 367434
rect 247918 360198 248154 360434
rect 247918 353198 248154 353434
rect 247918 346198 248154 346434
rect 247918 339198 248154 339434
rect 247918 332198 248154 332434
rect 247918 325198 248154 325434
rect 247918 318198 248154 318434
rect 247918 311198 248154 311434
rect 247918 304198 248154 304434
rect 247918 297198 248154 297434
rect 247918 290198 248154 290434
rect 247918 283198 248154 283434
rect 247918 276198 248154 276434
rect 247918 269198 248154 269434
rect 247918 262198 248154 262434
rect 247918 255198 248154 255434
rect 247918 248198 248154 248434
rect 247918 241198 248154 241434
rect 247918 234198 248154 234434
rect 247918 227198 248154 227434
rect 247918 220198 248154 220434
rect 247918 213198 248154 213434
rect 247918 206198 248154 206434
rect 247918 199198 248154 199434
rect 247918 192198 248154 192434
rect 247918 185198 248154 185434
rect 247918 178198 248154 178434
rect 247918 171198 248154 171434
rect 247918 164198 248154 164434
rect 247918 157198 248154 157434
rect 247918 150198 248154 150434
rect 247918 143198 248154 143434
rect 247918 136198 248154 136434
rect 247918 129198 248154 129434
rect 247918 122198 248154 122434
rect 247918 115198 248154 115434
rect 247918 108198 248154 108434
rect 247918 101198 248154 101434
rect 247918 94198 248154 94434
rect 247918 87198 248154 87434
rect 247918 80198 248154 80434
rect 247918 73198 248154 73434
rect 247918 66198 248154 66434
rect 247918 59198 248154 59434
rect 247918 52198 248154 52434
rect 247918 45198 248154 45434
rect 247918 38198 248154 38434
rect 247918 31198 248154 31434
rect 247918 24198 248154 24434
rect 247918 17198 248154 17434
rect 247918 10198 248154 10434
rect 247918 3198 248154 3434
rect 247918 -1942 248154 -1706
rect 247918 -2262 248154 -2026
rect 253186 705002 253422 705238
rect 253186 704682 253422 704918
rect 253186 695258 253422 695494
rect 253186 688258 253422 688494
rect 253186 681258 253422 681494
rect 253186 674258 253422 674494
rect 253186 667258 253422 667494
rect 253186 660258 253422 660494
rect 253186 653258 253422 653494
rect 253186 646258 253422 646494
rect 253186 639258 253422 639494
rect 253186 632258 253422 632494
rect 253186 625258 253422 625494
rect 253186 618258 253422 618494
rect 253186 611258 253422 611494
rect 253186 604258 253422 604494
rect 253186 597258 253422 597494
rect 253186 590258 253422 590494
rect 253186 583258 253422 583494
rect 253186 576258 253422 576494
rect 253186 569258 253422 569494
rect 253186 562258 253422 562494
rect 253186 555258 253422 555494
rect 253186 548258 253422 548494
rect 253186 541258 253422 541494
rect 253186 534258 253422 534494
rect 253186 527258 253422 527494
rect 253186 520258 253422 520494
rect 253186 513258 253422 513494
rect 253186 506258 253422 506494
rect 253186 499258 253422 499494
rect 253186 492258 253422 492494
rect 253186 485258 253422 485494
rect 253186 478258 253422 478494
rect 253186 471258 253422 471494
rect 253186 464258 253422 464494
rect 253186 457258 253422 457494
rect 253186 450258 253422 450494
rect 253186 443258 253422 443494
rect 253186 436258 253422 436494
rect 253186 429258 253422 429494
rect 253186 422258 253422 422494
rect 253186 415258 253422 415494
rect 253186 408258 253422 408494
rect 253186 401258 253422 401494
rect 253186 394258 253422 394494
rect 253186 387258 253422 387494
rect 253186 380258 253422 380494
rect 253186 373258 253422 373494
rect 253186 366258 253422 366494
rect 253186 359258 253422 359494
rect 253186 352258 253422 352494
rect 253186 345258 253422 345494
rect 253186 338258 253422 338494
rect 253186 331258 253422 331494
rect 253186 324258 253422 324494
rect 253186 317258 253422 317494
rect 253186 310258 253422 310494
rect 253186 303258 253422 303494
rect 253186 296258 253422 296494
rect 253186 289258 253422 289494
rect 253186 282258 253422 282494
rect 253186 275258 253422 275494
rect 253186 268258 253422 268494
rect 253186 261258 253422 261494
rect 253186 254258 253422 254494
rect 253186 247258 253422 247494
rect 253186 240258 253422 240494
rect 253186 233258 253422 233494
rect 253186 226258 253422 226494
rect 253186 219258 253422 219494
rect 253186 212258 253422 212494
rect 253186 205258 253422 205494
rect 253186 198258 253422 198494
rect 253186 191258 253422 191494
rect 253186 184258 253422 184494
rect 253186 177258 253422 177494
rect 253186 170258 253422 170494
rect 253186 163258 253422 163494
rect 253186 156258 253422 156494
rect 253186 149258 253422 149494
rect 253186 142258 253422 142494
rect 253186 135258 253422 135494
rect 253186 128258 253422 128494
rect 253186 121258 253422 121494
rect 253186 114258 253422 114494
rect 253186 107258 253422 107494
rect 253186 100258 253422 100494
rect 253186 93258 253422 93494
rect 253186 86258 253422 86494
rect 253186 79258 253422 79494
rect 253186 72258 253422 72494
rect 253186 65258 253422 65494
rect 253186 58258 253422 58494
rect 253186 51258 253422 51494
rect 253186 44258 253422 44494
rect 253186 37258 253422 37494
rect 253186 30258 253422 30494
rect 253186 23258 253422 23494
rect 253186 16258 253422 16494
rect 253186 9258 253422 9494
rect 253186 2258 253422 2494
rect 253186 -982 253422 -746
rect 253186 -1302 253422 -1066
rect 254918 705962 255154 706198
rect 254918 705642 255154 705878
rect 254918 696198 255154 696434
rect 254918 689198 255154 689434
rect 254918 682198 255154 682434
rect 254918 675198 255154 675434
rect 254918 668198 255154 668434
rect 254918 661198 255154 661434
rect 254918 654198 255154 654434
rect 254918 647198 255154 647434
rect 254918 640198 255154 640434
rect 254918 633198 255154 633434
rect 254918 626198 255154 626434
rect 254918 619198 255154 619434
rect 254918 612198 255154 612434
rect 254918 605198 255154 605434
rect 254918 598198 255154 598434
rect 254918 591198 255154 591434
rect 254918 584198 255154 584434
rect 254918 577198 255154 577434
rect 254918 570198 255154 570434
rect 254918 563198 255154 563434
rect 254918 556198 255154 556434
rect 254918 549198 255154 549434
rect 254918 542198 255154 542434
rect 254918 535198 255154 535434
rect 254918 528198 255154 528434
rect 254918 521198 255154 521434
rect 254918 514198 255154 514434
rect 254918 507198 255154 507434
rect 254918 500198 255154 500434
rect 254918 493198 255154 493434
rect 254918 486198 255154 486434
rect 254918 479198 255154 479434
rect 254918 472198 255154 472434
rect 254918 465198 255154 465434
rect 254918 458198 255154 458434
rect 254918 451198 255154 451434
rect 254918 444198 255154 444434
rect 254918 437198 255154 437434
rect 254918 430198 255154 430434
rect 254918 423198 255154 423434
rect 254918 416198 255154 416434
rect 254918 409198 255154 409434
rect 254918 402198 255154 402434
rect 254918 395198 255154 395434
rect 254918 388198 255154 388434
rect 254918 381198 255154 381434
rect 254918 374198 255154 374434
rect 254918 367198 255154 367434
rect 254918 360198 255154 360434
rect 254918 353198 255154 353434
rect 254918 346198 255154 346434
rect 254918 339198 255154 339434
rect 254918 332198 255154 332434
rect 254918 325198 255154 325434
rect 254918 318198 255154 318434
rect 254918 311198 255154 311434
rect 254918 304198 255154 304434
rect 254918 297198 255154 297434
rect 254918 290198 255154 290434
rect 254918 283198 255154 283434
rect 254918 276198 255154 276434
rect 254918 269198 255154 269434
rect 254918 262198 255154 262434
rect 254918 255198 255154 255434
rect 254918 248198 255154 248434
rect 254918 241198 255154 241434
rect 254918 234198 255154 234434
rect 254918 227198 255154 227434
rect 254918 220198 255154 220434
rect 254918 213198 255154 213434
rect 254918 206198 255154 206434
rect 254918 199198 255154 199434
rect 254918 192198 255154 192434
rect 254918 185198 255154 185434
rect 254918 178198 255154 178434
rect 254918 171198 255154 171434
rect 254918 164198 255154 164434
rect 254918 157198 255154 157434
rect 254918 150198 255154 150434
rect 254918 143198 255154 143434
rect 254918 136198 255154 136434
rect 254918 129198 255154 129434
rect 254918 122198 255154 122434
rect 254918 115198 255154 115434
rect 254918 108198 255154 108434
rect 254918 101198 255154 101434
rect 254918 94198 255154 94434
rect 254918 87198 255154 87434
rect 254918 80198 255154 80434
rect 254918 73198 255154 73434
rect 254918 66198 255154 66434
rect 254918 59198 255154 59434
rect 254918 52198 255154 52434
rect 254918 45198 255154 45434
rect 254918 38198 255154 38434
rect 254918 31198 255154 31434
rect 254918 24198 255154 24434
rect 254918 17198 255154 17434
rect 254918 10198 255154 10434
rect 254918 3198 255154 3434
rect 254918 -1942 255154 -1706
rect 254918 -2262 255154 -2026
rect 260186 705002 260422 705238
rect 260186 704682 260422 704918
rect 260186 695258 260422 695494
rect 260186 688258 260422 688494
rect 260186 681258 260422 681494
rect 260186 674258 260422 674494
rect 260186 667258 260422 667494
rect 260186 660258 260422 660494
rect 260186 653258 260422 653494
rect 260186 646258 260422 646494
rect 260186 639258 260422 639494
rect 260186 632258 260422 632494
rect 260186 625258 260422 625494
rect 260186 618258 260422 618494
rect 260186 611258 260422 611494
rect 260186 604258 260422 604494
rect 260186 597258 260422 597494
rect 260186 590258 260422 590494
rect 260186 583258 260422 583494
rect 260186 576258 260422 576494
rect 260186 569258 260422 569494
rect 260186 562258 260422 562494
rect 260186 555258 260422 555494
rect 260186 548258 260422 548494
rect 260186 541258 260422 541494
rect 260186 534258 260422 534494
rect 260186 527258 260422 527494
rect 260186 520258 260422 520494
rect 260186 513258 260422 513494
rect 260186 506258 260422 506494
rect 260186 499258 260422 499494
rect 260186 492258 260422 492494
rect 260186 485258 260422 485494
rect 260186 478258 260422 478494
rect 260186 471258 260422 471494
rect 260186 464258 260422 464494
rect 260186 457258 260422 457494
rect 260186 450258 260422 450494
rect 260186 443258 260422 443494
rect 260186 436258 260422 436494
rect 260186 429258 260422 429494
rect 260186 422258 260422 422494
rect 260186 415258 260422 415494
rect 260186 408258 260422 408494
rect 260186 401258 260422 401494
rect 260186 394258 260422 394494
rect 260186 387258 260422 387494
rect 260186 380258 260422 380494
rect 260186 373258 260422 373494
rect 260186 366258 260422 366494
rect 260186 359258 260422 359494
rect 260186 352258 260422 352494
rect 260186 345258 260422 345494
rect 260186 338258 260422 338494
rect 260186 331258 260422 331494
rect 260186 324258 260422 324494
rect 260186 317258 260422 317494
rect 260186 310258 260422 310494
rect 260186 303258 260422 303494
rect 260186 296258 260422 296494
rect 260186 289258 260422 289494
rect 260186 282258 260422 282494
rect 260186 275258 260422 275494
rect 260186 268258 260422 268494
rect 260186 261258 260422 261494
rect 260186 254258 260422 254494
rect 260186 247258 260422 247494
rect 260186 240258 260422 240494
rect 260186 233258 260422 233494
rect 260186 226258 260422 226494
rect 260186 219258 260422 219494
rect 260186 212258 260422 212494
rect 260186 205258 260422 205494
rect 260186 198258 260422 198494
rect 260186 191258 260422 191494
rect 260186 184258 260422 184494
rect 260186 177258 260422 177494
rect 260186 170258 260422 170494
rect 260186 163258 260422 163494
rect 260186 156258 260422 156494
rect 260186 149258 260422 149494
rect 260186 142258 260422 142494
rect 260186 135258 260422 135494
rect 260186 128258 260422 128494
rect 260186 121258 260422 121494
rect 260186 114258 260422 114494
rect 260186 107258 260422 107494
rect 260186 100258 260422 100494
rect 260186 93258 260422 93494
rect 260186 86258 260422 86494
rect 260186 79258 260422 79494
rect 260186 72258 260422 72494
rect 260186 65258 260422 65494
rect 260186 58258 260422 58494
rect 260186 51258 260422 51494
rect 260186 44258 260422 44494
rect 260186 37258 260422 37494
rect 260186 30258 260422 30494
rect 260186 23258 260422 23494
rect 260186 16258 260422 16494
rect 260186 9258 260422 9494
rect 260186 2258 260422 2494
rect 260186 -982 260422 -746
rect 260186 -1302 260422 -1066
rect 261918 705962 262154 706198
rect 261918 705642 262154 705878
rect 261918 696198 262154 696434
rect 261918 689198 262154 689434
rect 261918 682198 262154 682434
rect 261918 675198 262154 675434
rect 261918 668198 262154 668434
rect 261918 661198 262154 661434
rect 261918 654198 262154 654434
rect 261918 647198 262154 647434
rect 261918 640198 262154 640434
rect 261918 633198 262154 633434
rect 261918 626198 262154 626434
rect 261918 619198 262154 619434
rect 261918 612198 262154 612434
rect 261918 605198 262154 605434
rect 261918 598198 262154 598434
rect 261918 591198 262154 591434
rect 261918 584198 262154 584434
rect 261918 577198 262154 577434
rect 261918 570198 262154 570434
rect 261918 563198 262154 563434
rect 261918 556198 262154 556434
rect 261918 549198 262154 549434
rect 261918 542198 262154 542434
rect 261918 535198 262154 535434
rect 261918 528198 262154 528434
rect 261918 521198 262154 521434
rect 261918 514198 262154 514434
rect 261918 507198 262154 507434
rect 261918 500198 262154 500434
rect 261918 493198 262154 493434
rect 261918 486198 262154 486434
rect 261918 479198 262154 479434
rect 261918 472198 262154 472434
rect 261918 465198 262154 465434
rect 261918 458198 262154 458434
rect 261918 451198 262154 451434
rect 261918 444198 262154 444434
rect 261918 437198 262154 437434
rect 261918 430198 262154 430434
rect 261918 423198 262154 423434
rect 261918 416198 262154 416434
rect 261918 409198 262154 409434
rect 261918 402198 262154 402434
rect 261918 395198 262154 395434
rect 261918 388198 262154 388434
rect 261918 381198 262154 381434
rect 261918 374198 262154 374434
rect 261918 367198 262154 367434
rect 261918 360198 262154 360434
rect 261918 353198 262154 353434
rect 261918 346198 262154 346434
rect 261918 339198 262154 339434
rect 261918 332198 262154 332434
rect 261918 325198 262154 325434
rect 261918 318198 262154 318434
rect 261918 311198 262154 311434
rect 261918 304198 262154 304434
rect 261918 297198 262154 297434
rect 261918 290198 262154 290434
rect 261918 283198 262154 283434
rect 261918 276198 262154 276434
rect 261918 269198 262154 269434
rect 261918 262198 262154 262434
rect 261918 255198 262154 255434
rect 261918 248198 262154 248434
rect 261918 241198 262154 241434
rect 261918 234198 262154 234434
rect 261918 227198 262154 227434
rect 261918 220198 262154 220434
rect 261918 213198 262154 213434
rect 261918 206198 262154 206434
rect 261918 199198 262154 199434
rect 261918 192198 262154 192434
rect 261918 185198 262154 185434
rect 261918 178198 262154 178434
rect 261918 171198 262154 171434
rect 261918 164198 262154 164434
rect 261918 157198 262154 157434
rect 261918 150198 262154 150434
rect 261918 143198 262154 143434
rect 261918 136198 262154 136434
rect 261918 129198 262154 129434
rect 261918 122198 262154 122434
rect 261918 115198 262154 115434
rect 261918 108198 262154 108434
rect 261918 101198 262154 101434
rect 261918 94198 262154 94434
rect 261918 87198 262154 87434
rect 261918 80198 262154 80434
rect 261918 73198 262154 73434
rect 261918 66198 262154 66434
rect 261918 59198 262154 59434
rect 261918 52198 262154 52434
rect 261918 45198 262154 45434
rect 261918 38198 262154 38434
rect 261918 31198 262154 31434
rect 261918 24198 262154 24434
rect 261918 17198 262154 17434
rect 261918 10198 262154 10434
rect 261918 3198 262154 3434
rect 261918 -1942 262154 -1706
rect 261918 -2262 262154 -2026
rect 267186 705002 267422 705238
rect 267186 704682 267422 704918
rect 267186 695258 267422 695494
rect 267186 688258 267422 688494
rect 267186 681258 267422 681494
rect 267186 674258 267422 674494
rect 267186 667258 267422 667494
rect 267186 660258 267422 660494
rect 267186 653258 267422 653494
rect 267186 646258 267422 646494
rect 267186 639258 267422 639494
rect 267186 632258 267422 632494
rect 267186 625258 267422 625494
rect 267186 618258 267422 618494
rect 267186 611258 267422 611494
rect 267186 604258 267422 604494
rect 267186 597258 267422 597494
rect 267186 590258 267422 590494
rect 267186 583258 267422 583494
rect 267186 576258 267422 576494
rect 267186 569258 267422 569494
rect 267186 562258 267422 562494
rect 267186 555258 267422 555494
rect 267186 548258 267422 548494
rect 267186 541258 267422 541494
rect 267186 534258 267422 534494
rect 267186 527258 267422 527494
rect 267186 520258 267422 520494
rect 267186 513258 267422 513494
rect 267186 506258 267422 506494
rect 267186 499258 267422 499494
rect 267186 492258 267422 492494
rect 267186 485258 267422 485494
rect 267186 478258 267422 478494
rect 267186 471258 267422 471494
rect 267186 464258 267422 464494
rect 267186 457258 267422 457494
rect 267186 450258 267422 450494
rect 267186 443258 267422 443494
rect 267186 436258 267422 436494
rect 267186 429258 267422 429494
rect 267186 422258 267422 422494
rect 267186 415258 267422 415494
rect 267186 408258 267422 408494
rect 267186 401258 267422 401494
rect 267186 394258 267422 394494
rect 267186 387258 267422 387494
rect 267186 380258 267422 380494
rect 267186 373258 267422 373494
rect 267186 366258 267422 366494
rect 267186 359258 267422 359494
rect 267186 352258 267422 352494
rect 267186 345258 267422 345494
rect 267186 338258 267422 338494
rect 267186 331258 267422 331494
rect 267186 324258 267422 324494
rect 267186 317258 267422 317494
rect 267186 310258 267422 310494
rect 267186 303258 267422 303494
rect 267186 296258 267422 296494
rect 267186 289258 267422 289494
rect 267186 282258 267422 282494
rect 267186 275258 267422 275494
rect 267186 268258 267422 268494
rect 267186 261258 267422 261494
rect 267186 254258 267422 254494
rect 267186 247258 267422 247494
rect 267186 240258 267422 240494
rect 267186 233258 267422 233494
rect 267186 226258 267422 226494
rect 267186 219258 267422 219494
rect 267186 212258 267422 212494
rect 267186 205258 267422 205494
rect 267186 198258 267422 198494
rect 267186 191258 267422 191494
rect 267186 184258 267422 184494
rect 267186 177258 267422 177494
rect 267186 170258 267422 170494
rect 267186 163258 267422 163494
rect 267186 156258 267422 156494
rect 267186 149258 267422 149494
rect 267186 142258 267422 142494
rect 267186 135258 267422 135494
rect 267186 128258 267422 128494
rect 267186 121258 267422 121494
rect 267186 114258 267422 114494
rect 267186 107258 267422 107494
rect 267186 100258 267422 100494
rect 267186 93258 267422 93494
rect 267186 86258 267422 86494
rect 267186 79258 267422 79494
rect 267186 72258 267422 72494
rect 267186 65258 267422 65494
rect 267186 58258 267422 58494
rect 267186 51258 267422 51494
rect 267186 44258 267422 44494
rect 267186 37258 267422 37494
rect 267186 30258 267422 30494
rect 267186 23258 267422 23494
rect 267186 16258 267422 16494
rect 267186 9258 267422 9494
rect 267186 2258 267422 2494
rect 267186 -982 267422 -746
rect 267186 -1302 267422 -1066
rect 268918 705962 269154 706198
rect 268918 705642 269154 705878
rect 268918 696198 269154 696434
rect 268918 689198 269154 689434
rect 268918 682198 269154 682434
rect 268918 675198 269154 675434
rect 268918 668198 269154 668434
rect 268918 661198 269154 661434
rect 268918 654198 269154 654434
rect 268918 647198 269154 647434
rect 268918 640198 269154 640434
rect 268918 633198 269154 633434
rect 268918 626198 269154 626434
rect 268918 619198 269154 619434
rect 268918 612198 269154 612434
rect 268918 605198 269154 605434
rect 268918 598198 269154 598434
rect 268918 591198 269154 591434
rect 268918 584198 269154 584434
rect 268918 577198 269154 577434
rect 268918 570198 269154 570434
rect 268918 563198 269154 563434
rect 268918 556198 269154 556434
rect 268918 549198 269154 549434
rect 268918 542198 269154 542434
rect 268918 535198 269154 535434
rect 268918 528198 269154 528434
rect 268918 521198 269154 521434
rect 268918 514198 269154 514434
rect 268918 507198 269154 507434
rect 268918 500198 269154 500434
rect 268918 493198 269154 493434
rect 268918 486198 269154 486434
rect 268918 479198 269154 479434
rect 268918 472198 269154 472434
rect 268918 465198 269154 465434
rect 268918 458198 269154 458434
rect 268918 451198 269154 451434
rect 268918 444198 269154 444434
rect 268918 437198 269154 437434
rect 268918 430198 269154 430434
rect 268918 423198 269154 423434
rect 268918 416198 269154 416434
rect 268918 409198 269154 409434
rect 268918 402198 269154 402434
rect 268918 395198 269154 395434
rect 268918 388198 269154 388434
rect 268918 381198 269154 381434
rect 268918 374198 269154 374434
rect 268918 367198 269154 367434
rect 268918 360198 269154 360434
rect 268918 353198 269154 353434
rect 268918 346198 269154 346434
rect 268918 339198 269154 339434
rect 268918 332198 269154 332434
rect 268918 325198 269154 325434
rect 268918 318198 269154 318434
rect 268918 311198 269154 311434
rect 268918 304198 269154 304434
rect 268918 297198 269154 297434
rect 268918 290198 269154 290434
rect 268918 283198 269154 283434
rect 268918 276198 269154 276434
rect 268918 269198 269154 269434
rect 268918 262198 269154 262434
rect 268918 255198 269154 255434
rect 268918 248198 269154 248434
rect 268918 241198 269154 241434
rect 268918 234198 269154 234434
rect 268918 227198 269154 227434
rect 268918 220198 269154 220434
rect 268918 213198 269154 213434
rect 268918 206198 269154 206434
rect 268918 199198 269154 199434
rect 268918 192198 269154 192434
rect 268918 185198 269154 185434
rect 268918 178198 269154 178434
rect 268918 171198 269154 171434
rect 268918 164198 269154 164434
rect 268918 157198 269154 157434
rect 268918 150198 269154 150434
rect 268918 143198 269154 143434
rect 268918 136198 269154 136434
rect 268918 129198 269154 129434
rect 268918 122198 269154 122434
rect 268918 115198 269154 115434
rect 268918 108198 269154 108434
rect 268918 101198 269154 101434
rect 268918 94198 269154 94434
rect 268918 87198 269154 87434
rect 268918 80198 269154 80434
rect 268918 73198 269154 73434
rect 268918 66198 269154 66434
rect 268918 59198 269154 59434
rect 268918 52198 269154 52434
rect 268918 45198 269154 45434
rect 268918 38198 269154 38434
rect 268918 31198 269154 31434
rect 268918 24198 269154 24434
rect 268918 17198 269154 17434
rect 268918 10198 269154 10434
rect 268918 3198 269154 3434
rect 268918 -1942 269154 -1706
rect 268918 -2262 269154 -2026
rect 274186 705002 274422 705238
rect 274186 704682 274422 704918
rect 274186 695258 274422 695494
rect 274186 688258 274422 688494
rect 274186 681258 274422 681494
rect 274186 674258 274422 674494
rect 274186 667258 274422 667494
rect 274186 660258 274422 660494
rect 274186 653258 274422 653494
rect 274186 646258 274422 646494
rect 274186 639258 274422 639494
rect 274186 632258 274422 632494
rect 274186 625258 274422 625494
rect 274186 618258 274422 618494
rect 274186 611258 274422 611494
rect 274186 604258 274422 604494
rect 274186 597258 274422 597494
rect 274186 590258 274422 590494
rect 274186 583258 274422 583494
rect 274186 576258 274422 576494
rect 274186 569258 274422 569494
rect 274186 562258 274422 562494
rect 274186 555258 274422 555494
rect 274186 548258 274422 548494
rect 274186 541258 274422 541494
rect 274186 534258 274422 534494
rect 274186 527258 274422 527494
rect 274186 520258 274422 520494
rect 274186 513258 274422 513494
rect 274186 506258 274422 506494
rect 274186 499258 274422 499494
rect 274186 492258 274422 492494
rect 274186 485258 274422 485494
rect 274186 478258 274422 478494
rect 274186 471258 274422 471494
rect 274186 464258 274422 464494
rect 274186 457258 274422 457494
rect 274186 450258 274422 450494
rect 274186 443258 274422 443494
rect 274186 436258 274422 436494
rect 274186 429258 274422 429494
rect 274186 422258 274422 422494
rect 274186 415258 274422 415494
rect 274186 408258 274422 408494
rect 274186 401258 274422 401494
rect 274186 394258 274422 394494
rect 274186 387258 274422 387494
rect 274186 380258 274422 380494
rect 274186 373258 274422 373494
rect 274186 366258 274422 366494
rect 274186 359258 274422 359494
rect 274186 352258 274422 352494
rect 274186 345258 274422 345494
rect 274186 338258 274422 338494
rect 274186 331258 274422 331494
rect 274186 324258 274422 324494
rect 274186 317258 274422 317494
rect 274186 310258 274422 310494
rect 274186 303258 274422 303494
rect 274186 296258 274422 296494
rect 274186 289258 274422 289494
rect 274186 282258 274422 282494
rect 274186 275258 274422 275494
rect 274186 268258 274422 268494
rect 274186 261258 274422 261494
rect 274186 254258 274422 254494
rect 274186 247258 274422 247494
rect 274186 240258 274422 240494
rect 274186 233258 274422 233494
rect 274186 226258 274422 226494
rect 274186 219258 274422 219494
rect 274186 212258 274422 212494
rect 274186 205258 274422 205494
rect 274186 198258 274422 198494
rect 274186 191258 274422 191494
rect 274186 184258 274422 184494
rect 274186 177258 274422 177494
rect 274186 170258 274422 170494
rect 274186 163258 274422 163494
rect 274186 156258 274422 156494
rect 274186 149258 274422 149494
rect 274186 142258 274422 142494
rect 274186 135258 274422 135494
rect 274186 128258 274422 128494
rect 274186 121258 274422 121494
rect 274186 114258 274422 114494
rect 274186 107258 274422 107494
rect 274186 100258 274422 100494
rect 274186 93258 274422 93494
rect 274186 86258 274422 86494
rect 274186 79258 274422 79494
rect 274186 72258 274422 72494
rect 274186 65258 274422 65494
rect 274186 58258 274422 58494
rect 274186 51258 274422 51494
rect 274186 44258 274422 44494
rect 274186 37258 274422 37494
rect 274186 30258 274422 30494
rect 274186 23258 274422 23494
rect 274186 16258 274422 16494
rect 274186 9258 274422 9494
rect 274186 2258 274422 2494
rect 274186 -982 274422 -746
rect 274186 -1302 274422 -1066
rect 275918 705962 276154 706198
rect 275918 705642 276154 705878
rect 275918 696198 276154 696434
rect 275918 689198 276154 689434
rect 275918 682198 276154 682434
rect 275918 675198 276154 675434
rect 275918 668198 276154 668434
rect 275918 661198 276154 661434
rect 275918 654198 276154 654434
rect 275918 647198 276154 647434
rect 275918 640198 276154 640434
rect 275918 633198 276154 633434
rect 275918 626198 276154 626434
rect 275918 619198 276154 619434
rect 275918 612198 276154 612434
rect 275918 605198 276154 605434
rect 275918 598198 276154 598434
rect 275918 591198 276154 591434
rect 275918 584198 276154 584434
rect 275918 577198 276154 577434
rect 275918 570198 276154 570434
rect 275918 563198 276154 563434
rect 275918 556198 276154 556434
rect 275918 549198 276154 549434
rect 275918 542198 276154 542434
rect 275918 535198 276154 535434
rect 275918 528198 276154 528434
rect 275918 521198 276154 521434
rect 275918 514198 276154 514434
rect 275918 507198 276154 507434
rect 275918 500198 276154 500434
rect 275918 493198 276154 493434
rect 275918 486198 276154 486434
rect 275918 479198 276154 479434
rect 275918 472198 276154 472434
rect 275918 465198 276154 465434
rect 275918 458198 276154 458434
rect 275918 451198 276154 451434
rect 275918 444198 276154 444434
rect 275918 437198 276154 437434
rect 275918 430198 276154 430434
rect 275918 423198 276154 423434
rect 275918 416198 276154 416434
rect 275918 409198 276154 409434
rect 275918 402198 276154 402434
rect 275918 395198 276154 395434
rect 275918 388198 276154 388434
rect 275918 381198 276154 381434
rect 275918 374198 276154 374434
rect 275918 367198 276154 367434
rect 275918 360198 276154 360434
rect 275918 353198 276154 353434
rect 275918 346198 276154 346434
rect 275918 339198 276154 339434
rect 275918 332198 276154 332434
rect 275918 325198 276154 325434
rect 275918 318198 276154 318434
rect 275918 311198 276154 311434
rect 275918 304198 276154 304434
rect 275918 297198 276154 297434
rect 275918 290198 276154 290434
rect 275918 283198 276154 283434
rect 275918 276198 276154 276434
rect 275918 269198 276154 269434
rect 275918 262198 276154 262434
rect 275918 255198 276154 255434
rect 275918 248198 276154 248434
rect 275918 241198 276154 241434
rect 275918 234198 276154 234434
rect 275918 227198 276154 227434
rect 275918 220198 276154 220434
rect 275918 213198 276154 213434
rect 275918 206198 276154 206434
rect 275918 199198 276154 199434
rect 275918 192198 276154 192434
rect 275918 185198 276154 185434
rect 275918 178198 276154 178434
rect 275918 171198 276154 171434
rect 275918 164198 276154 164434
rect 275918 157198 276154 157434
rect 275918 150198 276154 150434
rect 275918 143198 276154 143434
rect 275918 136198 276154 136434
rect 275918 129198 276154 129434
rect 275918 122198 276154 122434
rect 275918 115198 276154 115434
rect 275918 108198 276154 108434
rect 275918 101198 276154 101434
rect 275918 94198 276154 94434
rect 275918 87198 276154 87434
rect 275918 80198 276154 80434
rect 275918 73198 276154 73434
rect 275918 66198 276154 66434
rect 275918 59198 276154 59434
rect 275918 52198 276154 52434
rect 275918 45198 276154 45434
rect 275918 38198 276154 38434
rect 275918 31198 276154 31434
rect 275918 24198 276154 24434
rect 275918 17198 276154 17434
rect 275918 10198 276154 10434
rect 275918 3198 276154 3434
rect 275918 -1942 276154 -1706
rect 275918 -2262 276154 -2026
rect 281186 705002 281422 705238
rect 281186 704682 281422 704918
rect 281186 695258 281422 695494
rect 281186 688258 281422 688494
rect 281186 681258 281422 681494
rect 281186 674258 281422 674494
rect 281186 667258 281422 667494
rect 281186 660258 281422 660494
rect 281186 653258 281422 653494
rect 281186 646258 281422 646494
rect 281186 639258 281422 639494
rect 281186 632258 281422 632494
rect 281186 625258 281422 625494
rect 281186 618258 281422 618494
rect 281186 611258 281422 611494
rect 281186 604258 281422 604494
rect 281186 597258 281422 597494
rect 281186 590258 281422 590494
rect 281186 583258 281422 583494
rect 281186 576258 281422 576494
rect 281186 569258 281422 569494
rect 281186 562258 281422 562494
rect 281186 555258 281422 555494
rect 281186 548258 281422 548494
rect 281186 541258 281422 541494
rect 281186 534258 281422 534494
rect 281186 527258 281422 527494
rect 281186 520258 281422 520494
rect 281186 513258 281422 513494
rect 281186 506258 281422 506494
rect 281186 499258 281422 499494
rect 281186 492258 281422 492494
rect 281186 485258 281422 485494
rect 281186 478258 281422 478494
rect 281186 471258 281422 471494
rect 281186 464258 281422 464494
rect 281186 457258 281422 457494
rect 281186 450258 281422 450494
rect 281186 443258 281422 443494
rect 281186 436258 281422 436494
rect 281186 429258 281422 429494
rect 281186 422258 281422 422494
rect 281186 415258 281422 415494
rect 281186 408258 281422 408494
rect 281186 401258 281422 401494
rect 281186 394258 281422 394494
rect 281186 387258 281422 387494
rect 281186 380258 281422 380494
rect 281186 373258 281422 373494
rect 281186 366258 281422 366494
rect 281186 359258 281422 359494
rect 281186 352258 281422 352494
rect 281186 345258 281422 345494
rect 281186 338258 281422 338494
rect 281186 331258 281422 331494
rect 281186 324258 281422 324494
rect 281186 317258 281422 317494
rect 281186 310258 281422 310494
rect 281186 303258 281422 303494
rect 281186 296258 281422 296494
rect 281186 289258 281422 289494
rect 281186 282258 281422 282494
rect 281186 275258 281422 275494
rect 281186 268258 281422 268494
rect 281186 261258 281422 261494
rect 281186 254258 281422 254494
rect 281186 247258 281422 247494
rect 281186 240258 281422 240494
rect 281186 233258 281422 233494
rect 281186 226258 281422 226494
rect 281186 219258 281422 219494
rect 281186 212258 281422 212494
rect 281186 205258 281422 205494
rect 281186 198258 281422 198494
rect 281186 191258 281422 191494
rect 281186 184258 281422 184494
rect 281186 177258 281422 177494
rect 281186 170258 281422 170494
rect 281186 163258 281422 163494
rect 281186 156258 281422 156494
rect 281186 149258 281422 149494
rect 281186 142258 281422 142494
rect 281186 135258 281422 135494
rect 281186 128258 281422 128494
rect 281186 121258 281422 121494
rect 281186 114258 281422 114494
rect 281186 107258 281422 107494
rect 281186 100258 281422 100494
rect 281186 93258 281422 93494
rect 281186 86258 281422 86494
rect 281186 79258 281422 79494
rect 281186 72258 281422 72494
rect 281186 65258 281422 65494
rect 281186 58258 281422 58494
rect 281186 51258 281422 51494
rect 281186 44258 281422 44494
rect 281186 37258 281422 37494
rect 281186 30258 281422 30494
rect 281186 23258 281422 23494
rect 281186 16258 281422 16494
rect 281186 9258 281422 9494
rect 281186 2258 281422 2494
rect 281186 -982 281422 -746
rect 281186 -1302 281422 -1066
rect 282918 705962 283154 706198
rect 282918 705642 283154 705878
rect 282918 696198 283154 696434
rect 282918 689198 283154 689434
rect 282918 682198 283154 682434
rect 282918 675198 283154 675434
rect 282918 668198 283154 668434
rect 282918 661198 283154 661434
rect 282918 654198 283154 654434
rect 282918 647198 283154 647434
rect 282918 640198 283154 640434
rect 282918 633198 283154 633434
rect 282918 626198 283154 626434
rect 282918 619198 283154 619434
rect 282918 612198 283154 612434
rect 282918 605198 283154 605434
rect 282918 598198 283154 598434
rect 282918 591198 283154 591434
rect 282918 584198 283154 584434
rect 282918 577198 283154 577434
rect 282918 570198 283154 570434
rect 282918 563198 283154 563434
rect 282918 556198 283154 556434
rect 282918 549198 283154 549434
rect 282918 542198 283154 542434
rect 282918 535198 283154 535434
rect 282918 528198 283154 528434
rect 282918 521198 283154 521434
rect 282918 514198 283154 514434
rect 282918 507198 283154 507434
rect 282918 500198 283154 500434
rect 282918 493198 283154 493434
rect 282918 486198 283154 486434
rect 282918 479198 283154 479434
rect 282918 472198 283154 472434
rect 282918 465198 283154 465434
rect 282918 458198 283154 458434
rect 282918 451198 283154 451434
rect 282918 444198 283154 444434
rect 282918 437198 283154 437434
rect 282918 430198 283154 430434
rect 282918 423198 283154 423434
rect 282918 416198 283154 416434
rect 282918 409198 283154 409434
rect 282918 402198 283154 402434
rect 282918 395198 283154 395434
rect 282918 388198 283154 388434
rect 282918 381198 283154 381434
rect 282918 374198 283154 374434
rect 282918 367198 283154 367434
rect 282918 360198 283154 360434
rect 282918 353198 283154 353434
rect 282918 346198 283154 346434
rect 282918 339198 283154 339434
rect 282918 332198 283154 332434
rect 282918 325198 283154 325434
rect 282918 318198 283154 318434
rect 282918 311198 283154 311434
rect 282918 304198 283154 304434
rect 282918 297198 283154 297434
rect 282918 290198 283154 290434
rect 282918 283198 283154 283434
rect 282918 276198 283154 276434
rect 282918 269198 283154 269434
rect 282918 262198 283154 262434
rect 282918 255198 283154 255434
rect 282918 248198 283154 248434
rect 282918 241198 283154 241434
rect 282918 234198 283154 234434
rect 282918 227198 283154 227434
rect 282918 220198 283154 220434
rect 282918 213198 283154 213434
rect 282918 206198 283154 206434
rect 282918 199198 283154 199434
rect 282918 192198 283154 192434
rect 282918 185198 283154 185434
rect 282918 178198 283154 178434
rect 282918 171198 283154 171434
rect 282918 164198 283154 164434
rect 282918 157198 283154 157434
rect 282918 150198 283154 150434
rect 282918 143198 283154 143434
rect 282918 136198 283154 136434
rect 282918 129198 283154 129434
rect 282918 122198 283154 122434
rect 282918 115198 283154 115434
rect 282918 108198 283154 108434
rect 282918 101198 283154 101434
rect 282918 94198 283154 94434
rect 282918 87198 283154 87434
rect 282918 80198 283154 80434
rect 282918 73198 283154 73434
rect 282918 66198 283154 66434
rect 282918 59198 283154 59434
rect 282918 52198 283154 52434
rect 282918 45198 283154 45434
rect 282918 38198 283154 38434
rect 282918 31198 283154 31434
rect 282918 24198 283154 24434
rect 282918 17198 283154 17434
rect 282918 10198 283154 10434
rect 282918 3198 283154 3434
rect 282918 -1942 283154 -1706
rect 282918 -2262 283154 -2026
rect 288186 705002 288422 705238
rect 288186 704682 288422 704918
rect 288186 695258 288422 695494
rect 288186 688258 288422 688494
rect 288186 681258 288422 681494
rect 288186 674258 288422 674494
rect 288186 667258 288422 667494
rect 288186 660258 288422 660494
rect 288186 653258 288422 653494
rect 288186 646258 288422 646494
rect 288186 639258 288422 639494
rect 288186 632258 288422 632494
rect 288186 625258 288422 625494
rect 288186 618258 288422 618494
rect 288186 611258 288422 611494
rect 288186 604258 288422 604494
rect 288186 597258 288422 597494
rect 288186 590258 288422 590494
rect 288186 583258 288422 583494
rect 288186 576258 288422 576494
rect 288186 569258 288422 569494
rect 288186 562258 288422 562494
rect 288186 555258 288422 555494
rect 288186 548258 288422 548494
rect 288186 541258 288422 541494
rect 288186 534258 288422 534494
rect 288186 527258 288422 527494
rect 288186 520258 288422 520494
rect 288186 513258 288422 513494
rect 288186 506258 288422 506494
rect 288186 499258 288422 499494
rect 288186 492258 288422 492494
rect 288186 485258 288422 485494
rect 288186 478258 288422 478494
rect 288186 471258 288422 471494
rect 288186 464258 288422 464494
rect 288186 457258 288422 457494
rect 288186 450258 288422 450494
rect 288186 443258 288422 443494
rect 288186 436258 288422 436494
rect 288186 429258 288422 429494
rect 288186 422258 288422 422494
rect 288186 415258 288422 415494
rect 288186 408258 288422 408494
rect 288186 401258 288422 401494
rect 288186 394258 288422 394494
rect 288186 387258 288422 387494
rect 288186 380258 288422 380494
rect 288186 373258 288422 373494
rect 288186 366258 288422 366494
rect 288186 359258 288422 359494
rect 288186 352258 288422 352494
rect 288186 345258 288422 345494
rect 288186 338258 288422 338494
rect 288186 331258 288422 331494
rect 288186 324258 288422 324494
rect 288186 317258 288422 317494
rect 288186 310258 288422 310494
rect 288186 303258 288422 303494
rect 288186 296258 288422 296494
rect 288186 289258 288422 289494
rect 288186 282258 288422 282494
rect 288186 275258 288422 275494
rect 288186 268258 288422 268494
rect 288186 261258 288422 261494
rect 288186 254258 288422 254494
rect 288186 247258 288422 247494
rect 288186 240258 288422 240494
rect 288186 233258 288422 233494
rect 288186 226258 288422 226494
rect 288186 219258 288422 219494
rect 288186 212258 288422 212494
rect 288186 205258 288422 205494
rect 288186 198258 288422 198494
rect 288186 191258 288422 191494
rect 288186 184258 288422 184494
rect 288186 177258 288422 177494
rect 288186 170258 288422 170494
rect 288186 163258 288422 163494
rect 288186 156258 288422 156494
rect 288186 149258 288422 149494
rect 288186 142258 288422 142494
rect 288186 135258 288422 135494
rect 288186 128258 288422 128494
rect 288186 121258 288422 121494
rect 288186 114258 288422 114494
rect 288186 107258 288422 107494
rect 288186 100258 288422 100494
rect 288186 93258 288422 93494
rect 288186 86258 288422 86494
rect 288186 79258 288422 79494
rect 288186 72258 288422 72494
rect 288186 65258 288422 65494
rect 288186 58258 288422 58494
rect 288186 51258 288422 51494
rect 288186 44258 288422 44494
rect 288186 37258 288422 37494
rect 288186 30258 288422 30494
rect 288186 23258 288422 23494
rect 288186 16258 288422 16494
rect 288186 9258 288422 9494
rect 288186 2258 288422 2494
rect 288186 -982 288422 -746
rect 288186 -1302 288422 -1066
rect 289918 705962 290154 706198
rect 289918 705642 290154 705878
rect 289918 696198 290154 696434
rect 289918 689198 290154 689434
rect 289918 682198 290154 682434
rect 289918 675198 290154 675434
rect 289918 668198 290154 668434
rect 289918 661198 290154 661434
rect 289918 654198 290154 654434
rect 289918 647198 290154 647434
rect 289918 640198 290154 640434
rect 289918 633198 290154 633434
rect 289918 626198 290154 626434
rect 289918 619198 290154 619434
rect 289918 612198 290154 612434
rect 289918 605198 290154 605434
rect 289918 598198 290154 598434
rect 289918 591198 290154 591434
rect 289918 584198 290154 584434
rect 289918 577198 290154 577434
rect 289918 570198 290154 570434
rect 289918 563198 290154 563434
rect 289918 556198 290154 556434
rect 289918 549198 290154 549434
rect 289918 542198 290154 542434
rect 289918 535198 290154 535434
rect 289918 528198 290154 528434
rect 289918 521198 290154 521434
rect 289918 514198 290154 514434
rect 289918 507198 290154 507434
rect 289918 500198 290154 500434
rect 289918 493198 290154 493434
rect 289918 486198 290154 486434
rect 289918 479198 290154 479434
rect 289918 472198 290154 472434
rect 289918 465198 290154 465434
rect 289918 458198 290154 458434
rect 289918 451198 290154 451434
rect 289918 444198 290154 444434
rect 289918 437198 290154 437434
rect 289918 430198 290154 430434
rect 289918 423198 290154 423434
rect 289918 416198 290154 416434
rect 289918 409198 290154 409434
rect 289918 402198 290154 402434
rect 289918 395198 290154 395434
rect 289918 388198 290154 388434
rect 289918 381198 290154 381434
rect 289918 374198 290154 374434
rect 295186 705002 295422 705238
rect 295186 704682 295422 704918
rect 295186 695258 295422 695494
rect 295186 688258 295422 688494
rect 295186 681258 295422 681494
rect 295186 674258 295422 674494
rect 295186 667258 295422 667494
rect 295186 660258 295422 660494
rect 295186 653258 295422 653494
rect 295186 646258 295422 646494
rect 295186 639258 295422 639494
rect 295186 632258 295422 632494
rect 295186 625258 295422 625494
rect 295186 618258 295422 618494
rect 295186 611258 295422 611494
rect 295186 604258 295422 604494
rect 295186 597258 295422 597494
rect 295186 590258 295422 590494
rect 295186 583258 295422 583494
rect 295186 576258 295422 576494
rect 295186 569258 295422 569494
rect 295186 562258 295422 562494
rect 295186 555258 295422 555494
rect 295186 548258 295422 548494
rect 295186 541258 295422 541494
rect 295186 534258 295422 534494
rect 295186 527258 295422 527494
rect 295186 520258 295422 520494
rect 295186 513258 295422 513494
rect 295186 506258 295422 506494
rect 295186 499258 295422 499494
rect 295186 492258 295422 492494
rect 295186 485258 295422 485494
rect 295186 478258 295422 478494
rect 295186 471258 295422 471494
rect 295186 464258 295422 464494
rect 295186 457258 295422 457494
rect 295186 450258 295422 450494
rect 295186 443258 295422 443494
rect 295186 436258 295422 436494
rect 295186 429258 295422 429494
rect 295186 422258 295422 422494
rect 295186 415258 295422 415494
rect 295186 408258 295422 408494
rect 295186 401258 295422 401494
rect 295186 394258 295422 394494
rect 295186 387258 295422 387494
rect 295186 380258 295422 380494
rect 295186 373258 295422 373494
rect 296918 705962 297154 706198
rect 296918 705642 297154 705878
rect 296918 696198 297154 696434
rect 296918 689198 297154 689434
rect 296918 682198 297154 682434
rect 296918 675198 297154 675434
rect 296918 668198 297154 668434
rect 296918 661198 297154 661434
rect 296918 654198 297154 654434
rect 296918 647198 297154 647434
rect 296918 640198 297154 640434
rect 296918 633198 297154 633434
rect 296918 626198 297154 626434
rect 296918 619198 297154 619434
rect 296918 612198 297154 612434
rect 296918 605198 297154 605434
rect 296918 598198 297154 598434
rect 296918 591198 297154 591434
rect 296918 584198 297154 584434
rect 296918 577198 297154 577434
rect 296918 570198 297154 570434
rect 296918 563198 297154 563434
rect 296918 556198 297154 556434
rect 296918 549198 297154 549434
rect 296918 542198 297154 542434
rect 296918 535198 297154 535434
rect 296918 528198 297154 528434
rect 296918 521198 297154 521434
rect 296918 514198 297154 514434
rect 296918 507198 297154 507434
rect 296918 500198 297154 500434
rect 296918 493198 297154 493434
rect 296918 486198 297154 486434
rect 296918 479198 297154 479434
rect 296918 472198 297154 472434
rect 296918 465198 297154 465434
rect 296918 458198 297154 458434
rect 296918 451198 297154 451434
rect 296918 444198 297154 444434
rect 296918 437198 297154 437434
rect 296918 430198 297154 430434
rect 296918 423198 297154 423434
rect 296918 416198 297154 416434
rect 296918 409198 297154 409434
rect 296918 402198 297154 402434
rect 296918 395198 297154 395434
rect 296918 388198 297154 388434
rect 296918 381198 297154 381434
rect 296918 374198 297154 374434
rect 302186 705002 302422 705238
rect 302186 704682 302422 704918
rect 302186 695258 302422 695494
rect 302186 688258 302422 688494
rect 302186 681258 302422 681494
rect 302186 674258 302422 674494
rect 302186 667258 302422 667494
rect 302186 660258 302422 660494
rect 302186 653258 302422 653494
rect 302186 646258 302422 646494
rect 302186 639258 302422 639494
rect 302186 632258 302422 632494
rect 302186 625258 302422 625494
rect 302186 618258 302422 618494
rect 302186 611258 302422 611494
rect 302186 604258 302422 604494
rect 302186 597258 302422 597494
rect 302186 590258 302422 590494
rect 302186 583258 302422 583494
rect 302186 576258 302422 576494
rect 302186 569258 302422 569494
rect 302186 562258 302422 562494
rect 302186 555258 302422 555494
rect 302186 548258 302422 548494
rect 302186 541258 302422 541494
rect 302186 534258 302422 534494
rect 302186 527258 302422 527494
rect 302186 520258 302422 520494
rect 302186 513258 302422 513494
rect 302186 506258 302422 506494
rect 302186 499258 302422 499494
rect 302186 492258 302422 492494
rect 302186 485258 302422 485494
rect 302186 478258 302422 478494
rect 302186 471258 302422 471494
rect 302186 464258 302422 464494
rect 302186 457258 302422 457494
rect 302186 450258 302422 450494
rect 302186 443258 302422 443494
rect 302186 436258 302422 436494
rect 302186 429258 302422 429494
rect 302186 422258 302422 422494
rect 302186 415258 302422 415494
rect 302186 408258 302422 408494
rect 302186 401258 302422 401494
rect 302186 394258 302422 394494
rect 302186 387258 302422 387494
rect 302186 380258 302422 380494
rect 302186 373258 302422 373494
rect 303918 705962 304154 706198
rect 303918 705642 304154 705878
rect 303918 696198 304154 696434
rect 303918 689198 304154 689434
rect 303918 682198 304154 682434
rect 303918 675198 304154 675434
rect 303918 668198 304154 668434
rect 303918 661198 304154 661434
rect 303918 654198 304154 654434
rect 303918 647198 304154 647434
rect 303918 640198 304154 640434
rect 303918 633198 304154 633434
rect 303918 626198 304154 626434
rect 303918 619198 304154 619434
rect 303918 612198 304154 612434
rect 303918 605198 304154 605434
rect 303918 598198 304154 598434
rect 303918 591198 304154 591434
rect 303918 584198 304154 584434
rect 303918 577198 304154 577434
rect 303918 570198 304154 570434
rect 303918 563198 304154 563434
rect 303918 556198 304154 556434
rect 303918 549198 304154 549434
rect 303918 542198 304154 542434
rect 303918 535198 304154 535434
rect 303918 528198 304154 528434
rect 303918 521198 304154 521434
rect 303918 514198 304154 514434
rect 303918 507198 304154 507434
rect 303918 500198 304154 500434
rect 303918 493198 304154 493434
rect 303918 486198 304154 486434
rect 303918 479198 304154 479434
rect 303918 472198 304154 472434
rect 303918 465198 304154 465434
rect 303918 458198 304154 458434
rect 303918 451198 304154 451434
rect 303918 444198 304154 444434
rect 303918 437198 304154 437434
rect 303918 430198 304154 430434
rect 303918 423198 304154 423434
rect 303918 416198 304154 416434
rect 303918 409198 304154 409434
rect 303918 402198 304154 402434
rect 303918 395198 304154 395434
rect 303918 388198 304154 388434
rect 303918 381198 304154 381434
rect 303918 374198 304154 374434
rect 309186 705002 309422 705238
rect 309186 704682 309422 704918
rect 309186 695258 309422 695494
rect 309186 688258 309422 688494
rect 309186 681258 309422 681494
rect 309186 674258 309422 674494
rect 309186 667258 309422 667494
rect 309186 660258 309422 660494
rect 309186 653258 309422 653494
rect 309186 646258 309422 646494
rect 309186 639258 309422 639494
rect 309186 632258 309422 632494
rect 309186 625258 309422 625494
rect 309186 618258 309422 618494
rect 309186 611258 309422 611494
rect 309186 604258 309422 604494
rect 309186 597258 309422 597494
rect 309186 590258 309422 590494
rect 309186 583258 309422 583494
rect 309186 576258 309422 576494
rect 309186 569258 309422 569494
rect 309186 562258 309422 562494
rect 309186 555258 309422 555494
rect 309186 548258 309422 548494
rect 309186 541258 309422 541494
rect 309186 534258 309422 534494
rect 309186 527258 309422 527494
rect 309186 520258 309422 520494
rect 309186 513258 309422 513494
rect 309186 506258 309422 506494
rect 309186 499258 309422 499494
rect 309186 492258 309422 492494
rect 309186 485258 309422 485494
rect 309186 478258 309422 478494
rect 309186 471258 309422 471494
rect 309186 464258 309422 464494
rect 309186 457258 309422 457494
rect 309186 450258 309422 450494
rect 309186 443258 309422 443494
rect 309186 436258 309422 436494
rect 309186 429258 309422 429494
rect 309186 422258 309422 422494
rect 309186 415258 309422 415494
rect 309186 408258 309422 408494
rect 309186 401258 309422 401494
rect 309186 394258 309422 394494
rect 309186 387258 309422 387494
rect 309186 380258 309422 380494
rect 309186 373258 309422 373494
rect 289918 367198 290154 367434
rect 309186 366258 309422 366494
rect 289918 360198 290154 360434
rect 289918 353198 290154 353434
rect 289918 346198 290154 346434
rect 289918 339198 290154 339434
rect 289918 332198 290154 332434
rect 289918 325198 290154 325434
rect 289918 318198 290154 318434
rect 289918 311198 290154 311434
rect 289918 304198 290154 304434
rect 289918 297198 290154 297434
rect 289918 290198 290154 290434
rect 289918 283198 290154 283434
rect 289918 276198 290154 276434
rect 289918 269198 290154 269434
rect 289918 262198 290154 262434
rect 289918 255198 290154 255434
rect 289918 248198 290154 248434
rect 289918 241198 290154 241434
rect 289918 234198 290154 234434
rect 289918 227198 290154 227434
rect 289918 220198 290154 220434
rect 289918 213198 290154 213434
rect 289918 206198 290154 206434
rect 295186 359258 295422 359494
rect 295186 352258 295422 352494
rect 295186 345258 295422 345494
rect 295186 338258 295422 338494
rect 295186 331258 295422 331494
rect 295186 324258 295422 324494
rect 295186 317258 295422 317494
rect 295186 310258 295422 310494
rect 295186 303258 295422 303494
rect 295186 296258 295422 296494
rect 295186 289258 295422 289494
rect 295186 282258 295422 282494
rect 295186 275258 295422 275494
rect 295186 268258 295422 268494
rect 295186 261258 295422 261494
rect 295186 254258 295422 254494
rect 295186 247258 295422 247494
rect 295186 240258 295422 240494
rect 295186 233258 295422 233494
rect 295186 226258 295422 226494
rect 295186 219258 295422 219494
rect 295186 212258 295422 212494
rect 295186 205258 295422 205494
rect 296918 360198 297154 360434
rect 296918 353198 297154 353434
rect 296918 346198 297154 346434
rect 296918 339198 297154 339434
rect 296918 332198 297154 332434
rect 296918 325198 297154 325434
rect 296918 318198 297154 318434
rect 296918 311198 297154 311434
rect 296918 304198 297154 304434
rect 296918 297198 297154 297434
rect 296918 290198 297154 290434
rect 296918 283198 297154 283434
rect 296918 276198 297154 276434
rect 296918 269198 297154 269434
rect 296918 262198 297154 262434
rect 296918 255198 297154 255434
rect 296918 248198 297154 248434
rect 296918 241198 297154 241434
rect 296918 234198 297154 234434
rect 296918 227198 297154 227434
rect 296918 220198 297154 220434
rect 296918 213198 297154 213434
rect 296918 206198 297154 206434
rect 302186 359258 302422 359494
rect 302186 352258 302422 352494
rect 302186 345258 302422 345494
rect 302186 338258 302422 338494
rect 302186 331258 302422 331494
rect 302186 324258 302422 324494
rect 302186 317258 302422 317494
rect 302186 310258 302422 310494
rect 302186 303258 302422 303494
rect 302186 296258 302422 296494
rect 302186 289258 302422 289494
rect 302186 282258 302422 282494
rect 302186 275258 302422 275494
rect 302186 268258 302422 268494
rect 302186 261258 302422 261494
rect 302186 254258 302422 254494
rect 302186 247258 302422 247494
rect 302186 240258 302422 240494
rect 302186 233258 302422 233494
rect 302186 226258 302422 226494
rect 302186 219258 302422 219494
rect 302186 212258 302422 212494
rect 302186 205258 302422 205494
rect 303918 360198 304154 360434
rect 303918 353198 304154 353434
rect 303918 346198 304154 346434
rect 303918 339198 304154 339434
rect 303918 332198 304154 332434
rect 303918 325198 304154 325434
rect 303918 318198 304154 318434
rect 303918 311198 304154 311434
rect 303918 304198 304154 304434
rect 303918 297198 304154 297434
rect 303918 290198 304154 290434
rect 303918 283198 304154 283434
rect 303918 276198 304154 276434
rect 303918 269198 304154 269434
rect 303918 262198 304154 262434
rect 303918 255198 304154 255434
rect 303918 248198 304154 248434
rect 303918 241198 304154 241434
rect 303918 234198 304154 234434
rect 303918 227198 304154 227434
rect 303918 220198 304154 220434
rect 303918 213198 304154 213434
rect 303918 206198 304154 206434
rect 309186 359258 309422 359494
rect 309186 352258 309422 352494
rect 309186 345258 309422 345494
rect 309186 338258 309422 338494
rect 309186 331258 309422 331494
rect 309186 324258 309422 324494
rect 309186 317258 309422 317494
rect 309186 310258 309422 310494
rect 309186 303258 309422 303494
rect 309186 296258 309422 296494
rect 309186 289258 309422 289494
rect 309186 282258 309422 282494
rect 309186 275258 309422 275494
rect 309186 268258 309422 268494
rect 309186 261258 309422 261494
rect 309186 254258 309422 254494
rect 309186 247258 309422 247494
rect 309186 240258 309422 240494
rect 309186 233258 309422 233494
rect 309186 226258 309422 226494
rect 309186 219258 309422 219494
rect 309186 212258 309422 212494
rect 309186 205258 309422 205494
rect 289918 199198 290154 199434
rect 309186 198258 309422 198494
rect 289918 192198 290154 192434
rect 289918 185198 290154 185434
rect 289918 178198 290154 178434
rect 289918 171198 290154 171434
rect 289918 164198 290154 164434
rect 289918 157198 290154 157434
rect 289918 150198 290154 150434
rect 289918 143198 290154 143434
rect 289918 136198 290154 136434
rect 289918 129198 290154 129434
rect 289918 122198 290154 122434
rect 289918 115198 290154 115434
rect 289918 108198 290154 108434
rect 289918 101198 290154 101434
rect 289918 94198 290154 94434
rect 289918 87198 290154 87434
rect 289918 80198 290154 80434
rect 289918 73198 290154 73434
rect 289918 66198 290154 66434
rect 289918 59198 290154 59434
rect 289918 52198 290154 52434
rect 289918 45198 290154 45434
rect 289918 38198 290154 38434
rect 289918 31198 290154 31434
rect 289918 24198 290154 24434
rect 289918 17198 290154 17434
rect 289918 10198 290154 10434
rect 289918 3198 290154 3434
rect 289918 -1942 290154 -1706
rect 289918 -2262 290154 -2026
rect 295186 191258 295422 191494
rect 295186 184258 295422 184494
rect 295186 177258 295422 177494
rect 295186 170258 295422 170494
rect 295186 163258 295422 163494
rect 295186 156258 295422 156494
rect 295186 149258 295422 149494
rect 295186 142258 295422 142494
rect 295186 135258 295422 135494
rect 295186 128258 295422 128494
rect 295186 121258 295422 121494
rect 295186 114258 295422 114494
rect 295186 107258 295422 107494
rect 295186 100258 295422 100494
rect 295186 93258 295422 93494
rect 295186 86258 295422 86494
rect 295186 79258 295422 79494
rect 295186 72258 295422 72494
rect 295186 65258 295422 65494
rect 295186 58258 295422 58494
rect 295186 51258 295422 51494
rect 295186 44258 295422 44494
rect 295186 37258 295422 37494
rect 295186 30258 295422 30494
rect 295186 23258 295422 23494
rect 295186 16258 295422 16494
rect 295186 9258 295422 9494
rect 295186 2258 295422 2494
rect 295186 -982 295422 -746
rect 295186 -1302 295422 -1066
rect 296918 192198 297154 192434
rect 296918 185198 297154 185434
rect 296918 178198 297154 178434
rect 296918 171198 297154 171434
rect 296918 164198 297154 164434
rect 296918 157198 297154 157434
rect 296918 150198 297154 150434
rect 296918 143198 297154 143434
rect 296918 136198 297154 136434
rect 296918 129198 297154 129434
rect 296918 122198 297154 122434
rect 296918 115198 297154 115434
rect 296918 108198 297154 108434
rect 296918 101198 297154 101434
rect 296918 94198 297154 94434
rect 296918 87198 297154 87434
rect 296918 80198 297154 80434
rect 296918 73198 297154 73434
rect 296918 66198 297154 66434
rect 296918 59198 297154 59434
rect 296918 52198 297154 52434
rect 296918 45198 297154 45434
rect 296918 38198 297154 38434
rect 296918 31198 297154 31434
rect 296918 24198 297154 24434
rect 296918 17198 297154 17434
rect 296918 10198 297154 10434
rect 296918 3198 297154 3434
rect 296918 -1942 297154 -1706
rect 296918 -2262 297154 -2026
rect 302186 191258 302422 191494
rect 302186 184258 302422 184494
rect 302186 177258 302422 177494
rect 302186 170258 302422 170494
rect 302186 163258 302422 163494
rect 302186 156258 302422 156494
rect 302186 149258 302422 149494
rect 302186 142258 302422 142494
rect 302186 135258 302422 135494
rect 302186 128258 302422 128494
rect 302186 121258 302422 121494
rect 302186 114258 302422 114494
rect 302186 107258 302422 107494
rect 302186 100258 302422 100494
rect 302186 93258 302422 93494
rect 302186 86258 302422 86494
rect 302186 79258 302422 79494
rect 302186 72258 302422 72494
rect 302186 65258 302422 65494
rect 302186 58258 302422 58494
rect 302186 51258 302422 51494
rect 302186 44258 302422 44494
rect 302186 37258 302422 37494
rect 302186 30258 302422 30494
rect 302186 23258 302422 23494
rect 302186 16258 302422 16494
rect 302186 9258 302422 9494
rect 302186 2258 302422 2494
rect 302186 -982 302422 -746
rect 302186 -1302 302422 -1066
rect 303918 192198 304154 192434
rect 303918 185198 304154 185434
rect 303918 178198 304154 178434
rect 303918 171198 304154 171434
rect 303918 164198 304154 164434
rect 303918 157198 304154 157434
rect 303918 150198 304154 150434
rect 303918 143198 304154 143434
rect 303918 136198 304154 136434
rect 303918 129198 304154 129434
rect 303918 122198 304154 122434
rect 303918 115198 304154 115434
rect 303918 108198 304154 108434
rect 303918 101198 304154 101434
rect 303918 94198 304154 94434
rect 303918 87198 304154 87434
rect 303918 80198 304154 80434
rect 303918 73198 304154 73434
rect 303918 66198 304154 66434
rect 303918 59198 304154 59434
rect 303918 52198 304154 52434
rect 303918 45198 304154 45434
rect 303918 38198 304154 38434
rect 303918 31198 304154 31434
rect 303918 24198 304154 24434
rect 303918 17198 304154 17434
rect 303918 10198 304154 10434
rect 303918 3198 304154 3434
rect 303918 -1942 304154 -1706
rect 303918 -2262 304154 -2026
rect 309186 191258 309422 191494
rect 309186 184258 309422 184494
rect 309186 177258 309422 177494
rect 309186 170258 309422 170494
rect 309186 163258 309422 163494
rect 309186 156258 309422 156494
rect 309186 149258 309422 149494
rect 309186 142258 309422 142494
rect 309186 135258 309422 135494
rect 309186 128258 309422 128494
rect 309186 121258 309422 121494
rect 309186 114258 309422 114494
rect 309186 107258 309422 107494
rect 309186 100258 309422 100494
rect 309186 93258 309422 93494
rect 309186 86258 309422 86494
rect 309186 79258 309422 79494
rect 309186 72258 309422 72494
rect 309186 65258 309422 65494
rect 309186 58258 309422 58494
rect 309186 51258 309422 51494
rect 309186 44258 309422 44494
rect 309186 37258 309422 37494
rect 309186 30258 309422 30494
rect 309186 23258 309422 23494
rect 309186 16258 309422 16494
rect 309186 9258 309422 9494
rect 309186 2258 309422 2494
rect 309186 -982 309422 -746
rect 309186 -1302 309422 -1066
rect 310918 705962 311154 706198
rect 310918 705642 311154 705878
rect 310918 696198 311154 696434
rect 310918 689198 311154 689434
rect 310918 682198 311154 682434
rect 310918 675198 311154 675434
rect 310918 668198 311154 668434
rect 310918 661198 311154 661434
rect 310918 654198 311154 654434
rect 310918 647198 311154 647434
rect 310918 640198 311154 640434
rect 310918 633198 311154 633434
rect 310918 626198 311154 626434
rect 310918 619198 311154 619434
rect 310918 612198 311154 612434
rect 310918 605198 311154 605434
rect 310918 598198 311154 598434
rect 310918 591198 311154 591434
rect 310918 584198 311154 584434
rect 310918 577198 311154 577434
rect 310918 570198 311154 570434
rect 310918 563198 311154 563434
rect 310918 556198 311154 556434
rect 310918 549198 311154 549434
rect 310918 542198 311154 542434
rect 310918 535198 311154 535434
rect 310918 528198 311154 528434
rect 310918 521198 311154 521434
rect 310918 514198 311154 514434
rect 310918 507198 311154 507434
rect 310918 500198 311154 500434
rect 310918 493198 311154 493434
rect 310918 486198 311154 486434
rect 310918 479198 311154 479434
rect 310918 472198 311154 472434
rect 310918 465198 311154 465434
rect 310918 458198 311154 458434
rect 310918 451198 311154 451434
rect 310918 444198 311154 444434
rect 310918 437198 311154 437434
rect 310918 430198 311154 430434
rect 310918 423198 311154 423434
rect 310918 416198 311154 416434
rect 310918 409198 311154 409434
rect 310918 402198 311154 402434
rect 310918 395198 311154 395434
rect 310918 388198 311154 388434
rect 310918 381198 311154 381434
rect 310918 374198 311154 374434
rect 310918 367198 311154 367434
rect 310918 360198 311154 360434
rect 310918 353198 311154 353434
rect 310918 346198 311154 346434
rect 310918 339198 311154 339434
rect 310918 332198 311154 332434
rect 310918 325198 311154 325434
rect 310918 318198 311154 318434
rect 310918 311198 311154 311434
rect 310918 304198 311154 304434
rect 310918 297198 311154 297434
rect 310918 290198 311154 290434
rect 310918 283198 311154 283434
rect 310918 276198 311154 276434
rect 310918 269198 311154 269434
rect 310918 262198 311154 262434
rect 310918 255198 311154 255434
rect 310918 248198 311154 248434
rect 310918 241198 311154 241434
rect 310918 234198 311154 234434
rect 310918 227198 311154 227434
rect 310918 220198 311154 220434
rect 310918 213198 311154 213434
rect 310918 206198 311154 206434
rect 310918 199198 311154 199434
rect 310918 192198 311154 192434
rect 310918 185198 311154 185434
rect 310918 178198 311154 178434
rect 310918 171198 311154 171434
rect 310918 164198 311154 164434
rect 310918 157198 311154 157434
rect 310918 150198 311154 150434
rect 310918 143198 311154 143434
rect 310918 136198 311154 136434
rect 310918 129198 311154 129434
rect 310918 122198 311154 122434
rect 310918 115198 311154 115434
rect 310918 108198 311154 108434
rect 310918 101198 311154 101434
rect 310918 94198 311154 94434
rect 310918 87198 311154 87434
rect 310918 80198 311154 80434
rect 310918 73198 311154 73434
rect 310918 66198 311154 66434
rect 310918 59198 311154 59434
rect 310918 52198 311154 52434
rect 310918 45198 311154 45434
rect 310918 38198 311154 38434
rect 310918 31198 311154 31434
rect 310918 24198 311154 24434
rect 310918 17198 311154 17434
rect 310918 10198 311154 10434
rect 310918 3198 311154 3434
rect 310918 -1942 311154 -1706
rect 310918 -2262 311154 -2026
rect 316186 705002 316422 705238
rect 316186 704682 316422 704918
rect 316186 695258 316422 695494
rect 316186 688258 316422 688494
rect 316186 681258 316422 681494
rect 316186 674258 316422 674494
rect 316186 667258 316422 667494
rect 316186 660258 316422 660494
rect 316186 653258 316422 653494
rect 316186 646258 316422 646494
rect 316186 639258 316422 639494
rect 316186 632258 316422 632494
rect 316186 625258 316422 625494
rect 316186 618258 316422 618494
rect 316186 611258 316422 611494
rect 316186 604258 316422 604494
rect 316186 597258 316422 597494
rect 316186 590258 316422 590494
rect 316186 583258 316422 583494
rect 316186 576258 316422 576494
rect 316186 569258 316422 569494
rect 316186 562258 316422 562494
rect 316186 555258 316422 555494
rect 316186 548258 316422 548494
rect 316186 541258 316422 541494
rect 316186 534258 316422 534494
rect 316186 527258 316422 527494
rect 316186 520258 316422 520494
rect 316186 513258 316422 513494
rect 316186 506258 316422 506494
rect 316186 499258 316422 499494
rect 316186 492258 316422 492494
rect 316186 485258 316422 485494
rect 316186 478258 316422 478494
rect 316186 471258 316422 471494
rect 316186 464258 316422 464494
rect 316186 457258 316422 457494
rect 316186 450258 316422 450494
rect 316186 443258 316422 443494
rect 316186 436258 316422 436494
rect 316186 429258 316422 429494
rect 316186 422258 316422 422494
rect 316186 415258 316422 415494
rect 316186 408258 316422 408494
rect 316186 401258 316422 401494
rect 316186 394258 316422 394494
rect 316186 387258 316422 387494
rect 316186 380258 316422 380494
rect 316186 373258 316422 373494
rect 316186 366258 316422 366494
rect 316186 359258 316422 359494
rect 316186 352258 316422 352494
rect 316186 345258 316422 345494
rect 316186 338258 316422 338494
rect 316186 331258 316422 331494
rect 316186 324258 316422 324494
rect 316186 317258 316422 317494
rect 316186 310258 316422 310494
rect 316186 303258 316422 303494
rect 316186 296258 316422 296494
rect 316186 289258 316422 289494
rect 316186 282258 316422 282494
rect 316186 275258 316422 275494
rect 316186 268258 316422 268494
rect 316186 261258 316422 261494
rect 316186 254258 316422 254494
rect 316186 247258 316422 247494
rect 316186 240258 316422 240494
rect 316186 233258 316422 233494
rect 316186 226258 316422 226494
rect 316186 219258 316422 219494
rect 316186 212258 316422 212494
rect 316186 205258 316422 205494
rect 316186 198258 316422 198494
rect 316186 191258 316422 191494
rect 316186 184258 316422 184494
rect 316186 177258 316422 177494
rect 316186 170258 316422 170494
rect 316186 163258 316422 163494
rect 316186 156258 316422 156494
rect 316186 149258 316422 149494
rect 316186 142258 316422 142494
rect 316186 135258 316422 135494
rect 316186 128258 316422 128494
rect 316186 121258 316422 121494
rect 316186 114258 316422 114494
rect 316186 107258 316422 107494
rect 316186 100258 316422 100494
rect 316186 93258 316422 93494
rect 316186 86258 316422 86494
rect 316186 79258 316422 79494
rect 316186 72258 316422 72494
rect 316186 65258 316422 65494
rect 316186 58258 316422 58494
rect 316186 51258 316422 51494
rect 316186 44258 316422 44494
rect 316186 37258 316422 37494
rect 316186 30258 316422 30494
rect 316186 23258 316422 23494
rect 316186 16258 316422 16494
rect 316186 9258 316422 9494
rect 316186 2258 316422 2494
rect 316186 -982 316422 -746
rect 316186 -1302 316422 -1066
rect 317918 705962 318154 706198
rect 317918 705642 318154 705878
rect 317918 696198 318154 696434
rect 317918 689198 318154 689434
rect 317918 682198 318154 682434
rect 317918 675198 318154 675434
rect 317918 668198 318154 668434
rect 317918 661198 318154 661434
rect 317918 654198 318154 654434
rect 317918 647198 318154 647434
rect 317918 640198 318154 640434
rect 317918 633198 318154 633434
rect 317918 626198 318154 626434
rect 317918 619198 318154 619434
rect 317918 612198 318154 612434
rect 317918 605198 318154 605434
rect 317918 598198 318154 598434
rect 317918 591198 318154 591434
rect 317918 584198 318154 584434
rect 317918 577198 318154 577434
rect 317918 570198 318154 570434
rect 317918 563198 318154 563434
rect 317918 556198 318154 556434
rect 317918 549198 318154 549434
rect 317918 542198 318154 542434
rect 317918 535198 318154 535434
rect 317918 528198 318154 528434
rect 317918 521198 318154 521434
rect 317918 514198 318154 514434
rect 317918 507198 318154 507434
rect 317918 500198 318154 500434
rect 317918 493198 318154 493434
rect 317918 486198 318154 486434
rect 317918 479198 318154 479434
rect 317918 472198 318154 472434
rect 317918 465198 318154 465434
rect 317918 458198 318154 458434
rect 317918 451198 318154 451434
rect 317918 444198 318154 444434
rect 317918 437198 318154 437434
rect 317918 430198 318154 430434
rect 317918 423198 318154 423434
rect 317918 416198 318154 416434
rect 317918 409198 318154 409434
rect 317918 402198 318154 402434
rect 317918 395198 318154 395434
rect 317918 388198 318154 388434
rect 317918 381198 318154 381434
rect 317918 374198 318154 374434
rect 317918 367198 318154 367434
rect 317918 360198 318154 360434
rect 317918 353198 318154 353434
rect 317918 346198 318154 346434
rect 317918 339198 318154 339434
rect 317918 332198 318154 332434
rect 317918 325198 318154 325434
rect 317918 318198 318154 318434
rect 317918 311198 318154 311434
rect 317918 304198 318154 304434
rect 317918 297198 318154 297434
rect 317918 290198 318154 290434
rect 317918 283198 318154 283434
rect 317918 276198 318154 276434
rect 317918 269198 318154 269434
rect 317918 262198 318154 262434
rect 317918 255198 318154 255434
rect 317918 248198 318154 248434
rect 317918 241198 318154 241434
rect 317918 234198 318154 234434
rect 317918 227198 318154 227434
rect 317918 220198 318154 220434
rect 317918 213198 318154 213434
rect 317918 206198 318154 206434
rect 317918 199198 318154 199434
rect 317918 192198 318154 192434
rect 317918 185198 318154 185434
rect 317918 178198 318154 178434
rect 317918 171198 318154 171434
rect 317918 164198 318154 164434
rect 317918 157198 318154 157434
rect 317918 150198 318154 150434
rect 317918 143198 318154 143434
rect 317918 136198 318154 136434
rect 317918 129198 318154 129434
rect 317918 122198 318154 122434
rect 317918 115198 318154 115434
rect 317918 108198 318154 108434
rect 317918 101198 318154 101434
rect 317918 94198 318154 94434
rect 317918 87198 318154 87434
rect 317918 80198 318154 80434
rect 317918 73198 318154 73434
rect 317918 66198 318154 66434
rect 317918 59198 318154 59434
rect 317918 52198 318154 52434
rect 317918 45198 318154 45434
rect 317918 38198 318154 38434
rect 317918 31198 318154 31434
rect 317918 24198 318154 24434
rect 317918 17198 318154 17434
rect 317918 10198 318154 10434
rect 317918 3198 318154 3434
rect 317918 -1942 318154 -1706
rect 317918 -2262 318154 -2026
rect 323186 705002 323422 705238
rect 323186 704682 323422 704918
rect 323186 695258 323422 695494
rect 323186 688258 323422 688494
rect 323186 681258 323422 681494
rect 323186 674258 323422 674494
rect 323186 667258 323422 667494
rect 323186 660258 323422 660494
rect 323186 653258 323422 653494
rect 323186 646258 323422 646494
rect 323186 639258 323422 639494
rect 323186 632258 323422 632494
rect 323186 625258 323422 625494
rect 323186 618258 323422 618494
rect 323186 611258 323422 611494
rect 323186 604258 323422 604494
rect 323186 597258 323422 597494
rect 323186 590258 323422 590494
rect 323186 583258 323422 583494
rect 323186 576258 323422 576494
rect 323186 569258 323422 569494
rect 323186 562258 323422 562494
rect 323186 555258 323422 555494
rect 323186 548258 323422 548494
rect 323186 541258 323422 541494
rect 323186 534258 323422 534494
rect 323186 527258 323422 527494
rect 323186 520258 323422 520494
rect 323186 513258 323422 513494
rect 323186 506258 323422 506494
rect 323186 499258 323422 499494
rect 323186 492258 323422 492494
rect 323186 485258 323422 485494
rect 323186 478258 323422 478494
rect 323186 471258 323422 471494
rect 323186 464258 323422 464494
rect 323186 457258 323422 457494
rect 323186 450258 323422 450494
rect 323186 443258 323422 443494
rect 323186 436258 323422 436494
rect 323186 429258 323422 429494
rect 323186 422258 323422 422494
rect 323186 415258 323422 415494
rect 323186 408258 323422 408494
rect 323186 401258 323422 401494
rect 323186 394258 323422 394494
rect 323186 387258 323422 387494
rect 323186 380258 323422 380494
rect 323186 373258 323422 373494
rect 323186 366258 323422 366494
rect 323186 359258 323422 359494
rect 323186 352258 323422 352494
rect 323186 345258 323422 345494
rect 323186 338258 323422 338494
rect 323186 331258 323422 331494
rect 323186 324258 323422 324494
rect 323186 317258 323422 317494
rect 323186 310258 323422 310494
rect 323186 303258 323422 303494
rect 323186 296258 323422 296494
rect 323186 289258 323422 289494
rect 323186 282258 323422 282494
rect 323186 275258 323422 275494
rect 323186 268258 323422 268494
rect 323186 261258 323422 261494
rect 323186 254258 323422 254494
rect 323186 247258 323422 247494
rect 323186 240258 323422 240494
rect 323186 233258 323422 233494
rect 323186 226258 323422 226494
rect 323186 219258 323422 219494
rect 323186 212258 323422 212494
rect 323186 205258 323422 205494
rect 323186 198258 323422 198494
rect 323186 191258 323422 191494
rect 323186 184258 323422 184494
rect 323186 177258 323422 177494
rect 323186 170258 323422 170494
rect 323186 163258 323422 163494
rect 323186 156258 323422 156494
rect 323186 149258 323422 149494
rect 323186 142258 323422 142494
rect 323186 135258 323422 135494
rect 323186 128258 323422 128494
rect 323186 121258 323422 121494
rect 323186 114258 323422 114494
rect 323186 107258 323422 107494
rect 323186 100258 323422 100494
rect 323186 93258 323422 93494
rect 323186 86258 323422 86494
rect 323186 79258 323422 79494
rect 323186 72258 323422 72494
rect 323186 65258 323422 65494
rect 323186 58258 323422 58494
rect 323186 51258 323422 51494
rect 323186 44258 323422 44494
rect 323186 37258 323422 37494
rect 323186 30258 323422 30494
rect 323186 23258 323422 23494
rect 323186 16258 323422 16494
rect 323186 9258 323422 9494
rect 323186 2258 323422 2494
rect 323186 -982 323422 -746
rect 323186 -1302 323422 -1066
rect 324918 705962 325154 706198
rect 324918 705642 325154 705878
rect 324918 696198 325154 696434
rect 324918 689198 325154 689434
rect 324918 682198 325154 682434
rect 324918 675198 325154 675434
rect 324918 668198 325154 668434
rect 324918 661198 325154 661434
rect 324918 654198 325154 654434
rect 324918 647198 325154 647434
rect 324918 640198 325154 640434
rect 324918 633198 325154 633434
rect 324918 626198 325154 626434
rect 324918 619198 325154 619434
rect 324918 612198 325154 612434
rect 324918 605198 325154 605434
rect 324918 598198 325154 598434
rect 324918 591198 325154 591434
rect 324918 584198 325154 584434
rect 324918 577198 325154 577434
rect 324918 570198 325154 570434
rect 324918 563198 325154 563434
rect 324918 556198 325154 556434
rect 324918 549198 325154 549434
rect 324918 542198 325154 542434
rect 324918 535198 325154 535434
rect 324918 528198 325154 528434
rect 324918 521198 325154 521434
rect 324918 514198 325154 514434
rect 324918 507198 325154 507434
rect 324918 500198 325154 500434
rect 324918 493198 325154 493434
rect 324918 486198 325154 486434
rect 324918 479198 325154 479434
rect 324918 472198 325154 472434
rect 324918 465198 325154 465434
rect 324918 458198 325154 458434
rect 324918 451198 325154 451434
rect 324918 444198 325154 444434
rect 324918 437198 325154 437434
rect 324918 430198 325154 430434
rect 324918 423198 325154 423434
rect 324918 416198 325154 416434
rect 324918 409198 325154 409434
rect 324918 402198 325154 402434
rect 324918 395198 325154 395434
rect 324918 388198 325154 388434
rect 324918 381198 325154 381434
rect 324918 374198 325154 374434
rect 324918 367198 325154 367434
rect 324918 360198 325154 360434
rect 324918 353198 325154 353434
rect 324918 346198 325154 346434
rect 324918 339198 325154 339434
rect 324918 332198 325154 332434
rect 324918 325198 325154 325434
rect 324918 318198 325154 318434
rect 324918 311198 325154 311434
rect 324918 304198 325154 304434
rect 324918 297198 325154 297434
rect 324918 290198 325154 290434
rect 324918 283198 325154 283434
rect 324918 276198 325154 276434
rect 324918 269198 325154 269434
rect 324918 262198 325154 262434
rect 324918 255198 325154 255434
rect 324918 248198 325154 248434
rect 324918 241198 325154 241434
rect 324918 234198 325154 234434
rect 324918 227198 325154 227434
rect 324918 220198 325154 220434
rect 324918 213198 325154 213434
rect 324918 206198 325154 206434
rect 324918 199198 325154 199434
rect 324918 192198 325154 192434
rect 324918 185198 325154 185434
rect 324918 178198 325154 178434
rect 324918 171198 325154 171434
rect 324918 164198 325154 164434
rect 324918 157198 325154 157434
rect 324918 150198 325154 150434
rect 324918 143198 325154 143434
rect 324918 136198 325154 136434
rect 324918 129198 325154 129434
rect 324918 122198 325154 122434
rect 324918 115198 325154 115434
rect 324918 108198 325154 108434
rect 324918 101198 325154 101434
rect 324918 94198 325154 94434
rect 324918 87198 325154 87434
rect 324918 80198 325154 80434
rect 324918 73198 325154 73434
rect 324918 66198 325154 66434
rect 324918 59198 325154 59434
rect 324918 52198 325154 52434
rect 324918 45198 325154 45434
rect 324918 38198 325154 38434
rect 324918 31198 325154 31434
rect 324918 24198 325154 24434
rect 324918 17198 325154 17434
rect 324918 10198 325154 10434
rect 324918 3198 325154 3434
rect 324918 -1942 325154 -1706
rect 324918 -2262 325154 -2026
rect 330186 705002 330422 705238
rect 330186 704682 330422 704918
rect 330186 695258 330422 695494
rect 330186 688258 330422 688494
rect 330186 681258 330422 681494
rect 330186 674258 330422 674494
rect 330186 667258 330422 667494
rect 330186 660258 330422 660494
rect 330186 653258 330422 653494
rect 330186 646258 330422 646494
rect 330186 639258 330422 639494
rect 330186 632258 330422 632494
rect 330186 625258 330422 625494
rect 330186 618258 330422 618494
rect 330186 611258 330422 611494
rect 330186 604258 330422 604494
rect 330186 597258 330422 597494
rect 330186 590258 330422 590494
rect 330186 583258 330422 583494
rect 330186 576258 330422 576494
rect 330186 569258 330422 569494
rect 330186 562258 330422 562494
rect 330186 555258 330422 555494
rect 330186 548258 330422 548494
rect 330186 541258 330422 541494
rect 330186 534258 330422 534494
rect 330186 527258 330422 527494
rect 330186 520258 330422 520494
rect 330186 513258 330422 513494
rect 330186 506258 330422 506494
rect 330186 499258 330422 499494
rect 330186 492258 330422 492494
rect 330186 485258 330422 485494
rect 330186 478258 330422 478494
rect 330186 471258 330422 471494
rect 330186 464258 330422 464494
rect 330186 457258 330422 457494
rect 330186 450258 330422 450494
rect 330186 443258 330422 443494
rect 330186 436258 330422 436494
rect 330186 429258 330422 429494
rect 330186 422258 330422 422494
rect 330186 415258 330422 415494
rect 330186 408258 330422 408494
rect 330186 401258 330422 401494
rect 330186 394258 330422 394494
rect 330186 387258 330422 387494
rect 330186 380258 330422 380494
rect 330186 373258 330422 373494
rect 330186 366258 330422 366494
rect 330186 359258 330422 359494
rect 330186 352258 330422 352494
rect 330186 345258 330422 345494
rect 330186 338258 330422 338494
rect 330186 331258 330422 331494
rect 330186 324258 330422 324494
rect 330186 317258 330422 317494
rect 330186 310258 330422 310494
rect 330186 303258 330422 303494
rect 330186 296258 330422 296494
rect 330186 289258 330422 289494
rect 330186 282258 330422 282494
rect 330186 275258 330422 275494
rect 330186 268258 330422 268494
rect 330186 261258 330422 261494
rect 330186 254258 330422 254494
rect 330186 247258 330422 247494
rect 330186 240258 330422 240494
rect 330186 233258 330422 233494
rect 330186 226258 330422 226494
rect 330186 219258 330422 219494
rect 330186 212258 330422 212494
rect 330186 205258 330422 205494
rect 330186 198258 330422 198494
rect 330186 191258 330422 191494
rect 330186 184258 330422 184494
rect 330186 177258 330422 177494
rect 330186 170258 330422 170494
rect 330186 163258 330422 163494
rect 330186 156258 330422 156494
rect 330186 149258 330422 149494
rect 330186 142258 330422 142494
rect 330186 135258 330422 135494
rect 330186 128258 330422 128494
rect 330186 121258 330422 121494
rect 330186 114258 330422 114494
rect 330186 107258 330422 107494
rect 330186 100258 330422 100494
rect 330186 93258 330422 93494
rect 330186 86258 330422 86494
rect 330186 79258 330422 79494
rect 330186 72258 330422 72494
rect 330186 65258 330422 65494
rect 330186 58258 330422 58494
rect 330186 51258 330422 51494
rect 330186 44258 330422 44494
rect 330186 37258 330422 37494
rect 330186 30258 330422 30494
rect 330186 23258 330422 23494
rect 330186 16258 330422 16494
rect 330186 9258 330422 9494
rect 330186 2258 330422 2494
rect 330186 -982 330422 -746
rect 330186 -1302 330422 -1066
rect 331918 705962 332154 706198
rect 331918 705642 332154 705878
rect 331918 696198 332154 696434
rect 331918 689198 332154 689434
rect 331918 682198 332154 682434
rect 331918 675198 332154 675434
rect 331918 668198 332154 668434
rect 331918 661198 332154 661434
rect 331918 654198 332154 654434
rect 331918 647198 332154 647434
rect 331918 640198 332154 640434
rect 331918 633198 332154 633434
rect 331918 626198 332154 626434
rect 331918 619198 332154 619434
rect 331918 612198 332154 612434
rect 331918 605198 332154 605434
rect 331918 598198 332154 598434
rect 331918 591198 332154 591434
rect 331918 584198 332154 584434
rect 331918 577198 332154 577434
rect 331918 570198 332154 570434
rect 331918 563198 332154 563434
rect 331918 556198 332154 556434
rect 331918 549198 332154 549434
rect 331918 542198 332154 542434
rect 331918 535198 332154 535434
rect 331918 528198 332154 528434
rect 331918 521198 332154 521434
rect 331918 514198 332154 514434
rect 331918 507198 332154 507434
rect 331918 500198 332154 500434
rect 331918 493198 332154 493434
rect 331918 486198 332154 486434
rect 331918 479198 332154 479434
rect 331918 472198 332154 472434
rect 331918 465198 332154 465434
rect 331918 458198 332154 458434
rect 331918 451198 332154 451434
rect 331918 444198 332154 444434
rect 331918 437198 332154 437434
rect 331918 430198 332154 430434
rect 331918 423198 332154 423434
rect 331918 416198 332154 416434
rect 331918 409198 332154 409434
rect 331918 402198 332154 402434
rect 331918 395198 332154 395434
rect 331918 388198 332154 388434
rect 331918 381198 332154 381434
rect 331918 374198 332154 374434
rect 331918 367198 332154 367434
rect 331918 360198 332154 360434
rect 331918 353198 332154 353434
rect 331918 346198 332154 346434
rect 331918 339198 332154 339434
rect 331918 332198 332154 332434
rect 331918 325198 332154 325434
rect 331918 318198 332154 318434
rect 331918 311198 332154 311434
rect 331918 304198 332154 304434
rect 331918 297198 332154 297434
rect 331918 290198 332154 290434
rect 331918 283198 332154 283434
rect 331918 276198 332154 276434
rect 331918 269198 332154 269434
rect 331918 262198 332154 262434
rect 331918 255198 332154 255434
rect 331918 248198 332154 248434
rect 331918 241198 332154 241434
rect 331918 234198 332154 234434
rect 331918 227198 332154 227434
rect 331918 220198 332154 220434
rect 331918 213198 332154 213434
rect 331918 206198 332154 206434
rect 331918 199198 332154 199434
rect 331918 192198 332154 192434
rect 331918 185198 332154 185434
rect 331918 178198 332154 178434
rect 331918 171198 332154 171434
rect 331918 164198 332154 164434
rect 331918 157198 332154 157434
rect 331918 150198 332154 150434
rect 331918 143198 332154 143434
rect 331918 136198 332154 136434
rect 331918 129198 332154 129434
rect 331918 122198 332154 122434
rect 331918 115198 332154 115434
rect 331918 108198 332154 108434
rect 331918 101198 332154 101434
rect 331918 94198 332154 94434
rect 331918 87198 332154 87434
rect 331918 80198 332154 80434
rect 331918 73198 332154 73434
rect 331918 66198 332154 66434
rect 331918 59198 332154 59434
rect 331918 52198 332154 52434
rect 331918 45198 332154 45434
rect 331918 38198 332154 38434
rect 331918 31198 332154 31434
rect 331918 24198 332154 24434
rect 331918 17198 332154 17434
rect 331918 10198 332154 10434
rect 331918 3198 332154 3434
rect 331918 -1942 332154 -1706
rect 331918 -2262 332154 -2026
rect 337186 705002 337422 705238
rect 337186 704682 337422 704918
rect 337186 695258 337422 695494
rect 337186 688258 337422 688494
rect 337186 681258 337422 681494
rect 337186 674258 337422 674494
rect 337186 667258 337422 667494
rect 337186 660258 337422 660494
rect 337186 653258 337422 653494
rect 337186 646258 337422 646494
rect 337186 639258 337422 639494
rect 337186 632258 337422 632494
rect 337186 625258 337422 625494
rect 337186 618258 337422 618494
rect 337186 611258 337422 611494
rect 337186 604258 337422 604494
rect 337186 597258 337422 597494
rect 337186 590258 337422 590494
rect 337186 583258 337422 583494
rect 337186 576258 337422 576494
rect 337186 569258 337422 569494
rect 337186 562258 337422 562494
rect 337186 555258 337422 555494
rect 337186 548258 337422 548494
rect 337186 541258 337422 541494
rect 337186 534258 337422 534494
rect 337186 527258 337422 527494
rect 337186 520258 337422 520494
rect 337186 513258 337422 513494
rect 337186 506258 337422 506494
rect 337186 499258 337422 499494
rect 337186 492258 337422 492494
rect 337186 485258 337422 485494
rect 337186 478258 337422 478494
rect 337186 471258 337422 471494
rect 337186 464258 337422 464494
rect 337186 457258 337422 457494
rect 337186 450258 337422 450494
rect 337186 443258 337422 443494
rect 337186 436258 337422 436494
rect 337186 429258 337422 429494
rect 337186 422258 337422 422494
rect 337186 415258 337422 415494
rect 337186 408258 337422 408494
rect 337186 401258 337422 401494
rect 337186 394258 337422 394494
rect 337186 387258 337422 387494
rect 337186 380258 337422 380494
rect 337186 373258 337422 373494
rect 337186 366258 337422 366494
rect 337186 359258 337422 359494
rect 337186 352258 337422 352494
rect 337186 345258 337422 345494
rect 337186 338258 337422 338494
rect 337186 331258 337422 331494
rect 337186 324258 337422 324494
rect 337186 317258 337422 317494
rect 337186 310258 337422 310494
rect 337186 303258 337422 303494
rect 337186 296258 337422 296494
rect 337186 289258 337422 289494
rect 337186 282258 337422 282494
rect 337186 275258 337422 275494
rect 337186 268258 337422 268494
rect 337186 261258 337422 261494
rect 337186 254258 337422 254494
rect 337186 247258 337422 247494
rect 337186 240258 337422 240494
rect 337186 233258 337422 233494
rect 337186 226258 337422 226494
rect 337186 219258 337422 219494
rect 337186 212258 337422 212494
rect 337186 205258 337422 205494
rect 337186 198258 337422 198494
rect 337186 191258 337422 191494
rect 337186 184258 337422 184494
rect 337186 177258 337422 177494
rect 337186 170258 337422 170494
rect 337186 163258 337422 163494
rect 337186 156258 337422 156494
rect 337186 149258 337422 149494
rect 337186 142258 337422 142494
rect 337186 135258 337422 135494
rect 337186 128258 337422 128494
rect 337186 121258 337422 121494
rect 337186 114258 337422 114494
rect 337186 107258 337422 107494
rect 337186 100258 337422 100494
rect 337186 93258 337422 93494
rect 337186 86258 337422 86494
rect 337186 79258 337422 79494
rect 337186 72258 337422 72494
rect 337186 65258 337422 65494
rect 337186 58258 337422 58494
rect 337186 51258 337422 51494
rect 337186 44258 337422 44494
rect 337186 37258 337422 37494
rect 337186 30258 337422 30494
rect 337186 23258 337422 23494
rect 337186 16258 337422 16494
rect 337186 9258 337422 9494
rect 337186 2258 337422 2494
rect 337186 -982 337422 -746
rect 337186 -1302 337422 -1066
rect 338918 705962 339154 706198
rect 338918 705642 339154 705878
rect 338918 696198 339154 696434
rect 338918 689198 339154 689434
rect 338918 682198 339154 682434
rect 338918 675198 339154 675434
rect 338918 668198 339154 668434
rect 338918 661198 339154 661434
rect 338918 654198 339154 654434
rect 338918 647198 339154 647434
rect 338918 640198 339154 640434
rect 338918 633198 339154 633434
rect 338918 626198 339154 626434
rect 338918 619198 339154 619434
rect 338918 612198 339154 612434
rect 338918 605198 339154 605434
rect 338918 598198 339154 598434
rect 338918 591198 339154 591434
rect 338918 584198 339154 584434
rect 338918 577198 339154 577434
rect 338918 570198 339154 570434
rect 338918 563198 339154 563434
rect 338918 556198 339154 556434
rect 338918 549198 339154 549434
rect 338918 542198 339154 542434
rect 338918 535198 339154 535434
rect 338918 528198 339154 528434
rect 338918 521198 339154 521434
rect 338918 514198 339154 514434
rect 338918 507198 339154 507434
rect 338918 500198 339154 500434
rect 338918 493198 339154 493434
rect 338918 486198 339154 486434
rect 338918 479198 339154 479434
rect 338918 472198 339154 472434
rect 338918 465198 339154 465434
rect 338918 458198 339154 458434
rect 338918 451198 339154 451434
rect 338918 444198 339154 444434
rect 338918 437198 339154 437434
rect 338918 430198 339154 430434
rect 338918 423198 339154 423434
rect 338918 416198 339154 416434
rect 338918 409198 339154 409434
rect 338918 402198 339154 402434
rect 338918 395198 339154 395434
rect 338918 388198 339154 388434
rect 338918 381198 339154 381434
rect 338918 374198 339154 374434
rect 338918 367198 339154 367434
rect 338918 360198 339154 360434
rect 338918 353198 339154 353434
rect 338918 346198 339154 346434
rect 338918 339198 339154 339434
rect 338918 332198 339154 332434
rect 338918 325198 339154 325434
rect 338918 318198 339154 318434
rect 338918 311198 339154 311434
rect 338918 304198 339154 304434
rect 338918 297198 339154 297434
rect 338918 290198 339154 290434
rect 338918 283198 339154 283434
rect 338918 276198 339154 276434
rect 338918 269198 339154 269434
rect 338918 262198 339154 262434
rect 338918 255198 339154 255434
rect 338918 248198 339154 248434
rect 338918 241198 339154 241434
rect 338918 234198 339154 234434
rect 338918 227198 339154 227434
rect 338918 220198 339154 220434
rect 338918 213198 339154 213434
rect 338918 206198 339154 206434
rect 338918 199198 339154 199434
rect 338918 192198 339154 192434
rect 338918 185198 339154 185434
rect 338918 178198 339154 178434
rect 338918 171198 339154 171434
rect 338918 164198 339154 164434
rect 338918 157198 339154 157434
rect 338918 150198 339154 150434
rect 338918 143198 339154 143434
rect 338918 136198 339154 136434
rect 338918 129198 339154 129434
rect 338918 122198 339154 122434
rect 338918 115198 339154 115434
rect 338918 108198 339154 108434
rect 338918 101198 339154 101434
rect 338918 94198 339154 94434
rect 338918 87198 339154 87434
rect 338918 80198 339154 80434
rect 338918 73198 339154 73434
rect 338918 66198 339154 66434
rect 338918 59198 339154 59434
rect 338918 52198 339154 52434
rect 338918 45198 339154 45434
rect 338918 38198 339154 38434
rect 338918 31198 339154 31434
rect 338918 24198 339154 24434
rect 338918 17198 339154 17434
rect 338918 10198 339154 10434
rect 338918 3198 339154 3434
rect 338918 -1942 339154 -1706
rect 338918 -2262 339154 -2026
rect 344186 705002 344422 705238
rect 344186 704682 344422 704918
rect 344186 695258 344422 695494
rect 344186 688258 344422 688494
rect 344186 681258 344422 681494
rect 344186 674258 344422 674494
rect 344186 667258 344422 667494
rect 344186 660258 344422 660494
rect 344186 653258 344422 653494
rect 344186 646258 344422 646494
rect 344186 639258 344422 639494
rect 344186 632258 344422 632494
rect 344186 625258 344422 625494
rect 344186 618258 344422 618494
rect 344186 611258 344422 611494
rect 344186 604258 344422 604494
rect 344186 597258 344422 597494
rect 344186 590258 344422 590494
rect 344186 583258 344422 583494
rect 344186 576258 344422 576494
rect 344186 569258 344422 569494
rect 344186 562258 344422 562494
rect 344186 555258 344422 555494
rect 344186 548258 344422 548494
rect 344186 541258 344422 541494
rect 344186 534258 344422 534494
rect 344186 527258 344422 527494
rect 344186 520258 344422 520494
rect 344186 513258 344422 513494
rect 344186 506258 344422 506494
rect 344186 499258 344422 499494
rect 344186 492258 344422 492494
rect 344186 485258 344422 485494
rect 344186 478258 344422 478494
rect 344186 471258 344422 471494
rect 344186 464258 344422 464494
rect 344186 457258 344422 457494
rect 344186 450258 344422 450494
rect 344186 443258 344422 443494
rect 344186 436258 344422 436494
rect 344186 429258 344422 429494
rect 344186 422258 344422 422494
rect 344186 415258 344422 415494
rect 344186 408258 344422 408494
rect 344186 401258 344422 401494
rect 344186 394258 344422 394494
rect 344186 387258 344422 387494
rect 344186 380258 344422 380494
rect 344186 373258 344422 373494
rect 344186 366258 344422 366494
rect 344186 359258 344422 359494
rect 344186 352258 344422 352494
rect 344186 345258 344422 345494
rect 344186 338258 344422 338494
rect 344186 331258 344422 331494
rect 344186 324258 344422 324494
rect 344186 317258 344422 317494
rect 344186 310258 344422 310494
rect 344186 303258 344422 303494
rect 344186 296258 344422 296494
rect 344186 289258 344422 289494
rect 344186 282258 344422 282494
rect 344186 275258 344422 275494
rect 344186 268258 344422 268494
rect 344186 261258 344422 261494
rect 344186 254258 344422 254494
rect 344186 247258 344422 247494
rect 344186 240258 344422 240494
rect 344186 233258 344422 233494
rect 344186 226258 344422 226494
rect 344186 219258 344422 219494
rect 344186 212258 344422 212494
rect 344186 205258 344422 205494
rect 344186 198258 344422 198494
rect 344186 191258 344422 191494
rect 344186 184258 344422 184494
rect 344186 177258 344422 177494
rect 344186 170258 344422 170494
rect 344186 163258 344422 163494
rect 344186 156258 344422 156494
rect 344186 149258 344422 149494
rect 344186 142258 344422 142494
rect 344186 135258 344422 135494
rect 344186 128258 344422 128494
rect 344186 121258 344422 121494
rect 344186 114258 344422 114494
rect 344186 107258 344422 107494
rect 344186 100258 344422 100494
rect 344186 93258 344422 93494
rect 344186 86258 344422 86494
rect 344186 79258 344422 79494
rect 344186 72258 344422 72494
rect 344186 65258 344422 65494
rect 344186 58258 344422 58494
rect 344186 51258 344422 51494
rect 344186 44258 344422 44494
rect 344186 37258 344422 37494
rect 344186 30258 344422 30494
rect 344186 23258 344422 23494
rect 344186 16258 344422 16494
rect 344186 9258 344422 9494
rect 344186 2258 344422 2494
rect 344186 -982 344422 -746
rect 344186 -1302 344422 -1066
rect 345918 705962 346154 706198
rect 345918 705642 346154 705878
rect 345918 696198 346154 696434
rect 345918 689198 346154 689434
rect 345918 682198 346154 682434
rect 345918 675198 346154 675434
rect 345918 668198 346154 668434
rect 345918 661198 346154 661434
rect 345918 654198 346154 654434
rect 345918 647198 346154 647434
rect 345918 640198 346154 640434
rect 345918 633198 346154 633434
rect 345918 626198 346154 626434
rect 345918 619198 346154 619434
rect 345918 612198 346154 612434
rect 345918 605198 346154 605434
rect 345918 598198 346154 598434
rect 345918 591198 346154 591434
rect 345918 584198 346154 584434
rect 345918 577198 346154 577434
rect 345918 570198 346154 570434
rect 345918 563198 346154 563434
rect 345918 556198 346154 556434
rect 345918 549198 346154 549434
rect 345918 542198 346154 542434
rect 345918 535198 346154 535434
rect 345918 528198 346154 528434
rect 345918 521198 346154 521434
rect 345918 514198 346154 514434
rect 345918 507198 346154 507434
rect 345918 500198 346154 500434
rect 345918 493198 346154 493434
rect 345918 486198 346154 486434
rect 345918 479198 346154 479434
rect 345918 472198 346154 472434
rect 345918 465198 346154 465434
rect 345918 458198 346154 458434
rect 345918 451198 346154 451434
rect 345918 444198 346154 444434
rect 345918 437198 346154 437434
rect 345918 430198 346154 430434
rect 345918 423198 346154 423434
rect 345918 416198 346154 416434
rect 345918 409198 346154 409434
rect 345918 402198 346154 402434
rect 345918 395198 346154 395434
rect 345918 388198 346154 388434
rect 345918 381198 346154 381434
rect 345918 374198 346154 374434
rect 345918 367198 346154 367434
rect 345918 360198 346154 360434
rect 345918 353198 346154 353434
rect 345918 346198 346154 346434
rect 345918 339198 346154 339434
rect 345918 332198 346154 332434
rect 345918 325198 346154 325434
rect 345918 318198 346154 318434
rect 345918 311198 346154 311434
rect 345918 304198 346154 304434
rect 345918 297198 346154 297434
rect 345918 290198 346154 290434
rect 345918 283198 346154 283434
rect 345918 276198 346154 276434
rect 345918 269198 346154 269434
rect 345918 262198 346154 262434
rect 345918 255198 346154 255434
rect 345918 248198 346154 248434
rect 345918 241198 346154 241434
rect 345918 234198 346154 234434
rect 345918 227198 346154 227434
rect 345918 220198 346154 220434
rect 345918 213198 346154 213434
rect 345918 206198 346154 206434
rect 345918 199198 346154 199434
rect 345918 192198 346154 192434
rect 345918 185198 346154 185434
rect 345918 178198 346154 178434
rect 345918 171198 346154 171434
rect 345918 164198 346154 164434
rect 345918 157198 346154 157434
rect 345918 150198 346154 150434
rect 345918 143198 346154 143434
rect 345918 136198 346154 136434
rect 345918 129198 346154 129434
rect 345918 122198 346154 122434
rect 345918 115198 346154 115434
rect 345918 108198 346154 108434
rect 345918 101198 346154 101434
rect 345918 94198 346154 94434
rect 345918 87198 346154 87434
rect 345918 80198 346154 80434
rect 345918 73198 346154 73434
rect 345918 66198 346154 66434
rect 345918 59198 346154 59434
rect 345918 52198 346154 52434
rect 345918 45198 346154 45434
rect 345918 38198 346154 38434
rect 345918 31198 346154 31434
rect 345918 24198 346154 24434
rect 345918 17198 346154 17434
rect 345918 10198 346154 10434
rect 345918 3198 346154 3434
rect 345918 -1942 346154 -1706
rect 345918 -2262 346154 -2026
rect 351186 705002 351422 705238
rect 351186 704682 351422 704918
rect 351186 695258 351422 695494
rect 351186 688258 351422 688494
rect 351186 681258 351422 681494
rect 351186 674258 351422 674494
rect 351186 667258 351422 667494
rect 351186 660258 351422 660494
rect 351186 653258 351422 653494
rect 351186 646258 351422 646494
rect 351186 639258 351422 639494
rect 351186 632258 351422 632494
rect 351186 625258 351422 625494
rect 351186 618258 351422 618494
rect 351186 611258 351422 611494
rect 351186 604258 351422 604494
rect 351186 597258 351422 597494
rect 351186 590258 351422 590494
rect 351186 583258 351422 583494
rect 351186 576258 351422 576494
rect 351186 569258 351422 569494
rect 351186 562258 351422 562494
rect 351186 555258 351422 555494
rect 351186 548258 351422 548494
rect 351186 541258 351422 541494
rect 351186 534258 351422 534494
rect 351186 527258 351422 527494
rect 351186 520258 351422 520494
rect 351186 513258 351422 513494
rect 351186 506258 351422 506494
rect 351186 499258 351422 499494
rect 351186 492258 351422 492494
rect 351186 485258 351422 485494
rect 351186 478258 351422 478494
rect 351186 471258 351422 471494
rect 351186 464258 351422 464494
rect 351186 457258 351422 457494
rect 351186 450258 351422 450494
rect 351186 443258 351422 443494
rect 351186 436258 351422 436494
rect 351186 429258 351422 429494
rect 351186 422258 351422 422494
rect 351186 415258 351422 415494
rect 351186 408258 351422 408494
rect 351186 401258 351422 401494
rect 351186 394258 351422 394494
rect 351186 387258 351422 387494
rect 351186 380258 351422 380494
rect 351186 373258 351422 373494
rect 351186 366258 351422 366494
rect 351186 359258 351422 359494
rect 351186 352258 351422 352494
rect 351186 345258 351422 345494
rect 351186 338258 351422 338494
rect 351186 331258 351422 331494
rect 351186 324258 351422 324494
rect 351186 317258 351422 317494
rect 351186 310258 351422 310494
rect 351186 303258 351422 303494
rect 351186 296258 351422 296494
rect 351186 289258 351422 289494
rect 351186 282258 351422 282494
rect 351186 275258 351422 275494
rect 351186 268258 351422 268494
rect 351186 261258 351422 261494
rect 351186 254258 351422 254494
rect 351186 247258 351422 247494
rect 351186 240258 351422 240494
rect 351186 233258 351422 233494
rect 351186 226258 351422 226494
rect 351186 219258 351422 219494
rect 351186 212258 351422 212494
rect 351186 205258 351422 205494
rect 351186 198258 351422 198494
rect 351186 191258 351422 191494
rect 351186 184258 351422 184494
rect 351186 177258 351422 177494
rect 351186 170258 351422 170494
rect 351186 163258 351422 163494
rect 351186 156258 351422 156494
rect 351186 149258 351422 149494
rect 351186 142258 351422 142494
rect 351186 135258 351422 135494
rect 351186 128258 351422 128494
rect 351186 121258 351422 121494
rect 351186 114258 351422 114494
rect 351186 107258 351422 107494
rect 351186 100258 351422 100494
rect 351186 93258 351422 93494
rect 351186 86258 351422 86494
rect 351186 79258 351422 79494
rect 351186 72258 351422 72494
rect 351186 65258 351422 65494
rect 351186 58258 351422 58494
rect 351186 51258 351422 51494
rect 351186 44258 351422 44494
rect 351186 37258 351422 37494
rect 351186 30258 351422 30494
rect 351186 23258 351422 23494
rect 351186 16258 351422 16494
rect 351186 9258 351422 9494
rect 351186 2258 351422 2494
rect 351186 -982 351422 -746
rect 351186 -1302 351422 -1066
rect 352918 705962 353154 706198
rect 352918 705642 353154 705878
rect 352918 696198 353154 696434
rect 352918 689198 353154 689434
rect 352918 682198 353154 682434
rect 352918 675198 353154 675434
rect 352918 668198 353154 668434
rect 352918 661198 353154 661434
rect 352918 654198 353154 654434
rect 352918 647198 353154 647434
rect 352918 640198 353154 640434
rect 352918 633198 353154 633434
rect 352918 626198 353154 626434
rect 352918 619198 353154 619434
rect 352918 612198 353154 612434
rect 352918 605198 353154 605434
rect 352918 598198 353154 598434
rect 352918 591198 353154 591434
rect 352918 584198 353154 584434
rect 352918 577198 353154 577434
rect 352918 570198 353154 570434
rect 352918 563198 353154 563434
rect 352918 556198 353154 556434
rect 352918 549198 353154 549434
rect 352918 542198 353154 542434
rect 352918 535198 353154 535434
rect 352918 528198 353154 528434
rect 352918 521198 353154 521434
rect 352918 514198 353154 514434
rect 352918 507198 353154 507434
rect 352918 500198 353154 500434
rect 352918 493198 353154 493434
rect 352918 486198 353154 486434
rect 352918 479198 353154 479434
rect 352918 472198 353154 472434
rect 352918 465198 353154 465434
rect 352918 458198 353154 458434
rect 352918 451198 353154 451434
rect 352918 444198 353154 444434
rect 352918 437198 353154 437434
rect 352918 430198 353154 430434
rect 352918 423198 353154 423434
rect 352918 416198 353154 416434
rect 352918 409198 353154 409434
rect 352918 402198 353154 402434
rect 352918 395198 353154 395434
rect 352918 388198 353154 388434
rect 352918 381198 353154 381434
rect 352918 374198 353154 374434
rect 352918 367198 353154 367434
rect 352918 360198 353154 360434
rect 352918 353198 353154 353434
rect 352918 346198 353154 346434
rect 352918 339198 353154 339434
rect 352918 332198 353154 332434
rect 352918 325198 353154 325434
rect 352918 318198 353154 318434
rect 352918 311198 353154 311434
rect 352918 304198 353154 304434
rect 352918 297198 353154 297434
rect 352918 290198 353154 290434
rect 352918 283198 353154 283434
rect 352918 276198 353154 276434
rect 352918 269198 353154 269434
rect 352918 262198 353154 262434
rect 352918 255198 353154 255434
rect 352918 248198 353154 248434
rect 352918 241198 353154 241434
rect 352918 234198 353154 234434
rect 352918 227198 353154 227434
rect 352918 220198 353154 220434
rect 352918 213198 353154 213434
rect 352918 206198 353154 206434
rect 352918 199198 353154 199434
rect 352918 192198 353154 192434
rect 352918 185198 353154 185434
rect 352918 178198 353154 178434
rect 352918 171198 353154 171434
rect 352918 164198 353154 164434
rect 352918 157198 353154 157434
rect 352918 150198 353154 150434
rect 352918 143198 353154 143434
rect 352918 136198 353154 136434
rect 352918 129198 353154 129434
rect 352918 122198 353154 122434
rect 352918 115198 353154 115434
rect 352918 108198 353154 108434
rect 352918 101198 353154 101434
rect 352918 94198 353154 94434
rect 352918 87198 353154 87434
rect 352918 80198 353154 80434
rect 352918 73198 353154 73434
rect 352918 66198 353154 66434
rect 352918 59198 353154 59434
rect 352918 52198 353154 52434
rect 352918 45198 353154 45434
rect 352918 38198 353154 38434
rect 352918 31198 353154 31434
rect 352918 24198 353154 24434
rect 352918 17198 353154 17434
rect 352918 10198 353154 10434
rect 352918 3198 353154 3434
rect 352918 -1942 353154 -1706
rect 352918 -2262 353154 -2026
rect 358186 705002 358422 705238
rect 358186 704682 358422 704918
rect 358186 695258 358422 695494
rect 358186 688258 358422 688494
rect 358186 681258 358422 681494
rect 358186 674258 358422 674494
rect 358186 667258 358422 667494
rect 358186 660258 358422 660494
rect 358186 653258 358422 653494
rect 358186 646258 358422 646494
rect 358186 639258 358422 639494
rect 358186 632258 358422 632494
rect 358186 625258 358422 625494
rect 358186 618258 358422 618494
rect 358186 611258 358422 611494
rect 358186 604258 358422 604494
rect 358186 597258 358422 597494
rect 358186 590258 358422 590494
rect 358186 583258 358422 583494
rect 358186 576258 358422 576494
rect 358186 569258 358422 569494
rect 358186 562258 358422 562494
rect 358186 555258 358422 555494
rect 358186 548258 358422 548494
rect 358186 541258 358422 541494
rect 358186 534258 358422 534494
rect 358186 527258 358422 527494
rect 358186 520258 358422 520494
rect 358186 513258 358422 513494
rect 358186 506258 358422 506494
rect 358186 499258 358422 499494
rect 358186 492258 358422 492494
rect 358186 485258 358422 485494
rect 358186 478258 358422 478494
rect 358186 471258 358422 471494
rect 358186 464258 358422 464494
rect 358186 457258 358422 457494
rect 358186 450258 358422 450494
rect 358186 443258 358422 443494
rect 358186 436258 358422 436494
rect 358186 429258 358422 429494
rect 358186 422258 358422 422494
rect 358186 415258 358422 415494
rect 358186 408258 358422 408494
rect 358186 401258 358422 401494
rect 358186 394258 358422 394494
rect 358186 387258 358422 387494
rect 358186 380258 358422 380494
rect 358186 373258 358422 373494
rect 358186 366258 358422 366494
rect 358186 359258 358422 359494
rect 358186 352258 358422 352494
rect 358186 345258 358422 345494
rect 358186 338258 358422 338494
rect 358186 331258 358422 331494
rect 358186 324258 358422 324494
rect 358186 317258 358422 317494
rect 358186 310258 358422 310494
rect 358186 303258 358422 303494
rect 358186 296258 358422 296494
rect 358186 289258 358422 289494
rect 358186 282258 358422 282494
rect 358186 275258 358422 275494
rect 358186 268258 358422 268494
rect 358186 261258 358422 261494
rect 358186 254258 358422 254494
rect 358186 247258 358422 247494
rect 358186 240258 358422 240494
rect 358186 233258 358422 233494
rect 358186 226258 358422 226494
rect 358186 219258 358422 219494
rect 358186 212258 358422 212494
rect 358186 205258 358422 205494
rect 358186 198258 358422 198494
rect 358186 191258 358422 191494
rect 358186 184258 358422 184494
rect 358186 177258 358422 177494
rect 358186 170258 358422 170494
rect 358186 163258 358422 163494
rect 358186 156258 358422 156494
rect 358186 149258 358422 149494
rect 358186 142258 358422 142494
rect 358186 135258 358422 135494
rect 358186 128258 358422 128494
rect 358186 121258 358422 121494
rect 358186 114258 358422 114494
rect 358186 107258 358422 107494
rect 358186 100258 358422 100494
rect 358186 93258 358422 93494
rect 358186 86258 358422 86494
rect 358186 79258 358422 79494
rect 358186 72258 358422 72494
rect 358186 65258 358422 65494
rect 358186 58258 358422 58494
rect 358186 51258 358422 51494
rect 358186 44258 358422 44494
rect 358186 37258 358422 37494
rect 358186 30258 358422 30494
rect 358186 23258 358422 23494
rect 358186 16258 358422 16494
rect 358186 9258 358422 9494
rect 358186 2258 358422 2494
rect 358186 -982 358422 -746
rect 358186 -1302 358422 -1066
rect 359918 705962 360154 706198
rect 359918 705642 360154 705878
rect 359918 696198 360154 696434
rect 359918 689198 360154 689434
rect 359918 682198 360154 682434
rect 359918 675198 360154 675434
rect 359918 668198 360154 668434
rect 359918 661198 360154 661434
rect 359918 654198 360154 654434
rect 359918 647198 360154 647434
rect 359918 640198 360154 640434
rect 359918 633198 360154 633434
rect 359918 626198 360154 626434
rect 359918 619198 360154 619434
rect 359918 612198 360154 612434
rect 359918 605198 360154 605434
rect 359918 598198 360154 598434
rect 359918 591198 360154 591434
rect 359918 584198 360154 584434
rect 359918 577198 360154 577434
rect 359918 570198 360154 570434
rect 359918 563198 360154 563434
rect 359918 556198 360154 556434
rect 359918 549198 360154 549434
rect 359918 542198 360154 542434
rect 359918 535198 360154 535434
rect 359918 528198 360154 528434
rect 359918 521198 360154 521434
rect 359918 514198 360154 514434
rect 359918 507198 360154 507434
rect 359918 500198 360154 500434
rect 359918 493198 360154 493434
rect 359918 486198 360154 486434
rect 359918 479198 360154 479434
rect 359918 472198 360154 472434
rect 359918 465198 360154 465434
rect 359918 458198 360154 458434
rect 359918 451198 360154 451434
rect 359918 444198 360154 444434
rect 359918 437198 360154 437434
rect 359918 430198 360154 430434
rect 359918 423198 360154 423434
rect 359918 416198 360154 416434
rect 359918 409198 360154 409434
rect 359918 402198 360154 402434
rect 359918 395198 360154 395434
rect 359918 388198 360154 388434
rect 359918 381198 360154 381434
rect 359918 374198 360154 374434
rect 359918 367198 360154 367434
rect 359918 360198 360154 360434
rect 359918 353198 360154 353434
rect 359918 346198 360154 346434
rect 359918 339198 360154 339434
rect 359918 332198 360154 332434
rect 359918 325198 360154 325434
rect 359918 318198 360154 318434
rect 359918 311198 360154 311434
rect 359918 304198 360154 304434
rect 359918 297198 360154 297434
rect 359918 290198 360154 290434
rect 359918 283198 360154 283434
rect 359918 276198 360154 276434
rect 359918 269198 360154 269434
rect 359918 262198 360154 262434
rect 359918 255198 360154 255434
rect 359918 248198 360154 248434
rect 359918 241198 360154 241434
rect 359918 234198 360154 234434
rect 359918 227198 360154 227434
rect 359918 220198 360154 220434
rect 359918 213198 360154 213434
rect 359918 206198 360154 206434
rect 359918 199198 360154 199434
rect 359918 192198 360154 192434
rect 359918 185198 360154 185434
rect 359918 178198 360154 178434
rect 359918 171198 360154 171434
rect 359918 164198 360154 164434
rect 359918 157198 360154 157434
rect 359918 150198 360154 150434
rect 359918 143198 360154 143434
rect 359918 136198 360154 136434
rect 359918 129198 360154 129434
rect 359918 122198 360154 122434
rect 359918 115198 360154 115434
rect 359918 108198 360154 108434
rect 359918 101198 360154 101434
rect 359918 94198 360154 94434
rect 359918 87198 360154 87434
rect 359918 80198 360154 80434
rect 359918 73198 360154 73434
rect 359918 66198 360154 66434
rect 359918 59198 360154 59434
rect 359918 52198 360154 52434
rect 359918 45198 360154 45434
rect 359918 38198 360154 38434
rect 359918 31198 360154 31434
rect 359918 24198 360154 24434
rect 359918 17198 360154 17434
rect 359918 10198 360154 10434
rect 359918 3198 360154 3434
rect 359918 -1942 360154 -1706
rect 359918 -2262 360154 -2026
rect 365186 705002 365422 705238
rect 365186 704682 365422 704918
rect 365186 695258 365422 695494
rect 365186 688258 365422 688494
rect 365186 681258 365422 681494
rect 365186 674258 365422 674494
rect 365186 667258 365422 667494
rect 365186 660258 365422 660494
rect 365186 653258 365422 653494
rect 365186 646258 365422 646494
rect 365186 639258 365422 639494
rect 365186 632258 365422 632494
rect 365186 625258 365422 625494
rect 365186 618258 365422 618494
rect 365186 611258 365422 611494
rect 365186 604258 365422 604494
rect 365186 597258 365422 597494
rect 365186 590258 365422 590494
rect 365186 583258 365422 583494
rect 365186 576258 365422 576494
rect 365186 569258 365422 569494
rect 365186 562258 365422 562494
rect 365186 555258 365422 555494
rect 365186 548258 365422 548494
rect 365186 541258 365422 541494
rect 365186 534258 365422 534494
rect 365186 527258 365422 527494
rect 365186 520258 365422 520494
rect 365186 513258 365422 513494
rect 365186 506258 365422 506494
rect 365186 499258 365422 499494
rect 365186 492258 365422 492494
rect 365186 485258 365422 485494
rect 365186 478258 365422 478494
rect 365186 471258 365422 471494
rect 365186 464258 365422 464494
rect 365186 457258 365422 457494
rect 365186 450258 365422 450494
rect 365186 443258 365422 443494
rect 365186 436258 365422 436494
rect 365186 429258 365422 429494
rect 365186 422258 365422 422494
rect 365186 415258 365422 415494
rect 365186 408258 365422 408494
rect 365186 401258 365422 401494
rect 365186 394258 365422 394494
rect 365186 387258 365422 387494
rect 365186 380258 365422 380494
rect 365186 373258 365422 373494
rect 365186 366258 365422 366494
rect 365186 359258 365422 359494
rect 365186 352258 365422 352494
rect 365186 345258 365422 345494
rect 365186 338258 365422 338494
rect 365186 331258 365422 331494
rect 365186 324258 365422 324494
rect 365186 317258 365422 317494
rect 365186 310258 365422 310494
rect 365186 303258 365422 303494
rect 365186 296258 365422 296494
rect 365186 289258 365422 289494
rect 365186 282258 365422 282494
rect 365186 275258 365422 275494
rect 365186 268258 365422 268494
rect 365186 261258 365422 261494
rect 365186 254258 365422 254494
rect 365186 247258 365422 247494
rect 365186 240258 365422 240494
rect 365186 233258 365422 233494
rect 365186 226258 365422 226494
rect 365186 219258 365422 219494
rect 365186 212258 365422 212494
rect 365186 205258 365422 205494
rect 365186 198258 365422 198494
rect 365186 191258 365422 191494
rect 365186 184258 365422 184494
rect 365186 177258 365422 177494
rect 365186 170258 365422 170494
rect 365186 163258 365422 163494
rect 365186 156258 365422 156494
rect 365186 149258 365422 149494
rect 365186 142258 365422 142494
rect 365186 135258 365422 135494
rect 365186 128258 365422 128494
rect 365186 121258 365422 121494
rect 365186 114258 365422 114494
rect 365186 107258 365422 107494
rect 365186 100258 365422 100494
rect 365186 93258 365422 93494
rect 365186 86258 365422 86494
rect 365186 79258 365422 79494
rect 365186 72258 365422 72494
rect 365186 65258 365422 65494
rect 365186 58258 365422 58494
rect 365186 51258 365422 51494
rect 365186 44258 365422 44494
rect 365186 37258 365422 37494
rect 365186 30258 365422 30494
rect 365186 23258 365422 23494
rect 365186 16258 365422 16494
rect 365186 9258 365422 9494
rect 365186 2258 365422 2494
rect 365186 -982 365422 -746
rect 365186 -1302 365422 -1066
rect 366918 705962 367154 706198
rect 366918 705642 367154 705878
rect 366918 696198 367154 696434
rect 366918 689198 367154 689434
rect 366918 682198 367154 682434
rect 366918 675198 367154 675434
rect 366918 668198 367154 668434
rect 366918 661198 367154 661434
rect 366918 654198 367154 654434
rect 366918 647198 367154 647434
rect 366918 640198 367154 640434
rect 366918 633198 367154 633434
rect 366918 626198 367154 626434
rect 366918 619198 367154 619434
rect 366918 612198 367154 612434
rect 366918 605198 367154 605434
rect 366918 598198 367154 598434
rect 366918 591198 367154 591434
rect 366918 584198 367154 584434
rect 366918 577198 367154 577434
rect 366918 570198 367154 570434
rect 366918 563198 367154 563434
rect 366918 556198 367154 556434
rect 366918 549198 367154 549434
rect 366918 542198 367154 542434
rect 366918 535198 367154 535434
rect 366918 528198 367154 528434
rect 366918 521198 367154 521434
rect 366918 514198 367154 514434
rect 366918 507198 367154 507434
rect 366918 500198 367154 500434
rect 366918 493198 367154 493434
rect 366918 486198 367154 486434
rect 366918 479198 367154 479434
rect 366918 472198 367154 472434
rect 366918 465198 367154 465434
rect 366918 458198 367154 458434
rect 366918 451198 367154 451434
rect 366918 444198 367154 444434
rect 366918 437198 367154 437434
rect 366918 430198 367154 430434
rect 366918 423198 367154 423434
rect 366918 416198 367154 416434
rect 366918 409198 367154 409434
rect 366918 402198 367154 402434
rect 366918 395198 367154 395434
rect 366918 388198 367154 388434
rect 366918 381198 367154 381434
rect 366918 374198 367154 374434
rect 366918 367198 367154 367434
rect 366918 360198 367154 360434
rect 366918 353198 367154 353434
rect 366918 346198 367154 346434
rect 366918 339198 367154 339434
rect 366918 332198 367154 332434
rect 366918 325198 367154 325434
rect 366918 318198 367154 318434
rect 366918 311198 367154 311434
rect 366918 304198 367154 304434
rect 366918 297198 367154 297434
rect 366918 290198 367154 290434
rect 366918 283198 367154 283434
rect 366918 276198 367154 276434
rect 366918 269198 367154 269434
rect 366918 262198 367154 262434
rect 366918 255198 367154 255434
rect 366918 248198 367154 248434
rect 366918 241198 367154 241434
rect 366918 234198 367154 234434
rect 366918 227198 367154 227434
rect 366918 220198 367154 220434
rect 366918 213198 367154 213434
rect 366918 206198 367154 206434
rect 366918 199198 367154 199434
rect 366918 192198 367154 192434
rect 366918 185198 367154 185434
rect 366918 178198 367154 178434
rect 366918 171198 367154 171434
rect 366918 164198 367154 164434
rect 366918 157198 367154 157434
rect 366918 150198 367154 150434
rect 366918 143198 367154 143434
rect 366918 136198 367154 136434
rect 366918 129198 367154 129434
rect 366918 122198 367154 122434
rect 366918 115198 367154 115434
rect 366918 108198 367154 108434
rect 366918 101198 367154 101434
rect 366918 94198 367154 94434
rect 366918 87198 367154 87434
rect 366918 80198 367154 80434
rect 366918 73198 367154 73434
rect 366918 66198 367154 66434
rect 366918 59198 367154 59434
rect 366918 52198 367154 52434
rect 366918 45198 367154 45434
rect 366918 38198 367154 38434
rect 366918 31198 367154 31434
rect 366918 24198 367154 24434
rect 366918 17198 367154 17434
rect 366918 10198 367154 10434
rect 366918 3198 367154 3434
rect 366918 -1942 367154 -1706
rect 366918 -2262 367154 -2026
rect 372186 705002 372422 705238
rect 372186 704682 372422 704918
rect 372186 695258 372422 695494
rect 372186 688258 372422 688494
rect 372186 681258 372422 681494
rect 372186 674258 372422 674494
rect 372186 667258 372422 667494
rect 372186 660258 372422 660494
rect 372186 653258 372422 653494
rect 372186 646258 372422 646494
rect 372186 639258 372422 639494
rect 372186 632258 372422 632494
rect 372186 625258 372422 625494
rect 372186 618258 372422 618494
rect 372186 611258 372422 611494
rect 372186 604258 372422 604494
rect 372186 597258 372422 597494
rect 372186 590258 372422 590494
rect 372186 583258 372422 583494
rect 372186 576258 372422 576494
rect 372186 569258 372422 569494
rect 372186 562258 372422 562494
rect 372186 555258 372422 555494
rect 372186 548258 372422 548494
rect 372186 541258 372422 541494
rect 372186 534258 372422 534494
rect 372186 527258 372422 527494
rect 372186 520258 372422 520494
rect 372186 513258 372422 513494
rect 372186 506258 372422 506494
rect 372186 499258 372422 499494
rect 372186 492258 372422 492494
rect 372186 485258 372422 485494
rect 372186 478258 372422 478494
rect 372186 471258 372422 471494
rect 372186 464258 372422 464494
rect 372186 457258 372422 457494
rect 372186 450258 372422 450494
rect 372186 443258 372422 443494
rect 372186 436258 372422 436494
rect 372186 429258 372422 429494
rect 372186 422258 372422 422494
rect 372186 415258 372422 415494
rect 372186 408258 372422 408494
rect 372186 401258 372422 401494
rect 372186 394258 372422 394494
rect 372186 387258 372422 387494
rect 372186 380258 372422 380494
rect 372186 373258 372422 373494
rect 372186 366258 372422 366494
rect 372186 359258 372422 359494
rect 372186 352258 372422 352494
rect 372186 345258 372422 345494
rect 372186 338258 372422 338494
rect 372186 331258 372422 331494
rect 372186 324258 372422 324494
rect 372186 317258 372422 317494
rect 372186 310258 372422 310494
rect 372186 303258 372422 303494
rect 372186 296258 372422 296494
rect 372186 289258 372422 289494
rect 372186 282258 372422 282494
rect 372186 275258 372422 275494
rect 372186 268258 372422 268494
rect 372186 261258 372422 261494
rect 372186 254258 372422 254494
rect 372186 247258 372422 247494
rect 372186 240258 372422 240494
rect 372186 233258 372422 233494
rect 372186 226258 372422 226494
rect 372186 219258 372422 219494
rect 372186 212258 372422 212494
rect 372186 205258 372422 205494
rect 372186 198258 372422 198494
rect 372186 191258 372422 191494
rect 372186 184258 372422 184494
rect 372186 177258 372422 177494
rect 372186 170258 372422 170494
rect 372186 163258 372422 163494
rect 372186 156258 372422 156494
rect 372186 149258 372422 149494
rect 372186 142258 372422 142494
rect 372186 135258 372422 135494
rect 372186 128258 372422 128494
rect 372186 121258 372422 121494
rect 372186 114258 372422 114494
rect 372186 107258 372422 107494
rect 372186 100258 372422 100494
rect 372186 93258 372422 93494
rect 372186 86258 372422 86494
rect 372186 79258 372422 79494
rect 372186 72258 372422 72494
rect 372186 65258 372422 65494
rect 372186 58258 372422 58494
rect 372186 51258 372422 51494
rect 372186 44258 372422 44494
rect 372186 37258 372422 37494
rect 372186 30258 372422 30494
rect 372186 23258 372422 23494
rect 372186 16258 372422 16494
rect 372186 9258 372422 9494
rect 372186 2258 372422 2494
rect 372186 -982 372422 -746
rect 372186 -1302 372422 -1066
rect 373918 705962 374154 706198
rect 373918 705642 374154 705878
rect 373918 696198 374154 696434
rect 373918 689198 374154 689434
rect 373918 682198 374154 682434
rect 373918 675198 374154 675434
rect 373918 668198 374154 668434
rect 373918 661198 374154 661434
rect 373918 654198 374154 654434
rect 373918 647198 374154 647434
rect 373918 640198 374154 640434
rect 373918 633198 374154 633434
rect 373918 626198 374154 626434
rect 373918 619198 374154 619434
rect 373918 612198 374154 612434
rect 373918 605198 374154 605434
rect 373918 598198 374154 598434
rect 373918 591198 374154 591434
rect 373918 584198 374154 584434
rect 373918 577198 374154 577434
rect 373918 570198 374154 570434
rect 373918 563198 374154 563434
rect 373918 556198 374154 556434
rect 373918 549198 374154 549434
rect 373918 542198 374154 542434
rect 373918 535198 374154 535434
rect 373918 528198 374154 528434
rect 373918 521198 374154 521434
rect 373918 514198 374154 514434
rect 373918 507198 374154 507434
rect 373918 500198 374154 500434
rect 373918 493198 374154 493434
rect 373918 486198 374154 486434
rect 373918 479198 374154 479434
rect 373918 472198 374154 472434
rect 373918 465198 374154 465434
rect 373918 458198 374154 458434
rect 373918 451198 374154 451434
rect 373918 444198 374154 444434
rect 373918 437198 374154 437434
rect 373918 430198 374154 430434
rect 373918 423198 374154 423434
rect 373918 416198 374154 416434
rect 373918 409198 374154 409434
rect 373918 402198 374154 402434
rect 373918 395198 374154 395434
rect 373918 388198 374154 388434
rect 373918 381198 374154 381434
rect 373918 374198 374154 374434
rect 373918 367198 374154 367434
rect 373918 360198 374154 360434
rect 373918 353198 374154 353434
rect 373918 346198 374154 346434
rect 373918 339198 374154 339434
rect 373918 332198 374154 332434
rect 373918 325198 374154 325434
rect 373918 318198 374154 318434
rect 373918 311198 374154 311434
rect 373918 304198 374154 304434
rect 373918 297198 374154 297434
rect 373918 290198 374154 290434
rect 373918 283198 374154 283434
rect 373918 276198 374154 276434
rect 373918 269198 374154 269434
rect 373918 262198 374154 262434
rect 373918 255198 374154 255434
rect 373918 248198 374154 248434
rect 373918 241198 374154 241434
rect 373918 234198 374154 234434
rect 373918 227198 374154 227434
rect 373918 220198 374154 220434
rect 373918 213198 374154 213434
rect 373918 206198 374154 206434
rect 373918 199198 374154 199434
rect 373918 192198 374154 192434
rect 373918 185198 374154 185434
rect 373918 178198 374154 178434
rect 373918 171198 374154 171434
rect 373918 164198 374154 164434
rect 373918 157198 374154 157434
rect 373918 150198 374154 150434
rect 373918 143198 374154 143434
rect 373918 136198 374154 136434
rect 373918 129198 374154 129434
rect 373918 122198 374154 122434
rect 373918 115198 374154 115434
rect 373918 108198 374154 108434
rect 373918 101198 374154 101434
rect 373918 94198 374154 94434
rect 373918 87198 374154 87434
rect 373918 80198 374154 80434
rect 373918 73198 374154 73434
rect 373918 66198 374154 66434
rect 373918 59198 374154 59434
rect 373918 52198 374154 52434
rect 373918 45198 374154 45434
rect 373918 38198 374154 38434
rect 373918 31198 374154 31434
rect 373918 24198 374154 24434
rect 373918 17198 374154 17434
rect 373918 10198 374154 10434
rect 373918 3198 374154 3434
rect 373918 -1942 374154 -1706
rect 373918 -2262 374154 -2026
rect 379186 705002 379422 705238
rect 379186 704682 379422 704918
rect 379186 695258 379422 695494
rect 379186 688258 379422 688494
rect 379186 681258 379422 681494
rect 379186 674258 379422 674494
rect 379186 667258 379422 667494
rect 379186 660258 379422 660494
rect 379186 653258 379422 653494
rect 379186 646258 379422 646494
rect 379186 639258 379422 639494
rect 379186 632258 379422 632494
rect 379186 625258 379422 625494
rect 379186 618258 379422 618494
rect 379186 611258 379422 611494
rect 379186 604258 379422 604494
rect 379186 597258 379422 597494
rect 379186 590258 379422 590494
rect 379186 583258 379422 583494
rect 379186 576258 379422 576494
rect 379186 569258 379422 569494
rect 379186 562258 379422 562494
rect 379186 555258 379422 555494
rect 379186 548258 379422 548494
rect 379186 541258 379422 541494
rect 379186 534258 379422 534494
rect 379186 527258 379422 527494
rect 379186 520258 379422 520494
rect 379186 513258 379422 513494
rect 379186 506258 379422 506494
rect 379186 499258 379422 499494
rect 379186 492258 379422 492494
rect 379186 485258 379422 485494
rect 379186 478258 379422 478494
rect 379186 471258 379422 471494
rect 379186 464258 379422 464494
rect 379186 457258 379422 457494
rect 379186 450258 379422 450494
rect 379186 443258 379422 443494
rect 379186 436258 379422 436494
rect 379186 429258 379422 429494
rect 379186 422258 379422 422494
rect 379186 415258 379422 415494
rect 379186 408258 379422 408494
rect 379186 401258 379422 401494
rect 379186 394258 379422 394494
rect 379186 387258 379422 387494
rect 379186 380258 379422 380494
rect 379186 373258 379422 373494
rect 379186 366258 379422 366494
rect 379186 359258 379422 359494
rect 379186 352258 379422 352494
rect 379186 345258 379422 345494
rect 379186 338258 379422 338494
rect 379186 331258 379422 331494
rect 379186 324258 379422 324494
rect 379186 317258 379422 317494
rect 379186 310258 379422 310494
rect 379186 303258 379422 303494
rect 379186 296258 379422 296494
rect 379186 289258 379422 289494
rect 379186 282258 379422 282494
rect 379186 275258 379422 275494
rect 379186 268258 379422 268494
rect 379186 261258 379422 261494
rect 379186 254258 379422 254494
rect 379186 247258 379422 247494
rect 379186 240258 379422 240494
rect 379186 233258 379422 233494
rect 379186 226258 379422 226494
rect 379186 219258 379422 219494
rect 379186 212258 379422 212494
rect 379186 205258 379422 205494
rect 379186 198258 379422 198494
rect 379186 191258 379422 191494
rect 379186 184258 379422 184494
rect 379186 177258 379422 177494
rect 379186 170258 379422 170494
rect 379186 163258 379422 163494
rect 379186 156258 379422 156494
rect 379186 149258 379422 149494
rect 379186 142258 379422 142494
rect 379186 135258 379422 135494
rect 379186 128258 379422 128494
rect 379186 121258 379422 121494
rect 379186 114258 379422 114494
rect 379186 107258 379422 107494
rect 379186 100258 379422 100494
rect 379186 93258 379422 93494
rect 379186 86258 379422 86494
rect 379186 79258 379422 79494
rect 379186 72258 379422 72494
rect 379186 65258 379422 65494
rect 379186 58258 379422 58494
rect 379186 51258 379422 51494
rect 379186 44258 379422 44494
rect 379186 37258 379422 37494
rect 379186 30258 379422 30494
rect 379186 23258 379422 23494
rect 379186 16258 379422 16494
rect 379186 9258 379422 9494
rect 379186 2258 379422 2494
rect 379186 -982 379422 -746
rect 379186 -1302 379422 -1066
rect 380918 705962 381154 706198
rect 380918 705642 381154 705878
rect 380918 696198 381154 696434
rect 380918 689198 381154 689434
rect 380918 682198 381154 682434
rect 380918 675198 381154 675434
rect 380918 668198 381154 668434
rect 380918 661198 381154 661434
rect 380918 654198 381154 654434
rect 380918 647198 381154 647434
rect 380918 640198 381154 640434
rect 380918 633198 381154 633434
rect 380918 626198 381154 626434
rect 380918 619198 381154 619434
rect 380918 612198 381154 612434
rect 380918 605198 381154 605434
rect 380918 598198 381154 598434
rect 380918 591198 381154 591434
rect 380918 584198 381154 584434
rect 380918 577198 381154 577434
rect 380918 570198 381154 570434
rect 380918 563198 381154 563434
rect 380918 556198 381154 556434
rect 380918 549198 381154 549434
rect 380918 542198 381154 542434
rect 380918 535198 381154 535434
rect 380918 528198 381154 528434
rect 380918 521198 381154 521434
rect 380918 514198 381154 514434
rect 380918 507198 381154 507434
rect 380918 500198 381154 500434
rect 380918 493198 381154 493434
rect 380918 486198 381154 486434
rect 380918 479198 381154 479434
rect 380918 472198 381154 472434
rect 380918 465198 381154 465434
rect 380918 458198 381154 458434
rect 380918 451198 381154 451434
rect 380918 444198 381154 444434
rect 380918 437198 381154 437434
rect 380918 430198 381154 430434
rect 380918 423198 381154 423434
rect 380918 416198 381154 416434
rect 380918 409198 381154 409434
rect 380918 402198 381154 402434
rect 380918 395198 381154 395434
rect 380918 388198 381154 388434
rect 380918 381198 381154 381434
rect 380918 374198 381154 374434
rect 380918 367198 381154 367434
rect 380918 360198 381154 360434
rect 380918 353198 381154 353434
rect 380918 346198 381154 346434
rect 380918 339198 381154 339434
rect 380918 332198 381154 332434
rect 380918 325198 381154 325434
rect 380918 318198 381154 318434
rect 380918 311198 381154 311434
rect 380918 304198 381154 304434
rect 380918 297198 381154 297434
rect 380918 290198 381154 290434
rect 380918 283198 381154 283434
rect 380918 276198 381154 276434
rect 380918 269198 381154 269434
rect 380918 262198 381154 262434
rect 380918 255198 381154 255434
rect 380918 248198 381154 248434
rect 380918 241198 381154 241434
rect 380918 234198 381154 234434
rect 380918 227198 381154 227434
rect 380918 220198 381154 220434
rect 380918 213198 381154 213434
rect 380918 206198 381154 206434
rect 380918 199198 381154 199434
rect 380918 192198 381154 192434
rect 380918 185198 381154 185434
rect 380918 178198 381154 178434
rect 380918 171198 381154 171434
rect 380918 164198 381154 164434
rect 380918 157198 381154 157434
rect 380918 150198 381154 150434
rect 380918 143198 381154 143434
rect 380918 136198 381154 136434
rect 380918 129198 381154 129434
rect 380918 122198 381154 122434
rect 380918 115198 381154 115434
rect 380918 108198 381154 108434
rect 380918 101198 381154 101434
rect 380918 94198 381154 94434
rect 380918 87198 381154 87434
rect 380918 80198 381154 80434
rect 380918 73198 381154 73434
rect 380918 66198 381154 66434
rect 380918 59198 381154 59434
rect 380918 52198 381154 52434
rect 380918 45198 381154 45434
rect 380918 38198 381154 38434
rect 380918 31198 381154 31434
rect 380918 24198 381154 24434
rect 380918 17198 381154 17434
rect 380918 10198 381154 10434
rect 380918 3198 381154 3434
rect 380918 -1942 381154 -1706
rect 380918 -2262 381154 -2026
rect 386186 705002 386422 705238
rect 386186 704682 386422 704918
rect 386186 695258 386422 695494
rect 386186 688258 386422 688494
rect 386186 681258 386422 681494
rect 386186 674258 386422 674494
rect 386186 667258 386422 667494
rect 386186 660258 386422 660494
rect 386186 653258 386422 653494
rect 386186 646258 386422 646494
rect 386186 639258 386422 639494
rect 386186 632258 386422 632494
rect 386186 625258 386422 625494
rect 386186 618258 386422 618494
rect 386186 611258 386422 611494
rect 386186 604258 386422 604494
rect 386186 597258 386422 597494
rect 386186 590258 386422 590494
rect 386186 583258 386422 583494
rect 386186 576258 386422 576494
rect 386186 569258 386422 569494
rect 386186 562258 386422 562494
rect 386186 555258 386422 555494
rect 386186 548258 386422 548494
rect 386186 541258 386422 541494
rect 386186 534258 386422 534494
rect 386186 527258 386422 527494
rect 386186 520258 386422 520494
rect 386186 513258 386422 513494
rect 386186 506258 386422 506494
rect 386186 499258 386422 499494
rect 386186 492258 386422 492494
rect 386186 485258 386422 485494
rect 386186 478258 386422 478494
rect 386186 471258 386422 471494
rect 386186 464258 386422 464494
rect 386186 457258 386422 457494
rect 386186 450258 386422 450494
rect 386186 443258 386422 443494
rect 386186 436258 386422 436494
rect 386186 429258 386422 429494
rect 386186 422258 386422 422494
rect 386186 415258 386422 415494
rect 386186 408258 386422 408494
rect 386186 401258 386422 401494
rect 386186 394258 386422 394494
rect 386186 387258 386422 387494
rect 386186 380258 386422 380494
rect 386186 373258 386422 373494
rect 386186 366258 386422 366494
rect 386186 359258 386422 359494
rect 386186 352258 386422 352494
rect 386186 345258 386422 345494
rect 386186 338258 386422 338494
rect 386186 331258 386422 331494
rect 386186 324258 386422 324494
rect 386186 317258 386422 317494
rect 386186 310258 386422 310494
rect 386186 303258 386422 303494
rect 386186 296258 386422 296494
rect 386186 289258 386422 289494
rect 386186 282258 386422 282494
rect 386186 275258 386422 275494
rect 386186 268258 386422 268494
rect 386186 261258 386422 261494
rect 386186 254258 386422 254494
rect 386186 247258 386422 247494
rect 386186 240258 386422 240494
rect 386186 233258 386422 233494
rect 386186 226258 386422 226494
rect 386186 219258 386422 219494
rect 386186 212258 386422 212494
rect 386186 205258 386422 205494
rect 386186 198258 386422 198494
rect 386186 191258 386422 191494
rect 386186 184258 386422 184494
rect 386186 177258 386422 177494
rect 386186 170258 386422 170494
rect 386186 163258 386422 163494
rect 386186 156258 386422 156494
rect 386186 149258 386422 149494
rect 386186 142258 386422 142494
rect 386186 135258 386422 135494
rect 386186 128258 386422 128494
rect 386186 121258 386422 121494
rect 386186 114258 386422 114494
rect 386186 107258 386422 107494
rect 386186 100258 386422 100494
rect 386186 93258 386422 93494
rect 386186 86258 386422 86494
rect 386186 79258 386422 79494
rect 386186 72258 386422 72494
rect 386186 65258 386422 65494
rect 386186 58258 386422 58494
rect 386186 51258 386422 51494
rect 386186 44258 386422 44494
rect 386186 37258 386422 37494
rect 386186 30258 386422 30494
rect 386186 23258 386422 23494
rect 386186 16258 386422 16494
rect 386186 9258 386422 9494
rect 386186 2258 386422 2494
rect 386186 -982 386422 -746
rect 386186 -1302 386422 -1066
rect 387918 705962 388154 706198
rect 387918 705642 388154 705878
rect 387918 696198 388154 696434
rect 387918 689198 388154 689434
rect 387918 682198 388154 682434
rect 387918 675198 388154 675434
rect 387918 668198 388154 668434
rect 387918 661198 388154 661434
rect 387918 654198 388154 654434
rect 387918 647198 388154 647434
rect 387918 640198 388154 640434
rect 387918 633198 388154 633434
rect 387918 626198 388154 626434
rect 387918 619198 388154 619434
rect 387918 612198 388154 612434
rect 387918 605198 388154 605434
rect 387918 598198 388154 598434
rect 387918 591198 388154 591434
rect 387918 584198 388154 584434
rect 387918 577198 388154 577434
rect 387918 570198 388154 570434
rect 387918 563198 388154 563434
rect 387918 556198 388154 556434
rect 387918 549198 388154 549434
rect 387918 542198 388154 542434
rect 387918 535198 388154 535434
rect 387918 528198 388154 528434
rect 387918 521198 388154 521434
rect 387918 514198 388154 514434
rect 387918 507198 388154 507434
rect 387918 500198 388154 500434
rect 387918 493198 388154 493434
rect 387918 486198 388154 486434
rect 387918 479198 388154 479434
rect 387918 472198 388154 472434
rect 387918 465198 388154 465434
rect 387918 458198 388154 458434
rect 387918 451198 388154 451434
rect 387918 444198 388154 444434
rect 387918 437198 388154 437434
rect 387918 430198 388154 430434
rect 387918 423198 388154 423434
rect 387918 416198 388154 416434
rect 387918 409198 388154 409434
rect 387918 402198 388154 402434
rect 387918 395198 388154 395434
rect 387918 388198 388154 388434
rect 387918 381198 388154 381434
rect 387918 374198 388154 374434
rect 387918 367198 388154 367434
rect 387918 360198 388154 360434
rect 387918 353198 388154 353434
rect 387918 346198 388154 346434
rect 387918 339198 388154 339434
rect 387918 332198 388154 332434
rect 387918 325198 388154 325434
rect 387918 318198 388154 318434
rect 387918 311198 388154 311434
rect 387918 304198 388154 304434
rect 387918 297198 388154 297434
rect 387918 290198 388154 290434
rect 387918 283198 388154 283434
rect 387918 276198 388154 276434
rect 387918 269198 388154 269434
rect 387918 262198 388154 262434
rect 387918 255198 388154 255434
rect 387918 248198 388154 248434
rect 387918 241198 388154 241434
rect 387918 234198 388154 234434
rect 387918 227198 388154 227434
rect 387918 220198 388154 220434
rect 387918 213198 388154 213434
rect 387918 206198 388154 206434
rect 387918 199198 388154 199434
rect 387918 192198 388154 192434
rect 387918 185198 388154 185434
rect 387918 178198 388154 178434
rect 387918 171198 388154 171434
rect 387918 164198 388154 164434
rect 387918 157198 388154 157434
rect 387918 150198 388154 150434
rect 387918 143198 388154 143434
rect 387918 136198 388154 136434
rect 387918 129198 388154 129434
rect 387918 122198 388154 122434
rect 387918 115198 388154 115434
rect 387918 108198 388154 108434
rect 387918 101198 388154 101434
rect 387918 94198 388154 94434
rect 387918 87198 388154 87434
rect 387918 80198 388154 80434
rect 387918 73198 388154 73434
rect 387918 66198 388154 66434
rect 387918 59198 388154 59434
rect 387918 52198 388154 52434
rect 387918 45198 388154 45434
rect 387918 38198 388154 38434
rect 387918 31198 388154 31434
rect 387918 24198 388154 24434
rect 387918 17198 388154 17434
rect 387918 10198 388154 10434
rect 387918 3198 388154 3434
rect 387918 -1942 388154 -1706
rect 387918 -2262 388154 -2026
rect 393186 705002 393422 705238
rect 393186 704682 393422 704918
rect 393186 695258 393422 695494
rect 393186 688258 393422 688494
rect 393186 681258 393422 681494
rect 393186 674258 393422 674494
rect 393186 667258 393422 667494
rect 393186 660258 393422 660494
rect 393186 653258 393422 653494
rect 393186 646258 393422 646494
rect 393186 639258 393422 639494
rect 393186 632258 393422 632494
rect 393186 625258 393422 625494
rect 393186 618258 393422 618494
rect 393186 611258 393422 611494
rect 393186 604258 393422 604494
rect 393186 597258 393422 597494
rect 393186 590258 393422 590494
rect 393186 583258 393422 583494
rect 393186 576258 393422 576494
rect 393186 569258 393422 569494
rect 393186 562258 393422 562494
rect 393186 555258 393422 555494
rect 393186 548258 393422 548494
rect 393186 541258 393422 541494
rect 393186 534258 393422 534494
rect 393186 527258 393422 527494
rect 393186 520258 393422 520494
rect 393186 513258 393422 513494
rect 393186 506258 393422 506494
rect 393186 499258 393422 499494
rect 393186 492258 393422 492494
rect 393186 485258 393422 485494
rect 393186 478258 393422 478494
rect 393186 471258 393422 471494
rect 393186 464258 393422 464494
rect 393186 457258 393422 457494
rect 393186 450258 393422 450494
rect 393186 443258 393422 443494
rect 393186 436258 393422 436494
rect 393186 429258 393422 429494
rect 393186 422258 393422 422494
rect 393186 415258 393422 415494
rect 393186 408258 393422 408494
rect 393186 401258 393422 401494
rect 393186 394258 393422 394494
rect 393186 387258 393422 387494
rect 393186 380258 393422 380494
rect 393186 373258 393422 373494
rect 393186 366258 393422 366494
rect 393186 359258 393422 359494
rect 393186 352258 393422 352494
rect 393186 345258 393422 345494
rect 393186 338258 393422 338494
rect 393186 331258 393422 331494
rect 393186 324258 393422 324494
rect 393186 317258 393422 317494
rect 393186 310258 393422 310494
rect 393186 303258 393422 303494
rect 393186 296258 393422 296494
rect 393186 289258 393422 289494
rect 393186 282258 393422 282494
rect 393186 275258 393422 275494
rect 393186 268258 393422 268494
rect 393186 261258 393422 261494
rect 393186 254258 393422 254494
rect 393186 247258 393422 247494
rect 393186 240258 393422 240494
rect 393186 233258 393422 233494
rect 393186 226258 393422 226494
rect 393186 219258 393422 219494
rect 393186 212258 393422 212494
rect 393186 205258 393422 205494
rect 393186 198258 393422 198494
rect 393186 191258 393422 191494
rect 393186 184258 393422 184494
rect 393186 177258 393422 177494
rect 393186 170258 393422 170494
rect 393186 163258 393422 163494
rect 393186 156258 393422 156494
rect 393186 149258 393422 149494
rect 393186 142258 393422 142494
rect 393186 135258 393422 135494
rect 393186 128258 393422 128494
rect 393186 121258 393422 121494
rect 393186 114258 393422 114494
rect 393186 107258 393422 107494
rect 393186 100258 393422 100494
rect 393186 93258 393422 93494
rect 393186 86258 393422 86494
rect 393186 79258 393422 79494
rect 393186 72258 393422 72494
rect 393186 65258 393422 65494
rect 393186 58258 393422 58494
rect 393186 51258 393422 51494
rect 393186 44258 393422 44494
rect 393186 37258 393422 37494
rect 393186 30258 393422 30494
rect 393186 23258 393422 23494
rect 393186 16258 393422 16494
rect 393186 9258 393422 9494
rect 393186 2258 393422 2494
rect 393186 -982 393422 -746
rect 393186 -1302 393422 -1066
rect 394918 705962 395154 706198
rect 394918 705642 395154 705878
rect 394918 696198 395154 696434
rect 394918 689198 395154 689434
rect 394918 682198 395154 682434
rect 394918 675198 395154 675434
rect 394918 668198 395154 668434
rect 394918 661198 395154 661434
rect 394918 654198 395154 654434
rect 394918 647198 395154 647434
rect 394918 640198 395154 640434
rect 394918 633198 395154 633434
rect 394918 626198 395154 626434
rect 394918 619198 395154 619434
rect 394918 612198 395154 612434
rect 394918 605198 395154 605434
rect 394918 598198 395154 598434
rect 394918 591198 395154 591434
rect 394918 584198 395154 584434
rect 394918 577198 395154 577434
rect 394918 570198 395154 570434
rect 394918 563198 395154 563434
rect 394918 556198 395154 556434
rect 394918 549198 395154 549434
rect 394918 542198 395154 542434
rect 394918 535198 395154 535434
rect 394918 528198 395154 528434
rect 394918 521198 395154 521434
rect 394918 514198 395154 514434
rect 394918 507198 395154 507434
rect 394918 500198 395154 500434
rect 394918 493198 395154 493434
rect 394918 486198 395154 486434
rect 394918 479198 395154 479434
rect 394918 472198 395154 472434
rect 394918 465198 395154 465434
rect 394918 458198 395154 458434
rect 394918 451198 395154 451434
rect 394918 444198 395154 444434
rect 394918 437198 395154 437434
rect 394918 430198 395154 430434
rect 394918 423198 395154 423434
rect 394918 416198 395154 416434
rect 394918 409198 395154 409434
rect 394918 402198 395154 402434
rect 394918 395198 395154 395434
rect 394918 388198 395154 388434
rect 394918 381198 395154 381434
rect 394918 374198 395154 374434
rect 394918 367198 395154 367434
rect 394918 360198 395154 360434
rect 394918 353198 395154 353434
rect 394918 346198 395154 346434
rect 394918 339198 395154 339434
rect 394918 332198 395154 332434
rect 394918 325198 395154 325434
rect 394918 318198 395154 318434
rect 394918 311198 395154 311434
rect 394918 304198 395154 304434
rect 394918 297198 395154 297434
rect 394918 290198 395154 290434
rect 394918 283198 395154 283434
rect 394918 276198 395154 276434
rect 394918 269198 395154 269434
rect 394918 262198 395154 262434
rect 394918 255198 395154 255434
rect 394918 248198 395154 248434
rect 394918 241198 395154 241434
rect 394918 234198 395154 234434
rect 394918 227198 395154 227434
rect 394918 220198 395154 220434
rect 394918 213198 395154 213434
rect 394918 206198 395154 206434
rect 394918 199198 395154 199434
rect 394918 192198 395154 192434
rect 394918 185198 395154 185434
rect 394918 178198 395154 178434
rect 394918 171198 395154 171434
rect 394918 164198 395154 164434
rect 394918 157198 395154 157434
rect 394918 150198 395154 150434
rect 394918 143198 395154 143434
rect 394918 136198 395154 136434
rect 394918 129198 395154 129434
rect 394918 122198 395154 122434
rect 394918 115198 395154 115434
rect 394918 108198 395154 108434
rect 394918 101198 395154 101434
rect 394918 94198 395154 94434
rect 394918 87198 395154 87434
rect 394918 80198 395154 80434
rect 394918 73198 395154 73434
rect 394918 66198 395154 66434
rect 394918 59198 395154 59434
rect 394918 52198 395154 52434
rect 394918 45198 395154 45434
rect 394918 38198 395154 38434
rect 394918 31198 395154 31434
rect 394918 24198 395154 24434
rect 394918 17198 395154 17434
rect 394918 10198 395154 10434
rect 394918 3198 395154 3434
rect 394918 -1942 395154 -1706
rect 394918 -2262 395154 -2026
rect 400186 705002 400422 705238
rect 400186 704682 400422 704918
rect 400186 695258 400422 695494
rect 400186 688258 400422 688494
rect 400186 681258 400422 681494
rect 400186 674258 400422 674494
rect 400186 667258 400422 667494
rect 400186 660258 400422 660494
rect 400186 653258 400422 653494
rect 400186 646258 400422 646494
rect 400186 639258 400422 639494
rect 400186 632258 400422 632494
rect 400186 625258 400422 625494
rect 400186 618258 400422 618494
rect 400186 611258 400422 611494
rect 400186 604258 400422 604494
rect 400186 597258 400422 597494
rect 400186 590258 400422 590494
rect 400186 583258 400422 583494
rect 400186 576258 400422 576494
rect 400186 569258 400422 569494
rect 400186 562258 400422 562494
rect 400186 555258 400422 555494
rect 400186 548258 400422 548494
rect 400186 541258 400422 541494
rect 400186 534258 400422 534494
rect 400186 527258 400422 527494
rect 400186 520258 400422 520494
rect 400186 513258 400422 513494
rect 400186 506258 400422 506494
rect 400186 499258 400422 499494
rect 400186 492258 400422 492494
rect 400186 485258 400422 485494
rect 400186 478258 400422 478494
rect 400186 471258 400422 471494
rect 400186 464258 400422 464494
rect 400186 457258 400422 457494
rect 400186 450258 400422 450494
rect 400186 443258 400422 443494
rect 400186 436258 400422 436494
rect 400186 429258 400422 429494
rect 400186 422258 400422 422494
rect 400186 415258 400422 415494
rect 400186 408258 400422 408494
rect 400186 401258 400422 401494
rect 400186 394258 400422 394494
rect 400186 387258 400422 387494
rect 400186 380258 400422 380494
rect 400186 373258 400422 373494
rect 400186 366258 400422 366494
rect 400186 359258 400422 359494
rect 400186 352258 400422 352494
rect 400186 345258 400422 345494
rect 400186 338258 400422 338494
rect 400186 331258 400422 331494
rect 400186 324258 400422 324494
rect 400186 317258 400422 317494
rect 400186 310258 400422 310494
rect 400186 303258 400422 303494
rect 400186 296258 400422 296494
rect 400186 289258 400422 289494
rect 400186 282258 400422 282494
rect 400186 275258 400422 275494
rect 400186 268258 400422 268494
rect 400186 261258 400422 261494
rect 400186 254258 400422 254494
rect 400186 247258 400422 247494
rect 400186 240258 400422 240494
rect 400186 233258 400422 233494
rect 400186 226258 400422 226494
rect 400186 219258 400422 219494
rect 400186 212258 400422 212494
rect 400186 205258 400422 205494
rect 400186 198258 400422 198494
rect 400186 191258 400422 191494
rect 400186 184258 400422 184494
rect 400186 177258 400422 177494
rect 400186 170258 400422 170494
rect 400186 163258 400422 163494
rect 400186 156258 400422 156494
rect 400186 149258 400422 149494
rect 400186 142258 400422 142494
rect 400186 135258 400422 135494
rect 400186 128258 400422 128494
rect 400186 121258 400422 121494
rect 400186 114258 400422 114494
rect 400186 107258 400422 107494
rect 400186 100258 400422 100494
rect 400186 93258 400422 93494
rect 400186 86258 400422 86494
rect 400186 79258 400422 79494
rect 400186 72258 400422 72494
rect 400186 65258 400422 65494
rect 400186 58258 400422 58494
rect 400186 51258 400422 51494
rect 400186 44258 400422 44494
rect 400186 37258 400422 37494
rect 400186 30258 400422 30494
rect 400186 23258 400422 23494
rect 400186 16258 400422 16494
rect 400186 9258 400422 9494
rect 400186 2258 400422 2494
rect 400186 -982 400422 -746
rect 400186 -1302 400422 -1066
rect 401918 705962 402154 706198
rect 401918 705642 402154 705878
rect 401918 696198 402154 696434
rect 401918 689198 402154 689434
rect 401918 682198 402154 682434
rect 401918 675198 402154 675434
rect 401918 668198 402154 668434
rect 401918 661198 402154 661434
rect 401918 654198 402154 654434
rect 401918 647198 402154 647434
rect 401918 640198 402154 640434
rect 401918 633198 402154 633434
rect 401918 626198 402154 626434
rect 401918 619198 402154 619434
rect 401918 612198 402154 612434
rect 401918 605198 402154 605434
rect 401918 598198 402154 598434
rect 401918 591198 402154 591434
rect 401918 584198 402154 584434
rect 401918 577198 402154 577434
rect 401918 570198 402154 570434
rect 401918 563198 402154 563434
rect 401918 556198 402154 556434
rect 401918 549198 402154 549434
rect 401918 542198 402154 542434
rect 401918 535198 402154 535434
rect 401918 528198 402154 528434
rect 401918 521198 402154 521434
rect 401918 514198 402154 514434
rect 401918 507198 402154 507434
rect 401918 500198 402154 500434
rect 401918 493198 402154 493434
rect 401918 486198 402154 486434
rect 401918 479198 402154 479434
rect 401918 472198 402154 472434
rect 401918 465198 402154 465434
rect 401918 458198 402154 458434
rect 401918 451198 402154 451434
rect 401918 444198 402154 444434
rect 401918 437198 402154 437434
rect 401918 430198 402154 430434
rect 401918 423198 402154 423434
rect 401918 416198 402154 416434
rect 401918 409198 402154 409434
rect 401918 402198 402154 402434
rect 401918 395198 402154 395434
rect 401918 388198 402154 388434
rect 401918 381198 402154 381434
rect 401918 374198 402154 374434
rect 401918 367198 402154 367434
rect 401918 360198 402154 360434
rect 401918 353198 402154 353434
rect 401918 346198 402154 346434
rect 401918 339198 402154 339434
rect 401918 332198 402154 332434
rect 401918 325198 402154 325434
rect 401918 318198 402154 318434
rect 401918 311198 402154 311434
rect 401918 304198 402154 304434
rect 401918 297198 402154 297434
rect 401918 290198 402154 290434
rect 401918 283198 402154 283434
rect 401918 276198 402154 276434
rect 401918 269198 402154 269434
rect 401918 262198 402154 262434
rect 401918 255198 402154 255434
rect 401918 248198 402154 248434
rect 401918 241198 402154 241434
rect 401918 234198 402154 234434
rect 401918 227198 402154 227434
rect 401918 220198 402154 220434
rect 401918 213198 402154 213434
rect 401918 206198 402154 206434
rect 401918 199198 402154 199434
rect 401918 192198 402154 192434
rect 401918 185198 402154 185434
rect 401918 178198 402154 178434
rect 401918 171198 402154 171434
rect 401918 164198 402154 164434
rect 401918 157198 402154 157434
rect 401918 150198 402154 150434
rect 401918 143198 402154 143434
rect 401918 136198 402154 136434
rect 401918 129198 402154 129434
rect 401918 122198 402154 122434
rect 401918 115198 402154 115434
rect 401918 108198 402154 108434
rect 401918 101198 402154 101434
rect 401918 94198 402154 94434
rect 401918 87198 402154 87434
rect 401918 80198 402154 80434
rect 401918 73198 402154 73434
rect 401918 66198 402154 66434
rect 401918 59198 402154 59434
rect 401918 52198 402154 52434
rect 401918 45198 402154 45434
rect 401918 38198 402154 38434
rect 401918 31198 402154 31434
rect 401918 24198 402154 24434
rect 401918 17198 402154 17434
rect 401918 10198 402154 10434
rect 401918 3198 402154 3434
rect 401918 -1942 402154 -1706
rect 401918 -2262 402154 -2026
rect 407186 705002 407422 705238
rect 407186 704682 407422 704918
rect 407186 695258 407422 695494
rect 407186 688258 407422 688494
rect 407186 681258 407422 681494
rect 407186 674258 407422 674494
rect 407186 667258 407422 667494
rect 407186 660258 407422 660494
rect 407186 653258 407422 653494
rect 407186 646258 407422 646494
rect 407186 639258 407422 639494
rect 407186 632258 407422 632494
rect 407186 625258 407422 625494
rect 407186 618258 407422 618494
rect 407186 611258 407422 611494
rect 407186 604258 407422 604494
rect 407186 597258 407422 597494
rect 407186 590258 407422 590494
rect 407186 583258 407422 583494
rect 407186 576258 407422 576494
rect 407186 569258 407422 569494
rect 407186 562258 407422 562494
rect 407186 555258 407422 555494
rect 407186 548258 407422 548494
rect 407186 541258 407422 541494
rect 407186 534258 407422 534494
rect 407186 527258 407422 527494
rect 407186 520258 407422 520494
rect 407186 513258 407422 513494
rect 407186 506258 407422 506494
rect 407186 499258 407422 499494
rect 407186 492258 407422 492494
rect 407186 485258 407422 485494
rect 407186 478258 407422 478494
rect 407186 471258 407422 471494
rect 407186 464258 407422 464494
rect 407186 457258 407422 457494
rect 407186 450258 407422 450494
rect 407186 443258 407422 443494
rect 407186 436258 407422 436494
rect 407186 429258 407422 429494
rect 407186 422258 407422 422494
rect 407186 415258 407422 415494
rect 407186 408258 407422 408494
rect 407186 401258 407422 401494
rect 407186 394258 407422 394494
rect 407186 387258 407422 387494
rect 407186 380258 407422 380494
rect 407186 373258 407422 373494
rect 407186 366258 407422 366494
rect 407186 359258 407422 359494
rect 407186 352258 407422 352494
rect 407186 345258 407422 345494
rect 407186 338258 407422 338494
rect 407186 331258 407422 331494
rect 407186 324258 407422 324494
rect 407186 317258 407422 317494
rect 407186 310258 407422 310494
rect 407186 303258 407422 303494
rect 407186 296258 407422 296494
rect 407186 289258 407422 289494
rect 407186 282258 407422 282494
rect 407186 275258 407422 275494
rect 407186 268258 407422 268494
rect 407186 261258 407422 261494
rect 407186 254258 407422 254494
rect 407186 247258 407422 247494
rect 407186 240258 407422 240494
rect 407186 233258 407422 233494
rect 407186 226258 407422 226494
rect 407186 219258 407422 219494
rect 407186 212258 407422 212494
rect 407186 205258 407422 205494
rect 407186 198258 407422 198494
rect 407186 191258 407422 191494
rect 407186 184258 407422 184494
rect 407186 177258 407422 177494
rect 407186 170258 407422 170494
rect 407186 163258 407422 163494
rect 407186 156258 407422 156494
rect 407186 149258 407422 149494
rect 407186 142258 407422 142494
rect 407186 135258 407422 135494
rect 407186 128258 407422 128494
rect 407186 121258 407422 121494
rect 407186 114258 407422 114494
rect 407186 107258 407422 107494
rect 407186 100258 407422 100494
rect 407186 93258 407422 93494
rect 407186 86258 407422 86494
rect 407186 79258 407422 79494
rect 407186 72258 407422 72494
rect 407186 65258 407422 65494
rect 407186 58258 407422 58494
rect 407186 51258 407422 51494
rect 407186 44258 407422 44494
rect 407186 37258 407422 37494
rect 407186 30258 407422 30494
rect 407186 23258 407422 23494
rect 407186 16258 407422 16494
rect 407186 9258 407422 9494
rect 407186 2258 407422 2494
rect 407186 -982 407422 -746
rect 407186 -1302 407422 -1066
rect 408918 705962 409154 706198
rect 408918 705642 409154 705878
rect 408918 696198 409154 696434
rect 408918 689198 409154 689434
rect 408918 682198 409154 682434
rect 408918 675198 409154 675434
rect 408918 668198 409154 668434
rect 408918 661198 409154 661434
rect 408918 654198 409154 654434
rect 408918 647198 409154 647434
rect 408918 640198 409154 640434
rect 408918 633198 409154 633434
rect 408918 626198 409154 626434
rect 408918 619198 409154 619434
rect 408918 612198 409154 612434
rect 408918 605198 409154 605434
rect 408918 598198 409154 598434
rect 408918 591198 409154 591434
rect 408918 584198 409154 584434
rect 408918 577198 409154 577434
rect 408918 570198 409154 570434
rect 408918 563198 409154 563434
rect 408918 556198 409154 556434
rect 408918 549198 409154 549434
rect 408918 542198 409154 542434
rect 408918 535198 409154 535434
rect 408918 528198 409154 528434
rect 408918 521198 409154 521434
rect 408918 514198 409154 514434
rect 408918 507198 409154 507434
rect 408918 500198 409154 500434
rect 408918 493198 409154 493434
rect 408918 486198 409154 486434
rect 408918 479198 409154 479434
rect 408918 472198 409154 472434
rect 408918 465198 409154 465434
rect 408918 458198 409154 458434
rect 408918 451198 409154 451434
rect 408918 444198 409154 444434
rect 408918 437198 409154 437434
rect 408918 430198 409154 430434
rect 408918 423198 409154 423434
rect 408918 416198 409154 416434
rect 408918 409198 409154 409434
rect 408918 402198 409154 402434
rect 408918 395198 409154 395434
rect 408918 388198 409154 388434
rect 408918 381198 409154 381434
rect 408918 374198 409154 374434
rect 408918 367198 409154 367434
rect 408918 360198 409154 360434
rect 408918 353198 409154 353434
rect 408918 346198 409154 346434
rect 408918 339198 409154 339434
rect 408918 332198 409154 332434
rect 408918 325198 409154 325434
rect 408918 318198 409154 318434
rect 408918 311198 409154 311434
rect 408918 304198 409154 304434
rect 408918 297198 409154 297434
rect 408918 290198 409154 290434
rect 408918 283198 409154 283434
rect 408918 276198 409154 276434
rect 408918 269198 409154 269434
rect 408918 262198 409154 262434
rect 408918 255198 409154 255434
rect 408918 248198 409154 248434
rect 408918 241198 409154 241434
rect 408918 234198 409154 234434
rect 408918 227198 409154 227434
rect 408918 220198 409154 220434
rect 408918 213198 409154 213434
rect 408918 206198 409154 206434
rect 408918 199198 409154 199434
rect 408918 192198 409154 192434
rect 408918 185198 409154 185434
rect 408918 178198 409154 178434
rect 408918 171198 409154 171434
rect 408918 164198 409154 164434
rect 408918 157198 409154 157434
rect 408918 150198 409154 150434
rect 408918 143198 409154 143434
rect 408918 136198 409154 136434
rect 408918 129198 409154 129434
rect 408918 122198 409154 122434
rect 408918 115198 409154 115434
rect 408918 108198 409154 108434
rect 408918 101198 409154 101434
rect 408918 94198 409154 94434
rect 408918 87198 409154 87434
rect 408918 80198 409154 80434
rect 408918 73198 409154 73434
rect 408918 66198 409154 66434
rect 408918 59198 409154 59434
rect 408918 52198 409154 52434
rect 408918 45198 409154 45434
rect 408918 38198 409154 38434
rect 408918 31198 409154 31434
rect 408918 24198 409154 24434
rect 408918 17198 409154 17434
rect 408918 10198 409154 10434
rect 408918 3198 409154 3434
rect 408918 -1942 409154 -1706
rect 408918 -2262 409154 -2026
rect 414186 705002 414422 705238
rect 414186 704682 414422 704918
rect 414186 695258 414422 695494
rect 414186 688258 414422 688494
rect 414186 681258 414422 681494
rect 414186 674258 414422 674494
rect 414186 667258 414422 667494
rect 414186 660258 414422 660494
rect 414186 653258 414422 653494
rect 414186 646258 414422 646494
rect 414186 639258 414422 639494
rect 414186 632258 414422 632494
rect 414186 625258 414422 625494
rect 414186 618258 414422 618494
rect 414186 611258 414422 611494
rect 414186 604258 414422 604494
rect 414186 597258 414422 597494
rect 414186 590258 414422 590494
rect 414186 583258 414422 583494
rect 414186 576258 414422 576494
rect 414186 569258 414422 569494
rect 414186 562258 414422 562494
rect 414186 555258 414422 555494
rect 414186 548258 414422 548494
rect 414186 541258 414422 541494
rect 414186 534258 414422 534494
rect 414186 527258 414422 527494
rect 414186 520258 414422 520494
rect 414186 513258 414422 513494
rect 414186 506258 414422 506494
rect 414186 499258 414422 499494
rect 414186 492258 414422 492494
rect 414186 485258 414422 485494
rect 414186 478258 414422 478494
rect 414186 471258 414422 471494
rect 414186 464258 414422 464494
rect 414186 457258 414422 457494
rect 414186 450258 414422 450494
rect 414186 443258 414422 443494
rect 414186 436258 414422 436494
rect 414186 429258 414422 429494
rect 414186 422258 414422 422494
rect 414186 415258 414422 415494
rect 414186 408258 414422 408494
rect 414186 401258 414422 401494
rect 414186 394258 414422 394494
rect 414186 387258 414422 387494
rect 414186 380258 414422 380494
rect 414186 373258 414422 373494
rect 414186 366258 414422 366494
rect 414186 359258 414422 359494
rect 414186 352258 414422 352494
rect 414186 345258 414422 345494
rect 414186 338258 414422 338494
rect 414186 331258 414422 331494
rect 414186 324258 414422 324494
rect 414186 317258 414422 317494
rect 414186 310258 414422 310494
rect 414186 303258 414422 303494
rect 414186 296258 414422 296494
rect 414186 289258 414422 289494
rect 414186 282258 414422 282494
rect 414186 275258 414422 275494
rect 414186 268258 414422 268494
rect 414186 261258 414422 261494
rect 414186 254258 414422 254494
rect 414186 247258 414422 247494
rect 414186 240258 414422 240494
rect 414186 233258 414422 233494
rect 414186 226258 414422 226494
rect 414186 219258 414422 219494
rect 414186 212258 414422 212494
rect 414186 205258 414422 205494
rect 414186 198258 414422 198494
rect 414186 191258 414422 191494
rect 414186 184258 414422 184494
rect 414186 177258 414422 177494
rect 414186 170258 414422 170494
rect 414186 163258 414422 163494
rect 414186 156258 414422 156494
rect 414186 149258 414422 149494
rect 414186 142258 414422 142494
rect 414186 135258 414422 135494
rect 414186 128258 414422 128494
rect 414186 121258 414422 121494
rect 414186 114258 414422 114494
rect 414186 107258 414422 107494
rect 414186 100258 414422 100494
rect 414186 93258 414422 93494
rect 414186 86258 414422 86494
rect 414186 79258 414422 79494
rect 414186 72258 414422 72494
rect 414186 65258 414422 65494
rect 414186 58258 414422 58494
rect 414186 51258 414422 51494
rect 414186 44258 414422 44494
rect 414186 37258 414422 37494
rect 414186 30258 414422 30494
rect 414186 23258 414422 23494
rect 414186 16258 414422 16494
rect 414186 9258 414422 9494
rect 414186 2258 414422 2494
rect 414186 -982 414422 -746
rect 414186 -1302 414422 -1066
rect 415918 705962 416154 706198
rect 415918 705642 416154 705878
rect 415918 696198 416154 696434
rect 415918 689198 416154 689434
rect 415918 682198 416154 682434
rect 415918 675198 416154 675434
rect 415918 668198 416154 668434
rect 415918 661198 416154 661434
rect 415918 654198 416154 654434
rect 415918 647198 416154 647434
rect 415918 640198 416154 640434
rect 415918 633198 416154 633434
rect 415918 626198 416154 626434
rect 415918 619198 416154 619434
rect 415918 612198 416154 612434
rect 415918 605198 416154 605434
rect 415918 598198 416154 598434
rect 415918 591198 416154 591434
rect 415918 584198 416154 584434
rect 415918 577198 416154 577434
rect 415918 570198 416154 570434
rect 415918 563198 416154 563434
rect 415918 556198 416154 556434
rect 415918 549198 416154 549434
rect 415918 542198 416154 542434
rect 415918 535198 416154 535434
rect 415918 528198 416154 528434
rect 415918 521198 416154 521434
rect 415918 514198 416154 514434
rect 415918 507198 416154 507434
rect 415918 500198 416154 500434
rect 415918 493198 416154 493434
rect 415918 486198 416154 486434
rect 415918 479198 416154 479434
rect 415918 472198 416154 472434
rect 415918 465198 416154 465434
rect 415918 458198 416154 458434
rect 415918 451198 416154 451434
rect 415918 444198 416154 444434
rect 415918 437198 416154 437434
rect 415918 430198 416154 430434
rect 415918 423198 416154 423434
rect 415918 416198 416154 416434
rect 415918 409198 416154 409434
rect 415918 402198 416154 402434
rect 415918 395198 416154 395434
rect 415918 388198 416154 388434
rect 415918 381198 416154 381434
rect 415918 374198 416154 374434
rect 415918 367198 416154 367434
rect 415918 360198 416154 360434
rect 415918 353198 416154 353434
rect 415918 346198 416154 346434
rect 415918 339198 416154 339434
rect 415918 332198 416154 332434
rect 415918 325198 416154 325434
rect 415918 318198 416154 318434
rect 415918 311198 416154 311434
rect 415918 304198 416154 304434
rect 415918 297198 416154 297434
rect 415918 290198 416154 290434
rect 415918 283198 416154 283434
rect 415918 276198 416154 276434
rect 415918 269198 416154 269434
rect 415918 262198 416154 262434
rect 415918 255198 416154 255434
rect 415918 248198 416154 248434
rect 415918 241198 416154 241434
rect 415918 234198 416154 234434
rect 415918 227198 416154 227434
rect 415918 220198 416154 220434
rect 415918 213198 416154 213434
rect 415918 206198 416154 206434
rect 415918 199198 416154 199434
rect 415918 192198 416154 192434
rect 415918 185198 416154 185434
rect 415918 178198 416154 178434
rect 415918 171198 416154 171434
rect 415918 164198 416154 164434
rect 415918 157198 416154 157434
rect 415918 150198 416154 150434
rect 415918 143198 416154 143434
rect 415918 136198 416154 136434
rect 415918 129198 416154 129434
rect 415918 122198 416154 122434
rect 415918 115198 416154 115434
rect 415918 108198 416154 108434
rect 415918 101198 416154 101434
rect 415918 94198 416154 94434
rect 415918 87198 416154 87434
rect 415918 80198 416154 80434
rect 415918 73198 416154 73434
rect 415918 66198 416154 66434
rect 415918 59198 416154 59434
rect 415918 52198 416154 52434
rect 415918 45198 416154 45434
rect 415918 38198 416154 38434
rect 415918 31198 416154 31434
rect 415918 24198 416154 24434
rect 415918 17198 416154 17434
rect 415918 10198 416154 10434
rect 415918 3198 416154 3434
rect 415918 -1942 416154 -1706
rect 415918 -2262 416154 -2026
rect 421186 705002 421422 705238
rect 421186 704682 421422 704918
rect 421186 695258 421422 695494
rect 421186 688258 421422 688494
rect 421186 681258 421422 681494
rect 421186 674258 421422 674494
rect 421186 667258 421422 667494
rect 421186 660258 421422 660494
rect 421186 653258 421422 653494
rect 421186 646258 421422 646494
rect 421186 639258 421422 639494
rect 421186 632258 421422 632494
rect 421186 625258 421422 625494
rect 421186 618258 421422 618494
rect 421186 611258 421422 611494
rect 421186 604258 421422 604494
rect 421186 597258 421422 597494
rect 421186 590258 421422 590494
rect 421186 583258 421422 583494
rect 421186 576258 421422 576494
rect 421186 569258 421422 569494
rect 421186 562258 421422 562494
rect 421186 555258 421422 555494
rect 421186 548258 421422 548494
rect 421186 541258 421422 541494
rect 421186 534258 421422 534494
rect 421186 527258 421422 527494
rect 421186 520258 421422 520494
rect 421186 513258 421422 513494
rect 421186 506258 421422 506494
rect 421186 499258 421422 499494
rect 421186 492258 421422 492494
rect 421186 485258 421422 485494
rect 421186 478258 421422 478494
rect 421186 471258 421422 471494
rect 421186 464258 421422 464494
rect 421186 457258 421422 457494
rect 421186 450258 421422 450494
rect 421186 443258 421422 443494
rect 421186 436258 421422 436494
rect 421186 429258 421422 429494
rect 421186 422258 421422 422494
rect 421186 415258 421422 415494
rect 421186 408258 421422 408494
rect 421186 401258 421422 401494
rect 421186 394258 421422 394494
rect 421186 387258 421422 387494
rect 421186 380258 421422 380494
rect 421186 373258 421422 373494
rect 421186 366258 421422 366494
rect 421186 359258 421422 359494
rect 421186 352258 421422 352494
rect 421186 345258 421422 345494
rect 421186 338258 421422 338494
rect 421186 331258 421422 331494
rect 421186 324258 421422 324494
rect 421186 317258 421422 317494
rect 421186 310258 421422 310494
rect 421186 303258 421422 303494
rect 421186 296258 421422 296494
rect 421186 289258 421422 289494
rect 421186 282258 421422 282494
rect 421186 275258 421422 275494
rect 421186 268258 421422 268494
rect 421186 261258 421422 261494
rect 421186 254258 421422 254494
rect 421186 247258 421422 247494
rect 421186 240258 421422 240494
rect 421186 233258 421422 233494
rect 421186 226258 421422 226494
rect 421186 219258 421422 219494
rect 421186 212258 421422 212494
rect 421186 205258 421422 205494
rect 421186 198258 421422 198494
rect 421186 191258 421422 191494
rect 421186 184258 421422 184494
rect 421186 177258 421422 177494
rect 421186 170258 421422 170494
rect 421186 163258 421422 163494
rect 421186 156258 421422 156494
rect 421186 149258 421422 149494
rect 421186 142258 421422 142494
rect 421186 135258 421422 135494
rect 421186 128258 421422 128494
rect 421186 121258 421422 121494
rect 421186 114258 421422 114494
rect 421186 107258 421422 107494
rect 421186 100258 421422 100494
rect 421186 93258 421422 93494
rect 421186 86258 421422 86494
rect 421186 79258 421422 79494
rect 421186 72258 421422 72494
rect 421186 65258 421422 65494
rect 421186 58258 421422 58494
rect 421186 51258 421422 51494
rect 421186 44258 421422 44494
rect 421186 37258 421422 37494
rect 421186 30258 421422 30494
rect 421186 23258 421422 23494
rect 421186 16258 421422 16494
rect 421186 9258 421422 9494
rect 421186 2258 421422 2494
rect 421186 -982 421422 -746
rect 421186 -1302 421422 -1066
rect 422918 705962 423154 706198
rect 422918 705642 423154 705878
rect 422918 696198 423154 696434
rect 422918 689198 423154 689434
rect 422918 682198 423154 682434
rect 422918 675198 423154 675434
rect 422918 668198 423154 668434
rect 422918 661198 423154 661434
rect 422918 654198 423154 654434
rect 422918 647198 423154 647434
rect 422918 640198 423154 640434
rect 422918 633198 423154 633434
rect 422918 626198 423154 626434
rect 422918 619198 423154 619434
rect 422918 612198 423154 612434
rect 422918 605198 423154 605434
rect 422918 598198 423154 598434
rect 422918 591198 423154 591434
rect 422918 584198 423154 584434
rect 422918 577198 423154 577434
rect 422918 570198 423154 570434
rect 422918 563198 423154 563434
rect 422918 556198 423154 556434
rect 422918 549198 423154 549434
rect 422918 542198 423154 542434
rect 422918 535198 423154 535434
rect 422918 528198 423154 528434
rect 422918 521198 423154 521434
rect 422918 514198 423154 514434
rect 422918 507198 423154 507434
rect 422918 500198 423154 500434
rect 422918 493198 423154 493434
rect 422918 486198 423154 486434
rect 422918 479198 423154 479434
rect 422918 472198 423154 472434
rect 422918 465198 423154 465434
rect 422918 458198 423154 458434
rect 422918 451198 423154 451434
rect 422918 444198 423154 444434
rect 422918 437198 423154 437434
rect 422918 430198 423154 430434
rect 422918 423198 423154 423434
rect 422918 416198 423154 416434
rect 422918 409198 423154 409434
rect 422918 402198 423154 402434
rect 422918 395198 423154 395434
rect 422918 388198 423154 388434
rect 422918 381198 423154 381434
rect 422918 374198 423154 374434
rect 422918 367198 423154 367434
rect 422918 360198 423154 360434
rect 422918 353198 423154 353434
rect 422918 346198 423154 346434
rect 422918 339198 423154 339434
rect 422918 332198 423154 332434
rect 422918 325198 423154 325434
rect 422918 318198 423154 318434
rect 422918 311198 423154 311434
rect 422918 304198 423154 304434
rect 422918 297198 423154 297434
rect 422918 290198 423154 290434
rect 422918 283198 423154 283434
rect 422918 276198 423154 276434
rect 422918 269198 423154 269434
rect 422918 262198 423154 262434
rect 422918 255198 423154 255434
rect 422918 248198 423154 248434
rect 422918 241198 423154 241434
rect 422918 234198 423154 234434
rect 422918 227198 423154 227434
rect 422918 220198 423154 220434
rect 422918 213198 423154 213434
rect 422918 206198 423154 206434
rect 422918 199198 423154 199434
rect 422918 192198 423154 192434
rect 422918 185198 423154 185434
rect 422918 178198 423154 178434
rect 422918 171198 423154 171434
rect 422918 164198 423154 164434
rect 422918 157198 423154 157434
rect 422918 150198 423154 150434
rect 422918 143198 423154 143434
rect 422918 136198 423154 136434
rect 422918 129198 423154 129434
rect 422918 122198 423154 122434
rect 422918 115198 423154 115434
rect 422918 108198 423154 108434
rect 422918 101198 423154 101434
rect 422918 94198 423154 94434
rect 422918 87198 423154 87434
rect 422918 80198 423154 80434
rect 422918 73198 423154 73434
rect 422918 66198 423154 66434
rect 422918 59198 423154 59434
rect 422918 52198 423154 52434
rect 422918 45198 423154 45434
rect 422918 38198 423154 38434
rect 422918 31198 423154 31434
rect 422918 24198 423154 24434
rect 422918 17198 423154 17434
rect 422918 10198 423154 10434
rect 422918 3198 423154 3434
rect 422918 -1942 423154 -1706
rect 422918 -2262 423154 -2026
rect 428186 705002 428422 705238
rect 428186 704682 428422 704918
rect 428186 695258 428422 695494
rect 428186 688258 428422 688494
rect 428186 681258 428422 681494
rect 428186 674258 428422 674494
rect 428186 667258 428422 667494
rect 428186 660258 428422 660494
rect 428186 653258 428422 653494
rect 428186 646258 428422 646494
rect 428186 639258 428422 639494
rect 428186 632258 428422 632494
rect 428186 625258 428422 625494
rect 428186 618258 428422 618494
rect 428186 611258 428422 611494
rect 428186 604258 428422 604494
rect 428186 597258 428422 597494
rect 428186 590258 428422 590494
rect 428186 583258 428422 583494
rect 428186 576258 428422 576494
rect 428186 569258 428422 569494
rect 428186 562258 428422 562494
rect 428186 555258 428422 555494
rect 428186 548258 428422 548494
rect 428186 541258 428422 541494
rect 428186 534258 428422 534494
rect 428186 527258 428422 527494
rect 428186 520258 428422 520494
rect 428186 513258 428422 513494
rect 428186 506258 428422 506494
rect 428186 499258 428422 499494
rect 428186 492258 428422 492494
rect 428186 485258 428422 485494
rect 428186 478258 428422 478494
rect 428186 471258 428422 471494
rect 428186 464258 428422 464494
rect 428186 457258 428422 457494
rect 428186 450258 428422 450494
rect 428186 443258 428422 443494
rect 428186 436258 428422 436494
rect 428186 429258 428422 429494
rect 428186 422258 428422 422494
rect 428186 415258 428422 415494
rect 428186 408258 428422 408494
rect 428186 401258 428422 401494
rect 428186 394258 428422 394494
rect 428186 387258 428422 387494
rect 428186 380258 428422 380494
rect 428186 373258 428422 373494
rect 428186 366258 428422 366494
rect 428186 359258 428422 359494
rect 428186 352258 428422 352494
rect 428186 345258 428422 345494
rect 428186 338258 428422 338494
rect 428186 331258 428422 331494
rect 428186 324258 428422 324494
rect 428186 317258 428422 317494
rect 428186 310258 428422 310494
rect 428186 303258 428422 303494
rect 428186 296258 428422 296494
rect 428186 289258 428422 289494
rect 428186 282258 428422 282494
rect 428186 275258 428422 275494
rect 428186 268258 428422 268494
rect 428186 261258 428422 261494
rect 428186 254258 428422 254494
rect 428186 247258 428422 247494
rect 428186 240258 428422 240494
rect 428186 233258 428422 233494
rect 428186 226258 428422 226494
rect 428186 219258 428422 219494
rect 428186 212258 428422 212494
rect 428186 205258 428422 205494
rect 428186 198258 428422 198494
rect 428186 191258 428422 191494
rect 428186 184258 428422 184494
rect 428186 177258 428422 177494
rect 428186 170258 428422 170494
rect 428186 163258 428422 163494
rect 428186 156258 428422 156494
rect 428186 149258 428422 149494
rect 428186 142258 428422 142494
rect 428186 135258 428422 135494
rect 428186 128258 428422 128494
rect 428186 121258 428422 121494
rect 428186 114258 428422 114494
rect 428186 107258 428422 107494
rect 428186 100258 428422 100494
rect 428186 93258 428422 93494
rect 428186 86258 428422 86494
rect 428186 79258 428422 79494
rect 428186 72258 428422 72494
rect 428186 65258 428422 65494
rect 428186 58258 428422 58494
rect 428186 51258 428422 51494
rect 428186 44258 428422 44494
rect 428186 37258 428422 37494
rect 428186 30258 428422 30494
rect 428186 23258 428422 23494
rect 428186 16258 428422 16494
rect 428186 9258 428422 9494
rect 428186 2258 428422 2494
rect 428186 -982 428422 -746
rect 428186 -1302 428422 -1066
rect 429918 705962 430154 706198
rect 429918 705642 430154 705878
rect 429918 696198 430154 696434
rect 429918 689198 430154 689434
rect 429918 682198 430154 682434
rect 429918 675198 430154 675434
rect 429918 668198 430154 668434
rect 429918 661198 430154 661434
rect 429918 654198 430154 654434
rect 429918 647198 430154 647434
rect 429918 640198 430154 640434
rect 429918 633198 430154 633434
rect 429918 626198 430154 626434
rect 429918 619198 430154 619434
rect 429918 612198 430154 612434
rect 429918 605198 430154 605434
rect 429918 598198 430154 598434
rect 429918 591198 430154 591434
rect 429918 584198 430154 584434
rect 429918 577198 430154 577434
rect 429918 570198 430154 570434
rect 429918 563198 430154 563434
rect 429918 556198 430154 556434
rect 429918 549198 430154 549434
rect 429918 542198 430154 542434
rect 429918 535198 430154 535434
rect 429918 528198 430154 528434
rect 429918 521198 430154 521434
rect 429918 514198 430154 514434
rect 429918 507198 430154 507434
rect 429918 500198 430154 500434
rect 429918 493198 430154 493434
rect 429918 486198 430154 486434
rect 429918 479198 430154 479434
rect 429918 472198 430154 472434
rect 429918 465198 430154 465434
rect 429918 458198 430154 458434
rect 429918 451198 430154 451434
rect 429918 444198 430154 444434
rect 429918 437198 430154 437434
rect 429918 430198 430154 430434
rect 429918 423198 430154 423434
rect 429918 416198 430154 416434
rect 429918 409198 430154 409434
rect 429918 402198 430154 402434
rect 429918 395198 430154 395434
rect 429918 388198 430154 388434
rect 429918 381198 430154 381434
rect 429918 374198 430154 374434
rect 429918 367198 430154 367434
rect 429918 360198 430154 360434
rect 429918 353198 430154 353434
rect 429918 346198 430154 346434
rect 429918 339198 430154 339434
rect 429918 332198 430154 332434
rect 429918 325198 430154 325434
rect 429918 318198 430154 318434
rect 429918 311198 430154 311434
rect 429918 304198 430154 304434
rect 429918 297198 430154 297434
rect 429918 290198 430154 290434
rect 429918 283198 430154 283434
rect 429918 276198 430154 276434
rect 429918 269198 430154 269434
rect 429918 262198 430154 262434
rect 429918 255198 430154 255434
rect 429918 248198 430154 248434
rect 429918 241198 430154 241434
rect 429918 234198 430154 234434
rect 429918 227198 430154 227434
rect 429918 220198 430154 220434
rect 429918 213198 430154 213434
rect 429918 206198 430154 206434
rect 429918 199198 430154 199434
rect 429918 192198 430154 192434
rect 429918 185198 430154 185434
rect 429918 178198 430154 178434
rect 429918 171198 430154 171434
rect 429918 164198 430154 164434
rect 429918 157198 430154 157434
rect 429918 150198 430154 150434
rect 429918 143198 430154 143434
rect 429918 136198 430154 136434
rect 429918 129198 430154 129434
rect 429918 122198 430154 122434
rect 429918 115198 430154 115434
rect 429918 108198 430154 108434
rect 429918 101198 430154 101434
rect 429918 94198 430154 94434
rect 429918 87198 430154 87434
rect 429918 80198 430154 80434
rect 429918 73198 430154 73434
rect 429918 66198 430154 66434
rect 429918 59198 430154 59434
rect 429918 52198 430154 52434
rect 429918 45198 430154 45434
rect 429918 38198 430154 38434
rect 429918 31198 430154 31434
rect 429918 24198 430154 24434
rect 429918 17198 430154 17434
rect 429918 10198 430154 10434
rect 429918 3198 430154 3434
rect 429918 -1942 430154 -1706
rect 429918 -2262 430154 -2026
rect 435186 705002 435422 705238
rect 435186 704682 435422 704918
rect 435186 695258 435422 695494
rect 435186 688258 435422 688494
rect 435186 681258 435422 681494
rect 435186 674258 435422 674494
rect 435186 667258 435422 667494
rect 435186 660258 435422 660494
rect 435186 653258 435422 653494
rect 435186 646258 435422 646494
rect 435186 639258 435422 639494
rect 435186 632258 435422 632494
rect 435186 625258 435422 625494
rect 435186 618258 435422 618494
rect 435186 611258 435422 611494
rect 435186 604258 435422 604494
rect 435186 597258 435422 597494
rect 435186 590258 435422 590494
rect 435186 583258 435422 583494
rect 435186 576258 435422 576494
rect 435186 569258 435422 569494
rect 435186 562258 435422 562494
rect 435186 555258 435422 555494
rect 435186 548258 435422 548494
rect 435186 541258 435422 541494
rect 435186 534258 435422 534494
rect 435186 527258 435422 527494
rect 435186 520258 435422 520494
rect 435186 513258 435422 513494
rect 435186 506258 435422 506494
rect 435186 499258 435422 499494
rect 435186 492258 435422 492494
rect 435186 485258 435422 485494
rect 435186 478258 435422 478494
rect 435186 471258 435422 471494
rect 435186 464258 435422 464494
rect 435186 457258 435422 457494
rect 435186 450258 435422 450494
rect 435186 443258 435422 443494
rect 435186 436258 435422 436494
rect 435186 429258 435422 429494
rect 435186 422258 435422 422494
rect 435186 415258 435422 415494
rect 435186 408258 435422 408494
rect 435186 401258 435422 401494
rect 435186 394258 435422 394494
rect 435186 387258 435422 387494
rect 435186 380258 435422 380494
rect 435186 373258 435422 373494
rect 435186 366258 435422 366494
rect 435186 359258 435422 359494
rect 435186 352258 435422 352494
rect 435186 345258 435422 345494
rect 435186 338258 435422 338494
rect 435186 331258 435422 331494
rect 435186 324258 435422 324494
rect 435186 317258 435422 317494
rect 435186 310258 435422 310494
rect 435186 303258 435422 303494
rect 435186 296258 435422 296494
rect 435186 289258 435422 289494
rect 435186 282258 435422 282494
rect 435186 275258 435422 275494
rect 435186 268258 435422 268494
rect 435186 261258 435422 261494
rect 435186 254258 435422 254494
rect 435186 247258 435422 247494
rect 435186 240258 435422 240494
rect 435186 233258 435422 233494
rect 435186 226258 435422 226494
rect 435186 219258 435422 219494
rect 435186 212258 435422 212494
rect 435186 205258 435422 205494
rect 435186 198258 435422 198494
rect 435186 191258 435422 191494
rect 435186 184258 435422 184494
rect 435186 177258 435422 177494
rect 435186 170258 435422 170494
rect 435186 163258 435422 163494
rect 435186 156258 435422 156494
rect 435186 149258 435422 149494
rect 435186 142258 435422 142494
rect 435186 135258 435422 135494
rect 435186 128258 435422 128494
rect 435186 121258 435422 121494
rect 435186 114258 435422 114494
rect 435186 107258 435422 107494
rect 435186 100258 435422 100494
rect 435186 93258 435422 93494
rect 435186 86258 435422 86494
rect 435186 79258 435422 79494
rect 435186 72258 435422 72494
rect 435186 65258 435422 65494
rect 435186 58258 435422 58494
rect 435186 51258 435422 51494
rect 435186 44258 435422 44494
rect 435186 37258 435422 37494
rect 435186 30258 435422 30494
rect 435186 23258 435422 23494
rect 435186 16258 435422 16494
rect 435186 9258 435422 9494
rect 435186 2258 435422 2494
rect 435186 -982 435422 -746
rect 435186 -1302 435422 -1066
rect 436918 705962 437154 706198
rect 436918 705642 437154 705878
rect 436918 696198 437154 696434
rect 436918 689198 437154 689434
rect 436918 682198 437154 682434
rect 436918 675198 437154 675434
rect 436918 668198 437154 668434
rect 436918 661198 437154 661434
rect 436918 654198 437154 654434
rect 436918 647198 437154 647434
rect 436918 640198 437154 640434
rect 436918 633198 437154 633434
rect 436918 626198 437154 626434
rect 436918 619198 437154 619434
rect 436918 612198 437154 612434
rect 436918 605198 437154 605434
rect 436918 598198 437154 598434
rect 436918 591198 437154 591434
rect 436918 584198 437154 584434
rect 436918 577198 437154 577434
rect 436918 570198 437154 570434
rect 436918 563198 437154 563434
rect 436918 556198 437154 556434
rect 436918 549198 437154 549434
rect 436918 542198 437154 542434
rect 436918 535198 437154 535434
rect 436918 528198 437154 528434
rect 436918 521198 437154 521434
rect 436918 514198 437154 514434
rect 436918 507198 437154 507434
rect 436918 500198 437154 500434
rect 436918 493198 437154 493434
rect 436918 486198 437154 486434
rect 436918 479198 437154 479434
rect 436918 472198 437154 472434
rect 436918 465198 437154 465434
rect 436918 458198 437154 458434
rect 436918 451198 437154 451434
rect 436918 444198 437154 444434
rect 436918 437198 437154 437434
rect 436918 430198 437154 430434
rect 436918 423198 437154 423434
rect 436918 416198 437154 416434
rect 436918 409198 437154 409434
rect 436918 402198 437154 402434
rect 436918 395198 437154 395434
rect 436918 388198 437154 388434
rect 436918 381198 437154 381434
rect 436918 374198 437154 374434
rect 436918 367198 437154 367434
rect 436918 360198 437154 360434
rect 436918 353198 437154 353434
rect 436918 346198 437154 346434
rect 436918 339198 437154 339434
rect 436918 332198 437154 332434
rect 436918 325198 437154 325434
rect 436918 318198 437154 318434
rect 436918 311198 437154 311434
rect 436918 304198 437154 304434
rect 436918 297198 437154 297434
rect 436918 290198 437154 290434
rect 436918 283198 437154 283434
rect 436918 276198 437154 276434
rect 436918 269198 437154 269434
rect 436918 262198 437154 262434
rect 436918 255198 437154 255434
rect 436918 248198 437154 248434
rect 436918 241198 437154 241434
rect 436918 234198 437154 234434
rect 436918 227198 437154 227434
rect 436918 220198 437154 220434
rect 436918 213198 437154 213434
rect 436918 206198 437154 206434
rect 436918 199198 437154 199434
rect 436918 192198 437154 192434
rect 436918 185198 437154 185434
rect 436918 178198 437154 178434
rect 436918 171198 437154 171434
rect 436918 164198 437154 164434
rect 436918 157198 437154 157434
rect 436918 150198 437154 150434
rect 436918 143198 437154 143434
rect 436918 136198 437154 136434
rect 436918 129198 437154 129434
rect 436918 122198 437154 122434
rect 436918 115198 437154 115434
rect 436918 108198 437154 108434
rect 436918 101198 437154 101434
rect 436918 94198 437154 94434
rect 436918 87198 437154 87434
rect 436918 80198 437154 80434
rect 436918 73198 437154 73434
rect 436918 66198 437154 66434
rect 436918 59198 437154 59434
rect 436918 52198 437154 52434
rect 436918 45198 437154 45434
rect 436918 38198 437154 38434
rect 436918 31198 437154 31434
rect 436918 24198 437154 24434
rect 436918 17198 437154 17434
rect 436918 10198 437154 10434
rect 436918 3198 437154 3434
rect 436918 -1942 437154 -1706
rect 436918 -2262 437154 -2026
rect 442186 705002 442422 705238
rect 442186 704682 442422 704918
rect 442186 695258 442422 695494
rect 442186 688258 442422 688494
rect 442186 681258 442422 681494
rect 442186 674258 442422 674494
rect 442186 667258 442422 667494
rect 442186 660258 442422 660494
rect 442186 653258 442422 653494
rect 442186 646258 442422 646494
rect 442186 639258 442422 639494
rect 442186 632258 442422 632494
rect 442186 625258 442422 625494
rect 442186 618258 442422 618494
rect 442186 611258 442422 611494
rect 442186 604258 442422 604494
rect 442186 597258 442422 597494
rect 442186 590258 442422 590494
rect 442186 583258 442422 583494
rect 442186 576258 442422 576494
rect 442186 569258 442422 569494
rect 442186 562258 442422 562494
rect 442186 555258 442422 555494
rect 442186 548258 442422 548494
rect 442186 541258 442422 541494
rect 442186 534258 442422 534494
rect 442186 527258 442422 527494
rect 442186 520258 442422 520494
rect 442186 513258 442422 513494
rect 442186 506258 442422 506494
rect 442186 499258 442422 499494
rect 442186 492258 442422 492494
rect 442186 485258 442422 485494
rect 442186 478258 442422 478494
rect 442186 471258 442422 471494
rect 442186 464258 442422 464494
rect 442186 457258 442422 457494
rect 442186 450258 442422 450494
rect 442186 443258 442422 443494
rect 442186 436258 442422 436494
rect 442186 429258 442422 429494
rect 442186 422258 442422 422494
rect 442186 415258 442422 415494
rect 442186 408258 442422 408494
rect 442186 401258 442422 401494
rect 442186 394258 442422 394494
rect 442186 387258 442422 387494
rect 442186 380258 442422 380494
rect 442186 373258 442422 373494
rect 442186 366258 442422 366494
rect 442186 359258 442422 359494
rect 442186 352258 442422 352494
rect 442186 345258 442422 345494
rect 442186 338258 442422 338494
rect 442186 331258 442422 331494
rect 442186 324258 442422 324494
rect 442186 317258 442422 317494
rect 442186 310258 442422 310494
rect 442186 303258 442422 303494
rect 442186 296258 442422 296494
rect 442186 289258 442422 289494
rect 442186 282258 442422 282494
rect 442186 275258 442422 275494
rect 442186 268258 442422 268494
rect 442186 261258 442422 261494
rect 442186 254258 442422 254494
rect 442186 247258 442422 247494
rect 442186 240258 442422 240494
rect 442186 233258 442422 233494
rect 442186 226258 442422 226494
rect 442186 219258 442422 219494
rect 442186 212258 442422 212494
rect 442186 205258 442422 205494
rect 442186 198258 442422 198494
rect 442186 191258 442422 191494
rect 442186 184258 442422 184494
rect 442186 177258 442422 177494
rect 442186 170258 442422 170494
rect 442186 163258 442422 163494
rect 442186 156258 442422 156494
rect 442186 149258 442422 149494
rect 442186 142258 442422 142494
rect 442186 135258 442422 135494
rect 442186 128258 442422 128494
rect 442186 121258 442422 121494
rect 442186 114258 442422 114494
rect 442186 107258 442422 107494
rect 442186 100258 442422 100494
rect 442186 93258 442422 93494
rect 442186 86258 442422 86494
rect 442186 79258 442422 79494
rect 442186 72258 442422 72494
rect 442186 65258 442422 65494
rect 442186 58258 442422 58494
rect 442186 51258 442422 51494
rect 442186 44258 442422 44494
rect 442186 37258 442422 37494
rect 442186 30258 442422 30494
rect 442186 23258 442422 23494
rect 442186 16258 442422 16494
rect 442186 9258 442422 9494
rect 442186 2258 442422 2494
rect 442186 -982 442422 -746
rect 442186 -1302 442422 -1066
rect 443918 705962 444154 706198
rect 443918 705642 444154 705878
rect 443918 696198 444154 696434
rect 443918 689198 444154 689434
rect 443918 682198 444154 682434
rect 443918 675198 444154 675434
rect 443918 668198 444154 668434
rect 443918 661198 444154 661434
rect 443918 654198 444154 654434
rect 443918 647198 444154 647434
rect 443918 640198 444154 640434
rect 443918 633198 444154 633434
rect 443918 626198 444154 626434
rect 443918 619198 444154 619434
rect 443918 612198 444154 612434
rect 443918 605198 444154 605434
rect 443918 598198 444154 598434
rect 443918 591198 444154 591434
rect 443918 584198 444154 584434
rect 443918 577198 444154 577434
rect 443918 570198 444154 570434
rect 443918 563198 444154 563434
rect 443918 556198 444154 556434
rect 443918 549198 444154 549434
rect 443918 542198 444154 542434
rect 443918 535198 444154 535434
rect 443918 528198 444154 528434
rect 443918 521198 444154 521434
rect 443918 514198 444154 514434
rect 443918 507198 444154 507434
rect 443918 500198 444154 500434
rect 443918 493198 444154 493434
rect 443918 486198 444154 486434
rect 443918 479198 444154 479434
rect 443918 472198 444154 472434
rect 443918 465198 444154 465434
rect 443918 458198 444154 458434
rect 443918 451198 444154 451434
rect 443918 444198 444154 444434
rect 443918 437198 444154 437434
rect 443918 430198 444154 430434
rect 443918 423198 444154 423434
rect 443918 416198 444154 416434
rect 443918 409198 444154 409434
rect 443918 402198 444154 402434
rect 443918 395198 444154 395434
rect 443918 388198 444154 388434
rect 443918 381198 444154 381434
rect 443918 374198 444154 374434
rect 443918 367198 444154 367434
rect 443918 360198 444154 360434
rect 443918 353198 444154 353434
rect 443918 346198 444154 346434
rect 443918 339198 444154 339434
rect 443918 332198 444154 332434
rect 443918 325198 444154 325434
rect 443918 318198 444154 318434
rect 443918 311198 444154 311434
rect 443918 304198 444154 304434
rect 443918 297198 444154 297434
rect 443918 290198 444154 290434
rect 443918 283198 444154 283434
rect 443918 276198 444154 276434
rect 443918 269198 444154 269434
rect 443918 262198 444154 262434
rect 443918 255198 444154 255434
rect 443918 248198 444154 248434
rect 443918 241198 444154 241434
rect 443918 234198 444154 234434
rect 443918 227198 444154 227434
rect 443918 220198 444154 220434
rect 443918 213198 444154 213434
rect 443918 206198 444154 206434
rect 443918 199198 444154 199434
rect 443918 192198 444154 192434
rect 443918 185198 444154 185434
rect 443918 178198 444154 178434
rect 443918 171198 444154 171434
rect 443918 164198 444154 164434
rect 443918 157198 444154 157434
rect 443918 150198 444154 150434
rect 443918 143198 444154 143434
rect 443918 136198 444154 136434
rect 443918 129198 444154 129434
rect 443918 122198 444154 122434
rect 443918 115198 444154 115434
rect 443918 108198 444154 108434
rect 443918 101198 444154 101434
rect 443918 94198 444154 94434
rect 443918 87198 444154 87434
rect 443918 80198 444154 80434
rect 443918 73198 444154 73434
rect 443918 66198 444154 66434
rect 443918 59198 444154 59434
rect 443918 52198 444154 52434
rect 443918 45198 444154 45434
rect 443918 38198 444154 38434
rect 443918 31198 444154 31434
rect 443918 24198 444154 24434
rect 443918 17198 444154 17434
rect 443918 10198 444154 10434
rect 443918 3198 444154 3434
rect 443918 -1942 444154 -1706
rect 443918 -2262 444154 -2026
rect 449186 705002 449422 705238
rect 449186 704682 449422 704918
rect 449186 695258 449422 695494
rect 449186 688258 449422 688494
rect 449186 681258 449422 681494
rect 449186 674258 449422 674494
rect 449186 667258 449422 667494
rect 449186 660258 449422 660494
rect 449186 653258 449422 653494
rect 449186 646258 449422 646494
rect 449186 639258 449422 639494
rect 449186 632258 449422 632494
rect 449186 625258 449422 625494
rect 449186 618258 449422 618494
rect 449186 611258 449422 611494
rect 449186 604258 449422 604494
rect 449186 597258 449422 597494
rect 449186 590258 449422 590494
rect 449186 583258 449422 583494
rect 449186 576258 449422 576494
rect 449186 569258 449422 569494
rect 449186 562258 449422 562494
rect 449186 555258 449422 555494
rect 449186 548258 449422 548494
rect 449186 541258 449422 541494
rect 449186 534258 449422 534494
rect 449186 527258 449422 527494
rect 449186 520258 449422 520494
rect 449186 513258 449422 513494
rect 449186 506258 449422 506494
rect 449186 499258 449422 499494
rect 449186 492258 449422 492494
rect 449186 485258 449422 485494
rect 449186 478258 449422 478494
rect 449186 471258 449422 471494
rect 449186 464258 449422 464494
rect 449186 457258 449422 457494
rect 449186 450258 449422 450494
rect 449186 443258 449422 443494
rect 449186 436258 449422 436494
rect 449186 429258 449422 429494
rect 449186 422258 449422 422494
rect 449186 415258 449422 415494
rect 449186 408258 449422 408494
rect 449186 401258 449422 401494
rect 449186 394258 449422 394494
rect 449186 387258 449422 387494
rect 449186 380258 449422 380494
rect 449186 373258 449422 373494
rect 449186 366258 449422 366494
rect 449186 359258 449422 359494
rect 449186 352258 449422 352494
rect 449186 345258 449422 345494
rect 449186 338258 449422 338494
rect 449186 331258 449422 331494
rect 449186 324258 449422 324494
rect 449186 317258 449422 317494
rect 449186 310258 449422 310494
rect 449186 303258 449422 303494
rect 449186 296258 449422 296494
rect 449186 289258 449422 289494
rect 449186 282258 449422 282494
rect 449186 275258 449422 275494
rect 449186 268258 449422 268494
rect 449186 261258 449422 261494
rect 449186 254258 449422 254494
rect 449186 247258 449422 247494
rect 449186 240258 449422 240494
rect 449186 233258 449422 233494
rect 449186 226258 449422 226494
rect 449186 219258 449422 219494
rect 449186 212258 449422 212494
rect 449186 205258 449422 205494
rect 449186 198258 449422 198494
rect 449186 191258 449422 191494
rect 449186 184258 449422 184494
rect 449186 177258 449422 177494
rect 449186 170258 449422 170494
rect 449186 163258 449422 163494
rect 449186 156258 449422 156494
rect 449186 149258 449422 149494
rect 449186 142258 449422 142494
rect 449186 135258 449422 135494
rect 449186 128258 449422 128494
rect 449186 121258 449422 121494
rect 449186 114258 449422 114494
rect 449186 107258 449422 107494
rect 449186 100258 449422 100494
rect 449186 93258 449422 93494
rect 449186 86258 449422 86494
rect 449186 79258 449422 79494
rect 449186 72258 449422 72494
rect 449186 65258 449422 65494
rect 449186 58258 449422 58494
rect 449186 51258 449422 51494
rect 449186 44258 449422 44494
rect 449186 37258 449422 37494
rect 449186 30258 449422 30494
rect 449186 23258 449422 23494
rect 449186 16258 449422 16494
rect 449186 9258 449422 9494
rect 449186 2258 449422 2494
rect 449186 -982 449422 -746
rect 449186 -1302 449422 -1066
rect 450918 705962 451154 706198
rect 450918 705642 451154 705878
rect 450918 696198 451154 696434
rect 450918 689198 451154 689434
rect 450918 682198 451154 682434
rect 450918 675198 451154 675434
rect 450918 668198 451154 668434
rect 450918 661198 451154 661434
rect 450918 654198 451154 654434
rect 450918 647198 451154 647434
rect 450918 640198 451154 640434
rect 450918 633198 451154 633434
rect 450918 626198 451154 626434
rect 450918 619198 451154 619434
rect 450918 612198 451154 612434
rect 450918 605198 451154 605434
rect 450918 598198 451154 598434
rect 450918 591198 451154 591434
rect 450918 584198 451154 584434
rect 450918 577198 451154 577434
rect 450918 570198 451154 570434
rect 450918 563198 451154 563434
rect 450918 556198 451154 556434
rect 450918 549198 451154 549434
rect 450918 542198 451154 542434
rect 450918 535198 451154 535434
rect 450918 528198 451154 528434
rect 450918 521198 451154 521434
rect 450918 514198 451154 514434
rect 450918 507198 451154 507434
rect 450918 500198 451154 500434
rect 450918 493198 451154 493434
rect 450918 486198 451154 486434
rect 450918 479198 451154 479434
rect 450918 472198 451154 472434
rect 450918 465198 451154 465434
rect 450918 458198 451154 458434
rect 450918 451198 451154 451434
rect 450918 444198 451154 444434
rect 450918 437198 451154 437434
rect 450918 430198 451154 430434
rect 450918 423198 451154 423434
rect 450918 416198 451154 416434
rect 450918 409198 451154 409434
rect 450918 402198 451154 402434
rect 450918 395198 451154 395434
rect 450918 388198 451154 388434
rect 450918 381198 451154 381434
rect 450918 374198 451154 374434
rect 450918 367198 451154 367434
rect 450918 360198 451154 360434
rect 450918 353198 451154 353434
rect 450918 346198 451154 346434
rect 450918 339198 451154 339434
rect 450918 332198 451154 332434
rect 450918 325198 451154 325434
rect 450918 318198 451154 318434
rect 450918 311198 451154 311434
rect 450918 304198 451154 304434
rect 450918 297198 451154 297434
rect 450918 290198 451154 290434
rect 450918 283198 451154 283434
rect 450918 276198 451154 276434
rect 450918 269198 451154 269434
rect 450918 262198 451154 262434
rect 450918 255198 451154 255434
rect 450918 248198 451154 248434
rect 450918 241198 451154 241434
rect 450918 234198 451154 234434
rect 450918 227198 451154 227434
rect 450918 220198 451154 220434
rect 450918 213198 451154 213434
rect 450918 206198 451154 206434
rect 450918 199198 451154 199434
rect 450918 192198 451154 192434
rect 450918 185198 451154 185434
rect 450918 178198 451154 178434
rect 450918 171198 451154 171434
rect 450918 164198 451154 164434
rect 450918 157198 451154 157434
rect 450918 150198 451154 150434
rect 450918 143198 451154 143434
rect 450918 136198 451154 136434
rect 450918 129198 451154 129434
rect 450918 122198 451154 122434
rect 450918 115198 451154 115434
rect 450918 108198 451154 108434
rect 450918 101198 451154 101434
rect 450918 94198 451154 94434
rect 450918 87198 451154 87434
rect 450918 80198 451154 80434
rect 450918 73198 451154 73434
rect 450918 66198 451154 66434
rect 450918 59198 451154 59434
rect 450918 52198 451154 52434
rect 450918 45198 451154 45434
rect 450918 38198 451154 38434
rect 450918 31198 451154 31434
rect 450918 24198 451154 24434
rect 450918 17198 451154 17434
rect 450918 10198 451154 10434
rect 450918 3198 451154 3434
rect 450918 -1942 451154 -1706
rect 450918 -2262 451154 -2026
rect 456186 705002 456422 705238
rect 456186 704682 456422 704918
rect 456186 695258 456422 695494
rect 456186 688258 456422 688494
rect 456186 681258 456422 681494
rect 456186 674258 456422 674494
rect 456186 667258 456422 667494
rect 456186 660258 456422 660494
rect 456186 653258 456422 653494
rect 456186 646258 456422 646494
rect 456186 639258 456422 639494
rect 456186 632258 456422 632494
rect 456186 625258 456422 625494
rect 456186 618258 456422 618494
rect 456186 611258 456422 611494
rect 456186 604258 456422 604494
rect 456186 597258 456422 597494
rect 456186 590258 456422 590494
rect 456186 583258 456422 583494
rect 456186 576258 456422 576494
rect 456186 569258 456422 569494
rect 456186 562258 456422 562494
rect 456186 555258 456422 555494
rect 456186 548258 456422 548494
rect 456186 541258 456422 541494
rect 456186 534258 456422 534494
rect 456186 527258 456422 527494
rect 456186 520258 456422 520494
rect 456186 513258 456422 513494
rect 456186 506258 456422 506494
rect 456186 499258 456422 499494
rect 456186 492258 456422 492494
rect 456186 485258 456422 485494
rect 456186 478258 456422 478494
rect 456186 471258 456422 471494
rect 456186 464258 456422 464494
rect 456186 457258 456422 457494
rect 456186 450258 456422 450494
rect 456186 443258 456422 443494
rect 456186 436258 456422 436494
rect 456186 429258 456422 429494
rect 456186 422258 456422 422494
rect 456186 415258 456422 415494
rect 456186 408258 456422 408494
rect 456186 401258 456422 401494
rect 456186 394258 456422 394494
rect 456186 387258 456422 387494
rect 456186 380258 456422 380494
rect 456186 373258 456422 373494
rect 456186 366258 456422 366494
rect 456186 359258 456422 359494
rect 456186 352258 456422 352494
rect 456186 345258 456422 345494
rect 456186 338258 456422 338494
rect 456186 331258 456422 331494
rect 456186 324258 456422 324494
rect 456186 317258 456422 317494
rect 456186 310258 456422 310494
rect 456186 303258 456422 303494
rect 456186 296258 456422 296494
rect 456186 289258 456422 289494
rect 456186 282258 456422 282494
rect 456186 275258 456422 275494
rect 456186 268258 456422 268494
rect 456186 261258 456422 261494
rect 456186 254258 456422 254494
rect 456186 247258 456422 247494
rect 456186 240258 456422 240494
rect 456186 233258 456422 233494
rect 456186 226258 456422 226494
rect 456186 219258 456422 219494
rect 456186 212258 456422 212494
rect 456186 205258 456422 205494
rect 456186 198258 456422 198494
rect 456186 191258 456422 191494
rect 456186 184258 456422 184494
rect 456186 177258 456422 177494
rect 456186 170258 456422 170494
rect 456186 163258 456422 163494
rect 456186 156258 456422 156494
rect 456186 149258 456422 149494
rect 456186 142258 456422 142494
rect 456186 135258 456422 135494
rect 456186 128258 456422 128494
rect 456186 121258 456422 121494
rect 456186 114258 456422 114494
rect 456186 107258 456422 107494
rect 456186 100258 456422 100494
rect 456186 93258 456422 93494
rect 456186 86258 456422 86494
rect 456186 79258 456422 79494
rect 456186 72258 456422 72494
rect 456186 65258 456422 65494
rect 456186 58258 456422 58494
rect 456186 51258 456422 51494
rect 456186 44258 456422 44494
rect 456186 37258 456422 37494
rect 456186 30258 456422 30494
rect 456186 23258 456422 23494
rect 456186 16258 456422 16494
rect 456186 9258 456422 9494
rect 456186 2258 456422 2494
rect 456186 -982 456422 -746
rect 456186 -1302 456422 -1066
rect 457918 705962 458154 706198
rect 457918 705642 458154 705878
rect 457918 696198 458154 696434
rect 457918 689198 458154 689434
rect 457918 682198 458154 682434
rect 457918 675198 458154 675434
rect 457918 668198 458154 668434
rect 457918 661198 458154 661434
rect 457918 654198 458154 654434
rect 457918 647198 458154 647434
rect 457918 640198 458154 640434
rect 457918 633198 458154 633434
rect 457918 626198 458154 626434
rect 457918 619198 458154 619434
rect 457918 612198 458154 612434
rect 457918 605198 458154 605434
rect 457918 598198 458154 598434
rect 457918 591198 458154 591434
rect 457918 584198 458154 584434
rect 457918 577198 458154 577434
rect 457918 570198 458154 570434
rect 457918 563198 458154 563434
rect 457918 556198 458154 556434
rect 457918 549198 458154 549434
rect 457918 542198 458154 542434
rect 457918 535198 458154 535434
rect 457918 528198 458154 528434
rect 457918 521198 458154 521434
rect 457918 514198 458154 514434
rect 457918 507198 458154 507434
rect 457918 500198 458154 500434
rect 457918 493198 458154 493434
rect 457918 486198 458154 486434
rect 457918 479198 458154 479434
rect 457918 472198 458154 472434
rect 457918 465198 458154 465434
rect 457918 458198 458154 458434
rect 457918 451198 458154 451434
rect 457918 444198 458154 444434
rect 457918 437198 458154 437434
rect 457918 430198 458154 430434
rect 457918 423198 458154 423434
rect 457918 416198 458154 416434
rect 457918 409198 458154 409434
rect 457918 402198 458154 402434
rect 457918 395198 458154 395434
rect 457918 388198 458154 388434
rect 457918 381198 458154 381434
rect 457918 374198 458154 374434
rect 457918 367198 458154 367434
rect 457918 360198 458154 360434
rect 457918 353198 458154 353434
rect 457918 346198 458154 346434
rect 457918 339198 458154 339434
rect 457918 332198 458154 332434
rect 457918 325198 458154 325434
rect 457918 318198 458154 318434
rect 457918 311198 458154 311434
rect 457918 304198 458154 304434
rect 457918 297198 458154 297434
rect 457918 290198 458154 290434
rect 457918 283198 458154 283434
rect 457918 276198 458154 276434
rect 457918 269198 458154 269434
rect 457918 262198 458154 262434
rect 457918 255198 458154 255434
rect 457918 248198 458154 248434
rect 457918 241198 458154 241434
rect 457918 234198 458154 234434
rect 457918 227198 458154 227434
rect 457918 220198 458154 220434
rect 457918 213198 458154 213434
rect 457918 206198 458154 206434
rect 457918 199198 458154 199434
rect 457918 192198 458154 192434
rect 457918 185198 458154 185434
rect 457918 178198 458154 178434
rect 457918 171198 458154 171434
rect 457918 164198 458154 164434
rect 457918 157198 458154 157434
rect 457918 150198 458154 150434
rect 457918 143198 458154 143434
rect 457918 136198 458154 136434
rect 457918 129198 458154 129434
rect 457918 122198 458154 122434
rect 457918 115198 458154 115434
rect 457918 108198 458154 108434
rect 457918 101198 458154 101434
rect 457918 94198 458154 94434
rect 457918 87198 458154 87434
rect 457918 80198 458154 80434
rect 457918 73198 458154 73434
rect 457918 66198 458154 66434
rect 457918 59198 458154 59434
rect 457918 52198 458154 52434
rect 457918 45198 458154 45434
rect 457918 38198 458154 38434
rect 457918 31198 458154 31434
rect 457918 24198 458154 24434
rect 457918 17198 458154 17434
rect 457918 10198 458154 10434
rect 457918 3198 458154 3434
rect 457918 -1942 458154 -1706
rect 457918 -2262 458154 -2026
rect 463186 705002 463422 705238
rect 463186 704682 463422 704918
rect 463186 695258 463422 695494
rect 463186 688258 463422 688494
rect 463186 681258 463422 681494
rect 463186 674258 463422 674494
rect 463186 667258 463422 667494
rect 463186 660258 463422 660494
rect 463186 653258 463422 653494
rect 463186 646258 463422 646494
rect 463186 639258 463422 639494
rect 463186 632258 463422 632494
rect 463186 625258 463422 625494
rect 463186 618258 463422 618494
rect 463186 611258 463422 611494
rect 463186 604258 463422 604494
rect 463186 597258 463422 597494
rect 463186 590258 463422 590494
rect 463186 583258 463422 583494
rect 463186 576258 463422 576494
rect 463186 569258 463422 569494
rect 463186 562258 463422 562494
rect 463186 555258 463422 555494
rect 463186 548258 463422 548494
rect 463186 541258 463422 541494
rect 463186 534258 463422 534494
rect 463186 527258 463422 527494
rect 463186 520258 463422 520494
rect 463186 513258 463422 513494
rect 463186 506258 463422 506494
rect 463186 499258 463422 499494
rect 463186 492258 463422 492494
rect 463186 485258 463422 485494
rect 463186 478258 463422 478494
rect 463186 471258 463422 471494
rect 463186 464258 463422 464494
rect 463186 457258 463422 457494
rect 463186 450258 463422 450494
rect 463186 443258 463422 443494
rect 463186 436258 463422 436494
rect 463186 429258 463422 429494
rect 463186 422258 463422 422494
rect 463186 415258 463422 415494
rect 463186 408258 463422 408494
rect 463186 401258 463422 401494
rect 463186 394258 463422 394494
rect 463186 387258 463422 387494
rect 463186 380258 463422 380494
rect 463186 373258 463422 373494
rect 463186 366258 463422 366494
rect 463186 359258 463422 359494
rect 463186 352258 463422 352494
rect 463186 345258 463422 345494
rect 463186 338258 463422 338494
rect 463186 331258 463422 331494
rect 463186 324258 463422 324494
rect 463186 317258 463422 317494
rect 463186 310258 463422 310494
rect 463186 303258 463422 303494
rect 463186 296258 463422 296494
rect 463186 289258 463422 289494
rect 463186 282258 463422 282494
rect 463186 275258 463422 275494
rect 463186 268258 463422 268494
rect 463186 261258 463422 261494
rect 463186 254258 463422 254494
rect 463186 247258 463422 247494
rect 463186 240258 463422 240494
rect 463186 233258 463422 233494
rect 463186 226258 463422 226494
rect 463186 219258 463422 219494
rect 463186 212258 463422 212494
rect 463186 205258 463422 205494
rect 463186 198258 463422 198494
rect 463186 191258 463422 191494
rect 463186 184258 463422 184494
rect 463186 177258 463422 177494
rect 463186 170258 463422 170494
rect 463186 163258 463422 163494
rect 463186 156258 463422 156494
rect 463186 149258 463422 149494
rect 463186 142258 463422 142494
rect 463186 135258 463422 135494
rect 463186 128258 463422 128494
rect 463186 121258 463422 121494
rect 463186 114258 463422 114494
rect 463186 107258 463422 107494
rect 463186 100258 463422 100494
rect 463186 93258 463422 93494
rect 463186 86258 463422 86494
rect 463186 79258 463422 79494
rect 463186 72258 463422 72494
rect 463186 65258 463422 65494
rect 463186 58258 463422 58494
rect 463186 51258 463422 51494
rect 463186 44258 463422 44494
rect 463186 37258 463422 37494
rect 463186 30258 463422 30494
rect 463186 23258 463422 23494
rect 463186 16258 463422 16494
rect 463186 9258 463422 9494
rect 463186 2258 463422 2494
rect 463186 -982 463422 -746
rect 463186 -1302 463422 -1066
rect 464918 705962 465154 706198
rect 464918 705642 465154 705878
rect 464918 696198 465154 696434
rect 464918 689198 465154 689434
rect 464918 682198 465154 682434
rect 464918 675198 465154 675434
rect 464918 668198 465154 668434
rect 464918 661198 465154 661434
rect 464918 654198 465154 654434
rect 464918 647198 465154 647434
rect 464918 640198 465154 640434
rect 464918 633198 465154 633434
rect 464918 626198 465154 626434
rect 464918 619198 465154 619434
rect 464918 612198 465154 612434
rect 464918 605198 465154 605434
rect 464918 598198 465154 598434
rect 464918 591198 465154 591434
rect 464918 584198 465154 584434
rect 464918 577198 465154 577434
rect 464918 570198 465154 570434
rect 464918 563198 465154 563434
rect 464918 556198 465154 556434
rect 464918 549198 465154 549434
rect 464918 542198 465154 542434
rect 464918 535198 465154 535434
rect 464918 528198 465154 528434
rect 464918 521198 465154 521434
rect 464918 514198 465154 514434
rect 464918 507198 465154 507434
rect 464918 500198 465154 500434
rect 464918 493198 465154 493434
rect 464918 486198 465154 486434
rect 464918 479198 465154 479434
rect 464918 472198 465154 472434
rect 464918 465198 465154 465434
rect 464918 458198 465154 458434
rect 464918 451198 465154 451434
rect 464918 444198 465154 444434
rect 464918 437198 465154 437434
rect 464918 430198 465154 430434
rect 464918 423198 465154 423434
rect 464918 416198 465154 416434
rect 464918 409198 465154 409434
rect 464918 402198 465154 402434
rect 464918 395198 465154 395434
rect 464918 388198 465154 388434
rect 464918 381198 465154 381434
rect 464918 374198 465154 374434
rect 464918 367198 465154 367434
rect 464918 360198 465154 360434
rect 464918 353198 465154 353434
rect 464918 346198 465154 346434
rect 464918 339198 465154 339434
rect 464918 332198 465154 332434
rect 464918 325198 465154 325434
rect 464918 318198 465154 318434
rect 464918 311198 465154 311434
rect 464918 304198 465154 304434
rect 464918 297198 465154 297434
rect 464918 290198 465154 290434
rect 464918 283198 465154 283434
rect 464918 276198 465154 276434
rect 464918 269198 465154 269434
rect 464918 262198 465154 262434
rect 464918 255198 465154 255434
rect 464918 248198 465154 248434
rect 464918 241198 465154 241434
rect 464918 234198 465154 234434
rect 464918 227198 465154 227434
rect 464918 220198 465154 220434
rect 464918 213198 465154 213434
rect 464918 206198 465154 206434
rect 464918 199198 465154 199434
rect 464918 192198 465154 192434
rect 464918 185198 465154 185434
rect 464918 178198 465154 178434
rect 464918 171198 465154 171434
rect 464918 164198 465154 164434
rect 464918 157198 465154 157434
rect 464918 150198 465154 150434
rect 464918 143198 465154 143434
rect 464918 136198 465154 136434
rect 464918 129198 465154 129434
rect 464918 122198 465154 122434
rect 464918 115198 465154 115434
rect 464918 108198 465154 108434
rect 464918 101198 465154 101434
rect 464918 94198 465154 94434
rect 464918 87198 465154 87434
rect 464918 80198 465154 80434
rect 464918 73198 465154 73434
rect 464918 66198 465154 66434
rect 464918 59198 465154 59434
rect 464918 52198 465154 52434
rect 464918 45198 465154 45434
rect 464918 38198 465154 38434
rect 464918 31198 465154 31434
rect 464918 24198 465154 24434
rect 464918 17198 465154 17434
rect 464918 10198 465154 10434
rect 464918 3198 465154 3434
rect 464918 -1942 465154 -1706
rect 464918 -2262 465154 -2026
rect 470186 705002 470422 705238
rect 470186 704682 470422 704918
rect 470186 695258 470422 695494
rect 470186 688258 470422 688494
rect 470186 681258 470422 681494
rect 470186 674258 470422 674494
rect 470186 667258 470422 667494
rect 470186 660258 470422 660494
rect 470186 653258 470422 653494
rect 470186 646258 470422 646494
rect 470186 639258 470422 639494
rect 470186 632258 470422 632494
rect 470186 625258 470422 625494
rect 470186 618258 470422 618494
rect 470186 611258 470422 611494
rect 470186 604258 470422 604494
rect 470186 597258 470422 597494
rect 470186 590258 470422 590494
rect 470186 583258 470422 583494
rect 470186 576258 470422 576494
rect 470186 569258 470422 569494
rect 470186 562258 470422 562494
rect 470186 555258 470422 555494
rect 470186 548258 470422 548494
rect 470186 541258 470422 541494
rect 470186 534258 470422 534494
rect 470186 527258 470422 527494
rect 470186 520258 470422 520494
rect 470186 513258 470422 513494
rect 470186 506258 470422 506494
rect 470186 499258 470422 499494
rect 470186 492258 470422 492494
rect 470186 485258 470422 485494
rect 470186 478258 470422 478494
rect 470186 471258 470422 471494
rect 470186 464258 470422 464494
rect 470186 457258 470422 457494
rect 470186 450258 470422 450494
rect 470186 443258 470422 443494
rect 470186 436258 470422 436494
rect 470186 429258 470422 429494
rect 470186 422258 470422 422494
rect 470186 415258 470422 415494
rect 470186 408258 470422 408494
rect 470186 401258 470422 401494
rect 470186 394258 470422 394494
rect 470186 387258 470422 387494
rect 470186 380258 470422 380494
rect 470186 373258 470422 373494
rect 470186 366258 470422 366494
rect 470186 359258 470422 359494
rect 470186 352258 470422 352494
rect 470186 345258 470422 345494
rect 470186 338258 470422 338494
rect 470186 331258 470422 331494
rect 470186 324258 470422 324494
rect 470186 317258 470422 317494
rect 470186 310258 470422 310494
rect 470186 303258 470422 303494
rect 470186 296258 470422 296494
rect 470186 289258 470422 289494
rect 470186 282258 470422 282494
rect 470186 275258 470422 275494
rect 470186 268258 470422 268494
rect 470186 261258 470422 261494
rect 470186 254258 470422 254494
rect 470186 247258 470422 247494
rect 470186 240258 470422 240494
rect 470186 233258 470422 233494
rect 470186 226258 470422 226494
rect 470186 219258 470422 219494
rect 470186 212258 470422 212494
rect 470186 205258 470422 205494
rect 470186 198258 470422 198494
rect 470186 191258 470422 191494
rect 470186 184258 470422 184494
rect 470186 177258 470422 177494
rect 470186 170258 470422 170494
rect 470186 163258 470422 163494
rect 470186 156258 470422 156494
rect 470186 149258 470422 149494
rect 470186 142258 470422 142494
rect 470186 135258 470422 135494
rect 470186 128258 470422 128494
rect 470186 121258 470422 121494
rect 470186 114258 470422 114494
rect 470186 107258 470422 107494
rect 470186 100258 470422 100494
rect 470186 93258 470422 93494
rect 470186 86258 470422 86494
rect 470186 79258 470422 79494
rect 470186 72258 470422 72494
rect 470186 65258 470422 65494
rect 470186 58258 470422 58494
rect 470186 51258 470422 51494
rect 470186 44258 470422 44494
rect 470186 37258 470422 37494
rect 470186 30258 470422 30494
rect 470186 23258 470422 23494
rect 470186 16258 470422 16494
rect 470186 9258 470422 9494
rect 470186 2258 470422 2494
rect 470186 -982 470422 -746
rect 470186 -1302 470422 -1066
rect 471918 705962 472154 706198
rect 471918 705642 472154 705878
rect 471918 696198 472154 696434
rect 471918 689198 472154 689434
rect 471918 682198 472154 682434
rect 471918 675198 472154 675434
rect 471918 668198 472154 668434
rect 471918 661198 472154 661434
rect 471918 654198 472154 654434
rect 471918 647198 472154 647434
rect 471918 640198 472154 640434
rect 471918 633198 472154 633434
rect 471918 626198 472154 626434
rect 471918 619198 472154 619434
rect 471918 612198 472154 612434
rect 471918 605198 472154 605434
rect 471918 598198 472154 598434
rect 471918 591198 472154 591434
rect 471918 584198 472154 584434
rect 471918 577198 472154 577434
rect 471918 570198 472154 570434
rect 471918 563198 472154 563434
rect 471918 556198 472154 556434
rect 471918 549198 472154 549434
rect 471918 542198 472154 542434
rect 471918 535198 472154 535434
rect 471918 528198 472154 528434
rect 471918 521198 472154 521434
rect 471918 514198 472154 514434
rect 471918 507198 472154 507434
rect 471918 500198 472154 500434
rect 471918 493198 472154 493434
rect 471918 486198 472154 486434
rect 471918 479198 472154 479434
rect 471918 472198 472154 472434
rect 471918 465198 472154 465434
rect 471918 458198 472154 458434
rect 471918 451198 472154 451434
rect 471918 444198 472154 444434
rect 471918 437198 472154 437434
rect 471918 430198 472154 430434
rect 471918 423198 472154 423434
rect 471918 416198 472154 416434
rect 471918 409198 472154 409434
rect 471918 402198 472154 402434
rect 471918 395198 472154 395434
rect 471918 388198 472154 388434
rect 471918 381198 472154 381434
rect 471918 374198 472154 374434
rect 471918 367198 472154 367434
rect 471918 360198 472154 360434
rect 471918 353198 472154 353434
rect 471918 346198 472154 346434
rect 471918 339198 472154 339434
rect 471918 332198 472154 332434
rect 471918 325198 472154 325434
rect 471918 318198 472154 318434
rect 471918 311198 472154 311434
rect 471918 304198 472154 304434
rect 471918 297198 472154 297434
rect 471918 290198 472154 290434
rect 471918 283198 472154 283434
rect 471918 276198 472154 276434
rect 471918 269198 472154 269434
rect 471918 262198 472154 262434
rect 471918 255198 472154 255434
rect 471918 248198 472154 248434
rect 471918 241198 472154 241434
rect 471918 234198 472154 234434
rect 471918 227198 472154 227434
rect 471918 220198 472154 220434
rect 471918 213198 472154 213434
rect 471918 206198 472154 206434
rect 471918 199198 472154 199434
rect 471918 192198 472154 192434
rect 471918 185198 472154 185434
rect 471918 178198 472154 178434
rect 471918 171198 472154 171434
rect 471918 164198 472154 164434
rect 471918 157198 472154 157434
rect 471918 150198 472154 150434
rect 471918 143198 472154 143434
rect 471918 136198 472154 136434
rect 471918 129198 472154 129434
rect 471918 122198 472154 122434
rect 471918 115198 472154 115434
rect 471918 108198 472154 108434
rect 471918 101198 472154 101434
rect 471918 94198 472154 94434
rect 471918 87198 472154 87434
rect 471918 80198 472154 80434
rect 471918 73198 472154 73434
rect 471918 66198 472154 66434
rect 471918 59198 472154 59434
rect 471918 52198 472154 52434
rect 471918 45198 472154 45434
rect 471918 38198 472154 38434
rect 471918 31198 472154 31434
rect 471918 24198 472154 24434
rect 471918 17198 472154 17434
rect 471918 10198 472154 10434
rect 471918 3198 472154 3434
rect 471918 -1942 472154 -1706
rect 471918 -2262 472154 -2026
rect 477186 705002 477422 705238
rect 477186 704682 477422 704918
rect 477186 695258 477422 695494
rect 477186 688258 477422 688494
rect 477186 681258 477422 681494
rect 477186 674258 477422 674494
rect 477186 667258 477422 667494
rect 477186 660258 477422 660494
rect 477186 653258 477422 653494
rect 477186 646258 477422 646494
rect 477186 639258 477422 639494
rect 477186 632258 477422 632494
rect 477186 625258 477422 625494
rect 477186 618258 477422 618494
rect 477186 611258 477422 611494
rect 477186 604258 477422 604494
rect 477186 597258 477422 597494
rect 477186 590258 477422 590494
rect 477186 583258 477422 583494
rect 477186 576258 477422 576494
rect 477186 569258 477422 569494
rect 477186 562258 477422 562494
rect 477186 555258 477422 555494
rect 477186 548258 477422 548494
rect 477186 541258 477422 541494
rect 477186 534258 477422 534494
rect 477186 527258 477422 527494
rect 477186 520258 477422 520494
rect 477186 513258 477422 513494
rect 477186 506258 477422 506494
rect 477186 499258 477422 499494
rect 477186 492258 477422 492494
rect 477186 485258 477422 485494
rect 477186 478258 477422 478494
rect 477186 471258 477422 471494
rect 477186 464258 477422 464494
rect 477186 457258 477422 457494
rect 477186 450258 477422 450494
rect 477186 443258 477422 443494
rect 477186 436258 477422 436494
rect 477186 429258 477422 429494
rect 477186 422258 477422 422494
rect 477186 415258 477422 415494
rect 477186 408258 477422 408494
rect 477186 401258 477422 401494
rect 477186 394258 477422 394494
rect 477186 387258 477422 387494
rect 477186 380258 477422 380494
rect 477186 373258 477422 373494
rect 477186 366258 477422 366494
rect 477186 359258 477422 359494
rect 477186 352258 477422 352494
rect 477186 345258 477422 345494
rect 477186 338258 477422 338494
rect 477186 331258 477422 331494
rect 477186 324258 477422 324494
rect 477186 317258 477422 317494
rect 477186 310258 477422 310494
rect 477186 303258 477422 303494
rect 477186 296258 477422 296494
rect 477186 289258 477422 289494
rect 477186 282258 477422 282494
rect 477186 275258 477422 275494
rect 477186 268258 477422 268494
rect 477186 261258 477422 261494
rect 477186 254258 477422 254494
rect 477186 247258 477422 247494
rect 477186 240258 477422 240494
rect 477186 233258 477422 233494
rect 477186 226258 477422 226494
rect 477186 219258 477422 219494
rect 477186 212258 477422 212494
rect 477186 205258 477422 205494
rect 477186 198258 477422 198494
rect 477186 191258 477422 191494
rect 477186 184258 477422 184494
rect 477186 177258 477422 177494
rect 477186 170258 477422 170494
rect 477186 163258 477422 163494
rect 477186 156258 477422 156494
rect 477186 149258 477422 149494
rect 477186 142258 477422 142494
rect 477186 135258 477422 135494
rect 477186 128258 477422 128494
rect 477186 121258 477422 121494
rect 477186 114258 477422 114494
rect 477186 107258 477422 107494
rect 477186 100258 477422 100494
rect 477186 93258 477422 93494
rect 477186 86258 477422 86494
rect 477186 79258 477422 79494
rect 477186 72258 477422 72494
rect 477186 65258 477422 65494
rect 477186 58258 477422 58494
rect 477186 51258 477422 51494
rect 477186 44258 477422 44494
rect 477186 37258 477422 37494
rect 477186 30258 477422 30494
rect 477186 23258 477422 23494
rect 477186 16258 477422 16494
rect 477186 9258 477422 9494
rect 477186 2258 477422 2494
rect 477186 -982 477422 -746
rect 477186 -1302 477422 -1066
rect 478918 705962 479154 706198
rect 478918 705642 479154 705878
rect 478918 696198 479154 696434
rect 478918 689198 479154 689434
rect 478918 682198 479154 682434
rect 478918 675198 479154 675434
rect 478918 668198 479154 668434
rect 478918 661198 479154 661434
rect 478918 654198 479154 654434
rect 478918 647198 479154 647434
rect 478918 640198 479154 640434
rect 478918 633198 479154 633434
rect 478918 626198 479154 626434
rect 478918 619198 479154 619434
rect 478918 612198 479154 612434
rect 478918 605198 479154 605434
rect 478918 598198 479154 598434
rect 478918 591198 479154 591434
rect 478918 584198 479154 584434
rect 478918 577198 479154 577434
rect 478918 570198 479154 570434
rect 478918 563198 479154 563434
rect 478918 556198 479154 556434
rect 478918 549198 479154 549434
rect 478918 542198 479154 542434
rect 478918 535198 479154 535434
rect 478918 528198 479154 528434
rect 478918 521198 479154 521434
rect 478918 514198 479154 514434
rect 478918 507198 479154 507434
rect 478918 500198 479154 500434
rect 478918 493198 479154 493434
rect 478918 486198 479154 486434
rect 478918 479198 479154 479434
rect 478918 472198 479154 472434
rect 478918 465198 479154 465434
rect 478918 458198 479154 458434
rect 478918 451198 479154 451434
rect 478918 444198 479154 444434
rect 478918 437198 479154 437434
rect 478918 430198 479154 430434
rect 478918 423198 479154 423434
rect 478918 416198 479154 416434
rect 478918 409198 479154 409434
rect 478918 402198 479154 402434
rect 478918 395198 479154 395434
rect 478918 388198 479154 388434
rect 478918 381198 479154 381434
rect 478918 374198 479154 374434
rect 478918 367198 479154 367434
rect 478918 360198 479154 360434
rect 478918 353198 479154 353434
rect 478918 346198 479154 346434
rect 478918 339198 479154 339434
rect 478918 332198 479154 332434
rect 478918 325198 479154 325434
rect 478918 318198 479154 318434
rect 478918 311198 479154 311434
rect 478918 304198 479154 304434
rect 478918 297198 479154 297434
rect 478918 290198 479154 290434
rect 478918 283198 479154 283434
rect 478918 276198 479154 276434
rect 478918 269198 479154 269434
rect 478918 262198 479154 262434
rect 478918 255198 479154 255434
rect 478918 248198 479154 248434
rect 478918 241198 479154 241434
rect 478918 234198 479154 234434
rect 478918 227198 479154 227434
rect 478918 220198 479154 220434
rect 478918 213198 479154 213434
rect 478918 206198 479154 206434
rect 478918 199198 479154 199434
rect 478918 192198 479154 192434
rect 478918 185198 479154 185434
rect 478918 178198 479154 178434
rect 478918 171198 479154 171434
rect 478918 164198 479154 164434
rect 478918 157198 479154 157434
rect 478918 150198 479154 150434
rect 478918 143198 479154 143434
rect 478918 136198 479154 136434
rect 478918 129198 479154 129434
rect 478918 122198 479154 122434
rect 478918 115198 479154 115434
rect 478918 108198 479154 108434
rect 478918 101198 479154 101434
rect 478918 94198 479154 94434
rect 478918 87198 479154 87434
rect 478918 80198 479154 80434
rect 478918 73198 479154 73434
rect 478918 66198 479154 66434
rect 478918 59198 479154 59434
rect 478918 52198 479154 52434
rect 478918 45198 479154 45434
rect 478918 38198 479154 38434
rect 478918 31198 479154 31434
rect 478918 24198 479154 24434
rect 478918 17198 479154 17434
rect 478918 10198 479154 10434
rect 478918 3198 479154 3434
rect 478918 -1942 479154 -1706
rect 478918 -2262 479154 -2026
rect 484186 705002 484422 705238
rect 484186 704682 484422 704918
rect 484186 695258 484422 695494
rect 484186 688258 484422 688494
rect 484186 681258 484422 681494
rect 484186 674258 484422 674494
rect 484186 667258 484422 667494
rect 484186 660258 484422 660494
rect 484186 653258 484422 653494
rect 484186 646258 484422 646494
rect 484186 639258 484422 639494
rect 484186 632258 484422 632494
rect 484186 625258 484422 625494
rect 484186 618258 484422 618494
rect 484186 611258 484422 611494
rect 484186 604258 484422 604494
rect 484186 597258 484422 597494
rect 484186 590258 484422 590494
rect 484186 583258 484422 583494
rect 484186 576258 484422 576494
rect 484186 569258 484422 569494
rect 484186 562258 484422 562494
rect 484186 555258 484422 555494
rect 484186 548258 484422 548494
rect 484186 541258 484422 541494
rect 484186 534258 484422 534494
rect 484186 527258 484422 527494
rect 484186 520258 484422 520494
rect 484186 513258 484422 513494
rect 484186 506258 484422 506494
rect 484186 499258 484422 499494
rect 484186 492258 484422 492494
rect 484186 485258 484422 485494
rect 484186 478258 484422 478494
rect 484186 471258 484422 471494
rect 484186 464258 484422 464494
rect 484186 457258 484422 457494
rect 484186 450258 484422 450494
rect 484186 443258 484422 443494
rect 484186 436258 484422 436494
rect 484186 429258 484422 429494
rect 484186 422258 484422 422494
rect 484186 415258 484422 415494
rect 484186 408258 484422 408494
rect 484186 401258 484422 401494
rect 484186 394258 484422 394494
rect 484186 387258 484422 387494
rect 484186 380258 484422 380494
rect 484186 373258 484422 373494
rect 484186 366258 484422 366494
rect 484186 359258 484422 359494
rect 484186 352258 484422 352494
rect 484186 345258 484422 345494
rect 484186 338258 484422 338494
rect 484186 331258 484422 331494
rect 484186 324258 484422 324494
rect 484186 317258 484422 317494
rect 484186 310258 484422 310494
rect 484186 303258 484422 303494
rect 484186 296258 484422 296494
rect 484186 289258 484422 289494
rect 484186 282258 484422 282494
rect 484186 275258 484422 275494
rect 484186 268258 484422 268494
rect 484186 261258 484422 261494
rect 484186 254258 484422 254494
rect 484186 247258 484422 247494
rect 484186 240258 484422 240494
rect 484186 233258 484422 233494
rect 484186 226258 484422 226494
rect 484186 219258 484422 219494
rect 484186 212258 484422 212494
rect 484186 205258 484422 205494
rect 484186 198258 484422 198494
rect 484186 191258 484422 191494
rect 484186 184258 484422 184494
rect 484186 177258 484422 177494
rect 484186 170258 484422 170494
rect 484186 163258 484422 163494
rect 484186 156258 484422 156494
rect 484186 149258 484422 149494
rect 484186 142258 484422 142494
rect 484186 135258 484422 135494
rect 484186 128258 484422 128494
rect 484186 121258 484422 121494
rect 484186 114258 484422 114494
rect 484186 107258 484422 107494
rect 484186 100258 484422 100494
rect 484186 93258 484422 93494
rect 484186 86258 484422 86494
rect 484186 79258 484422 79494
rect 484186 72258 484422 72494
rect 484186 65258 484422 65494
rect 484186 58258 484422 58494
rect 484186 51258 484422 51494
rect 484186 44258 484422 44494
rect 484186 37258 484422 37494
rect 484186 30258 484422 30494
rect 484186 23258 484422 23494
rect 484186 16258 484422 16494
rect 484186 9258 484422 9494
rect 484186 2258 484422 2494
rect 484186 -982 484422 -746
rect 484186 -1302 484422 -1066
rect 485918 705962 486154 706198
rect 485918 705642 486154 705878
rect 485918 696198 486154 696434
rect 485918 689198 486154 689434
rect 485918 682198 486154 682434
rect 485918 675198 486154 675434
rect 485918 668198 486154 668434
rect 485918 661198 486154 661434
rect 485918 654198 486154 654434
rect 485918 647198 486154 647434
rect 485918 640198 486154 640434
rect 485918 633198 486154 633434
rect 485918 626198 486154 626434
rect 485918 619198 486154 619434
rect 485918 612198 486154 612434
rect 485918 605198 486154 605434
rect 485918 598198 486154 598434
rect 485918 591198 486154 591434
rect 485918 584198 486154 584434
rect 485918 577198 486154 577434
rect 485918 570198 486154 570434
rect 485918 563198 486154 563434
rect 485918 556198 486154 556434
rect 485918 549198 486154 549434
rect 485918 542198 486154 542434
rect 485918 535198 486154 535434
rect 485918 528198 486154 528434
rect 485918 521198 486154 521434
rect 485918 514198 486154 514434
rect 485918 507198 486154 507434
rect 485918 500198 486154 500434
rect 485918 493198 486154 493434
rect 485918 486198 486154 486434
rect 485918 479198 486154 479434
rect 485918 472198 486154 472434
rect 485918 465198 486154 465434
rect 485918 458198 486154 458434
rect 485918 451198 486154 451434
rect 485918 444198 486154 444434
rect 485918 437198 486154 437434
rect 485918 430198 486154 430434
rect 485918 423198 486154 423434
rect 485918 416198 486154 416434
rect 485918 409198 486154 409434
rect 485918 402198 486154 402434
rect 485918 395198 486154 395434
rect 485918 388198 486154 388434
rect 485918 381198 486154 381434
rect 485918 374198 486154 374434
rect 485918 367198 486154 367434
rect 485918 360198 486154 360434
rect 485918 353198 486154 353434
rect 485918 346198 486154 346434
rect 485918 339198 486154 339434
rect 485918 332198 486154 332434
rect 485918 325198 486154 325434
rect 485918 318198 486154 318434
rect 485918 311198 486154 311434
rect 485918 304198 486154 304434
rect 485918 297198 486154 297434
rect 485918 290198 486154 290434
rect 485918 283198 486154 283434
rect 485918 276198 486154 276434
rect 485918 269198 486154 269434
rect 485918 262198 486154 262434
rect 485918 255198 486154 255434
rect 485918 248198 486154 248434
rect 485918 241198 486154 241434
rect 485918 234198 486154 234434
rect 485918 227198 486154 227434
rect 485918 220198 486154 220434
rect 485918 213198 486154 213434
rect 485918 206198 486154 206434
rect 485918 199198 486154 199434
rect 485918 192198 486154 192434
rect 485918 185198 486154 185434
rect 485918 178198 486154 178434
rect 485918 171198 486154 171434
rect 485918 164198 486154 164434
rect 485918 157198 486154 157434
rect 485918 150198 486154 150434
rect 485918 143198 486154 143434
rect 485918 136198 486154 136434
rect 485918 129198 486154 129434
rect 485918 122198 486154 122434
rect 485918 115198 486154 115434
rect 485918 108198 486154 108434
rect 485918 101198 486154 101434
rect 485918 94198 486154 94434
rect 485918 87198 486154 87434
rect 485918 80198 486154 80434
rect 485918 73198 486154 73434
rect 485918 66198 486154 66434
rect 485918 59198 486154 59434
rect 485918 52198 486154 52434
rect 485918 45198 486154 45434
rect 485918 38198 486154 38434
rect 485918 31198 486154 31434
rect 485918 24198 486154 24434
rect 485918 17198 486154 17434
rect 485918 10198 486154 10434
rect 485918 3198 486154 3434
rect 485918 -1942 486154 -1706
rect 485918 -2262 486154 -2026
rect 491186 705002 491422 705238
rect 491186 704682 491422 704918
rect 491186 695258 491422 695494
rect 491186 688258 491422 688494
rect 491186 681258 491422 681494
rect 491186 674258 491422 674494
rect 491186 667258 491422 667494
rect 491186 660258 491422 660494
rect 491186 653258 491422 653494
rect 491186 646258 491422 646494
rect 491186 639258 491422 639494
rect 491186 632258 491422 632494
rect 491186 625258 491422 625494
rect 491186 618258 491422 618494
rect 491186 611258 491422 611494
rect 491186 604258 491422 604494
rect 491186 597258 491422 597494
rect 491186 590258 491422 590494
rect 491186 583258 491422 583494
rect 491186 576258 491422 576494
rect 491186 569258 491422 569494
rect 491186 562258 491422 562494
rect 491186 555258 491422 555494
rect 491186 548258 491422 548494
rect 491186 541258 491422 541494
rect 491186 534258 491422 534494
rect 491186 527258 491422 527494
rect 491186 520258 491422 520494
rect 491186 513258 491422 513494
rect 491186 506258 491422 506494
rect 491186 499258 491422 499494
rect 491186 492258 491422 492494
rect 491186 485258 491422 485494
rect 491186 478258 491422 478494
rect 491186 471258 491422 471494
rect 491186 464258 491422 464494
rect 491186 457258 491422 457494
rect 491186 450258 491422 450494
rect 491186 443258 491422 443494
rect 491186 436258 491422 436494
rect 491186 429258 491422 429494
rect 491186 422258 491422 422494
rect 491186 415258 491422 415494
rect 491186 408258 491422 408494
rect 491186 401258 491422 401494
rect 491186 394258 491422 394494
rect 491186 387258 491422 387494
rect 491186 380258 491422 380494
rect 491186 373258 491422 373494
rect 491186 366258 491422 366494
rect 491186 359258 491422 359494
rect 491186 352258 491422 352494
rect 491186 345258 491422 345494
rect 491186 338258 491422 338494
rect 491186 331258 491422 331494
rect 491186 324258 491422 324494
rect 491186 317258 491422 317494
rect 491186 310258 491422 310494
rect 491186 303258 491422 303494
rect 491186 296258 491422 296494
rect 491186 289258 491422 289494
rect 491186 282258 491422 282494
rect 491186 275258 491422 275494
rect 491186 268258 491422 268494
rect 491186 261258 491422 261494
rect 491186 254258 491422 254494
rect 491186 247258 491422 247494
rect 491186 240258 491422 240494
rect 491186 233258 491422 233494
rect 491186 226258 491422 226494
rect 491186 219258 491422 219494
rect 491186 212258 491422 212494
rect 491186 205258 491422 205494
rect 491186 198258 491422 198494
rect 491186 191258 491422 191494
rect 491186 184258 491422 184494
rect 491186 177258 491422 177494
rect 491186 170258 491422 170494
rect 491186 163258 491422 163494
rect 491186 156258 491422 156494
rect 491186 149258 491422 149494
rect 491186 142258 491422 142494
rect 491186 135258 491422 135494
rect 491186 128258 491422 128494
rect 491186 121258 491422 121494
rect 491186 114258 491422 114494
rect 491186 107258 491422 107494
rect 491186 100258 491422 100494
rect 491186 93258 491422 93494
rect 491186 86258 491422 86494
rect 491186 79258 491422 79494
rect 491186 72258 491422 72494
rect 491186 65258 491422 65494
rect 491186 58258 491422 58494
rect 491186 51258 491422 51494
rect 491186 44258 491422 44494
rect 491186 37258 491422 37494
rect 491186 30258 491422 30494
rect 491186 23258 491422 23494
rect 491186 16258 491422 16494
rect 491186 9258 491422 9494
rect 491186 2258 491422 2494
rect 491186 -982 491422 -746
rect 491186 -1302 491422 -1066
rect 492918 705962 493154 706198
rect 492918 705642 493154 705878
rect 492918 696198 493154 696434
rect 492918 689198 493154 689434
rect 492918 682198 493154 682434
rect 492918 675198 493154 675434
rect 492918 668198 493154 668434
rect 492918 661198 493154 661434
rect 492918 654198 493154 654434
rect 492918 647198 493154 647434
rect 492918 640198 493154 640434
rect 492918 633198 493154 633434
rect 492918 626198 493154 626434
rect 492918 619198 493154 619434
rect 492918 612198 493154 612434
rect 492918 605198 493154 605434
rect 492918 598198 493154 598434
rect 492918 591198 493154 591434
rect 492918 584198 493154 584434
rect 492918 577198 493154 577434
rect 492918 570198 493154 570434
rect 492918 563198 493154 563434
rect 492918 556198 493154 556434
rect 492918 549198 493154 549434
rect 492918 542198 493154 542434
rect 492918 535198 493154 535434
rect 492918 528198 493154 528434
rect 492918 521198 493154 521434
rect 492918 514198 493154 514434
rect 492918 507198 493154 507434
rect 492918 500198 493154 500434
rect 492918 493198 493154 493434
rect 492918 486198 493154 486434
rect 492918 479198 493154 479434
rect 492918 472198 493154 472434
rect 492918 465198 493154 465434
rect 492918 458198 493154 458434
rect 492918 451198 493154 451434
rect 492918 444198 493154 444434
rect 492918 437198 493154 437434
rect 492918 430198 493154 430434
rect 492918 423198 493154 423434
rect 492918 416198 493154 416434
rect 492918 409198 493154 409434
rect 492918 402198 493154 402434
rect 492918 395198 493154 395434
rect 492918 388198 493154 388434
rect 492918 381198 493154 381434
rect 492918 374198 493154 374434
rect 492918 367198 493154 367434
rect 492918 360198 493154 360434
rect 492918 353198 493154 353434
rect 492918 346198 493154 346434
rect 492918 339198 493154 339434
rect 492918 332198 493154 332434
rect 492918 325198 493154 325434
rect 492918 318198 493154 318434
rect 492918 311198 493154 311434
rect 492918 304198 493154 304434
rect 492918 297198 493154 297434
rect 492918 290198 493154 290434
rect 492918 283198 493154 283434
rect 492918 276198 493154 276434
rect 492918 269198 493154 269434
rect 492918 262198 493154 262434
rect 492918 255198 493154 255434
rect 492918 248198 493154 248434
rect 492918 241198 493154 241434
rect 492918 234198 493154 234434
rect 492918 227198 493154 227434
rect 492918 220198 493154 220434
rect 492918 213198 493154 213434
rect 492918 206198 493154 206434
rect 492918 199198 493154 199434
rect 492918 192198 493154 192434
rect 492918 185198 493154 185434
rect 492918 178198 493154 178434
rect 492918 171198 493154 171434
rect 492918 164198 493154 164434
rect 492918 157198 493154 157434
rect 492918 150198 493154 150434
rect 492918 143198 493154 143434
rect 492918 136198 493154 136434
rect 492918 129198 493154 129434
rect 492918 122198 493154 122434
rect 492918 115198 493154 115434
rect 492918 108198 493154 108434
rect 492918 101198 493154 101434
rect 492918 94198 493154 94434
rect 492918 87198 493154 87434
rect 492918 80198 493154 80434
rect 492918 73198 493154 73434
rect 492918 66198 493154 66434
rect 492918 59198 493154 59434
rect 492918 52198 493154 52434
rect 492918 45198 493154 45434
rect 492918 38198 493154 38434
rect 492918 31198 493154 31434
rect 492918 24198 493154 24434
rect 492918 17198 493154 17434
rect 492918 10198 493154 10434
rect 492918 3198 493154 3434
rect 492918 -1942 493154 -1706
rect 492918 -2262 493154 -2026
rect 498186 705002 498422 705238
rect 498186 704682 498422 704918
rect 498186 695258 498422 695494
rect 498186 688258 498422 688494
rect 498186 681258 498422 681494
rect 498186 674258 498422 674494
rect 498186 667258 498422 667494
rect 498186 660258 498422 660494
rect 498186 653258 498422 653494
rect 498186 646258 498422 646494
rect 498186 639258 498422 639494
rect 498186 632258 498422 632494
rect 498186 625258 498422 625494
rect 498186 618258 498422 618494
rect 498186 611258 498422 611494
rect 498186 604258 498422 604494
rect 498186 597258 498422 597494
rect 498186 590258 498422 590494
rect 498186 583258 498422 583494
rect 498186 576258 498422 576494
rect 498186 569258 498422 569494
rect 498186 562258 498422 562494
rect 498186 555258 498422 555494
rect 498186 548258 498422 548494
rect 498186 541258 498422 541494
rect 498186 534258 498422 534494
rect 498186 527258 498422 527494
rect 498186 520258 498422 520494
rect 498186 513258 498422 513494
rect 498186 506258 498422 506494
rect 498186 499258 498422 499494
rect 498186 492258 498422 492494
rect 498186 485258 498422 485494
rect 498186 478258 498422 478494
rect 498186 471258 498422 471494
rect 498186 464258 498422 464494
rect 498186 457258 498422 457494
rect 498186 450258 498422 450494
rect 498186 443258 498422 443494
rect 498186 436258 498422 436494
rect 498186 429258 498422 429494
rect 498186 422258 498422 422494
rect 498186 415258 498422 415494
rect 498186 408258 498422 408494
rect 498186 401258 498422 401494
rect 498186 394258 498422 394494
rect 498186 387258 498422 387494
rect 498186 380258 498422 380494
rect 498186 373258 498422 373494
rect 498186 366258 498422 366494
rect 498186 359258 498422 359494
rect 498186 352258 498422 352494
rect 498186 345258 498422 345494
rect 498186 338258 498422 338494
rect 498186 331258 498422 331494
rect 498186 324258 498422 324494
rect 498186 317258 498422 317494
rect 498186 310258 498422 310494
rect 498186 303258 498422 303494
rect 498186 296258 498422 296494
rect 498186 289258 498422 289494
rect 498186 282258 498422 282494
rect 498186 275258 498422 275494
rect 498186 268258 498422 268494
rect 498186 261258 498422 261494
rect 498186 254258 498422 254494
rect 498186 247258 498422 247494
rect 498186 240258 498422 240494
rect 498186 233258 498422 233494
rect 498186 226258 498422 226494
rect 498186 219258 498422 219494
rect 498186 212258 498422 212494
rect 498186 205258 498422 205494
rect 498186 198258 498422 198494
rect 498186 191258 498422 191494
rect 498186 184258 498422 184494
rect 498186 177258 498422 177494
rect 498186 170258 498422 170494
rect 498186 163258 498422 163494
rect 498186 156258 498422 156494
rect 498186 149258 498422 149494
rect 498186 142258 498422 142494
rect 498186 135258 498422 135494
rect 498186 128258 498422 128494
rect 498186 121258 498422 121494
rect 498186 114258 498422 114494
rect 498186 107258 498422 107494
rect 498186 100258 498422 100494
rect 498186 93258 498422 93494
rect 498186 86258 498422 86494
rect 498186 79258 498422 79494
rect 498186 72258 498422 72494
rect 498186 65258 498422 65494
rect 498186 58258 498422 58494
rect 498186 51258 498422 51494
rect 498186 44258 498422 44494
rect 498186 37258 498422 37494
rect 498186 30258 498422 30494
rect 498186 23258 498422 23494
rect 498186 16258 498422 16494
rect 498186 9258 498422 9494
rect 498186 2258 498422 2494
rect 498186 -982 498422 -746
rect 498186 -1302 498422 -1066
rect 499918 705962 500154 706198
rect 499918 705642 500154 705878
rect 499918 696198 500154 696434
rect 499918 689198 500154 689434
rect 499918 682198 500154 682434
rect 499918 675198 500154 675434
rect 499918 668198 500154 668434
rect 499918 661198 500154 661434
rect 499918 654198 500154 654434
rect 499918 647198 500154 647434
rect 499918 640198 500154 640434
rect 499918 633198 500154 633434
rect 499918 626198 500154 626434
rect 499918 619198 500154 619434
rect 499918 612198 500154 612434
rect 499918 605198 500154 605434
rect 499918 598198 500154 598434
rect 499918 591198 500154 591434
rect 499918 584198 500154 584434
rect 499918 577198 500154 577434
rect 499918 570198 500154 570434
rect 499918 563198 500154 563434
rect 499918 556198 500154 556434
rect 499918 549198 500154 549434
rect 499918 542198 500154 542434
rect 499918 535198 500154 535434
rect 499918 528198 500154 528434
rect 499918 521198 500154 521434
rect 499918 514198 500154 514434
rect 499918 507198 500154 507434
rect 499918 500198 500154 500434
rect 499918 493198 500154 493434
rect 499918 486198 500154 486434
rect 499918 479198 500154 479434
rect 499918 472198 500154 472434
rect 499918 465198 500154 465434
rect 499918 458198 500154 458434
rect 499918 451198 500154 451434
rect 499918 444198 500154 444434
rect 499918 437198 500154 437434
rect 499918 430198 500154 430434
rect 499918 423198 500154 423434
rect 499918 416198 500154 416434
rect 499918 409198 500154 409434
rect 499918 402198 500154 402434
rect 499918 395198 500154 395434
rect 499918 388198 500154 388434
rect 499918 381198 500154 381434
rect 499918 374198 500154 374434
rect 499918 367198 500154 367434
rect 499918 360198 500154 360434
rect 499918 353198 500154 353434
rect 499918 346198 500154 346434
rect 499918 339198 500154 339434
rect 499918 332198 500154 332434
rect 499918 325198 500154 325434
rect 499918 318198 500154 318434
rect 499918 311198 500154 311434
rect 499918 304198 500154 304434
rect 499918 297198 500154 297434
rect 499918 290198 500154 290434
rect 499918 283198 500154 283434
rect 499918 276198 500154 276434
rect 499918 269198 500154 269434
rect 499918 262198 500154 262434
rect 499918 255198 500154 255434
rect 499918 248198 500154 248434
rect 499918 241198 500154 241434
rect 499918 234198 500154 234434
rect 499918 227198 500154 227434
rect 499918 220198 500154 220434
rect 499918 213198 500154 213434
rect 499918 206198 500154 206434
rect 499918 199198 500154 199434
rect 499918 192198 500154 192434
rect 499918 185198 500154 185434
rect 499918 178198 500154 178434
rect 499918 171198 500154 171434
rect 499918 164198 500154 164434
rect 499918 157198 500154 157434
rect 499918 150198 500154 150434
rect 499918 143198 500154 143434
rect 499918 136198 500154 136434
rect 499918 129198 500154 129434
rect 499918 122198 500154 122434
rect 499918 115198 500154 115434
rect 499918 108198 500154 108434
rect 499918 101198 500154 101434
rect 499918 94198 500154 94434
rect 499918 87198 500154 87434
rect 499918 80198 500154 80434
rect 499918 73198 500154 73434
rect 499918 66198 500154 66434
rect 499918 59198 500154 59434
rect 499918 52198 500154 52434
rect 499918 45198 500154 45434
rect 499918 38198 500154 38434
rect 499918 31198 500154 31434
rect 499918 24198 500154 24434
rect 499918 17198 500154 17434
rect 499918 10198 500154 10434
rect 499918 3198 500154 3434
rect 499918 -1942 500154 -1706
rect 499918 -2262 500154 -2026
rect 505186 705002 505422 705238
rect 505186 704682 505422 704918
rect 505186 695258 505422 695494
rect 505186 688258 505422 688494
rect 505186 681258 505422 681494
rect 505186 674258 505422 674494
rect 505186 667258 505422 667494
rect 505186 660258 505422 660494
rect 505186 653258 505422 653494
rect 505186 646258 505422 646494
rect 505186 639258 505422 639494
rect 505186 632258 505422 632494
rect 505186 625258 505422 625494
rect 505186 618258 505422 618494
rect 505186 611258 505422 611494
rect 505186 604258 505422 604494
rect 505186 597258 505422 597494
rect 505186 590258 505422 590494
rect 505186 583258 505422 583494
rect 505186 576258 505422 576494
rect 505186 569258 505422 569494
rect 505186 562258 505422 562494
rect 505186 555258 505422 555494
rect 505186 548258 505422 548494
rect 505186 541258 505422 541494
rect 505186 534258 505422 534494
rect 505186 527258 505422 527494
rect 505186 520258 505422 520494
rect 505186 513258 505422 513494
rect 505186 506258 505422 506494
rect 505186 499258 505422 499494
rect 505186 492258 505422 492494
rect 505186 485258 505422 485494
rect 505186 478258 505422 478494
rect 505186 471258 505422 471494
rect 505186 464258 505422 464494
rect 505186 457258 505422 457494
rect 505186 450258 505422 450494
rect 505186 443258 505422 443494
rect 505186 436258 505422 436494
rect 505186 429258 505422 429494
rect 505186 422258 505422 422494
rect 505186 415258 505422 415494
rect 505186 408258 505422 408494
rect 505186 401258 505422 401494
rect 505186 394258 505422 394494
rect 505186 387258 505422 387494
rect 505186 380258 505422 380494
rect 505186 373258 505422 373494
rect 505186 366258 505422 366494
rect 505186 359258 505422 359494
rect 505186 352258 505422 352494
rect 505186 345258 505422 345494
rect 505186 338258 505422 338494
rect 505186 331258 505422 331494
rect 505186 324258 505422 324494
rect 505186 317258 505422 317494
rect 505186 310258 505422 310494
rect 505186 303258 505422 303494
rect 505186 296258 505422 296494
rect 505186 289258 505422 289494
rect 505186 282258 505422 282494
rect 505186 275258 505422 275494
rect 505186 268258 505422 268494
rect 505186 261258 505422 261494
rect 505186 254258 505422 254494
rect 505186 247258 505422 247494
rect 505186 240258 505422 240494
rect 505186 233258 505422 233494
rect 505186 226258 505422 226494
rect 505186 219258 505422 219494
rect 505186 212258 505422 212494
rect 505186 205258 505422 205494
rect 505186 198258 505422 198494
rect 505186 191258 505422 191494
rect 505186 184258 505422 184494
rect 505186 177258 505422 177494
rect 505186 170258 505422 170494
rect 505186 163258 505422 163494
rect 505186 156258 505422 156494
rect 505186 149258 505422 149494
rect 505186 142258 505422 142494
rect 505186 135258 505422 135494
rect 505186 128258 505422 128494
rect 505186 121258 505422 121494
rect 505186 114258 505422 114494
rect 505186 107258 505422 107494
rect 505186 100258 505422 100494
rect 505186 93258 505422 93494
rect 505186 86258 505422 86494
rect 505186 79258 505422 79494
rect 505186 72258 505422 72494
rect 505186 65258 505422 65494
rect 505186 58258 505422 58494
rect 505186 51258 505422 51494
rect 505186 44258 505422 44494
rect 505186 37258 505422 37494
rect 505186 30258 505422 30494
rect 505186 23258 505422 23494
rect 505186 16258 505422 16494
rect 505186 9258 505422 9494
rect 505186 2258 505422 2494
rect 505186 -982 505422 -746
rect 505186 -1302 505422 -1066
rect 506918 705962 507154 706198
rect 506918 705642 507154 705878
rect 506918 696198 507154 696434
rect 506918 689198 507154 689434
rect 506918 682198 507154 682434
rect 506918 675198 507154 675434
rect 506918 668198 507154 668434
rect 506918 661198 507154 661434
rect 506918 654198 507154 654434
rect 506918 647198 507154 647434
rect 506918 640198 507154 640434
rect 506918 633198 507154 633434
rect 506918 626198 507154 626434
rect 506918 619198 507154 619434
rect 506918 612198 507154 612434
rect 506918 605198 507154 605434
rect 506918 598198 507154 598434
rect 506918 591198 507154 591434
rect 506918 584198 507154 584434
rect 506918 577198 507154 577434
rect 506918 570198 507154 570434
rect 506918 563198 507154 563434
rect 506918 556198 507154 556434
rect 506918 549198 507154 549434
rect 506918 542198 507154 542434
rect 506918 535198 507154 535434
rect 506918 528198 507154 528434
rect 506918 521198 507154 521434
rect 506918 514198 507154 514434
rect 506918 507198 507154 507434
rect 506918 500198 507154 500434
rect 506918 493198 507154 493434
rect 506918 486198 507154 486434
rect 506918 479198 507154 479434
rect 506918 472198 507154 472434
rect 506918 465198 507154 465434
rect 506918 458198 507154 458434
rect 506918 451198 507154 451434
rect 506918 444198 507154 444434
rect 506918 437198 507154 437434
rect 506918 430198 507154 430434
rect 506918 423198 507154 423434
rect 506918 416198 507154 416434
rect 506918 409198 507154 409434
rect 506918 402198 507154 402434
rect 506918 395198 507154 395434
rect 506918 388198 507154 388434
rect 506918 381198 507154 381434
rect 506918 374198 507154 374434
rect 506918 367198 507154 367434
rect 506918 360198 507154 360434
rect 506918 353198 507154 353434
rect 506918 346198 507154 346434
rect 506918 339198 507154 339434
rect 506918 332198 507154 332434
rect 506918 325198 507154 325434
rect 506918 318198 507154 318434
rect 506918 311198 507154 311434
rect 506918 304198 507154 304434
rect 506918 297198 507154 297434
rect 506918 290198 507154 290434
rect 506918 283198 507154 283434
rect 506918 276198 507154 276434
rect 506918 269198 507154 269434
rect 506918 262198 507154 262434
rect 506918 255198 507154 255434
rect 506918 248198 507154 248434
rect 506918 241198 507154 241434
rect 506918 234198 507154 234434
rect 506918 227198 507154 227434
rect 506918 220198 507154 220434
rect 506918 213198 507154 213434
rect 506918 206198 507154 206434
rect 506918 199198 507154 199434
rect 506918 192198 507154 192434
rect 506918 185198 507154 185434
rect 506918 178198 507154 178434
rect 506918 171198 507154 171434
rect 506918 164198 507154 164434
rect 506918 157198 507154 157434
rect 506918 150198 507154 150434
rect 506918 143198 507154 143434
rect 506918 136198 507154 136434
rect 506918 129198 507154 129434
rect 506918 122198 507154 122434
rect 506918 115198 507154 115434
rect 506918 108198 507154 108434
rect 506918 101198 507154 101434
rect 506918 94198 507154 94434
rect 506918 87198 507154 87434
rect 506918 80198 507154 80434
rect 506918 73198 507154 73434
rect 506918 66198 507154 66434
rect 506918 59198 507154 59434
rect 506918 52198 507154 52434
rect 506918 45198 507154 45434
rect 506918 38198 507154 38434
rect 506918 31198 507154 31434
rect 506918 24198 507154 24434
rect 506918 17198 507154 17434
rect 506918 10198 507154 10434
rect 506918 3198 507154 3434
rect 506918 -1942 507154 -1706
rect 506918 -2262 507154 -2026
rect 512186 705002 512422 705238
rect 512186 704682 512422 704918
rect 512186 695258 512422 695494
rect 512186 688258 512422 688494
rect 512186 681258 512422 681494
rect 512186 674258 512422 674494
rect 512186 667258 512422 667494
rect 512186 660258 512422 660494
rect 512186 653258 512422 653494
rect 512186 646258 512422 646494
rect 512186 639258 512422 639494
rect 512186 632258 512422 632494
rect 512186 625258 512422 625494
rect 512186 618258 512422 618494
rect 512186 611258 512422 611494
rect 512186 604258 512422 604494
rect 512186 597258 512422 597494
rect 512186 590258 512422 590494
rect 512186 583258 512422 583494
rect 512186 576258 512422 576494
rect 512186 569258 512422 569494
rect 512186 562258 512422 562494
rect 512186 555258 512422 555494
rect 512186 548258 512422 548494
rect 512186 541258 512422 541494
rect 512186 534258 512422 534494
rect 512186 527258 512422 527494
rect 512186 520258 512422 520494
rect 512186 513258 512422 513494
rect 512186 506258 512422 506494
rect 512186 499258 512422 499494
rect 512186 492258 512422 492494
rect 512186 485258 512422 485494
rect 512186 478258 512422 478494
rect 512186 471258 512422 471494
rect 512186 464258 512422 464494
rect 512186 457258 512422 457494
rect 512186 450258 512422 450494
rect 512186 443258 512422 443494
rect 512186 436258 512422 436494
rect 512186 429258 512422 429494
rect 512186 422258 512422 422494
rect 512186 415258 512422 415494
rect 512186 408258 512422 408494
rect 512186 401258 512422 401494
rect 512186 394258 512422 394494
rect 512186 387258 512422 387494
rect 512186 380258 512422 380494
rect 512186 373258 512422 373494
rect 512186 366258 512422 366494
rect 512186 359258 512422 359494
rect 512186 352258 512422 352494
rect 512186 345258 512422 345494
rect 512186 338258 512422 338494
rect 512186 331258 512422 331494
rect 512186 324258 512422 324494
rect 512186 317258 512422 317494
rect 512186 310258 512422 310494
rect 512186 303258 512422 303494
rect 512186 296258 512422 296494
rect 512186 289258 512422 289494
rect 512186 282258 512422 282494
rect 512186 275258 512422 275494
rect 512186 268258 512422 268494
rect 512186 261258 512422 261494
rect 512186 254258 512422 254494
rect 512186 247258 512422 247494
rect 512186 240258 512422 240494
rect 512186 233258 512422 233494
rect 512186 226258 512422 226494
rect 512186 219258 512422 219494
rect 512186 212258 512422 212494
rect 512186 205258 512422 205494
rect 512186 198258 512422 198494
rect 512186 191258 512422 191494
rect 512186 184258 512422 184494
rect 512186 177258 512422 177494
rect 512186 170258 512422 170494
rect 512186 163258 512422 163494
rect 512186 156258 512422 156494
rect 512186 149258 512422 149494
rect 512186 142258 512422 142494
rect 512186 135258 512422 135494
rect 512186 128258 512422 128494
rect 512186 121258 512422 121494
rect 512186 114258 512422 114494
rect 512186 107258 512422 107494
rect 512186 100258 512422 100494
rect 512186 93258 512422 93494
rect 512186 86258 512422 86494
rect 512186 79258 512422 79494
rect 512186 72258 512422 72494
rect 512186 65258 512422 65494
rect 512186 58258 512422 58494
rect 512186 51258 512422 51494
rect 512186 44258 512422 44494
rect 512186 37258 512422 37494
rect 512186 30258 512422 30494
rect 512186 23258 512422 23494
rect 512186 16258 512422 16494
rect 512186 9258 512422 9494
rect 512186 2258 512422 2494
rect 512186 -982 512422 -746
rect 512186 -1302 512422 -1066
rect 513918 705962 514154 706198
rect 513918 705642 514154 705878
rect 513918 696198 514154 696434
rect 513918 689198 514154 689434
rect 513918 682198 514154 682434
rect 513918 675198 514154 675434
rect 513918 668198 514154 668434
rect 513918 661198 514154 661434
rect 513918 654198 514154 654434
rect 513918 647198 514154 647434
rect 513918 640198 514154 640434
rect 513918 633198 514154 633434
rect 513918 626198 514154 626434
rect 513918 619198 514154 619434
rect 513918 612198 514154 612434
rect 513918 605198 514154 605434
rect 513918 598198 514154 598434
rect 513918 591198 514154 591434
rect 513918 584198 514154 584434
rect 513918 577198 514154 577434
rect 513918 570198 514154 570434
rect 513918 563198 514154 563434
rect 513918 556198 514154 556434
rect 513918 549198 514154 549434
rect 513918 542198 514154 542434
rect 513918 535198 514154 535434
rect 513918 528198 514154 528434
rect 513918 521198 514154 521434
rect 513918 514198 514154 514434
rect 513918 507198 514154 507434
rect 513918 500198 514154 500434
rect 513918 493198 514154 493434
rect 513918 486198 514154 486434
rect 513918 479198 514154 479434
rect 513918 472198 514154 472434
rect 513918 465198 514154 465434
rect 513918 458198 514154 458434
rect 513918 451198 514154 451434
rect 513918 444198 514154 444434
rect 513918 437198 514154 437434
rect 513918 430198 514154 430434
rect 513918 423198 514154 423434
rect 513918 416198 514154 416434
rect 513918 409198 514154 409434
rect 513918 402198 514154 402434
rect 513918 395198 514154 395434
rect 513918 388198 514154 388434
rect 513918 381198 514154 381434
rect 513918 374198 514154 374434
rect 513918 367198 514154 367434
rect 513918 360198 514154 360434
rect 513918 353198 514154 353434
rect 513918 346198 514154 346434
rect 513918 339198 514154 339434
rect 513918 332198 514154 332434
rect 513918 325198 514154 325434
rect 513918 318198 514154 318434
rect 513918 311198 514154 311434
rect 513918 304198 514154 304434
rect 513918 297198 514154 297434
rect 513918 290198 514154 290434
rect 513918 283198 514154 283434
rect 513918 276198 514154 276434
rect 513918 269198 514154 269434
rect 513918 262198 514154 262434
rect 513918 255198 514154 255434
rect 513918 248198 514154 248434
rect 513918 241198 514154 241434
rect 513918 234198 514154 234434
rect 513918 227198 514154 227434
rect 513918 220198 514154 220434
rect 513918 213198 514154 213434
rect 513918 206198 514154 206434
rect 513918 199198 514154 199434
rect 513918 192198 514154 192434
rect 513918 185198 514154 185434
rect 513918 178198 514154 178434
rect 513918 171198 514154 171434
rect 513918 164198 514154 164434
rect 513918 157198 514154 157434
rect 513918 150198 514154 150434
rect 513918 143198 514154 143434
rect 513918 136198 514154 136434
rect 513918 129198 514154 129434
rect 513918 122198 514154 122434
rect 513918 115198 514154 115434
rect 513918 108198 514154 108434
rect 513918 101198 514154 101434
rect 513918 94198 514154 94434
rect 513918 87198 514154 87434
rect 513918 80198 514154 80434
rect 513918 73198 514154 73434
rect 513918 66198 514154 66434
rect 513918 59198 514154 59434
rect 513918 52198 514154 52434
rect 513918 45198 514154 45434
rect 513918 38198 514154 38434
rect 513918 31198 514154 31434
rect 513918 24198 514154 24434
rect 513918 17198 514154 17434
rect 513918 10198 514154 10434
rect 513918 3198 514154 3434
rect 513918 -1942 514154 -1706
rect 513918 -2262 514154 -2026
rect 519186 705002 519422 705238
rect 519186 704682 519422 704918
rect 519186 695258 519422 695494
rect 519186 688258 519422 688494
rect 519186 681258 519422 681494
rect 519186 674258 519422 674494
rect 519186 667258 519422 667494
rect 519186 660258 519422 660494
rect 519186 653258 519422 653494
rect 519186 646258 519422 646494
rect 519186 639258 519422 639494
rect 519186 632258 519422 632494
rect 519186 625258 519422 625494
rect 519186 618258 519422 618494
rect 519186 611258 519422 611494
rect 519186 604258 519422 604494
rect 519186 597258 519422 597494
rect 519186 590258 519422 590494
rect 519186 583258 519422 583494
rect 519186 576258 519422 576494
rect 519186 569258 519422 569494
rect 519186 562258 519422 562494
rect 519186 555258 519422 555494
rect 519186 548258 519422 548494
rect 519186 541258 519422 541494
rect 519186 534258 519422 534494
rect 519186 527258 519422 527494
rect 519186 520258 519422 520494
rect 519186 513258 519422 513494
rect 519186 506258 519422 506494
rect 519186 499258 519422 499494
rect 519186 492258 519422 492494
rect 519186 485258 519422 485494
rect 519186 478258 519422 478494
rect 519186 471258 519422 471494
rect 519186 464258 519422 464494
rect 519186 457258 519422 457494
rect 519186 450258 519422 450494
rect 519186 443258 519422 443494
rect 519186 436258 519422 436494
rect 519186 429258 519422 429494
rect 519186 422258 519422 422494
rect 520918 705962 521154 706198
rect 520918 705642 521154 705878
rect 520918 696198 521154 696434
rect 520918 689198 521154 689434
rect 520918 682198 521154 682434
rect 520918 675198 521154 675434
rect 520918 668198 521154 668434
rect 520918 661198 521154 661434
rect 520918 654198 521154 654434
rect 520918 647198 521154 647434
rect 520918 640198 521154 640434
rect 520918 633198 521154 633434
rect 520918 626198 521154 626434
rect 520918 619198 521154 619434
rect 520918 612198 521154 612434
rect 520918 605198 521154 605434
rect 520918 598198 521154 598434
rect 520918 591198 521154 591434
rect 520918 584198 521154 584434
rect 520918 577198 521154 577434
rect 520918 570198 521154 570434
rect 520918 563198 521154 563434
rect 520918 556198 521154 556434
rect 520918 549198 521154 549434
rect 520918 542198 521154 542434
rect 520918 535198 521154 535434
rect 520918 528198 521154 528434
rect 520918 521198 521154 521434
rect 520918 514198 521154 514434
rect 520918 507198 521154 507434
rect 520918 500198 521154 500434
rect 520918 493198 521154 493434
rect 520918 486198 521154 486434
rect 520918 479198 521154 479434
rect 520918 472198 521154 472434
rect 520918 465198 521154 465434
rect 520918 458198 521154 458434
rect 520918 451198 521154 451434
rect 520918 444198 521154 444434
rect 520918 437198 521154 437434
rect 520918 430198 521154 430434
rect 520918 423198 521154 423434
rect 526186 705002 526422 705238
rect 526186 704682 526422 704918
rect 526186 695258 526422 695494
rect 526186 688258 526422 688494
rect 526186 681258 526422 681494
rect 526186 674258 526422 674494
rect 526186 667258 526422 667494
rect 526186 660258 526422 660494
rect 526186 653258 526422 653494
rect 526186 646258 526422 646494
rect 526186 639258 526422 639494
rect 526186 632258 526422 632494
rect 526186 625258 526422 625494
rect 526186 618258 526422 618494
rect 526186 611258 526422 611494
rect 526186 604258 526422 604494
rect 526186 597258 526422 597494
rect 526186 590258 526422 590494
rect 526186 583258 526422 583494
rect 526186 576258 526422 576494
rect 526186 569258 526422 569494
rect 526186 562258 526422 562494
rect 526186 555258 526422 555494
rect 526186 548258 526422 548494
rect 526186 541258 526422 541494
rect 526186 534258 526422 534494
rect 526186 527258 526422 527494
rect 526186 520258 526422 520494
rect 526186 513258 526422 513494
rect 526186 506258 526422 506494
rect 526186 499258 526422 499494
rect 526186 492258 526422 492494
rect 526186 485258 526422 485494
rect 526186 478258 526422 478494
rect 526186 471258 526422 471494
rect 526186 464258 526422 464494
rect 526186 457258 526422 457494
rect 526186 450258 526422 450494
rect 526186 443258 526422 443494
rect 526186 436258 526422 436494
rect 526186 429258 526422 429494
rect 526186 422258 526422 422494
rect 527918 705962 528154 706198
rect 527918 705642 528154 705878
rect 527918 696198 528154 696434
rect 527918 689198 528154 689434
rect 527918 682198 528154 682434
rect 527918 675198 528154 675434
rect 527918 668198 528154 668434
rect 527918 661198 528154 661434
rect 527918 654198 528154 654434
rect 527918 647198 528154 647434
rect 527918 640198 528154 640434
rect 527918 633198 528154 633434
rect 527918 626198 528154 626434
rect 527918 619198 528154 619434
rect 527918 612198 528154 612434
rect 527918 605198 528154 605434
rect 527918 598198 528154 598434
rect 527918 591198 528154 591434
rect 527918 584198 528154 584434
rect 527918 577198 528154 577434
rect 527918 570198 528154 570434
rect 527918 563198 528154 563434
rect 527918 556198 528154 556434
rect 527918 549198 528154 549434
rect 527918 542198 528154 542434
rect 527918 535198 528154 535434
rect 527918 528198 528154 528434
rect 527918 521198 528154 521434
rect 527918 514198 528154 514434
rect 527918 507198 528154 507434
rect 527918 500198 528154 500434
rect 527918 493198 528154 493434
rect 527918 486198 528154 486434
rect 527918 479198 528154 479434
rect 527918 472198 528154 472434
rect 527918 465198 528154 465434
rect 527918 458198 528154 458434
rect 527918 451198 528154 451434
rect 527918 444198 528154 444434
rect 527918 437198 528154 437434
rect 527918 430198 528154 430434
rect 527918 423198 528154 423434
rect 520918 416198 521154 416434
rect 522850 416198 523086 416434
rect 524782 416198 525018 416434
rect 526714 416198 526950 416434
rect 527918 416198 528154 416434
rect 519186 415258 519422 415494
rect 519952 415258 520188 415494
rect 521884 415258 522120 415494
rect 523816 415258 524052 415494
rect 525748 415258 525984 415494
rect 520918 409198 521154 409434
rect 522850 409198 523086 409434
rect 524782 409198 525018 409434
rect 526714 409198 526950 409434
rect 527918 409198 528154 409434
rect 519186 408258 519422 408494
rect 519952 408258 520188 408494
rect 521884 408258 522120 408494
rect 523816 408258 524052 408494
rect 525748 408258 525984 408494
rect 520918 402198 521154 402434
rect 522850 402198 523086 402434
rect 524782 402198 525018 402434
rect 526714 402198 526950 402434
rect 527918 402198 528154 402434
rect 519186 401258 519422 401494
rect 519186 394258 519422 394494
rect 519186 387258 519422 387494
rect 520918 395198 521154 395434
rect 520918 388198 521154 388434
rect 526186 394258 526422 394494
rect 526186 387258 526422 387494
rect 527918 395198 528154 395434
rect 527918 388198 528154 388434
rect 519186 380258 519422 380494
rect 527918 381198 528154 381434
rect 520918 374198 521154 374434
rect 522850 374198 523086 374434
rect 524782 374198 525018 374434
rect 526714 374198 526950 374434
rect 527918 374198 528154 374434
rect 519186 373258 519422 373494
rect 519952 373258 520188 373494
rect 521884 373258 522120 373494
rect 523816 373258 524052 373494
rect 525748 373258 525984 373494
rect 520918 367198 521154 367434
rect 522850 367198 523086 367434
rect 524782 367198 525018 367434
rect 526714 367198 526950 367434
rect 527918 367198 528154 367434
rect 519186 366258 519422 366494
rect 519952 366258 520188 366494
rect 521884 366258 522120 366494
rect 523816 366258 524052 366494
rect 525748 366258 525984 366494
rect 527918 360198 528154 360434
rect 519186 359258 519422 359494
rect 519186 352258 519422 352494
rect 519186 345258 519422 345494
rect 520918 353198 521154 353434
rect 520918 346198 521154 346434
rect 526186 359258 526422 359494
rect 526186 352258 526422 352494
rect 526186 345258 526422 345494
rect 527918 353198 528154 353434
rect 527918 346198 528154 346434
rect 520918 339198 521154 339434
rect 522850 339198 523086 339434
rect 524782 339198 525018 339434
rect 526714 339198 526950 339434
rect 527918 339198 528154 339434
rect 519186 338258 519422 338494
rect 519952 338258 520188 338494
rect 521884 338258 522120 338494
rect 523816 338258 524052 338494
rect 525748 338258 525984 338494
rect 520918 332198 521154 332434
rect 522850 332198 523086 332434
rect 524782 332198 525018 332434
rect 526714 332198 526950 332434
rect 527918 332198 528154 332434
rect 519186 331258 519422 331494
rect 519952 331258 520188 331494
rect 521884 331258 522120 331494
rect 523816 331258 524052 331494
rect 525748 331258 525984 331494
rect 520918 325198 521154 325434
rect 522850 325198 523086 325434
rect 524782 325198 525018 325434
rect 526714 325198 526950 325434
rect 527918 325198 528154 325434
rect 519186 324258 519422 324494
rect 519952 324258 520188 324494
rect 521884 324258 522120 324494
rect 523816 324258 524052 324494
rect 525748 324258 525984 324494
rect 519186 317258 519422 317494
rect 519186 310258 519422 310494
rect 519186 303258 519422 303494
rect 520918 318198 521154 318434
rect 520918 311198 521154 311434
rect 520918 304198 521154 304434
rect 526186 317258 526422 317494
rect 526186 310258 526422 310494
rect 526186 303258 526422 303494
rect 527918 318198 528154 318434
rect 527918 311198 528154 311434
rect 527918 304198 528154 304434
rect 520918 297198 521154 297434
rect 522850 297198 523086 297434
rect 524782 297198 525018 297434
rect 526714 297198 526950 297434
rect 527918 297198 528154 297434
rect 519186 296258 519422 296494
rect 519952 296258 520188 296494
rect 521884 296258 522120 296494
rect 523816 296258 524052 296494
rect 525748 296258 525984 296494
rect 520918 290198 521154 290434
rect 522850 290198 523086 290434
rect 524782 290198 525018 290434
rect 526714 290198 526950 290434
rect 527918 290198 528154 290434
rect 519186 289258 519422 289494
rect 519952 289258 520188 289494
rect 521884 289258 522120 289494
rect 523816 289258 524052 289494
rect 525748 289258 525984 289494
rect 520918 283198 521154 283434
rect 522850 283198 523086 283434
rect 524782 283198 525018 283434
rect 526714 283198 526950 283434
rect 527918 283198 528154 283434
rect 519186 282258 519422 282494
rect 519952 282258 520188 282494
rect 521884 282258 522120 282494
rect 523816 282258 524052 282494
rect 525748 282258 525984 282494
rect 519186 275258 519422 275494
rect 519186 268258 519422 268494
rect 520918 276198 521154 276434
rect 520918 269198 521154 269434
rect 520918 262198 521154 262434
rect 526186 275258 526422 275494
rect 526186 268258 526422 268494
rect 527918 276198 528154 276434
rect 527918 269198 528154 269434
rect 527918 262198 528154 262434
rect 519186 261258 519422 261494
rect 520918 255198 521154 255434
rect 522850 255198 523086 255434
rect 524782 255198 525018 255434
rect 526714 255198 526950 255434
rect 527918 255198 528154 255434
rect 519186 254258 519422 254494
rect 519952 254258 520188 254494
rect 521884 254258 522120 254494
rect 523816 254258 524052 254494
rect 525748 254258 525984 254494
rect 520918 248198 521154 248434
rect 522850 248198 523086 248434
rect 524782 248198 525018 248434
rect 526714 248198 526950 248434
rect 527918 248198 528154 248434
rect 519186 247258 519422 247494
rect 519952 247258 520188 247494
rect 521884 247258 522120 247494
rect 523816 247258 524052 247494
rect 525748 247258 525984 247494
rect 519186 240258 519422 240494
rect 527918 241198 528154 241434
rect 519186 233258 519422 233494
rect 519186 226258 519422 226494
rect 519186 219258 519422 219494
rect 519186 212258 519422 212494
rect 519186 205258 519422 205494
rect 519186 198258 519422 198494
rect 519186 191258 519422 191494
rect 519186 184258 519422 184494
rect 519186 177258 519422 177494
rect 519186 170258 519422 170494
rect 519186 163258 519422 163494
rect 519186 156258 519422 156494
rect 519186 149258 519422 149494
rect 519186 142258 519422 142494
rect 519186 135258 519422 135494
rect 519186 128258 519422 128494
rect 519186 121258 519422 121494
rect 519186 114258 519422 114494
rect 519186 107258 519422 107494
rect 519186 100258 519422 100494
rect 519186 93258 519422 93494
rect 519186 86258 519422 86494
rect 519186 79258 519422 79494
rect 519186 72258 519422 72494
rect 519186 65258 519422 65494
rect 519186 58258 519422 58494
rect 519186 51258 519422 51494
rect 519186 44258 519422 44494
rect 519186 37258 519422 37494
rect 519186 30258 519422 30494
rect 519186 23258 519422 23494
rect 519186 16258 519422 16494
rect 519186 9258 519422 9494
rect 519186 2258 519422 2494
rect 519186 -982 519422 -746
rect 519186 -1302 519422 -1066
rect 520918 234198 521154 234434
rect 520918 227198 521154 227434
rect 520918 220198 521154 220434
rect 520918 213198 521154 213434
rect 520918 206198 521154 206434
rect 520918 199198 521154 199434
rect 520918 192198 521154 192434
rect 520918 185198 521154 185434
rect 520918 178198 521154 178434
rect 520918 171198 521154 171434
rect 520918 164198 521154 164434
rect 520918 157198 521154 157434
rect 520918 150198 521154 150434
rect 520918 143198 521154 143434
rect 520918 136198 521154 136434
rect 520918 129198 521154 129434
rect 520918 122198 521154 122434
rect 520918 115198 521154 115434
rect 520918 108198 521154 108434
rect 520918 101198 521154 101434
rect 520918 94198 521154 94434
rect 520918 87198 521154 87434
rect 520918 80198 521154 80434
rect 520918 73198 521154 73434
rect 520918 66198 521154 66434
rect 520918 59198 521154 59434
rect 520918 52198 521154 52434
rect 520918 45198 521154 45434
rect 520918 38198 521154 38434
rect 520918 31198 521154 31434
rect 520918 24198 521154 24434
rect 520918 17198 521154 17434
rect 520918 10198 521154 10434
rect 520918 3198 521154 3434
rect 520918 -1942 521154 -1706
rect 520918 -2262 521154 -2026
rect 526186 233258 526422 233494
rect 526186 226258 526422 226494
rect 526186 219258 526422 219494
rect 526186 212258 526422 212494
rect 526186 205258 526422 205494
rect 526186 198258 526422 198494
rect 526186 191258 526422 191494
rect 526186 184258 526422 184494
rect 526186 177258 526422 177494
rect 526186 170258 526422 170494
rect 526186 163258 526422 163494
rect 526186 156258 526422 156494
rect 526186 149258 526422 149494
rect 526186 142258 526422 142494
rect 526186 135258 526422 135494
rect 526186 128258 526422 128494
rect 526186 121258 526422 121494
rect 526186 114258 526422 114494
rect 526186 107258 526422 107494
rect 526186 100258 526422 100494
rect 526186 93258 526422 93494
rect 526186 86258 526422 86494
rect 526186 79258 526422 79494
rect 526186 72258 526422 72494
rect 526186 65258 526422 65494
rect 526186 58258 526422 58494
rect 526186 51258 526422 51494
rect 526186 44258 526422 44494
rect 526186 37258 526422 37494
rect 526186 30258 526422 30494
rect 526186 23258 526422 23494
rect 526186 16258 526422 16494
rect 526186 9258 526422 9494
rect 526186 2258 526422 2494
rect 526186 -982 526422 -746
rect 526186 -1302 526422 -1066
rect 527918 234198 528154 234434
rect 527918 227198 528154 227434
rect 527918 220198 528154 220434
rect 527918 213198 528154 213434
rect 527918 206198 528154 206434
rect 527918 199198 528154 199434
rect 527918 192198 528154 192434
rect 527918 185198 528154 185434
rect 527918 178198 528154 178434
rect 527918 171198 528154 171434
rect 527918 164198 528154 164434
rect 527918 157198 528154 157434
rect 527918 150198 528154 150434
rect 527918 143198 528154 143434
rect 527918 136198 528154 136434
rect 527918 129198 528154 129434
rect 527918 122198 528154 122434
rect 527918 115198 528154 115434
rect 527918 108198 528154 108434
rect 527918 101198 528154 101434
rect 527918 94198 528154 94434
rect 527918 87198 528154 87434
rect 527918 80198 528154 80434
rect 527918 73198 528154 73434
rect 527918 66198 528154 66434
rect 527918 59198 528154 59434
rect 527918 52198 528154 52434
rect 527918 45198 528154 45434
rect 527918 38198 528154 38434
rect 527918 31198 528154 31434
rect 527918 24198 528154 24434
rect 527918 17198 528154 17434
rect 527918 10198 528154 10434
rect 527918 3198 528154 3434
rect 527918 -1942 528154 -1706
rect 527918 -2262 528154 -2026
rect 533186 705002 533422 705238
rect 533186 704682 533422 704918
rect 533186 695258 533422 695494
rect 533186 688258 533422 688494
rect 533186 681258 533422 681494
rect 533186 674258 533422 674494
rect 533186 667258 533422 667494
rect 533186 660258 533422 660494
rect 533186 653258 533422 653494
rect 533186 646258 533422 646494
rect 533186 639258 533422 639494
rect 533186 632258 533422 632494
rect 533186 625258 533422 625494
rect 533186 618258 533422 618494
rect 533186 611258 533422 611494
rect 533186 604258 533422 604494
rect 533186 597258 533422 597494
rect 533186 590258 533422 590494
rect 533186 583258 533422 583494
rect 533186 576258 533422 576494
rect 533186 569258 533422 569494
rect 533186 562258 533422 562494
rect 533186 555258 533422 555494
rect 533186 548258 533422 548494
rect 533186 541258 533422 541494
rect 533186 534258 533422 534494
rect 533186 527258 533422 527494
rect 533186 520258 533422 520494
rect 533186 513258 533422 513494
rect 533186 506258 533422 506494
rect 533186 499258 533422 499494
rect 533186 492258 533422 492494
rect 533186 485258 533422 485494
rect 533186 478258 533422 478494
rect 533186 471258 533422 471494
rect 533186 464258 533422 464494
rect 533186 457258 533422 457494
rect 533186 450258 533422 450494
rect 533186 443258 533422 443494
rect 533186 436258 533422 436494
rect 533186 429258 533422 429494
rect 533186 422258 533422 422494
rect 533186 415258 533422 415494
rect 533186 408258 533422 408494
rect 533186 401258 533422 401494
rect 533186 394258 533422 394494
rect 533186 387258 533422 387494
rect 533186 380258 533422 380494
rect 533186 373258 533422 373494
rect 533186 366258 533422 366494
rect 533186 359258 533422 359494
rect 533186 352258 533422 352494
rect 533186 345258 533422 345494
rect 533186 338258 533422 338494
rect 533186 331258 533422 331494
rect 533186 324258 533422 324494
rect 533186 317258 533422 317494
rect 533186 310258 533422 310494
rect 533186 303258 533422 303494
rect 533186 296258 533422 296494
rect 533186 289258 533422 289494
rect 533186 282258 533422 282494
rect 533186 275258 533422 275494
rect 533186 268258 533422 268494
rect 533186 261258 533422 261494
rect 533186 254258 533422 254494
rect 533186 247258 533422 247494
rect 533186 240258 533422 240494
rect 533186 233258 533422 233494
rect 533186 226258 533422 226494
rect 533186 219258 533422 219494
rect 533186 212258 533422 212494
rect 533186 205258 533422 205494
rect 533186 198258 533422 198494
rect 533186 191258 533422 191494
rect 533186 184258 533422 184494
rect 533186 177258 533422 177494
rect 533186 170258 533422 170494
rect 533186 163258 533422 163494
rect 533186 156258 533422 156494
rect 533186 149258 533422 149494
rect 533186 142258 533422 142494
rect 533186 135258 533422 135494
rect 533186 128258 533422 128494
rect 533186 121258 533422 121494
rect 533186 114258 533422 114494
rect 533186 107258 533422 107494
rect 533186 100258 533422 100494
rect 533186 93258 533422 93494
rect 533186 86258 533422 86494
rect 533186 79258 533422 79494
rect 533186 72258 533422 72494
rect 533186 65258 533422 65494
rect 533186 58258 533422 58494
rect 533186 51258 533422 51494
rect 533186 44258 533422 44494
rect 533186 37258 533422 37494
rect 533186 30258 533422 30494
rect 533186 23258 533422 23494
rect 533186 16258 533422 16494
rect 533186 9258 533422 9494
rect 533186 2258 533422 2494
rect 533186 -982 533422 -746
rect 533186 -1302 533422 -1066
rect 534918 705962 535154 706198
rect 534918 705642 535154 705878
rect 534918 696198 535154 696434
rect 534918 689198 535154 689434
rect 534918 682198 535154 682434
rect 534918 675198 535154 675434
rect 534918 668198 535154 668434
rect 534918 661198 535154 661434
rect 534918 654198 535154 654434
rect 534918 647198 535154 647434
rect 534918 640198 535154 640434
rect 534918 633198 535154 633434
rect 534918 626198 535154 626434
rect 534918 619198 535154 619434
rect 534918 612198 535154 612434
rect 534918 605198 535154 605434
rect 534918 598198 535154 598434
rect 534918 591198 535154 591434
rect 534918 584198 535154 584434
rect 534918 577198 535154 577434
rect 534918 570198 535154 570434
rect 534918 563198 535154 563434
rect 534918 556198 535154 556434
rect 534918 549198 535154 549434
rect 534918 542198 535154 542434
rect 534918 535198 535154 535434
rect 534918 528198 535154 528434
rect 534918 521198 535154 521434
rect 534918 514198 535154 514434
rect 534918 507198 535154 507434
rect 534918 500198 535154 500434
rect 534918 493198 535154 493434
rect 534918 486198 535154 486434
rect 534918 479198 535154 479434
rect 534918 472198 535154 472434
rect 534918 465198 535154 465434
rect 534918 458198 535154 458434
rect 534918 451198 535154 451434
rect 534918 444198 535154 444434
rect 534918 437198 535154 437434
rect 534918 430198 535154 430434
rect 534918 423198 535154 423434
rect 534918 416198 535154 416434
rect 534918 409198 535154 409434
rect 534918 402198 535154 402434
rect 534918 395198 535154 395434
rect 534918 388198 535154 388434
rect 534918 381198 535154 381434
rect 534918 374198 535154 374434
rect 534918 367198 535154 367434
rect 534918 360198 535154 360434
rect 534918 353198 535154 353434
rect 534918 346198 535154 346434
rect 534918 339198 535154 339434
rect 534918 332198 535154 332434
rect 534918 325198 535154 325434
rect 534918 318198 535154 318434
rect 534918 311198 535154 311434
rect 534918 304198 535154 304434
rect 534918 297198 535154 297434
rect 534918 290198 535154 290434
rect 534918 283198 535154 283434
rect 534918 276198 535154 276434
rect 534918 269198 535154 269434
rect 534918 262198 535154 262434
rect 534918 255198 535154 255434
rect 534918 248198 535154 248434
rect 534918 241198 535154 241434
rect 534918 234198 535154 234434
rect 534918 227198 535154 227434
rect 534918 220198 535154 220434
rect 534918 213198 535154 213434
rect 534918 206198 535154 206434
rect 534918 199198 535154 199434
rect 534918 192198 535154 192434
rect 534918 185198 535154 185434
rect 534918 178198 535154 178434
rect 534918 171198 535154 171434
rect 534918 164198 535154 164434
rect 534918 157198 535154 157434
rect 534918 150198 535154 150434
rect 534918 143198 535154 143434
rect 534918 136198 535154 136434
rect 534918 129198 535154 129434
rect 534918 122198 535154 122434
rect 534918 115198 535154 115434
rect 534918 108198 535154 108434
rect 534918 101198 535154 101434
rect 534918 94198 535154 94434
rect 534918 87198 535154 87434
rect 534918 80198 535154 80434
rect 534918 73198 535154 73434
rect 534918 66198 535154 66434
rect 534918 59198 535154 59434
rect 534918 52198 535154 52434
rect 534918 45198 535154 45434
rect 534918 38198 535154 38434
rect 534918 31198 535154 31434
rect 534918 24198 535154 24434
rect 534918 17198 535154 17434
rect 534918 10198 535154 10434
rect 534918 3198 535154 3434
rect 534918 -1942 535154 -1706
rect 534918 -2262 535154 -2026
rect 540186 705002 540422 705238
rect 540186 704682 540422 704918
rect 540186 695258 540422 695494
rect 540186 688258 540422 688494
rect 540186 681258 540422 681494
rect 540186 674258 540422 674494
rect 540186 667258 540422 667494
rect 540186 660258 540422 660494
rect 540186 653258 540422 653494
rect 540186 646258 540422 646494
rect 540186 639258 540422 639494
rect 540186 632258 540422 632494
rect 540186 625258 540422 625494
rect 540186 618258 540422 618494
rect 540186 611258 540422 611494
rect 540186 604258 540422 604494
rect 540186 597258 540422 597494
rect 540186 590258 540422 590494
rect 540186 583258 540422 583494
rect 540186 576258 540422 576494
rect 540186 569258 540422 569494
rect 540186 562258 540422 562494
rect 540186 555258 540422 555494
rect 540186 548258 540422 548494
rect 540186 541258 540422 541494
rect 540186 534258 540422 534494
rect 540186 527258 540422 527494
rect 540186 520258 540422 520494
rect 540186 513258 540422 513494
rect 540186 506258 540422 506494
rect 540186 499258 540422 499494
rect 540186 492258 540422 492494
rect 540186 485258 540422 485494
rect 540186 478258 540422 478494
rect 540186 471258 540422 471494
rect 540186 464258 540422 464494
rect 540186 457258 540422 457494
rect 540186 450258 540422 450494
rect 540186 443258 540422 443494
rect 540186 436258 540422 436494
rect 540186 429258 540422 429494
rect 540186 422258 540422 422494
rect 540186 415258 540422 415494
rect 540186 408258 540422 408494
rect 540186 401258 540422 401494
rect 540186 394258 540422 394494
rect 540186 387258 540422 387494
rect 540186 380258 540422 380494
rect 540186 373258 540422 373494
rect 540186 366258 540422 366494
rect 540186 359258 540422 359494
rect 540186 352258 540422 352494
rect 540186 345258 540422 345494
rect 540186 338258 540422 338494
rect 540186 331258 540422 331494
rect 540186 324258 540422 324494
rect 540186 317258 540422 317494
rect 540186 310258 540422 310494
rect 540186 303258 540422 303494
rect 540186 296258 540422 296494
rect 540186 289258 540422 289494
rect 540186 282258 540422 282494
rect 540186 275258 540422 275494
rect 540186 268258 540422 268494
rect 540186 261258 540422 261494
rect 540186 254258 540422 254494
rect 540186 247258 540422 247494
rect 540186 240258 540422 240494
rect 540186 233258 540422 233494
rect 540186 226258 540422 226494
rect 540186 219258 540422 219494
rect 540186 212258 540422 212494
rect 540186 205258 540422 205494
rect 540186 198258 540422 198494
rect 540186 191258 540422 191494
rect 540186 184258 540422 184494
rect 540186 177258 540422 177494
rect 540186 170258 540422 170494
rect 540186 163258 540422 163494
rect 540186 156258 540422 156494
rect 540186 149258 540422 149494
rect 540186 142258 540422 142494
rect 540186 135258 540422 135494
rect 540186 128258 540422 128494
rect 540186 121258 540422 121494
rect 540186 114258 540422 114494
rect 540186 107258 540422 107494
rect 540186 100258 540422 100494
rect 540186 93258 540422 93494
rect 540186 86258 540422 86494
rect 540186 79258 540422 79494
rect 540186 72258 540422 72494
rect 540186 65258 540422 65494
rect 540186 58258 540422 58494
rect 540186 51258 540422 51494
rect 540186 44258 540422 44494
rect 540186 37258 540422 37494
rect 540186 30258 540422 30494
rect 540186 23258 540422 23494
rect 540186 16258 540422 16494
rect 540186 9258 540422 9494
rect 540186 2258 540422 2494
rect 540186 -982 540422 -746
rect 540186 -1302 540422 -1066
rect 541918 705962 542154 706198
rect 541918 705642 542154 705878
rect 541918 696198 542154 696434
rect 541918 689198 542154 689434
rect 541918 682198 542154 682434
rect 541918 675198 542154 675434
rect 541918 668198 542154 668434
rect 541918 661198 542154 661434
rect 541918 654198 542154 654434
rect 541918 647198 542154 647434
rect 541918 640198 542154 640434
rect 541918 633198 542154 633434
rect 541918 626198 542154 626434
rect 541918 619198 542154 619434
rect 541918 612198 542154 612434
rect 541918 605198 542154 605434
rect 541918 598198 542154 598434
rect 541918 591198 542154 591434
rect 541918 584198 542154 584434
rect 541918 577198 542154 577434
rect 541918 570198 542154 570434
rect 541918 563198 542154 563434
rect 541918 556198 542154 556434
rect 541918 549198 542154 549434
rect 541918 542198 542154 542434
rect 541918 535198 542154 535434
rect 541918 528198 542154 528434
rect 541918 521198 542154 521434
rect 541918 514198 542154 514434
rect 541918 507198 542154 507434
rect 541918 500198 542154 500434
rect 541918 493198 542154 493434
rect 541918 486198 542154 486434
rect 541918 479198 542154 479434
rect 541918 472198 542154 472434
rect 541918 465198 542154 465434
rect 541918 458198 542154 458434
rect 541918 451198 542154 451434
rect 541918 444198 542154 444434
rect 541918 437198 542154 437434
rect 541918 430198 542154 430434
rect 541918 423198 542154 423434
rect 541918 416198 542154 416434
rect 541918 409198 542154 409434
rect 541918 402198 542154 402434
rect 541918 395198 542154 395434
rect 541918 388198 542154 388434
rect 541918 381198 542154 381434
rect 541918 374198 542154 374434
rect 541918 367198 542154 367434
rect 541918 360198 542154 360434
rect 541918 353198 542154 353434
rect 541918 346198 542154 346434
rect 541918 339198 542154 339434
rect 541918 332198 542154 332434
rect 541918 325198 542154 325434
rect 541918 318198 542154 318434
rect 541918 311198 542154 311434
rect 541918 304198 542154 304434
rect 541918 297198 542154 297434
rect 541918 290198 542154 290434
rect 541918 283198 542154 283434
rect 541918 276198 542154 276434
rect 541918 269198 542154 269434
rect 541918 262198 542154 262434
rect 541918 255198 542154 255434
rect 541918 248198 542154 248434
rect 541918 241198 542154 241434
rect 541918 234198 542154 234434
rect 541918 227198 542154 227434
rect 541918 220198 542154 220434
rect 541918 213198 542154 213434
rect 541918 206198 542154 206434
rect 541918 199198 542154 199434
rect 541918 192198 542154 192434
rect 541918 185198 542154 185434
rect 541918 178198 542154 178434
rect 541918 171198 542154 171434
rect 541918 164198 542154 164434
rect 541918 157198 542154 157434
rect 541918 150198 542154 150434
rect 541918 143198 542154 143434
rect 541918 136198 542154 136434
rect 541918 129198 542154 129434
rect 541918 122198 542154 122434
rect 541918 115198 542154 115434
rect 541918 108198 542154 108434
rect 541918 101198 542154 101434
rect 541918 94198 542154 94434
rect 541918 87198 542154 87434
rect 541918 80198 542154 80434
rect 541918 73198 542154 73434
rect 541918 66198 542154 66434
rect 541918 59198 542154 59434
rect 541918 52198 542154 52434
rect 541918 45198 542154 45434
rect 541918 38198 542154 38434
rect 541918 31198 542154 31434
rect 541918 24198 542154 24434
rect 541918 17198 542154 17434
rect 541918 10198 542154 10434
rect 541918 3198 542154 3434
rect 541918 -1942 542154 -1706
rect 541918 -2262 542154 -2026
rect 547186 705002 547422 705238
rect 547186 704682 547422 704918
rect 547186 695258 547422 695494
rect 547186 688258 547422 688494
rect 547186 681258 547422 681494
rect 547186 674258 547422 674494
rect 547186 667258 547422 667494
rect 547186 660258 547422 660494
rect 547186 653258 547422 653494
rect 547186 646258 547422 646494
rect 547186 639258 547422 639494
rect 547186 632258 547422 632494
rect 547186 625258 547422 625494
rect 547186 618258 547422 618494
rect 547186 611258 547422 611494
rect 547186 604258 547422 604494
rect 547186 597258 547422 597494
rect 547186 590258 547422 590494
rect 547186 583258 547422 583494
rect 547186 576258 547422 576494
rect 547186 569258 547422 569494
rect 547186 562258 547422 562494
rect 547186 555258 547422 555494
rect 547186 548258 547422 548494
rect 547186 541258 547422 541494
rect 547186 534258 547422 534494
rect 547186 527258 547422 527494
rect 547186 520258 547422 520494
rect 547186 513258 547422 513494
rect 547186 506258 547422 506494
rect 547186 499258 547422 499494
rect 547186 492258 547422 492494
rect 547186 485258 547422 485494
rect 547186 478258 547422 478494
rect 547186 471258 547422 471494
rect 547186 464258 547422 464494
rect 547186 457258 547422 457494
rect 547186 450258 547422 450494
rect 547186 443258 547422 443494
rect 547186 436258 547422 436494
rect 547186 429258 547422 429494
rect 547186 422258 547422 422494
rect 547186 415258 547422 415494
rect 547186 408258 547422 408494
rect 547186 401258 547422 401494
rect 547186 394258 547422 394494
rect 547186 387258 547422 387494
rect 547186 380258 547422 380494
rect 547186 373258 547422 373494
rect 547186 366258 547422 366494
rect 547186 359258 547422 359494
rect 547186 352258 547422 352494
rect 547186 345258 547422 345494
rect 547186 338258 547422 338494
rect 547186 331258 547422 331494
rect 547186 324258 547422 324494
rect 547186 317258 547422 317494
rect 547186 310258 547422 310494
rect 547186 303258 547422 303494
rect 547186 296258 547422 296494
rect 547186 289258 547422 289494
rect 547186 282258 547422 282494
rect 547186 275258 547422 275494
rect 547186 268258 547422 268494
rect 547186 261258 547422 261494
rect 547186 254258 547422 254494
rect 547186 247258 547422 247494
rect 547186 240258 547422 240494
rect 547186 233258 547422 233494
rect 547186 226258 547422 226494
rect 547186 219258 547422 219494
rect 547186 212258 547422 212494
rect 547186 205258 547422 205494
rect 547186 198258 547422 198494
rect 547186 191258 547422 191494
rect 547186 184258 547422 184494
rect 547186 177258 547422 177494
rect 547186 170258 547422 170494
rect 547186 163258 547422 163494
rect 547186 156258 547422 156494
rect 547186 149258 547422 149494
rect 547186 142258 547422 142494
rect 547186 135258 547422 135494
rect 547186 128258 547422 128494
rect 547186 121258 547422 121494
rect 547186 114258 547422 114494
rect 547186 107258 547422 107494
rect 547186 100258 547422 100494
rect 547186 93258 547422 93494
rect 547186 86258 547422 86494
rect 547186 79258 547422 79494
rect 547186 72258 547422 72494
rect 547186 65258 547422 65494
rect 547186 58258 547422 58494
rect 547186 51258 547422 51494
rect 547186 44258 547422 44494
rect 547186 37258 547422 37494
rect 547186 30258 547422 30494
rect 547186 23258 547422 23494
rect 547186 16258 547422 16494
rect 547186 9258 547422 9494
rect 547186 2258 547422 2494
rect 547186 -982 547422 -746
rect 547186 -1302 547422 -1066
rect 548918 705962 549154 706198
rect 548918 705642 549154 705878
rect 548918 696198 549154 696434
rect 548918 689198 549154 689434
rect 548918 682198 549154 682434
rect 548918 675198 549154 675434
rect 548918 668198 549154 668434
rect 548918 661198 549154 661434
rect 548918 654198 549154 654434
rect 548918 647198 549154 647434
rect 548918 640198 549154 640434
rect 548918 633198 549154 633434
rect 548918 626198 549154 626434
rect 548918 619198 549154 619434
rect 548918 612198 549154 612434
rect 548918 605198 549154 605434
rect 548918 598198 549154 598434
rect 548918 591198 549154 591434
rect 548918 584198 549154 584434
rect 548918 577198 549154 577434
rect 548918 570198 549154 570434
rect 548918 563198 549154 563434
rect 548918 556198 549154 556434
rect 548918 549198 549154 549434
rect 548918 542198 549154 542434
rect 548918 535198 549154 535434
rect 548918 528198 549154 528434
rect 548918 521198 549154 521434
rect 548918 514198 549154 514434
rect 548918 507198 549154 507434
rect 548918 500198 549154 500434
rect 548918 493198 549154 493434
rect 548918 486198 549154 486434
rect 548918 479198 549154 479434
rect 548918 472198 549154 472434
rect 548918 465198 549154 465434
rect 548918 458198 549154 458434
rect 548918 451198 549154 451434
rect 548918 444198 549154 444434
rect 548918 437198 549154 437434
rect 548918 430198 549154 430434
rect 548918 423198 549154 423434
rect 548918 416198 549154 416434
rect 548918 409198 549154 409434
rect 548918 402198 549154 402434
rect 548918 395198 549154 395434
rect 548918 388198 549154 388434
rect 548918 381198 549154 381434
rect 548918 374198 549154 374434
rect 548918 367198 549154 367434
rect 548918 360198 549154 360434
rect 548918 353198 549154 353434
rect 548918 346198 549154 346434
rect 548918 339198 549154 339434
rect 548918 332198 549154 332434
rect 548918 325198 549154 325434
rect 548918 318198 549154 318434
rect 548918 311198 549154 311434
rect 548918 304198 549154 304434
rect 548918 297198 549154 297434
rect 548918 290198 549154 290434
rect 548918 283198 549154 283434
rect 548918 276198 549154 276434
rect 548918 269198 549154 269434
rect 548918 262198 549154 262434
rect 548918 255198 549154 255434
rect 548918 248198 549154 248434
rect 548918 241198 549154 241434
rect 548918 234198 549154 234434
rect 548918 227198 549154 227434
rect 548918 220198 549154 220434
rect 548918 213198 549154 213434
rect 548918 206198 549154 206434
rect 548918 199198 549154 199434
rect 548918 192198 549154 192434
rect 548918 185198 549154 185434
rect 548918 178198 549154 178434
rect 548918 171198 549154 171434
rect 548918 164198 549154 164434
rect 548918 157198 549154 157434
rect 548918 150198 549154 150434
rect 548918 143198 549154 143434
rect 548918 136198 549154 136434
rect 548918 129198 549154 129434
rect 548918 122198 549154 122434
rect 548918 115198 549154 115434
rect 548918 108198 549154 108434
rect 548918 101198 549154 101434
rect 548918 94198 549154 94434
rect 548918 87198 549154 87434
rect 548918 80198 549154 80434
rect 548918 73198 549154 73434
rect 548918 66198 549154 66434
rect 548918 59198 549154 59434
rect 548918 52198 549154 52434
rect 548918 45198 549154 45434
rect 548918 38198 549154 38434
rect 548918 31198 549154 31434
rect 548918 24198 549154 24434
rect 548918 17198 549154 17434
rect 548918 10198 549154 10434
rect 548918 3198 549154 3434
rect 548918 -1942 549154 -1706
rect 548918 -2262 549154 -2026
rect 554186 705002 554422 705238
rect 554186 704682 554422 704918
rect 554186 695258 554422 695494
rect 554186 688258 554422 688494
rect 554186 681258 554422 681494
rect 554186 674258 554422 674494
rect 554186 667258 554422 667494
rect 554186 660258 554422 660494
rect 554186 653258 554422 653494
rect 554186 646258 554422 646494
rect 554186 639258 554422 639494
rect 554186 632258 554422 632494
rect 554186 625258 554422 625494
rect 554186 618258 554422 618494
rect 554186 611258 554422 611494
rect 554186 604258 554422 604494
rect 554186 597258 554422 597494
rect 554186 590258 554422 590494
rect 554186 583258 554422 583494
rect 554186 576258 554422 576494
rect 554186 569258 554422 569494
rect 554186 562258 554422 562494
rect 554186 555258 554422 555494
rect 554186 548258 554422 548494
rect 554186 541258 554422 541494
rect 554186 534258 554422 534494
rect 554186 527258 554422 527494
rect 554186 520258 554422 520494
rect 554186 513258 554422 513494
rect 554186 506258 554422 506494
rect 554186 499258 554422 499494
rect 554186 492258 554422 492494
rect 554186 485258 554422 485494
rect 554186 478258 554422 478494
rect 554186 471258 554422 471494
rect 554186 464258 554422 464494
rect 554186 457258 554422 457494
rect 554186 450258 554422 450494
rect 554186 443258 554422 443494
rect 554186 436258 554422 436494
rect 554186 429258 554422 429494
rect 554186 422258 554422 422494
rect 554186 415258 554422 415494
rect 554186 408258 554422 408494
rect 554186 401258 554422 401494
rect 554186 394258 554422 394494
rect 554186 387258 554422 387494
rect 554186 380258 554422 380494
rect 554186 373258 554422 373494
rect 554186 366258 554422 366494
rect 554186 359258 554422 359494
rect 554186 352258 554422 352494
rect 554186 345258 554422 345494
rect 554186 338258 554422 338494
rect 554186 331258 554422 331494
rect 554186 324258 554422 324494
rect 554186 317258 554422 317494
rect 554186 310258 554422 310494
rect 554186 303258 554422 303494
rect 554186 296258 554422 296494
rect 554186 289258 554422 289494
rect 554186 282258 554422 282494
rect 554186 275258 554422 275494
rect 554186 268258 554422 268494
rect 554186 261258 554422 261494
rect 554186 254258 554422 254494
rect 554186 247258 554422 247494
rect 554186 240258 554422 240494
rect 554186 233258 554422 233494
rect 554186 226258 554422 226494
rect 554186 219258 554422 219494
rect 554186 212258 554422 212494
rect 554186 205258 554422 205494
rect 554186 198258 554422 198494
rect 554186 191258 554422 191494
rect 554186 184258 554422 184494
rect 554186 177258 554422 177494
rect 554186 170258 554422 170494
rect 554186 163258 554422 163494
rect 554186 156258 554422 156494
rect 554186 149258 554422 149494
rect 554186 142258 554422 142494
rect 554186 135258 554422 135494
rect 554186 128258 554422 128494
rect 554186 121258 554422 121494
rect 554186 114258 554422 114494
rect 554186 107258 554422 107494
rect 554186 100258 554422 100494
rect 554186 93258 554422 93494
rect 554186 86258 554422 86494
rect 554186 79258 554422 79494
rect 554186 72258 554422 72494
rect 554186 65258 554422 65494
rect 554186 58258 554422 58494
rect 554186 51258 554422 51494
rect 554186 44258 554422 44494
rect 554186 37258 554422 37494
rect 554186 30258 554422 30494
rect 554186 23258 554422 23494
rect 554186 16258 554422 16494
rect 554186 9258 554422 9494
rect 554186 2258 554422 2494
rect 554186 -982 554422 -746
rect 554186 -1302 554422 -1066
rect 555918 705962 556154 706198
rect 555918 705642 556154 705878
rect 555918 696198 556154 696434
rect 555918 689198 556154 689434
rect 555918 682198 556154 682434
rect 555918 675198 556154 675434
rect 555918 668198 556154 668434
rect 555918 661198 556154 661434
rect 555918 654198 556154 654434
rect 555918 647198 556154 647434
rect 555918 640198 556154 640434
rect 555918 633198 556154 633434
rect 555918 626198 556154 626434
rect 555918 619198 556154 619434
rect 555918 612198 556154 612434
rect 555918 605198 556154 605434
rect 555918 598198 556154 598434
rect 555918 591198 556154 591434
rect 555918 584198 556154 584434
rect 555918 577198 556154 577434
rect 555918 570198 556154 570434
rect 555918 563198 556154 563434
rect 555918 556198 556154 556434
rect 555918 549198 556154 549434
rect 555918 542198 556154 542434
rect 555918 535198 556154 535434
rect 555918 528198 556154 528434
rect 555918 521198 556154 521434
rect 555918 514198 556154 514434
rect 555918 507198 556154 507434
rect 555918 500198 556154 500434
rect 555918 493198 556154 493434
rect 555918 486198 556154 486434
rect 555918 479198 556154 479434
rect 555918 472198 556154 472434
rect 555918 465198 556154 465434
rect 555918 458198 556154 458434
rect 555918 451198 556154 451434
rect 555918 444198 556154 444434
rect 555918 437198 556154 437434
rect 555918 430198 556154 430434
rect 555918 423198 556154 423434
rect 555918 416198 556154 416434
rect 555918 409198 556154 409434
rect 555918 402198 556154 402434
rect 555918 395198 556154 395434
rect 555918 388198 556154 388434
rect 555918 381198 556154 381434
rect 555918 374198 556154 374434
rect 555918 367198 556154 367434
rect 555918 360198 556154 360434
rect 555918 353198 556154 353434
rect 555918 346198 556154 346434
rect 555918 339198 556154 339434
rect 555918 332198 556154 332434
rect 555918 325198 556154 325434
rect 555918 318198 556154 318434
rect 555918 311198 556154 311434
rect 555918 304198 556154 304434
rect 555918 297198 556154 297434
rect 555918 290198 556154 290434
rect 555918 283198 556154 283434
rect 555918 276198 556154 276434
rect 555918 269198 556154 269434
rect 555918 262198 556154 262434
rect 555918 255198 556154 255434
rect 555918 248198 556154 248434
rect 555918 241198 556154 241434
rect 555918 234198 556154 234434
rect 555918 227198 556154 227434
rect 555918 220198 556154 220434
rect 555918 213198 556154 213434
rect 555918 206198 556154 206434
rect 555918 199198 556154 199434
rect 555918 192198 556154 192434
rect 555918 185198 556154 185434
rect 555918 178198 556154 178434
rect 555918 171198 556154 171434
rect 555918 164198 556154 164434
rect 555918 157198 556154 157434
rect 555918 150198 556154 150434
rect 555918 143198 556154 143434
rect 555918 136198 556154 136434
rect 555918 129198 556154 129434
rect 555918 122198 556154 122434
rect 555918 115198 556154 115434
rect 555918 108198 556154 108434
rect 555918 101198 556154 101434
rect 555918 94198 556154 94434
rect 555918 87198 556154 87434
rect 555918 80198 556154 80434
rect 555918 73198 556154 73434
rect 555918 66198 556154 66434
rect 555918 59198 556154 59434
rect 555918 52198 556154 52434
rect 555918 45198 556154 45434
rect 555918 38198 556154 38434
rect 555918 31198 556154 31434
rect 555918 24198 556154 24434
rect 555918 17198 556154 17434
rect 555918 10198 556154 10434
rect 555918 3198 556154 3434
rect 555918 -1942 556154 -1706
rect 555918 -2262 556154 -2026
rect 561186 705002 561422 705238
rect 561186 704682 561422 704918
rect 561186 695258 561422 695494
rect 561186 688258 561422 688494
rect 561186 681258 561422 681494
rect 561186 674258 561422 674494
rect 561186 667258 561422 667494
rect 561186 660258 561422 660494
rect 561186 653258 561422 653494
rect 561186 646258 561422 646494
rect 561186 639258 561422 639494
rect 561186 632258 561422 632494
rect 561186 625258 561422 625494
rect 561186 618258 561422 618494
rect 561186 611258 561422 611494
rect 561186 604258 561422 604494
rect 561186 597258 561422 597494
rect 561186 590258 561422 590494
rect 561186 583258 561422 583494
rect 561186 576258 561422 576494
rect 561186 569258 561422 569494
rect 561186 562258 561422 562494
rect 561186 555258 561422 555494
rect 561186 548258 561422 548494
rect 561186 541258 561422 541494
rect 561186 534258 561422 534494
rect 561186 527258 561422 527494
rect 561186 520258 561422 520494
rect 561186 513258 561422 513494
rect 561186 506258 561422 506494
rect 561186 499258 561422 499494
rect 561186 492258 561422 492494
rect 561186 485258 561422 485494
rect 561186 478258 561422 478494
rect 561186 471258 561422 471494
rect 561186 464258 561422 464494
rect 561186 457258 561422 457494
rect 561186 450258 561422 450494
rect 561186 443258 561422 443494
rect 561186 436258 561422 436494
rect 561186 429258 561422 429494
rect 561186 422258 561422 422494
rect 561186 415258 561422 415494
rect 561186 408258 561422 408494
rect 561186 401258 561422 401494
rect 561186 394258 561422 394494
rect 561186 387258 561422 387494
rect 561186 380258 561422 380494
rect 561186 373258 561422 373494
rect 561186 366258 561422 366494
rect 561186 359258 561422 359494
rect 561186 352258 561422 352494
rect 561186 345258 561422 345494
rect 561186 338258 561422 338494
rect 561186 331258 561422 331494
rect 561186 324258 561422 324494
rect 561186 317258 561422 317494
rect 561186 310258 561422 310494
rect 561186 303258 561422 303494
rect 561186 296258 561422 296494
rect 561186 289258 561422 289494
rect 561186 282258 561422 282494
rect 561186 275258 561422 275494
rect 561186 268258 561422 268494
rect 561186 261258 561422 261494
rect 561186 254258 561422 254494
rect 561186 247258 561422 247494
rect 561186 240258 561422 240494
rect 561186 233258 561422 233494
rect 561186 226258 561422 226494
rect 561186 219258 561422 219494
rect 561186 212258 561422 212494
rect 561186 205258 561422 205494
rect 561186 198258 561422 198494
rect 561186 191258 561422 191494
rect 561186 184258 561422 184494
rect 561186 177258 561422 177494
rect 561186 170258 561422 170494
rect 561186 163258 561422 163494
rect 561186 156258 561422 156494
rect 561186 149258 561422 149494
rect 561186 142258 561422 142494
rect 561186 135258 561422 135494
rect 561186 128258 561422 128494
rect 561186 121258 561422 121494
rect 561186 114258 561422 114494
rect 561186 107258 561422 107494
rect 561186 100258 561422 100494
rect 561186 93258 561422 93494
rect 561186 86258 561422 86494
rect 561186 79258 561422 79494
rect 561186 72258 561422 72494
rect 561186 65258 561422 65494
rect 561186 58258 561422 58494
rect 561186 51258 561422 51494
rect 561186 44258 561422 44494
rect 561186 37258 561422 37494
rect 561186 30258 561422 30494
rect 561186 23258 561422 23494
rect 561186 16258 561422 16494
rect 561186 9258 561422 9494
rect 561186 2258 561422 2494
rect 561186 -982 561422 -746
rect 561186 -1302 561422 -1066
rect 562918 705962 563154 706198
rect 562918 705642 563154 705878
rect 562918 696198 563154 696434
rect 562918 689198 563154 689434
rect 562918 682198 563154 682434
rect 562918 675198 563154 675434
rect 562918 668198 563154 668434
rect 562918 661198 563154 661434
rect 562918 654198 563154 654434
rect 562918 647198 563154 647434
rect 562918 640198 563154 640434
rect 562918 633198 563154 633434
rect 562918 626198 563154 626434
rect 562918 619198 563154 619434
rect 562918 612198 563154 612434
rect 562918 605198 563154 605434
rect 562918 598198 563154 598434
rect 562918 591198 563154 591434
rect 562918 584198 563154 584434
rect 562918 577198 563154 577434
rect 562918 570198 563154 570434
rect 562918 563198 563154 563434
rect 562918 556198 563154 556434
rect 562918 549198 563154 549434
rect 562918 542198 563154 542434
rect 562918 535198 563154 535434
rect 562918 528198 563154 528434
rect 562918 521198 563154 521434
rect 562918 514198 563154 514434
rect 562918 507198 563154 507434
rect 562918 500198 563154 500434
rect 562918 493198 563154 493434
rect 562918 486198 563154 486434
rect 562918 479198 563154 479434
rect 562918 472198 563154 472434
rect 562918 465198 563154 465434
rect 562918 458198 563154 458434
rect 562918 451198 563154 451434
rect 562918 444198 563154 444434
rect 562918 437198 563154 437434
rect 562918 430198 563154 430434
rect 562918 423198 563154 423434
rect 562918 416198 563154 416434
rect 562918 409198 563154 409434
rect 562918 402198 563154 402434
rect 562918 395198 563154 395434
rect 562918 388198 563154 388434
rect 562918 381198 563154 381434
rect 562918 374198 563154 374434
rect 562918 367198 563154 367434
rect 562918 360198 563154 360434
rect 562918 353198 563154 353434
rect 562918 346198 563154 346434
rect 562918 339198 563154 339434
rect 562918 332198 563154 332434
rect 562918 325198 563154 325434
rect 562918 318198 563154 318434
rect 562918 311198 563154 311434
rect 562918 304198 563154 304434
rect 562918 297198 563154 297434
rect 562918 290198 563154 290434
rect 562918 283198 563154 283434
rect 562918 276198 563154 276434
rect 562918 269198 563154 269434
rect 562918 262198 563154 262434
rect 562918 255198 563154 255434
rect 562918 248198 563154 248434
rect 562918 241198 563154 241434
rect 562918 234198 563154 234434
rect 562918 227198 563154 227434
rect 562918 220198 563154 220434
rect 562918 213198 563154 213434
rect 562918 206198 563154 206434
rect 562918 199198 563154 199434
rect 562918 192198 563154 192434
rect 562918 185198 563154 185434
rect 562918 178198 563154 178434
rect 562918 171198 563154 171434
rect 562918 164198 563154 164434
rect 562918 157198 563154 157434
rect 562918 150198 563154 150434
rect 562918 143198 563154 143434
rect 562918 136198 563154 136434
rect 562918 129198 563154 129434
rect 562918 122198 563154 122434
rect 562918 115198 563154 115434
rect 562918 108198 563154 108434
rect 562918 101198 563154 101434
rect 562918 94198 563154 94434
rect 562918 87198 563154 87434
rect 562918 80198 563154 80434
rect 562918 73198 563154 73434
rect 562918 66198 563154 66434
rect 562918 59198 563154 59434
rect 562918 52198 563154 52434
rect 562918 45198 563154 45434
rect 562918 38198 563154 38434
rect 562918 31198 563154 31434
rect 562918 24198 563154 24434
rect 562918 17198 563154 17434
rect 562918 10198 563154 10434
rect 562918 3198 563154 3434
rect 562918 -1942 563154 -1706
rect 562918 -2262 563154 -2026
rect 568186 705002 568422 705238
rect 568186 704682 568422 704918
rect 568186 695258 568422 695494
rect 568186 688258 568422 688494
rect 568186 681258 568422 681494
rect 568186 674258 568422 674494
rect 568186 667258 568422 667494
rect 568186 660258 568422 660494
rect 568186 653258 568422 653494
rect 568186 646258 568422 646494
rect 568186 639258 568422 639494
rect 568186 632258 568422 632494
rect 568186 625258 568422 625494
rect 568186 618258 568422 618494
rect 568186 611258 568422 611494
rect 568186 604258 568422 604494
rect 568186 597258 568422 597494
rect 568186 590258 568422 590494
rect 568186 583258 568422 583494
rect 568186 576258 568422 576494
rect 568186 569258 568422 569494
rect 568186 562258 568422 562494
rect 568186 555258 568422 555494
rect 568186 548258 568422 548494
rect 568186 541258 568422 541494
rect 568186 534258 568422 534494
rect 568186 527258 568422 527494
rect 568186 520258 568422 520494
rect 568186 513258 568422 513494
rect 568186 506258 568422 506494
rect 568186 499258 568422 499494
rect 568186 492258 568422 492494
rect 568186 485258 568422 485494
rect 568186 478258 568422 478494
rect 568186 471258 568422 471494
rect 568186 464258 568422 464494
rect 568186 457258 568422 457494
rect 568186 450258 568422 450494
rect 568186 443258 568422 443494
rect 568186 436258 568422 436494
rect 568186 429258 568422 429494
rect 568186 422258 568422 422494
rect 568186 415258 568422 415494
rect 568186 408258 568422 408494
rect 568186 401258 568422 401494
rect 568186 394258 568422 394494
rect 568186 387258 568422 387494
rect 568186 380258 568422 380494
rect 568186 373258 568422 373494
rect 568186 366258 568422 366494
rect 568186 359258 568422 359494
rect 568186 352258 568422 352494
rect 568186 345258 568422 345494
rect 568186 338258 568422 338494
rect 568186 331258 568422 331494
rect 568186 324258 568422 324494
rect 568186 317258 568422 317494
rect 568186 310258 568422 310494
rect 568186 303258 568422 303494
rect 568186 296258 568422 296494
rect 568186 289258 568422 289494
rect 568186 282258 568422 282494
rect 568186 275258 568422 275494
rect 568186 268258 568422 268494
rect 568186 261258 568422 261494
rect 568186 254258 568422 254494
rect 568186 247258 568422 247494
rect 568186 240258 568422 240494
rect 568186 233258 568422 233494
rect 568186 226258 568422 226494
rect 568186 219258 568422 219494
rect 568186 212258 568422 212494
rect 568186 205258 568422 205494
rect 568186 198258 568422 198494
rect 568186 191258 568422 191494
rect 568186 184258 568422 184494
rect 568186 177258 568422 177494
rect 568186 170258 568422 170494
rect 568186 163258 568422 163494
rect 568186 156258 568422 156494
rect 568186 149258 568422 149494
rect 568186 142258 568422 142494
rect 568186 135258 568422 135494
rect 568186 128258 568422 128494
rect 568186 121258 568422 121494
rect 568186 114258 568422 114494
rect 568186 107258 568422 107494
rect 568186 100258 568422 100494
rect 568186 93258 568422 93494
rect 568186 86258 568422 86494
rect 568186 79258 568422 79494
rect 568186 72258 568422 72494
rect 568186 65258 568422 65494
rect 568186 58258 568422 58494
rect 568186 51258 568422 51494
rect 568186 44258 568422 44494
rect 568186 37258 568422 37494
rect 568186 30258 568422 30494
rect 568186 23258 568422 23494
rect 568186 16258 568422 16494
rect 568186 9258 568422 9494
rect 568186 2258 568422 2494
rect 568186 -982 568422 -746
rect 568186 -1302 568422 -1066
rect 569918 705962 570154 706198
rect 569918 705642 570154 705878
rect 569918 696198 570154 696434
rect 569918 689198 570154 689434
rect 569918 682198 570154 682434
rect 569918 675198 570154 675434
rect 569918 668198 570154 668434
rect 569918 661198 570154 661434
rect 569918 654198 570154 654434
rect 569918 647198 570154 647434
rect 569918 640198 570154 640434
rect 569918 633198 570154 633434
rect 569918 626198 570154 626434
rect 569918 619198 570154 619434
rect 569918 612198 570154 612434
rect 569918 605198 570154 605434
rect 569918 598198 570154 598434
rect 569918 591198 570154 591434
rect 569918 584198 570154 584434
rect 569918 577198 570154 577434
rect 569918 570198 570154 570434
rect 569918 563198 570154 563434
rect 569918 556198 570154 556434
rect 569918 549198 570154 549434
rect 569918 542198 570154 542434
rect 569918 535198 570154 535434
rect 569918 528198 570154 528434
rect 569918 521198 570154 521434
rect 569918 514198 570154 514434
rect 569918 507198 570154 507434
rect 569918 500198 570154 500434
rect 569918 493198 570154 493434
rect 569918 486198 570154 486434
rect 569918 479198 570154 479434
rect 569918 472198 570154 472434
rect 569918 465198 570154 465434
rect 569918 458198 570154 458434
rect 569918 451198 570154 451434
rect 569918 444198 570154 444434
rect 569918 437198 570154 437434
rect 569918 430198 570154 430434
rect 569918 423198 570154 423434
rect 569918 416198 570154 416434
rect 569918 409198 570154 409434
rect 569918 402198 570154 402434
rect 569918 395198 570154 395434
rect 569918 388198 570154 388434
rect 569918 381198 570154 381434
rect 569918 374198 570154 374434
rect 569918 367198 570154 367434
rect 569918 360198 570154 360434
rect 569918 353198 570154 353434
rect 569918 346198 570154 346434
rect 569918 339198 570154 339434
rect 569918 332198 570154 332434
rect 569918 325198 570154 325434
rect 569918 318198 570154 318434
rect 569918 311198 570154 311434
rect 569918 304198 570154 304434
rect 569918 297198 570154 297434
rect 569918 290198 570154 290434
rect 569918 283198 570154 283434
rect 569918 276198 570154 276434
rect 569918 269198 570154 269434
rect 569918 262198 570154 262434
rect 569918 255198 570154 255434
rect 569918 248198 570154 248434
rect 569918 241198 570154 241434
rect 569918 234198 570154 234434
rect 569918 227198 570154 227434
rect 569918 220198 570154 220434
rect 569918 213198 570154 213434
rect 569918 206198 570154 206434
rect 569918 199198 570154 199434
rect 569918 192198 570154 192434
rect 569918 185198 570154 185434
rect 569918 178198 570154 178434
rect 569918 171198 570154 171434
rect 569918 164198 570154 164434
rect 569918 157198 570154 157434
rect 569918 150198 570154 150434
rect 569918 143198 570154 143434
rect 569918 136198 570154 136434
rect 569918 129198 570154 129434
rect 569918 122198 570154 122434
rect 569918 115198 570154 115434
rect 569918 108198 570154 108434
rect 569918 101198 570154 101434
rect 569918 94198 570154 94434
rect 569918 87198 570154 87434
rect 569918 80198 570154 80434
rect 569918 73198 570154 73434
rect 569918 66198 570154 66434
rect 569918 59198 570154 59434
rect 569918 52198 570154 52434
rect 569918 45198 570154 45434
rect 569918 38198 570154 38434
rect 569918 31198 570154 31434
rect 569918 24198 570154 24434
rect 569918 17198 570154 17434
rect 569918 10198 570154 10434
rect 569918 3198 570154 3434
rect 569918 -1942 570154 -1706
rect 569918 -2262 570154 -2026
rect 575186 705002 575422 705238
rect 575186 704682 575422 704918
rect 575186 695258 575422 695494
rect 575186 688258 575422 688494
rect 575186 681258 575422 681494
rect 575186 674258 575422 674494
rect 575186 667258 575422 667494
rect 575186 660258 575422 660494
rect 575186 653258 575422 653494
rect 575186 646258 575422 646494
rect 575186 639258 575422 639494
rect 575186 632258 575422 632494
rect 575186 625258 575422 625494
rect 575186 618258 575422 618494
rect 575186 611258 575422 611494
rect 575186 604258 575422 604494
rect 575186 597258 575422 597494
rect 575186 590258 575422 590494
rect 575186 583258 575422 583494
rect 575186 576258 575422 576494
rect 575186 569258 575422 569494
rect 575186 562258 575422 562494
rect 575186 555258 575422 555494
rect 575186 548258 575422 548494
rect 575186 541258 575422 541494
rect 575186 534258 575422 534494
rect 575186 527258 575422 527494
rect 575186 520258 575422 520494
rect 575186 513258 575422 513494
rect 575186 506258 575422 506494
rect 575186 499258 575422 499494
rect 575186 492258 575422 492494
rect 575186 485258 575422 485494
rect 575186 478258 575422 478494
rect 575186 471258 575422 471494
rect 575186 464258 575422 464494
rect 575186 457258 575422 457494
rect 575186 450258 575422 450494
rect 575186 443258 575422 443494
rect 575186 436258 575422 436494
rect 575186 429258 575422 429494
rect 575186 422258 575422 422494
rect 575186 415258 575422 415494
rect 575186 408258 575422 408494
rect 575186 401258 575422 401494
rect 575186 394258 575422 394494
rect 575186 387258 575422 387494
rect 575186 380258 575422 380494
rect 575186 373258 575422 373494
rect 575186 366258 575422 366494
rect 575186 359258 575422 359494
rect 575186 352258 575422 352494
rect 575186 345258 575422 345494
rect 575186 338258 575422 338494
rect 575186 331258 575422 331494
rect 575186 324258 575422 324494
rect 575186 317258 575422 317494
rect 575186 310258 575422 310494
rect 575186 303258 575422 303494
rect 575186 296258 575422 296494
rect 575186 289258 575422 289494
rect 575186 282258 575422 282494
rect 575186 275258 575422 275494
rect 575186 268258 575422 268494
rect 575186 261258 575422 261494
rect 575186 254258 575422 254494
rect 575186 247258 575422 247494
rect 575186 240258 575422 240494
rect 575186 233258 575422 233494
rect 575186 226258 575422 226494
rect 575186 219258 575422 219494
rect 575186 212258 575422 212494
rect 575186 205258 575422 205494
rect 575186 198258 575422 198494
rect 575186 191258 575422 191494
rect 575186 184258 575422 184494
rect 575186 177258 575422 177494
rect 575186 170258 575422 170494
rect 575186 163258 575422 163494
rect 575186 156258 575422 156494
rect 575186 149258 575422 149494
rect 575186 142258 575422 142494
rect 575186 135258 575422 135494
rect 575186 128258 575422 128494
rect 575186 121258 575422 121494
rect 575186 114258 575422 114494
rect 575186 107258 575422 107494
rect 575186 100258 575422 100494
rect 575186 93258 575422 93494
rect 575186 86258 575422 86494
rect 575186 79258 575422 79494
rect 575186 72258 575422 72494
rect 575186 65258 575422 65494
rect 575186 58258 575422 58494
rect 575186 51258 575422 51494
rect 575186 44258 575422 44494
rect 575186 37258 575422 37494
rect 575186 30258 575422 30494
rect 575186 23258 575422 23494
rect 575186 16258 575422 16494
rect 575186 9258 575422 9494
rect 575186 2258 575422 2494
rect 575186 -982 575422 -746
rect 575186 -1302 575422 -1066
rect 576918 705962 577154 706198
rect 576918 705642 577154 705878
rect 576918 696198 577154 696434
rect 576918 689198 577154 689434
rect 576918 682198 577154 682434
rect 576918 675198 577154 675434
rect 576918 668198 577154 668434
rect 576918 661198 577154 661434
rect 576918 654198 577154 654434
rect 576918 647198 577154 647434
rect 576918 640198 577154 640434
rect 576918 633198 577154 633434
rect 576918 626198 577154 626434
rect 576918 619198 577154 619434
rect 576918 612198 577154 612434
rect 576918 605198 577154 605434
rect 576918 598198 577154 598434
rect 576918 591198 577154 591434
rect 576918 584198 577154 584434
rect 576918 577198 577154 577434
rect 576918 570198 577154 570434
rect 576918 563198 577154 563434
rect 576918 556198 577154 556434
rect 576918 549198 577154 549434
rect 576918 542198 577154 542434
rect 576918 535198 577154 535434
rect 576918 528198 577154 528434
rect 576918 521198 577154 521434
rect 576918 514198 577154 514434
rect 576918 507198 577154 507434
rect 576918 500198 577154 500434
rect 576918 493198 577154 493434
rect 576918 486198 577154 486434
rect 576918 479198 577154 479434
rect 576918 472198 577154 472434
rect 576918 465198 577154 465434
rect 576918 458198 577154 458434
rect 576918 451198 577154 451434
rect 576918 444198 577154 444434
rect 576918 437198 577154 437434
rect 576918 430198 577154 430434
rect 576918 423198 577154 423434
rect 576918 416198 577154 416434
rect 576918 409198 577154 409434
rect 576918 402198 577154 402434
rect 576918 395198 577154 395434
rect 576918 388198 577154 388434
rect 576918 381198 577154 381434
rect 576918 374198 577154 374434
rect 576918 367198 577154 367434
rect 576918 360198 577154 360434
rect 576918 353198 577154 353434
rect 576918 346198 577154 346434
rect 576918 339198 577154 339434
rect 576918 332198 577154 332434
rect 576918 325198 577154 325434
rect 576918 318198 577154 318434
rect 576918 311198 577154 311434
rect 576918 304198 577154 304434
rect 576918 297198 577154 297434
rect 576918 290198 577154 290434
rect 576918 283198 577154 283434
rect 576918 276198 577154 276434
rect 576918 269198 577154 269434
rect 576918 262198 577154 262434
rect 576918 255198 577154 255434
rect 576918 248198 577154 248434
rect 576918 241198 577154 241434
rect 576918 234198 577154 234434
rect 576918 227198 577154 227434
rect 576918 220198 577154 220434
rect 576918 213198 577154 213434
rect 576918 206198 577154 206434
rect 576918 199198 577154 199434
rect 576918 192198 577154 192434
rect 576918 185198 577154 185434
rect 576918 178198 577154 178434
rect 576918 171198 577154 171434
rect 576918 164198 577154 164434
rect 576918 157198 577154 157434
rect 576918 150198 577154 150434
rect 576918 143198 577154 143434
rect 576918 136198 577154 136434
rect 576918 129198 577154 129434
rect 576918 122198 577154 122434
rect 576918 115198 577154 115434
rect 576918 108198 577154 108434
rect 576918 101198 577154 101434
rect 576918 94198 577154 94434
rect 576918 87198 577154 87434
rect 576918 80198 577154 80434
rect 576918 73198 577154 73434
rect 576918 66198 577154 66434
rect 576918 59198 577154 59434
rect 576918 52198 577154 52434
rect 576918 45198 577154 45434
rect 576918 38198 577154 38434
rect 576918 31198 577154 31434
rect 576918 24198 577154 24434
rect 576918 17198 577154 17434
rect 576918 10198 577154 10434
rect 576918 3198 577154 3434
rect 576918 -1942 577154 -1706
rect 576918 -2262 577154 -2026
rect 582186 705002 582422 705238
rect 582186 704682 582422 704918
rect 582186 695258 582422 695494
rect 582186 688258 582422 688494
rect 582186 681258 582422 681494
rect 582186 674258 582422 674494
rect 582186 667258 582422 667494
rect 582186 660258 582422 660494
rect 582186 653258 582422 653494
rect 582186 646258 582422 646494
rect 582186 639258 582422 639494
rect 582186 632258 582422 632494
rect 582186 625258 582422 625494
rect 582186 618258 582422 618494
rect 582186 611258 582422 611494
rect 582186 604258 582422 604494
rect 582186 597258 582422 597494
rect 582186 590258 582422 590494
rect 582186 583258 582422 583494
rect 582186 576258 582422 576494
rect 582186 569258 582422 569494
rect 582186 562258 582422 562494
rect 582186 555258 582422 555494
rect 582186 548258 582422 548494
rect 582186 541258 582422 541494
rect 582186 534258 582422 534494
rect 582186 527258 582422 527494
rect 582186 520258 582422 520494
rect 582186 513258 582422 513494
rect 582186 506258 582422 506494
rect 582186 499258 582422 499494
rect 582186 492258 582422 492494
rect 582186 485258 582422 485494
rect 582186 478258 582422 478494
rect 582186 471258 582422 471494
rect 582186 464258 582422 464494
rect 582186 457258 582422 457494
rect 582186 450258 582422 450494
rect 582186 443258 582422 443494
rect 582186 436258 582422 436494
rect 582186 429258 582422 429494
rect 582186 422258 582422 422494
rect 582186 415258 582422 415494
rect 582186 408258 582422 408494
rect 582186 401258 582422 401494
rect 582186 394258 582422 394494
rect 582186 387258 582422 387494
rect 582186 380258 582422 380494
rect 582186 373258 582422 373494
rect 582186 366258 582422 366494
rect 582186 359258 582422 359494
rect 582186 352258 582422 352494
rect 582186 345258 582422 345494
rect 582186 338258 582422 338494
rect 582186 331258 582422 331494
rect 582186 324258 582422 324494
rect 582186 317258 582422 317494
rect 582186 310258 582422 310494
rect 582186 303258 582422 303494
rect 582186 296258 582422 296494
rect 582186 289258 582422 289494
rect 582186 282258 582422 282494
rect 582186 275258 582422 275494
rect 582186 268258 582422 268494
rect 582186 261258 582422 261494
rect 582186 254258 582422 254494
rect 582186 247258 582422 247494
rect 582186 240258 582422 240494
rect 582186 233258 582422 233494
rect 582186 226258 582422 226494
rect 582186 219258 582422 219494
rect 582186 212258 582422 212494
rect 582186 205258 582422 205494
rect 582186 198258 582422 198494
rect 582186 191258 582422 191494
rect 582186 184258 582422 184494
rect 582186 177258 582422 177494
rect 582186 170258 582422 170494
rect 582186 163258 582422 163494
rect 582186 156258 582422 156494
rect 582186 149258 582422 149494
rect 582186 142258 582422 142494
rect 582186 135258 582422 135494
rect 582186 128258 582422 128494
rect 582186 121258 582422 121494
rect 582186 114258 582422 114494
rect 582186 107258 582422 107494
rect 582186 100258 582422 100494
rect 582186 93258 582422 93494
rect 582186 86258 582422 86494
rect 582186 79258 582422 79494
rect 582186 72258 582422 72494
rect 582186 65258 582422 65494
rect 582186 58258 582422 58494
rect 582186 51258 582422 51494
rect 582186 44258 582422 44494
rect 582186 37258 582422 37494
rect 582186 30258 582422 30494
rect 582186 23258 582422 23494
rect 582186 16258 582422 16494
rect 582186 9258 582422 9494
rect 582186 2258 582422 2494
rect 582186 -982 582422 -746
rect 582186 -1302 582422 -1066
rect 585818 705002 586054 705238
rect 586138 705002 586374 705238
rect 586458 705002 586694 705238
rect 586778 705002 587014 705238
rect 585818 704682 586054 704918
rect 586138 704682 586374 704918
rect 586458 704682 586694 704918
rect 586778 704682 587014 704918
rect 585818 695258 586054 695494
rect 586138 695258 586374 695494
rect 586458 695258 586694 695494
rect 586778 695258 587014 695494
rect 585818 688258 586054 688494
rect 586138 688258 586374 688494
rect 586458 688258 586694 688494
rect 586778 688258 587014 688494
rect 585818 681258 586054 681494
rect 586138 681258 586374 681494
rect 586458 681258 586694 681494
rect 586778 681258 587014 681494
rect 585818 674258 586054 674494
rect 586138 674258 586374 674494
rect 586458 674258 586694 674494
rect 586778 674258 587014 674494
rect 585818 667258 586054 667494
rect 586138 667258 586374 667494
rect 586458 667258 586694 667494
rect 586778 667258 587014 667494
rect 585818 660258 586054 660494
rect 586138 660258 586374 660494
rect 586458 660258 586694 660494
rect 586778 660258 587014 660494
rect 585818 653258 586054 653494
rect 586138 653258 586374 653494
rect 586458 653258 586694 653494
rect 586778 653258 587014 653494
rect 585818 646258 586054 646494
rect 586138 646258 586374 646494
rect 586458 646258 586694 646494
rect 586778 646258 587014 646494
rect 585818 639258 586054 639494
rect 586138 639258 586374 639494
rect 586458 639258 586694 639494
rect 586778 639258 587014 639494
rect 585818 632258 586054 632494
rect 586138 632258 586374 632494
rect 586458 632258 586694 632494
rect 586778 632258 587014 632494
rect 585818 625258 586054 625494
rect 586138 625258 586374 625494
rect 586458 625258 586694 625494
rect 586778 625258 587014 625494
rect 585818 618258 586054 618494
rect 586138 618258 586374 618494
rect 586458 618258 586694 618494
rect 586778 618258 587014 618494
rect 585818 611258 586054 611494
rect 586138 611258 586374 611494
rect 586458 611258 586694 611494
rect 586778 611258 587014 611494
rect 585818 604258 586054 604494
rect 586138 604258 586374 604494
rect 586458 604258 586694 604494
rect 586778 604258 587014 604494
rect 585818 597258 586054 597494
rect 586138 597258 586374 597494
rect 586458 597258 586694 597494
rect 586778 597258 587014 597494
rect 585818 590258 586054 590494
rect 586138 590258 586374 590494
rect 586458 590258 586694 590494
rect 586778 590258 587014 590494
rect 585818 583258 586054 583494
rect 586138 583258 586374 583494
rect 586458 583258 586694 583494
rect 586778 583258 587014 583494
rect 585818 576258 586054 576494
rect 586138 576258 586374 576494
rect 586458 576258 586694 576494
rect 586778 576258 587014 576494
rect 585818 569258 586054 569494
rect 586138 569258 586374 569494
rect 586458 569258 586694 569494
rect 586778 569258 587014 569494
rect 585818 562258 586054 562494
rect 586138 562258 586374 562494
rect 586458 562258 586694 562494
rect 586778 562258 587014 562494
rect 585818 555258 586054 555494
rect 586138 555258 586374 555494
rect 586458 555258 586694 555494
rect 586778 555258 587014 555494
rect 585818 548258 586054 548494
rect 586138 548258 586374 548494
rect 586458 548258 586694 548494
rect 586778 548258 587014 548494
rect 585818 541258 586054 541494
rect 586138 541258 586374 541494
rect 586458 541258 586694 541494
rect 586778 541258 587014 541494
rect 585818 534258 586054 534494
rect 586138 534258 586374 534494
rect 586458 534258 586694 534494
rect 586778 534258 587014 534494
rect 585818 527258 586054 527494
rect 586138 527258 586374 527494
rect 586458 527258 586694 527494
rect 586778 527258 587014 527494
rect 585818 520258 586054 520494
rect 586138 520258 586374 520494
rect 586458 520258 586694 520494
rect 586778 520258 587014 520494
rect 585818 513258 586054 513494
rect 586138 513258 586374 513494
rect 586458 513258 586694 513494
rect 586778 513258 587014 513494
rect 585818 506258 586054 506494
rect 586138 506258 586374 506494
rect 586458 506258 586694 506494
rect 586778 506258 587014 506494
rect 585818 499258 586054 499494
rect 586138 499258 586374 499494
rect 586458 499258 586694 499494
rect 586778 499258 587014 499494
rect 585818 492258 586054 492494
rect 586138 492258 586374 492494
rect 586458 492258 586694 492494
rect 586778 492258 587014 492494
rect 585818 485258 586054 485494
rect 586138 485258 586374 485494
rect 586458 485258 586694 485494
rect 586778 485258 587014 485494
rect 585818 478258 586054 478494
rect 586138 478258 586374 478494
rect 586458 478258 586694 478494
rect 586778 478258 587014 478494
rect 585818 471258 586054 471494
rect 586138 471258 586374 471494
rect 586458 471258 586694 471494
rect 586778 471258 587014 471494
rect 585818 464258 586054 464494
rect 586138 464258 586374 464494
rect 586458 464258 586694 464494
rect 586778 464258 587014 464494
rect 585818 457258 586054 457494
rect 586138 457258 586374 457494
rect 586458 457258 586694 457494
rect 586778 457258 587014 457494
rect 585818 450258 586054 450494
rect 586138 450258 586374 450494
rect 586458 450258 586694 450494
rect 586778 450258 587014 450494
rect 585818 443258 586054 443494
rect 586138 443258 586374 443494
rect 586458 443258 586694 443494
rect 586778 443258 587014 443494
rect 585818 436258 586054 436494
rect 586138 436258 586374 436494
rect 586458 436258 586694 436494
rect 586778 436258 587014 436494
rect 585818 429258 586054 429494
rect 586138 429258 586374 429494
rect 586458 429258 586694 429494
rect 586778 429258 587014 429494
rect 585818 422258 586054 422494
rect 586138 422258 586374 422494
rect 586458 422258 586694 422494
rect 586778 422258 587014 422494
rect 585818 415258 586054 415494
rect 586138 415258 586374 415494
rect 586458 415258 586694 415494
rect 586778 415258 587014 415494
rect 585818 408258 586054 408494
rect 586138 408258 586374 408494
rect 586458 408258 586694 408494
rect 586778 408258 587014 408494
rect 585818 401258 586054 401494
rect 586138 401258 586374 401494
rect 586458 401258 586694 401494
rect 586778 401258 587014 401494
rect 585818 394258 586054 394494
rect 586138 394258 586374 394494
rect 586458 394258 586694 394494
rect 586778 394258 587014 394494
rect 585818 387258 586054 387494
rect 586138 387258 586374 387494
rect 586458 387258 586694 387494
rect 586778 387258 587014 387494
rect 585818 380258 586054 380494
rect 586138 380258 586374 380494
rect 586458 380258 586694 380494
rect 586778 380258 587014 380494
rect 585818 373258 586054 373494
rect 586138 373258 586374 373494
rect 586458 373258 586694 373494
rect 586778 373258 587014 373494
rect 585818 366258 586054 366494
rect 586138 366258 586374 366494
rect 586458 366258 586694 366494
rect 586778 366258 587014 366494
rect 585818 359258 586054 359494
rect 586138 359258 586374 359494
rect 586458 359258 586694 359494
rect 586778 359258 587014 359494
rect 585818 352258 586054 352494
rect 586138 352258 586374 352494
rect 586458 352258 586694 352494
rect 586778 352258 587014 352494
rect 585818 345258 586054 345494
rect 586138 345258 586374 345494
rect 586458 345258 586694 345494
rect 586778 345258 587014 345494
rect 585818 338258 586054 338494
rect 586138 338258 586374 338494
rect 586458 338258 586694 338494
rect 586778 338258 587014 338494
rect 585818 331258 586054 331494
rect 586138 331258 586374 331494
rect 586458 331258 586694 331494
rect 586778 331258 587014 331494
rect 585818 324258 586054 324494
rect 586138 324258 586374 324494
rect 586458 324258 586694 324494
rect 586778 324258 587014 324494
rect 585818 317258 586054 317494
rect 586138 317258 586374 317494
rect 586458 317258 586694 317494
rect 586778 317258 587014 317494
rect 585818 310258 586054 310494
rect 586138 310258 586374 310494
rect 586458 310258 586694 310494
rect 586778 310258 587014 310494
rect 585818 303258 586054 303494
rect 586138 303258 586374 303494
rect 586458 303258 586694 303494
rect 586778 303258 587014 303494
rect 585818 296258 586054 296494
rect 586138 296258 586374 296494
rect 586458 296258 586694 296494
rect 586778 296258 587014 296494
rect 585818 289258 586054 289494
rect 586138 289258 586374 289494
rect 586458 289258 586694 289494
rect 586778 289258 587014 289494
rect 585818 282258 586054 282494
rect 586138 282258 586374 282494
rect 586458 282258 586694 282494
rect 586778 282258 587014 282494
rect 585818 275258 586054 275494
rect 586138 275258 586374 275494
rect 586458 275258 586694 275494
rect 586778 275258 587014 275494
rect 585818 268258 586054 268494
rect 586138 268258 586374 268494
rect 586458 268258 586694 268494
rect 586778 268258 587014 268494
rect 585818 261258 586054 261494
rect 586138 261258 586374 261494
rect 586458 261258 586694 261494
rect 586778 261258 587014 261494
rect 585818 254258 586054 254494
rect 586138 254258 586374 254494
rect 586458 254258 586694 254494
rect 586778 254258 587014 254494
rect 585818 247258 586054 247494
rect 586138 247258 586374 247494
rect 586458 247258 586694 247494
rect 586778 247258 587014 247494
rect 585818 240258 586054 240494
rect 586138 240258 586374 240494
rect 586458 240258 586694 240494
rect 586778 240258 587014 240494
rect 585818 233258 586054 233494
rect 586138 233258 586374 233494
rect 586458 233258 586694 233494
rect 586778 233258 587014 233494
rect 585818 226258 586054 226494
rect 586138 226258 586374 226494
rect 586458 226258 586694 226494
rect 586778 226258 587014 226494
rect 585818 219258 586054 219494
rect 586138 219258 586374 219494
rect 586458 219258 586694 219494
rect 586778 219258 587014 219494
rect 585818 212258 586054 212494
rect 586138 212258 586374 212494
rect 586458 212258 586694 212494
rect 586778 212258 587014 212494
rect 585818 205258 586054 205494
rect 586138 205258 586374 205494
rect 586458 205258 586694 205494
rect 586778 205258 587014 205494
rect 585818 198258 586054 198494
rect 586138 198258 586374 198494
rect 586458 198258 586694 198494
rect 586778 198258 587014 198494
rect 585818 191258 586054 191494
rect 586138 191258 586374 191494
rect 586458 191258 586694 191494
rect 586778 191258 587014 191494
rect 585818 184258 586054 184494
rect 586138 184258 586374 184494
rect 586458 184258 586694 184494
rect 586778 184258 587014 184494
rect 585818 177258 586054 177494
rect 586138 177258 586374 177494
rect 586458 177258 586694 177494
rect 586778 177258 587014 177494
rect 585818 170258 586054 170494
rect 586138 170258 586374 170494
rect 586458 170258 586694 170494
rect 586778 170258 587014 170494
rect 585818 163258 586054 163494
rect 586138 163258 586374 163494
rect 586458 163258 586694 163494
rect 586778 163258 587014 163494
rect 585818 156258 586054 156494
rect 586138 156258 586374 156494
rect 586458 156258 586694 156494
rect 586778 156258 587014 156494
rect 585818 149258 586054 149494
rect 586138 149258 586374 149494
rect 586458 149258 586694 149494
rect 586778 149258 587014 149494
rect 585818 142258 586054 142494
rect 586138 142258 586374 142494
rect 586458 142258 586694 142494
rect 586778 142258 587014 142494
rect 585818 135258 586054 135494
rect 586138 135258 586374 135494
rect 586458 135258 586694 135494
rect 586778 135258 587014 135494
rect 585818 128258 586054 128494
rect 586138 128258 586374 128494
rect 586458 128258 586694 128494
rect 586778 128258 587014 128494
rect 585818 121258 586054 121494
rect 586138 121258 586374 121494
rect 586458 121258 586694 121494
rect 586778 121258 587014 121494
rect 585818 114258 586054 114494
rect 586138 114258 586374 114494
rect 586458 114258 586694 114494
rect 586778 114258 587014 114494
rect 585818 107258 586054 107494
rect 586138 107258 586374 107494
rect 586458 107258 586694 107494
rect 586778 107258 587014 107494
rect 585818 100258 586054 100494
rect 586138 100258 586374 100494
rect 586458 100258 586694 100494
rect 586778 100258 587014 100494
rect 585818 93258 586054 93494
rect 586138 93258 586374 93494
rect 586458 93258 586694 93494
rect 586778 93258 587014 93494
rect 585818 86258 586054 86494
rect 586138 86258 586374 86494
rect 586458 86258 586694 86494
rect 586778 86258 587014 86494
rect 585818 79258 586054 79494
rect 586138 79258 586374 79494
rect 586458 79258 586694 79494
rect 586778 79258 587014 79494
rect 585818 72258 586054 72494
rect 586138 72258 586374 72494
rect 586458 72258 586694 72494
rect 586778 72258 587014 72494
rect 585818 65258 586054 65494
rect 586138 65258 586374 65494
rect 586458 65258 586694 65494
rect 586778 65258 587014 65494
rect 585818 58258 586054 58494
rect 586138 58258 586374 58494
rect 586458 58258 586694 58494
rect 586778 58258 587014 58494
rect 585818 51258 586054 51494
rect 586138 51258 586374 51494
rect 586458 51258 586694 51494
rect 586778 51258 587014 51494
rect 585818 44258 586054 44494
rect 586138 44258 586374 44494
rect 586458 44258 586694 44494
rect 586778 44258 587014 44494
rect 585818 37258 586054 37494
rect 586138 37258 586374 37494
rect 586458 37258 586694 37494
rect 586778 37258 587014 37494
rect 585818 30258 586054 30494
rect 586138 30258 586374 30494
rect 586458 30258 586694 30494
rect 586778 30258 587014 30494
rect 585818 23258 586054 23494
rect 586138 23258 586374 23494
rect 586458 23258 586694 23494
rect 586778 23258 587014 23494
rect 585818 16258 586054 16494
rect 586138 16258 586374 16494
rect 586458 16258 586694 16494
rect 586778 16258 587014 16494
rect 585818 9258 586054 9494
rect 586138 9258 586374 9494
rect 586458 9258 586694 9494
rect 586778 9258 587014 9494
rect 585818 2258 586054 2494
rect 586138 2258 586374 2494
rect 586458 2258 586694 2494
rect 586778 2258 587014 2494
rect 585818 -982 586054 -746
rect 586138 -982 586374 -746
rect 586458 -982 586694 -746
rect 586778 -982 587014 -746
rect 585818 -1302 586054 -1066
rect 586138 -1302 586374 -1066
rect 586458 -1302 586694 -1066
rect 586778 -1302 587014 -1066
rect 587570 696198 587806 696434
rect 587890 696198 588126 696434
rect 588210 696198 588446 696434
rect 588530 696198 588766 696434
rect 587570 689198 587806 689434
rect 587890 689198 588126 689434
rect 588210 689198 588446 689434
rect 588530 689198 588766 689434
rect 587570 682198 587806 682434
rect 587890 682198 588126 682434
rect 588210 682198 588446 682434
rect 588530 682198 588766 682434
rect 587570 675198 587806 675434
rect 587890 675198 588126 675434
rect 588210 675198 588446 675434
rect 588530 675198 588766 675434
rect 587570 668198 587806 668434
rect 587890 668198 588126 668434
rect 588210 668198 588446 668434
rect 588530 668198 588766 668434
rect 587570 661198 587806 661434
rect 587890 661198 588126 661434
rect 588210 661198 588446 661434
rect 588530 661198 588766 661434
rect 587570 654198 587806 654434
rect 587890 654198 588126 654434
rect 588210 654198 588446 654434
rect 588530 654198 588766 654434
rect 587570 647198 587806 647434
rect 587890 647198 588126 647434
rect 588210 647198 588446 647434
rect 588530 647198 588766 647434
rect 587570 640198 587806 640434
rect 587890 640198 588126 640434
rect 588210 640198 588446 640434
rect 588530 640198 588766 640434
rect 587570 633198 587806 633434
rect 587890 633198 588126 633434
rect 588210 633198 588446 633434
rect 588530 633198 588766 633434
rect 587570 626198 587806 626434
rect 587890 626198 588126 626434
rect 588210 626198 588446 626434
rect 588530 626198 588766 626434
rect 587570 619198 587806 619434
rect 587890 619198 588126 619434
rect 588210 619198 588446 619434
rect 588530 619198 588766 619434
rect 587570 612198 587806 612434
rect 587890 612198 588126 612434
rect 588210 612198 588446 612434
rect 588530 612198 588766 612434
rect 587570 605198 587806 605434
rect 587890 605198 588126 605434
rect 588210 605198 588446 605434
rect 588530 605198 588766 605434
rect 587570 598198 587806 598434
rect 587890 598198 588126 598434
rect 588210 598198 588446 598434
rect 588530 598198 588766 598434
rect 587570 591198 587806 591434
rect 587890 591198 588126 591434
rect 588210 591198 588446 591434
rect 588530 591198 588766 591434
rect 587570 584198 587806 584434
rect 587890 584198 588126 584434
rect 588210 584198 588446 584434
rect 588530 584198 588766 584434
rect 587570 577198 587806 577434
rect 587890 577198 588126 577434
rect 588210 577198 588446 577434
rect 588530 577198 588766 577434
rect 587570 570198 587806 570434
rect 587890 570198 588126 570434
rect 588210 570198 588446 570434
rect 588530 570198 588766 570434
rect 587570 563198 587806 563434
rect 587890 563198 588126 563434
rect 588210 563198 588446 563434
rect 588530 563198 588766 563434
rect 587570 556198 587806 556434
rect 587890 556198 588126 556434
rect 588210 556198 588446 556434
rect 588530 556198 588766 556434
rect 587570 549198 587806 549434
rect 587890 549198 588126 549434
rect 588210 549198 588446 549434
rect 588530 549198 588766 549434
rect 587570 542198 587806 542434
rect 587890 542198 588126 542434
rect 588210 542198 588446 542434
rect 588530 542198 588766 542434
rect 587570 535198 587806 535434
rect 587890 535198 588126 535434
rect 588210 535198 588446 535434
rect 588530 535198 588766 535434
rect 587570 528198 587806 528434
rect 587890 528198 588126 528434
rect 588210 528198 588446 528434
rect 588530 528198 588766 528434
rect 587570 521198 587806 521434
rect 587890 521198 588126 521434
rect 588210 521198 588446 521434
rect 588530 521198 588766 521434
rect 587570 514198 587806 514434
rect 587890 514198 588126 514434
rect 588210 514198 588446 514434
rect 588530 514198 588766 514434
rect 587570 507198 587806 507434
rect 587890 507198 588126 507434
rect 588210 507198 588446 507434
rect 588530 507198 588766 507434
rect 587570 500198 587806 500434
rect 587890 500198 588126 500434
rect 588210 500198 588446 500434
rect 588530 500198 588766 500434
rect 587570 493198 587806 493434
rect 587890 493198 588126 493434
rect 588210 493198 588446 493434
rect 588530 493198 588766 493434
rect 587570 486198 587806 486434
rect 587890 486198 588126 486434
rect 588210 486198 588446 486434
rect 588530 486198 588766 486434
rect 587570 479198 587806 479434
rect 587890 479198 588126 479434
rect 588210 479198 588446 479434
rect 588530 479198 588766 479434
rect 587570 472198 587806 472434
rect 587890 472198 588126 472434
rect 588210 472198 588446 472434
rect 588530 472198 588766 472434
rect 587570 465198 587806 465434
rect 587890 465198 588126 465434
rect 588210 465198 588446 465434
rect 588530 465198 588766 465434
rect 587570 458198 587806 458434
rect 587890 458198 588126 458434
rect 588210 458198 588446 458434
rect 588530 458198 588766 458434
rect 587570 451198 587806 451434
rect 587890 451198 588126 451434
rect 588210 451198 588446 451434
rect 588530 451198 588766 451434
rect 587570 444198 587806 444434
rect 587890 444198 588126 444434
rect 588210 444198 588446 444434
rect 588530 444198 588766 444434
rect 587570 437198 587806 437434
rect 587890 437198 588126 437434
rect 588210 437198 588446 437434
rect 588530 437198 588766 437434
rect 587570 430198 587806 430434
rect 587890 430198 588126 430434
rect 588210 430198 588446 430434
rect 588530 430198 588766 430434
rect 587570 423198 587806 423434
rect 587890 423198 588126 423434
rect 588210 423198 588446 423434
rect 588530 423198 588766 423434
rect 587570 416198 587806 416434
rect 587890 416198 588126 416434
rect 588210 416198 588446 416434
rect 588530 416198 588766 416434
rect 587570 409198 587806 409434
rect 587890 409198 588126 409434
rect 588210 409198 588446 409434
rect 588530 409198 588766 409434
rect 587570 402198 587806 402434
rect 587890 402198 588126 402434
rect 588210 402198 588446 402434
rect 588530 402198 588766 402434
rect 587570 395198 587806 395434
rect 587890 395198 588126 395434
rect 588210 395198 588446 395434
rect 588530 395198 588766 395434
rect 587570 388198 587806 388434
rect 587890 388198 588126 388434
rect 588210 388198 588446 388434
rect 588530 388198 588766 388434
rect 587570 381198 587806 381434
rect 587890 381198 588126 381434
rect 588210 381198 588446 381434
rect 588530 381198 588766 381434
rect 587570 374198 587806 374434
rect 587890 374198 588126 374434
rect 588210 374198 588446 374434
rect 588530 374198 588766 374434
rect 587570 367198 587806 367434
rect 587890 367198 588126 367434
rect 588210 367198 588446 367434
rect 588530 367198 588766 367434
rect 587570 360198 587806 360434
rect 587890 360198 588126 360434
rect 588210 360198 588446 360434
rect 588530 360198 588766 360434
rect 587570 353198 587806 353434
rect 587890 353198 588126 353434
rect 588210 353198 588446 353434
rect 588530 353198 588766 353434
rect 587570 346198 587806 346434
rect 587890 346198 588126 346434
rect 588210 346198 588446 346434
rect 588530 346198 588766 346434
rect 587570 339198 587806 339434
rect 587890 339198 588126 339434
rect 588210 339198 588446 339434
rect 588530 339198 588766 339434
rect 587570 332198 587806 332434
rect 587890 332198 588126 332434
rect 588210 332198 588446 332434
rect 588530 332198 588766 332434
rect 587570 325198 587806 325434
rect 587890 325198 588126 325434
rect 588210 325198 588446 325434
rect 588530 325198 588766 325434
rect 587570 318198 587806 318434
rect 587890 318198 588126 318434
rect 588210 318198 588446 318434
rect 588530 318198 588766 318434
rect 587570 311198 587806 311434
rect 587890 311198 588126 311434
rect 588210 311198 588446 311434
rect 588530 311198 588766 311434
rect 587570 304198 587806 304434
rect 587890 304198 588126 304434
rect 588210 304198 588446 304434
rect 588530 304198 588766 304434
rect 587570 297198 587806 297434
rect 587890 297198 588126 297434
rect 588210 297198 588446 297434
rect 588530 297198 588766 297434
rect 587570 290198 587806 290434
rect 587890 290198 588126 290434
rect 588210 290198 588446 290434
rect 588530 290198 588766 290434
rect 587570 283198 587806 283434
rect 587890 283198 588126 283434
rect 588210 283198 588446 283434
rect 588530 283198 588766 283434
rect 587570 276198 587806 276434
rect 587890 276198 588126 276434
rect 588210 276198 588446 276434
rect 588530 276198 588766 276434
rect 587570 269198 587806 269434
rect 587890 269198 588126 269434
rect 588210 269198 588446 269434
rect 588530 269198 588766 269434
rect 587570 262198 587806 262434
rect 587890 262198 588126 262434
rect 588210 262198 588446 262434
rect 588530 262198 588766 262434
rect 587570 255198 587806 255434
rect 587890 255198 588126 255434
rect 588210 255198 588446 255434
rect 588530 255198 588766 255434
rect 587570 248198 587806 248434
rect 587890 248198 588126 248434
rect 588210 248198 588446 248434
rect 588530 248198 588766 248434
rect 587570 241198 587806 241434
rect 587890 241198 588126 241434
rect 588210 241198 588446 241434
rect 588530 241198 588766 241434
rect 587570 234198 587806 234434
rect 587890 234198 588126 234434
rect 588210 234198 588446 234434
rect 588530 234198 588766 234434
rect 587570 227198 587806 227434
rect 587890 227198 588126 227434
rect 588210 227198 588446 227434
rect 588530 227198 588766 227434
rect 587570 220198 587806 220434
rect 587890 220198 588126 220434
rect 588210 220198 588446 220434
rect 588530 220198 588766 220434
rect 587570 213198 587806 213434
rect 587890 213198 588126 213434
rect 588210 213198 588446 213434
rect 588530 213198 588766 213434
rect 587570 206198 587806 206434
rect 587890 206198 588126 206434
rect 588210 206198 588446 206434
rect 588530 206198 588766 206434
rect 587570 199198 587806 199434
rect 587890 199198 588126 199434
rect 588210 199198 588446 199434
rect 588530 199198 588766 199434
rect 587570 192198 587806 192434
rect 587890 192198 588126 192434
rect 588210 192198 588446 192434
rect 588530 192198 588766 192434
rect 587570 185198 587806 185434
rect 587890 185198 588126 185434
rect 588210 185198 588446 185434
rect 588530 185198 588766 185434
rect 587570 178198 587806 178434
rect 587890 178198 588126 178434
rect 588210 178198 588446 178434
rect 588530 178198 588766 178434
rect 587570 171198 587806 171434
rect 587890 171198 588126 171434
rect 588210 171198 588446 171434
rect 588530 171198 588766 171434
rect 587570 164198 587806 164434
rect 587890 164198 588126 164434
rect 588210 164198 588446 164434
rect 588530 164198 588766 164434
rect 587570 157198 587806 157434
rect 587890 157198 588126 157434
rect 588210 157198 588446 157434
rect 588530 157198 588766 157434
rect 587570 150198 587806 150434
rect 587890 150198 588126 150434
rect 588210 150198 588446 150434
rect 588530 150198 588766 150434
rect 587570 143198 587806 143434
rect 587890 143198 588126 143434
rect 588210 143198 588446 143434
rect 588530 143198 588766 143434
rect 587570 136198 587806 136434
rect 587890 136198 588126 136434
rect 588210 136198 588446 136434
rect 588530 136198 588766 136434
rect 587570 129198 587806 129434
rect 587890 129198 588126 129434
rect 588210 129198 588446 129434
rect 588530 129198 588766 129434
rect 587570 122198 587806 122434
rect 587890 122198 588126 122434
rect 588210 122198 588446 122434
rect 588530 122198 588766 122434
rect 587570 115198 587806 115434
rect 587890 115198 588126 115434
rect 588210 115198 588446 115434
rect 588530 115198 588766 115434
rect 587570 108198 587806 108434
rect 587890 108198 588126 108434
rect 588210 108198 588446 108434
rect 588530 108198 588766 108434
rect 587570 101198 587806 101434
rect 587890 101198 588126 101434
rect 588210 101198 588446 101434
rect 588530 101198 588766 101434
rect 587570 94198 587806 94434
rect 587890 94198 588126 94434
rect 588210 94198 588446 94434
rect 588530 94198 588766 94434
rect 587570 87198 587806 87434
rect 587890 87198 588126 87434
rect 588210 87198 588446 87434
rect 588530 87198 588766 87434
rect 587570 80198 587806 80434
rect 587890 80198 588126 80434
rect 588210 80198 588446 80434
rect 588530 80198 588766 80434
rect 587570 73198 587806 73434
rect 587890 73198 588126 73434
rect 588210 73198 588446 73434
rect 588530 73198 588766 73434
rect 587570 66198 587806 66434
rect 587890 66198 588126 66434
rect 588210 66198 588446 66434
rect 588530 66198 588766 66434
rect 587570 59198 587806 59434
rect 587890 59198 588126 59434
rect 588210 59198 588446 59434
rect 588530 59198 588766 59434
rect 587570 52198 587806 52434
rect 587890 52198 588126 52434
rect 588210 52198 588446 52434
rect 588530 52198 588766 52434
rect 587570 45198 587806 45434
rect 587890 45198 588126 45434
rect 588210 45198 588446 45434
rect 588530 45198 588766 45434
rect 587570 38198 587806 38434
rect 587890 38198 588126 38434
rect 588210 38198 588446 38434
rect 588530 38198 588766 38434
rect 587570 31198 587806 31434
rect 587890 31198 588126 31434
rect 588210 31198 588446 31434
rect 588530 31198 588766 31434
rect 587570 24198 587806 24434
rect 587890 24198 588126 24434
rect 588210 24198 588446 24434
rect 588530 24198 588766 24434
rect 587570 17198 587806 17434
rect 587890 17198 588126 17434
rect 588210 17198 588446 17434
rect 588530 17198 588766 17434
rect 587570 10198 587806 10434
rect 587890 10198 588126 10434
rect 588210 10198 588446 10434
rect 588530 10198 588766 10434
rect 587570 3198 587806 3434
rect 587890 3198 588126 3434
rect 588210 3198 588446 3434
rect 588530 3198 588766 3434
<< metal5 >>
rect -3366 706198 587290 706230
rect -3366 705962 2918 706198
rect 3154 705962 9918 706198
rect 10154 705962 16918 706198
rect 17154 705962 23918 706198
rect 24154 705962 30918 706198
rect 31154 705962 37918 706198
rect 38154 705962 44918 706198
rect 45154 705962 51918 706198
rect 52154 705962 58918 706198
rect 59154 705962 65918 706198
rect 66154 705962 72918 706198
rect 73154 705962 79918 706198
rect 80154 705962 86918 706198
rect 87154 705962 93918 706198
rect 94154 705962 100918 706198
rect 101154 705962 107918 706198
rect 108154 705962 114918 706198
rect 115154 705962 121918 706198
rect 122154 705962 128918 706198
rect 129154 705962 135918 706198
rect 136154 705962 142918 706198
rect 143154 705962 149918 706198
rect 150154 705962 156918 706198
rect 157154 705962 163918 706198
rect 164154 705962 170918 706198
rect 171154 705962 177918 706198
rect 178154 705962 184918 706198
rect 185154 705962 191918 706198
rect 192154 705962 198918 706198
rect 199154 705962 205918 706198
rect 206154 705962 212918 706198
rect 213154 705962 219918 706198
rect 220154 705962 226918 706198
rect 227154 705962 233918 706198
rect 234154 705962 240918 706198
rect 241154 705962 247918 706198
rect 248154 705962 254918 706198
rect 255154 705962 261918 706198
rect 262154 705962 268918 706198
rect 269154 705962 275918 706198
rect 276154 705962 282918 706198
rect 283154 705962 289918 706198
rect 290154 705962 296918 706198
rect 297154 705962 303918 706198
rect 304154 705962 310918 706198
rect 311154 705962 317918 706198
rect 318154 705962 324918 706198
rect 325154 705962 331918 706198
rect 332154 705962 338918 706198
rect 339154 705962 345918 706198
rect 346154 705962 352918 706198
rect 353154 705962 359918 706198
rect 360154 705962 366918 706198
rect 367154 705962 373918 706198
rect 374154 705962 380918 706198
rect 381154 705962 387918 706198
rect 388154 705962 394918 706198
rect 395154 705962 401918 706198
rect 402154 705962 408918 706198
rect 409154 705962 415918 706198
rect 416154 705962 422918 706198
rect 423154 705962 429918 706198
rect 430154 705962 436918 706198
rect 437154 705962 443918 706198
rect 444154 705962 450918 706198
rect 451154 705962 457918 706198
rect 458154 705962 464918 706198
rect 465154 705962 471918 706198
rect 472154 705962 478918 706198
rect 479154 705962 485918 706198
rect 486154 705962 492918 706198
rect 493154 705962 499918 706198
rect 500154 705962 506918 706198
rect 507154 705962 513918 706198
rect 514154 705962 520918 706198
rect 521154 705962 527918 706198
rect 528154 705962 534918 706198
rect 535154 705962 541918 706198
rect 542154 705962 548918 706198
rect 549154 705962 555918 706198
rect 556154 705962 562918 706198
rect 563154 705962 569918 706198
rect 570154 705962 576918 706198
rect 577154 705962 587290 706198
rect -3366 705878 587290 705962
rect -3366 705642 2918 705878
rect 3154 705642 9918 705878
rect 10154 705642 16918 705878
rect 17154 705642 23918 705878
rect 24154 705642 30918 705878
rect 31154 705642 37918 705878
rect 38154 705642 44918 705878
rect 45154 705642 51918 705878
rect 52154 705642 58918 705878
rect 59154 705642 65918 705878
rect 66154 705642 72918 705878
rect 73154 705642 79918 705878
rect 80154 705642 86918 705878
rect 87154 705642 93918 705878
rect 94154 705642 100918 705878
rect 101154 705642 107918 705878
rect 108154 705642 114918 705878
rect 115154 705642 121918 705878
rect 122154 705642 128918 705878
rect 129154 705642 135918 705878
rect 136154 705642 142918 705878
rect 143154 705642 149918 705878
rect 150154 705642 156918 705878
rect 157154 705642 163918 705878
rect 164154 705642 170918 705878
rect 171154 705642 177918 705878
rect 178154 705642 184918 705878
rect 185154 705642 191918 705878
rect 192154 705642 198918 705878
rect 199154 705642 205918 705878
rect 206154 705642 212918 705878
rect 213154 705642 219918 705878
rect 220154 705642 226918 705878
rect 227154 705642 233918 705878
rect 234154 705642 240918 705878
rect 241154 705642 247918 705878
rect 248154 705642 254918 705878
rect 255154 705642 261918 705878
rect 262154 705642 268918 705878
rect 269154 705642 275918 705878
rect 276154 705642 282918 705878
rect 283154 705642 289918 705878
rect 290154 705642 296918 705878
rect 297154 705642 303918 705878
rect 304154 705642 310918 705878
rect 311154 705642 317918 705878
rect 318154 705642 324918 705878
rect 325154 705642 331918 705878
rect 332154 705642 338918 705878
rect 339154 705642 345918 705878
rect 346154 705642 352918 705878
rect 353154 705642 359918 705878
rect 360154 705642 366918 705878
rect 367154 705642 373918 705878
rect 374154 705642 380918 705878
rect 381154 705642 387918 705878
rect 388154 705642 394918 705878
rect 395154 705642 401918 705878
rect 402154 705642 408918 705878
rect 409154 705642 415918 705878
rect 416154 705642 422918 705878
rect 423154 705642 429918 705878
rect 430154 705642 436918 705878
rect 437154 705642 443918 705878
rect 444154 705642 450918 705878
rect 451154 705642 457918 705878
rect 458154 705642 464918 705878
rect 465154 705642 471918 705878
rect 472154 705642 478918 705878
rect 479154 705642 485918 705878
rect 486154 705642 492918 705878
rect 493154 705642 499918 705878
rect 500154 705642 506918 705878
rect 507154 705642 513918 705878
rect 514154 705642 520918 705878
rect 521154 705642 527918 705878
rect 528154 705642 534918 705878
rect 535154 705642 541918 705878
rect 542154 705642 548918 705878
rect 549154 705642 555918 705878
rect 556154 705642 562918 705878
rect 563154 705642 569918 705878
rect 570154 705642 576918 705878
rect 577154 705642 587290 705878
rect -3366 705610 587290 705642
rect -2406 705238 587122 705270
rect -2406 705002 -2374 705238
rect -2138 705002 -2054 705238
rect -1818 705002 1186 705238
rect 1422 705002 8186 705238
rect 8422 705002 15186 705238
rect 15422 705002 22186 705238
rect 22422 705002 29186 705238
rect 29422 705002 36186 705238
rect 36422 705002 43186 705238
rect 43422 705002 50186 705238
rect 50422 705002 57186 705238
rect 57422 705002 64186 705238
rect 64422 705002 71186 705238
rect 71422 705002 78186 705238
rect 78422 705002 85186 705238
rect 85422 705002 92186 705238
rect 92422 705002 99186 705238
rect 99422 705002 106186 705238
rect 106422 705002 113186 705238
rect 113422 705002 120186 705238
rect 120422 705002 127186 705238
rect 127422 705002 134186 705238
rect 134422 705002 141186 705238
rect 141422 705002 148186 705238
rect 148422 705002 155186 705238
rect 155422 705002 162186 705238
rect 162422 705002 169186 705238
rect 169422 705002 176186 705238
rect 176422 705002 183186 705238
rect 183422 705002 190186 705238
rect 190422 705002 197186 705238
rect 197422 705002 204186 705238
rect 204422 705002 211186 705238
rect 211422 705002 218186 705238
rect 218422 705002 225186 705238
rect 225422 705002 232186 705238
rect 232422 705002 239186 705238
rect 239422 705002 246186 705238
rect 246422 705002 253186 705238
rect 253422 705002 260186 705238
rect 260422 705002 267186 705238
rect 267422 705002 274186 705238
rect 274422 705002 281186 705238
rect 281422 705002 288186 705238
rect 288422 705002 295186 705238
rect 295422 705002 302186 705238
rect 302422 705002 309186 705238
rect 309422 705002 316186 705238
rect 316422 705002 323186 705238
rect 323422 705002 330186 705238
rect 330422 705002 337186 705238
rect 337422 705002 344186 705238
rect 344422 705002 351186 705238
rect 351422 705002 358186 705238
rect 358422 705002 365186 705238
rect 365422 705002 372186 705238
rect 372422 705002 379186 705238
rect 379422 705002 386186 705238
rect 386422 705002 393186 705238
rect 393422 705002 400186 705238
rect 400422 705002 407186 705238
rect 407422 705002 414186 705238
rect 414422 705002 421186 705238
rect 421422 705002 428186 705238
rect 428422 705002 435186 705238
rect 435422 705002 442186 705238
rect 442422 705002 449186 705238
rect 449422 705002 456186 705238
rect 456422 705002 463186 705238
rect 463422 705002 470186 705238
rect 470422 705002 477186 705238
rect 477422 705002 484186 705238
rect 484422 705002 491186 705238
rect 491422 705002 498186 705238
rect 498422 705002 505186 705238
rect 505422 705002 512186 705238
rect 512422 705002 519186 705238
rect 519422 705002 526186 705238
rect 526422 705002 533186 705238
rect 533422 705002 540186 705238
rect 540422 705002 547186 705238
rect 547422 705002 554186 705238
rect 554422 705002 561186 705238
rect 561422 705002 568186 705238
rect 568422 705002 575186 705238
rect 575422 705002 582186 705238
rect 582422 705002 585818 705238
rect 586054 705002 586138 705238
rect 586374 705002 586458 705238
rect 586694 705002 586778 705238
rect 587014 705002 587122 705238
rect -2406 704918 587122 705002
rect -2406 704682 -2374 704918
rect -2138 704682 -2054 704918
rect -1818 704682 1186 704918
rect 1422 704682 8186 704918
rect 8422 704682 15186 704918
rect 15422 704682 22186 704918
rect 22422 704682 29186 704918
rect 29422 704682 36186 704918
rect 36422 704682 43186 704918
rect 43422 704682 50186 704918
rect 50422 704682 57186 704918
rect 57422 704682 64186 704918
rect 64422 704682 71186 704918
rect 71422 704682 78186 704918
rect 78422 704682 85186 704918
rect 85422 704682 92186 704918
rect 92422 704682 99186 704918
rect 99422 704682 106186 704918
rect 106422 704682 113186 704918
rect 113422 704682 120186 704918
rect 120422 704682 127186 704918
rect 127422 704682 134186 704918
rect 134422 704682 141186 704918
rect 141422 704682 148186 704918
rect 148422 704682 155186 704918
rect 155422 704682 162186 704918
rect 162422 704682 169186 704918
rect 169422 704682 176186 704918
rect 176422 704682 183186 704918
rect 183422 704682 190186 704918
rect 190422 704682 197186 704918
rect 197422 704682 204186 704918
rect 204422 704682 211186 704918
rect 211422 704682 218186 704918
rect 218422 704682 225186 704918
rect 225422 704682 232186 704918
rect 232422 704682 239186 704918
rect 239422 704682 246186 704918
rect 246422 704682 253186 704918
rect 253422 704682 260186 704918
rect 260422 704682 267186 704918
rect 267422 704682 274186 704918
rect 274422 704682 281186 704918
rect 281422 704682 288186 704918
rect 288422 704682 295186 704918
rect 295422 704682 302186 704918
rect 302422 704682 309186 704918
rect 309422 704682 316186 704918
rect 316422 704682 323186 704918
rect 323422 704682 330186 704918
rect 330422 704682 337186 704918
rect 337422 704682 344186 704918
rect 344422 704682 351186 704918
rect 351422 704682 358186 704918
rect 358422 704682 365186 704918
rect 365422 704682 372186 704918
rect 372422 704682 379186 704918
rect 379422 704682 386186 704918
rect 386422 704682 393186 704918
rect 393422 704682 400186 704918
rect 400422 704682 407186 704918
rect 407422 704682 414186 704918
rect 414422 704682 421186 704918
rect 421422 704682 428186 704918
rect 428422 704682 435186 704918
rect 435422 704682 442186 704918
rect 442422 704682 449186 704918
rect 449422 704682 456186 704918
rect 456422 704682 463186 704918
rect 463422 704682 470186 704918
rect 470422 704682 477186 704918
rect 477422 704682 484186 704918
rect 484422 704682 491186 704918
rect 491422 704682 498186 704918
rect 498422 704682 505186 704918
rect 505422 704682 512186 704918
rect 512422 704682 519186 704918
rect 519422 704682 526186 704918
rect 526422 704682 533186 704918
rect 533422 704682 540186 704918
rect 540422 704682 547186 704918
rect 547422 704682 554186 704918
rect 554422 704682 561186 704918
rect 561422 704682 568186 704918
rect 568422 704682 575186 704918
rect 575422 704682 582186 704918
rect 582422 704682 585818 704918
rect 586054 704682 586138 704918
rect 586374 704682 586458 704918
rect 586694 704682 586778 704918
rect 587014 704682 587122 704918
rect -2406 704650 587122 704682
rect -4950 696434 588874 696476
rect -4950 696198 -4842 696434
rect -4606 696198 -4522 696434
rect -4286 696198 -4202 696434
rect -3966 696198 -3882 696434
rect -3646 696198 2918 696434
rect 3154 696198 9918 696434
rect 10154 696198 16918 696434
rect 17154 696198 23918 696434
rect 24154 696198 30918 696434
rect 31154 696198 37918 696434
rect 38154 696198 44918 696434
rect 45154 696198 51918 696434
rect 52154 696198 58918 696434
rect 59154 696198 65918 696434
rect 66154 696198 72918 696434
rect 73154 696198 79918 696434
rect 80154 696198 86918 696434
rect 87154 696198 93918 696434
rect 94154 696198 100918 696434
rect 101154 696198 107918 696434
rect 108154 696198 114918 696434
rect 115154 696198 121918 696434
rect 122154 696198 128918 696434
rect 129154 696198 135918 696434
rect 136154 696198 142918 696434
rect 143154 696198 149918 696434
rect 150154 696198 156918 696434
rect 157154 696198 163918 696434
rect 164154 696198 170918 696434
rect 171154 696198 177918 696434
rect 178154 696198 184918 696434
rect 185154 696198 191918 696434
rect 192154 696198 198918 696434
rect 199154 696198 205918 696434
rect 206154 696198 212918 696434
rect 213154 696198 219918 696434
rect 220154 696198 226918 696434
rect 227154 696198 233918 696434
rect 234154 696198 240918 696434
rect 241154 696198 247918 696434
rect 248154 696198 254918 696434
rect 255154 696198 261918 696434
rect 262154 696198 268918 696434
rect 269154 696198 275918 696434
rect 276154 696198 282918 696434
rect 283154 696198 289918 696434
rect 290154 696198 296918 696434
rect 297154 696198 303918 696434
rect 304154 696198 310918 696434
rect 311154 696198 317918 696434
rect 318154 696198 324918 696434
rect 325154 696198 331918 696434
rect 332154 696198 338918 696434
rect 339154 696198 345918 696434
rect 346154 696198 352918 696434
rect 353154 696198 359918 696434
rect 360154 696198 366918 696434
rect 367154 696198 373918 696434
rect 374154 696198 380918 696434
rect 381154 696198 387918 696434
rect 388154 696198 394918 696434
rect 395154 696198 401918 696434
rect 402154 696198 408918 696434
rect 409154 696198 415918 696434
rect 416154 696198 422918 696434
rect 423154 696198 429918 696434
rect 430154 696198 436918 696434
rect 437154 696198 443918 696434
rect 444154 696198 450918 696434
rect 451154 696198 457918 696434
rect 458154 696198 464918 696434
rect 465154 696198 471918 696434
rect 472154 696198 478918 696434
rect 479154 696198 485918 696434
rect 486154 696198 492918 696434
rect 493154 696198 499918 696434
rect 500154 696198 506918 696434
rect 507154 696198 513918 696434
rect 514154 696198 520918 696434
rect 521154 696198 527918 696434
rect 528154 696198 534918 696434
rect 535154 696198 541918 696434
rect 542154 696198 548918 696434
rect 549154 696198 555918 696434
rect 556154 696198 562918 696434
rect 563154 696198 569918 696434
rect 570154 696198 576918 696434
rect 577154 696198 587570 696434
rect 587806 696198 587890 696434
rect 588126 696198 588210 696434
rect 588446 696198 588530 696434
rect 588766 696198 588874 696434
rect -4950 696156 588874 696198
rect -4950 695494 588874 695536
rect -4950 695258 -3090 695494
rect -2854 695258 -2770 695494
rect -2534 695258 -2450 695494
rect -2214 695258 -2130 695494
rect -1894 695258 1186 695494
rect 1422 695258 8186 695494
rect 8422 695258 15186 695494
rect 15422 695258 22186 695494
rect 22422 695258 29186 695494
rect 29422 695258 36186 695494
rect 36422 695258 43186 695494
rect 43422 695258 50186 695494
rect 50422 695258 57186 695494
rect 57422 695258 64186 695494
rect 64422 695258 71186 695494
rect 71422 695258 78186 695494
rect 78422 695258 85186 695494
rect 85422 695258 92186 695494
rect 92422 695258 99186 695494
rect 99422 695258 106186 695494
rect 106422 695258 113186 695494
rect 113422 695258 120186 695494
rect 120422 695258 127186 695494
rect 127422 695258 134186 695494
rect 134422 695258 141186 695494
rect 141422 695258 148186 695494
rect 148422 695258 155186 695494
rect 155422 695258 162186 695494
rect 162422 695258 169186 695494
rect 169422 695258 176186 695494
rect 176422 695258 183186 695494
rect 183422 695258 190186 695494
rect 190422 695258 197186 695494
rect 197422 695258 204186 695494
rect 204422 695258 211186 695494
rect 211422 695258 218186 695494
rect 218422 695258 225186 695494
rect 225422 695258 232186 695494
rect 232422 695258 239186 695494
rect 239422 695258 246186 695494
rect 246422 695258 253186 695494
rect 253422 695258 260186 695494
rect 260422 695258 267186 695494
rect 267422 695258 274186 695494
rect 274422 695258 281186 695494
rect 281422 695258 288186 695494
rect 288422 695258 295186 695494
rect 295422 695258 302186 695494
rect 302422 695258 309186 695494
rect 309422 695258 316186 695494
rect 316422 695258 323186 695494
rect 323422 695258 330186 695494
rect 330422 695258 337186 695494
rect 337422 695258 344186 695494
rect 344422 695258 351186 695494
rect 351422 695258 358186 695494
rect 358422 695258 365186 695494
rect 365422 695258 372186 695494
rect 372422 695258 379186 695494
rect 379422 695258 386186 695494
rect 386422 695258 393186 695494
rect 393422 695258 400186 695494
rect 400422 695258 407186 695494
rect 407422 695258 414186 695494
rect 414422 695258 421186 695494
rect 421422 695258 428186 695494
rect 428422 695258 435186 695494
rect 435422 695258 442186 695494
rect 442422 695258 449186 695494
rect 449422 695258 456186 695494
rect 456422 695258 463186 695494
rect 463422 695258 470186 695494
rect 470422 695258 477186 695494
rect 477422 695258 484186 695494
rect 484422 695258 491186 695494
rect 491422 695258 498186 695494
rect 498422 695258 505186 695494
rect 505422 695258 512186 695494
rect 512422 695258 519186 695494
rect 519422 695258 526186 695494
rect 526422 695258 533186 695494
rect 533422 695258 540186 695494
rect 540422 695258 547186 695494
rect 547422 695258 554186 695494
rect 554422 695258 561186 695494
rect 561422 695258 568186 695494
rect 568422 695258 575186 695494
rect 575422 695258 582186 695494
rect 582422 695258 585818 695494
rect 586054 695258 586138 695494
rect 586374 695258 586458 695494
rect 586694 695258 586778 695494
rect 587014 695258 588874 695494
rect -4950 695216 588874 695258
rect -4950 689434 588874 689476
rect -4950 689198 -4842 689434
rect -4606 689198 -4522 689434
rect -4286 689198 -4202 689434
rect -3966 689198 -3882 689434
rect -3646 689198 2918 689434
rect 3154 689198 9918 689434
rect 10154 689198 16918 689434
rect 17154 689198 23918 689434
rect 24154 689198 30918 689434
rect 31154 689198 37918 689434
rect 38154 689198 44918 689434
rect 45154 689198 51918 689434
rect 52154 689198 58918 689434
rect 59154 689198 65918 689434
rect 66154 689198 72918 689434
rect 73154 689198 79918 689434
rect 80154 689198 86918 689434
rect 87154 689198 93918 689434
rect 94154 689198 100918 689434
rect 101154 689198 107918 689434
rect 108154 689198 114918 689434
rect 115154 689198 121918 689434
rect 122154 689198 128918 689434
rect 129154 689198 135918 689434
rect 136154 689198 142918 689434
rect 143154 689198 149918 689434
rect 150154 689198 156918 689434
rect 157154 689198 163918 689434
rect 164154 689198 170918 689434
rect 171154 689198 177918 689434
rect 178154 689198 184918 689434
rect 185154 689198 191918 689434
rect 192154 689198 198918 689434
rect 199154 689198 205918 689434
rect 206154 689198 212918 689434
rect 213154 689198 219918 689434
rect 220154 689198 226918 689434
rect 227154 689198 233918 689434
rect 234154 689198 240918 689434
rect 241154 689198 247918 689434
rect 248154 689198 254918 689434
rect 255154 689198 261918 689434
rect 262154 689198 268918 689434
rect 269154 689198 275918 689434
rect 276154 689198 282918 689434
rect 283154 689198 289918 689434
rect 290154 689198 296918 689434
rect 297154 689198 303918 689434
rect 304154 689198 310918 689434
rect 311154 689198 317918 689434
rect 318154 689198 324918 689434
rect 325154 689198 331918 689434
rect 332154 689198 338918 689434
rect 339154 689198 345918 689434
rect 346154 689198 352918 689434
rect 353154 689198 359918 689434
rect 360154 689198 366918 689434
rect 367154 689198 373918 689434
rect 374154 689198 380918 689434
rect 381154 689198 387918 689434
rect 388154 689198 394918 689434
rect 395154 689198 401918 689434
rect 402154 689198 408918 689434
rect 409154 689198 415918 689434
rect 416154 689198 422918 689434
rect 423154 689198 429918 689434
rect 430154 689198 436918 689434
rect 437154 689198 443918 689434
rect 444154 689198 450918 689434
rect 451154 689198 457918 689434
rect 458154 689198 464918 689434
rect 465154 689198 471918 689434
rect 472154 689198 478918 689434
rect 479154 689198 485918 689434
rect 486154 689198 492918 689434
rect 493154 689198 499918 689434
rect 500154 689198 506918 689434
rect 507154 689198 513918 689434
rect 514154 689198 520918 689434
rect 521154 689198 527918 689434
rect 528154 689198 534918 689434
rect 535154 689198 541918 689434
rect 542154 689198 548918 689434
rect 549154 689198 555918 689434
rect 556154 689198 562918 689434
rect 563154 689198 569918 689434
rect 570154 689198 576918 689434
rect 577154 689198 587570 689434
rect 587806 689198 587890 689434
rect 588126 689198 588210 689434
rect 588446 689198 588530 689434
rect 588766 689198 588874 689434
rect -4950 689156 588874 689198
rect -4950 688494 588874 688536
rect -4950 688258 -3090 688494
rect -2854 688258 -2770 688494
rect -2534 688258 -2450 688494
rect -2214 688258 -2130 688494
rect -1894 688258 1186 688494
rect 1422 688258 8186 688494
rect 8422 688258 15186 688494
rect 15422 688258 22186 688494
rect 22422 688258 29186 688494
rect 29422 688258 36186 688494
rect 36422 688258 43186 688494
rect 43422 688258 50186 688494
rect 50422 688258 57186 688494
rect 57422 688258 64186 688494
rect 64422 688258 71186 688494
rect 71422 688258 78186 688494
rect 78422 688258 85186 688494
rect 85422 688258 92186 688494
rect 92422 688258 99186 688494
rect 99422 688258 106186 688494
rect 106422 688258 113186 688494
rect 113422 688258 120186 688494
rect 120422 688258 127186 688494
rect 127422 688258 134186 688494
rect 134422 688258 141186 688494
rect 141422 688258 148186 688494
rect 148422 688258 155186 688494
rect 155422 688258 162186 688494
rect 162422 688258 169186 688494
rect 169422 688258 176186 688494
rect 176422 688258 183186 688494
rect 183422 688258 190186 688494
rect 190422 688258 197186 688494
rect 197422 688258 204186 688494
rect 204422 688258 211186 688494
rect 211422 688258 218186 688494
rect 218422 688258 225186 688494
rect 225422 688258 232186 688494
rect 232422 688258 239186 688494
rect 239422 688258 246186 688494
rect 246422 688258 253186 688494
rect 253422 688258 260186 688494
rect 260422 688258 267186 688494
rect 267422 688258 274186 688494
rect 274422 688258 281186 688494
rect 281422 688258 288186 688494
rect 288422 688258 295186 688494
rect 295422 688258 302186 688494
rect 302422 688258 309186 688494
rect 309422 688258 316186 688494
rect 316422 688258 323186 688494
rect 323422 688258 330186 688494
rect 330422 688258 337186 688494
rect 337422 688258 344186 688494
rect 344422 688258 351186 688494
rect 351422 688258 358186 688494
rect 358422 688258 365186 688494
rect 365422 688258 372186 688494
rect 372422 688258 379186 688494
rect 379422 688258 386186 688494
rect 386422 688258 393186 688494
rect 393422 688258 400186 688494
rect 400422 688258 407186 688494
rect 407422 688258 414186 688494
rect 414422 688258 421186 688494
rect 421422 688258 428186 688494
rect 428422 688258 435186 688494
rect 435422 688258 442186 688494
rect 442422 688258 449186 688494
rect 449422 688258 456186 688494
rect 456422 688258 463186 688494
rect 463422 688258 470186 688494
rect 470422 688258 477186 688494
rect 477422 688258 484186 688494
rect 484422 688258 491186 688494
rect 491422 688258 498186 688494
rect 498422 688258 505186 688494
rect 505422 688258 512186 688494
rect 512422 688258 519186 688494
rect 519422 688258 526186 688494
rect 526422 688258 533186 688494
rect 533422 688258 540186 688494
rect 540422 688258 547186 688494
rect 547422 688258 554186 688494
rect 554422 688258 561186 688494
rect 561422 688258 568186 688494
rect 568422 688258 575186 688494
rect 575422 688258 582186 688494
rect 582422 688258 585818 688494
rect 586054 688258 586138 688494
rect 586374 688258 586458 688494
rect 586694 688258 586778 688494
rect 587014 688258 588874 688494
rect -4950 688216 588874 688258
rect -4950 682434 588874 682476
rect -4950 682198 -4842 682434
rect -4606 682198 -4522 682434
rect -4286 682198 -4202 682434
rect -3966 682198 -3882 682434
rect -3646 682198 2918 682434
rect 3154 682198 9918 682434
rect 10154 682198 16918 682434
rect 17154 682198 23918 682434
rect 24154 682198 30918 682434
rect 31154 682198 37918 682434
rect 38154 682198 44918 682434
rect 45154 682198 51918 682434
rect 52154 682198 58918 682434
rect 59154 682198 65918 682434
rect 66154 682198 72918 682434
rect 73154 682198 79918 682434
rect 80154 682198 86918 682434
rect 87154 682198 93918 682434
rect 94154 682198 100918 682434
rect 101154 682198 107918 682434
rect 108154 682198 114918 682434
rect 115154 682198 121918 682434
rect 122154 682198 128918 682434
rect 129154 682198 135918 682434
rect 136154 682198 142918 682434
rect 143154 682198 149918 682434
rect 150154 682198 156918 682434
rect 157154 682198 163918 682434
rect 164154 682198 170918 682434
rect 171154 682198 177918 682434
rect 178154 682198 184918 682434
rect 185154 682198 191918 682434
rect 192154 682198 198918 682434
rect 199154 682198 205918 682434
rect 206154 682198 212918 682434
rect 213154 682198 219918 682434
rect 220154 682198 226918 682434
rect 227154 682198 233918 682434
rect 234154 682198 240918 682434
rect 241154 682198 247918 682434
rect 248154 682198 254918 682434
rect 255154 682198 261918 682434
rect 262154 682198 268918 682434
rect 269154 682198 275918 682434
rect 276154 682198 282918 682434
rect 283154 682198 289918 682434
rect 290154 682198 296918 682434
rect 297154 682198 303918 682434
rect 304154 682198 310918 682434
rect 311154 682198 317918 682434
rect 318154 682198 324918 682434
rect 325154 682198 331918 682434
rect 332154 682198 338918 682434
rect 339154 682198 345918 682434
rect 346154 682198 352918 682434
rect 353154 682198 359918 682434
rect 360154 682198 366918 682434
rect 367154 682198 373918 682434
rect 374154 682198 380918 682434
rect 381154 682198 387918 682434
rect 388154 682198 394918 682434
rect 395154 682198 401918 682434
rect 402154 682198 408918 682434
rect 409154 682198 415918 682434
rect 416154 682198 422918 682434
rect 423154 682198 429918 682434
rect 430154 682198 436918 682434
rect 437154 682198 443918 682434
rect 444154 682198 450918 682434
rect 451154 682198 457918 682434
rect 458154 682198 464918 682434
rect 465154 682198 471918 682434
rect 472154 682198 478918 682434
rect 479154 682198 485918 682434
rect 486154 682198 492918 682434
rect 493154 682198 499918 682434
rect 500154 682198 506918 682434
rect 507154 682198 513918 682434
rect 514154 682198 520918 682434
rect 521154 682198 527918 682434
rect 528154 682198 534918 682434
rect 535154 682198 541918 682434
rect 542154 682198 548918 682434
rect 549154 682198 555918 682434
rect 556154 682198 562918 682434
rect 563154 682198 569918 682434
rect 570154 682198 576918 682434
rect 577154 682198 587570 682434
rect 587806 682198 587890 682434
rect 588126 682198 588210 682434
rect 588446 682198 588530 682434
rect 588766 682198 588874 682434
rect -4950 682156 588874 682198
rect -4950 681494 588874 681536
rect -4950 681258 -3090 681494
rect -2854 681258 -2770 681494
rect -2534 681258 -2450 681494
rect -2214 681258 -2130 681494
rect -1894 681258 1186 681494
rect 1422 681258 8186 681494
rect 8422 681258 15186 681494
rect 15422 681258 22186 681494
rect 22422 681258 29186 681494
rect 29422 681258 36186 681494
rect 36422 681258 43186 681494
rect 43422 681258 50186 681494
rect 50422 681258 57186 681494
rect 57422 681258 64186 681494
rect 64422 681258 71186 681494
rect 71422 681258 78186 681494
rect 78422 681258 85186 681494
rect 85422 681258 92186 681494
rect 92422 681258 99186 681494
rect 99422 681258 106186 681494
rect 106422 681258 113186 681494
rect 113422 681258 120186 681494
rect 120422 681258 127186 681494
rect 127422 681258 134186 681494
rect 134422 681258 141186 681494
rect 141422 681258 148186 681494
rect 148422 681258 155186 681494
rect 155422 681258 162186 681494
rect 162422 681258 169186 681494
rect 169422 681258 176186 681494
rect 176422 681258 183186 681494
rect 183422 681258 190186 681494
rect 190422 681258 197186 681494
rect 197422 681258 204186 681494
rect 204422 681258 211186 681494
rect 211422 681258 218186 681494
rect 218422 681258 225186 681494
rect 225422 681258 232186 681494
rect 232422 681258 239186 681494
rect 239422 681258 246186 681494
rect 246422 681258 253186 681494
rect 253422 681258 260186 681494
rect 260422 681258 267186 681494
rect 267422 681258 274186 681494
rect 274422 681258 281186 681494
rect 281422 681258 288186 681494
rect 288422 681258 295186 681494
rect 295422 681258 302186 681494
rect 302422 681258 309186 681494
rect 309422 681258 316186 681494
rect 316422 681258 323186 681494
rect 323422 681258 330186 681494
rect 330422 681258 337186 681494
rect 337422 681258 344186 681494
rect 344422 681258 351186 681494
rect 351422 681258 358186 681494
rect 358422 681258 365186 681494
rect 365422 681258 372186 681494
rect 372422 681258 379186 681494
rect 379422 681258 386186 681494
rect 386422 681258 393186 681494
rect 393422 681258 400186 681494
rect 400422 681258 407186 681494
rect 407422 681258 414186 681494
rect 414422 681258 421186 681494
rect 421422 681258 428186 681494
rect 428422 681258 435186 681494
rect 435422 681258 442186 681494
rect 442422 681258 449186 681494
rect 449422 681258 456186 681494
rect 456422 681258 463186 681494
rect 463422 681258 470186 681494
rect 470422 681258 477186 681494
rect 477422 681258 484186 681494
rect 484422 681258 491186 681494
rect 491422 681258 498186 681494
rect 498422 681258 505186 681494
rect 505422 681258 512186 681494
rect 512422 681258 519186 681494
rect 519422 681258 526186 681494
rect 526422 681258 533186 681494
rect 533422 681258 540186 681494
rect 540422 681258 547186 681494
rect 547422 681258 554186 681494
rect 554422 681258 561186 681494
rect 561422 681258 568186 681494
rect 568422 681258 575186 681494
rect 575422 681258 582186 681494
rect 582422 681258 585818 681494
rect 586054 681258 586138 681494
rect 586374 681258 586458 681494
rect 586694 681258 586778 681494
rect 587014 681258 588874 681494
rect -4950 681216 588874 681258
rect -4950 675434 588874 675476
rect -4950 675198 -4842 675434
rect -4606 675198 -4522 675434
rect -4286 675198 -4202 675434
rect -3966 675198 -3882 675434
rect -3646 675198 2918 675434
rect 3154 675198 9918 675434
rect 10154 675198 16918 675434
rect 17154 675198 23918 675434
rect 24154 675198 30918 675434
rect 31154 675198 37918 675434
rect 38154 675198 44918 675434
rect 45154 675198 51918 675434
rect 52154 675198 58918 675434
rect 59154 675198 65918 675434
rect 66154 675198 72918 675434
rect 73154 675198 79918 675434
rect 80154 675198 86918 675434
rect 87154 675198 93918 675434
rect 94154 675198 100918 675434
rect 101154 675198 107918 675434
rect 108154 675198 114918 675434
rect 115154 675198 121918 675434
rect 122154 675198 128918 675434
rect 129154 675198 135918 675434
rect 136154 675198 142918 675434
rect 143154 675198 149918 675434
rect 150154 675198 156918 675434
rect 157154 675198 163918 675434
rect 164154 675198 170918 675434
rect 171154 675198 177918 675434
rect 178154 675198 184918 675434
rect 185154 675198 191918 675434
rect 192154 675198 198918 675434
rect 199154 675198 205918 675434
rect 206154 675198 212918 675434
rect 213154 675198 219918 675434
rect 220154 675198 226918 675434
rect 227154 675198 233918 675434
rect 234154 675198 240918 675434
rect 241154 675198 247918 675434
rect 248154 675198 254918 675434
rect 255154 675198 261918 675434
rect 262154 675198 268918 675434
rect 269154 675198 275918 675434
rect 276154 675198 282918 675434
rect 283154 675198 289918 675434
rect 290154 675198 296918 675434
rect 297154 675198 303918 675434
rect 304154 675198 310918 675434
rect 311154 675198 317918 675434
rect 318154 675198 324918 675434
rect 325154 675198 331918 675434
rect 332154 675198 338918 675434
rect 339154 675198 345918 675434
rect 346154 675198 352918 675434
rect 353154 675198 359918 675434
rect 360154 675198 366918 675434
rect 367154 675198 373918 675434
rect 374154 675198 380918 675434
rect 381154 675198 387918 675434
rect 388154 675198 394918 675434
rect 395154 675198 401918 675434
rect 402154 675198 408918 675434
rect 409154 675198 415918 675434
rect 416154 675198 422918 675434
rect 423154 675198 429918 675434
rect 430154 675198 436918 675434
rect 437154 675198 443918 675434
rect 444154 675198 450918 675434
rect 451154 675198 457918 675434
rect 458154 675198 464918 675434
rect 465154 675198 471918 675434
rect 472154 675198 478918 675434
rect 479154 675198 485918 675434
rect 486154 675198 492918 675434
rect 493154 675198 499918 675434
rect 500154 675198 506918 675434
rect 507154 675198 513918 675434
rect 514154 675198 520918 675434
rect 521154 675198 527918 675434
rect 528154 675198 534918 675434
rect 535154 675198 541918 675434
rect 542154 675198 548918 675434
rect 549154 675198 555918 675434
rect 556154 675198 562918 675434
rect 563154 675198 569918 675434
rect 570154 675198 576918 675434
rect 577154 675198 587570 675434
rect 587806 675198 587890 675434
rect 588126 675198 588210 675434
rect 588446 675198 588530 675434
rect 588766 675198 588874 675434
rect -4950 675156 588874 675198
rect -4950 674494 588874 674536
rect -4950 674258 -3090 674494
rect -2854 674258 -2770 674494
rect -2534 674258 -2450 674494
rect -2214 674258 -2130 674494
rect -1894 674258 1186 674494
rect 1422 674258 8186 674494
rect 8422 674258 15186 674494
rect 15422 674258 22186 674494
rect 22422 674258 29186 674494
rect 29422 674258 36186 674494
rect 36422 674258 43186 674494
rect 43422 674258 50186 674494
rect 50422 674258 57186 674494
rect 57422 674258 64186 674494
rect 64422 674258 71186 674494
rect 71422 674258 78186 674494
rect 78422 674258 85186 674494
rect 85422 674258 92186 674494
rect 92422 674258 99186 674494
rect 99422 674258 106186 674494
rect 106422 674258 113186 674494
rect 113422 674258 120186 674494
rect 120422 674258 127186 674494
rect 127422 674258 134186 674494
rect 134422 674258 141186 674494
rect 141422 674258 148186 674494
rect 148422 674258 155186 674494
rect 155422 674258 162186 674494
rect 162422 674258 169186 674494
rect 169422 674258 176186 674494
rect 176422 674258 183186 674494
rect 183422 674258 190186 674494
rect 190422 674258 197186 674494
rect 197422 674258 204186 674494
rect 204422 674258 211186 674494
rect 211422 674258 218186 674494
rect 218422 674258 225186 674494
rect 225422 674258 232186 674494
rect 232422 674258 239186 674494
rect 239422 674258 246186 674494
rect 246422 674258 253186 674494
rect 253422 674258 260186 674494
rect 260422 674258 267186 674494
rect 267422 674258 274186 674494
rect 274422 674258 281186 674494
rect 281422 674258 288186 674494
rect 288422 674258 295186 674494
rect 295422 674258 302186 674494
rect 302422 674258 309186 674494
rect 309422 674258 316186 674494
rect 316422 674258 323186 674494
rect 323422 674258 330186 674494
rect 330422 674258 337186 674494
rect 337422 674258 344186 674494
rect 344422 674258 351186 674494
rect 351422 674258 358186 674494
rect 358422 674258 365186 674494
rect 365422 674258 372186 674494
rect 372422 674258 379186 674494
rect 379422 674258 386186 674494
rect 386422 674258 393186 674494
rect 393422 674258 400186 674494
rect 400422 674258 407186 674494
rect 407422 674258 414186 674494
rect 414422 674258 421186 674494
rect 421422 674258 428186 674494
rect 428422 674258 435186 674494
rect 435422 674258 442186 674494
rect 442422 674258 449186 674494
rect 449422 674258 456186 674494
rect 456422 674258 463186 674494
rect 463422 674258 470186 674494
rect 470422 674258 477186 674494
rect 477422 674258 484186 674494
rect 484422 674258 491186 674494
rect 491422 674258 498186 674494
rect 498422 674258 505186 674494
rect 505422 674258 512186 674494
rect 512422 674258 519186 674494
rect 519422 674258 526186 674494
rect 526422 674258 533186 674494
rect 533422 674258 540186 674494
rect 540422 674258 547186 674494
rect 547422 674258 554186 674494
rect 554422 674258 561186 674494
rect 561422 674258 568186 674494
rect 568422 674258 575186 674494
rect 575422 674258 582186 674494
rect 582422 674258 585818 674494
rect 586054 674258 586138 674494
rect 586374 674258 586458 674494
rect 586694 674258 586778 674494
rect 587014 674258 588874 674494
rect -4950 674216 588874 674258
rect -4950 668434 588874 668476
rect -4950 668198 -4842 668434
rect -4606 668198 -4522 668434
rect -4286 668198 -4202 668434
rect -3966 668198 -3882 668434
rect -3646 668198 2918 668434
rect 3154 668198 9918 668434
rect 10154 668198 16918 668434
rect 17154 668198 23918 668434
rect 24154 668198 30918 668434
rect 31154 668198 37918 668434
rect 38154 668198 44918 668434
rect 45154 668198 51918 668434
rect 52154 668198 58918 668434
rect 59154 668198 65918 668434
rect 66154 668198 72918 668434
rect 73154 668198 79918 668434
rect 80154 668198 86918 668434
rect 87154 668198 93918 668434
rect 94154 668198 100918 668434
rect 101154 668198 107918 668434
rect 108154 668198 114918 668434
rect 115154 668198 121918 668434
rect 122154 668198 128918 668434
rect 129154 668198 135918 668434
rect 136154 668198 142918 668434
rect 143154 668198 149918 668434
rect 150154 668198 156918 668434
rect 157154 668198 163918 668434
rect 164154 668198 170918 668434
rect 171154 668198 177918 668434
rect 178154 668198 184918 668434
rect 185154 668198 191918 668434
rect 192154 668198 198918 668434
rect 199154 668198 205918 668434
rect 206154 668198 212918 668434
rect 213154 668198 219918 668434
rect 220154 668198 226918 668434
rect 227154 668198 233918 668434
rect 234154 668198 240918 668434
rect 241154 668198 247918 668434
rect 248154 668198 254918 668434
rect 255154 668198 261918 668434
rect 262154 668198 268918 668434
rect 269154 668198 275918 668434
rect 276154 668198 282918 668434
rect 283154 668198 289918 668434
rect 290154 668198 296918 668434
rect 297154 668198 303918 668434
rect 304154 668198 310918 668434
rect 311154 668198 317918 668434
rect 318154 668198 324918 668434
rect 325154 668198 331918 668434
rect 332154 668198 338918 668434
rect 339154 668198 345918 668434
rect 346154 668198 352918 668434
rect 353154 668198 359918 668434
rect 360154 668198 366918 668434
rect 367154 668198 373918 668434
rect 374154 668198 380918 668434
rect 381154 668198 387918 668434
rect 388154 668198 394918 668434
rect 395154 668198 401918 668434
rect 402154 668198 408918 668434
rect 409154 668198 415918 668434
rect 416154 668198 422918 668434
rect 423154 668198 429918 668434
rect 430154 668198 436918 668434
rect 437154 668198 443918 668434
rect 444154 668198 450918 668434
rect 451154 668198 457918 668434
rect 458154 668198 464918 668434
rect 465154 668198 471918 668434
rect 472154 668198 478918 668434
rect 479154 668198 485918 668434
rect 486154 668198 492918 668434
rect 493154 668198 499918 668434
rect 500154 668198 506918 668434
rect 507154 668198 513918 668434
rect 514154 668198 520918 668434
rect 521154 668198 527918 668434
rect 528154 668198 534918 668434
rect 535154 668198 541918 668434
rect 542154 668198 548918 668434
rect 549154 668198 555918 668434
rect 556154 668198 562918 668434
rect 563154 668198 569918 668434
rect 570154 668198 576918 668434
rect 577154 668198 587570 668434
rect 587806 668198 587890 668434
rect 588126 668198 588210 668434
rect 588446 668198 588530 668434
rect 588766 668198 588874 668434
rect -4950 668156 588874 668198
rect -4950 667494 588874 667536
rect -4950 667258 -3090 667494
rect -2854 667258 -2770 667494
rect -2534 667258 -2450 667494
rect -2214 667258 -2130 667494
rect -1894 667258 1186 667494
rect 1422 667258 8186 667494
rect 8422 667258 15186 667494
rect 15422 667258 22186 667494
rect 22422 667258 29186 667494
rect 29422 667258 36186 667494
rect 36422 667258 43186 667494
rect 43422 667258 50186 667494
rect 50422 667258 57186 667494
rect 57422 667258 64186 667494
rect 64422 667258 71186 667494
rect 71422 667258 78186 667494
rect 78422 667258 85186 667494
rect 85422 667258 92186 667494
rect 92422 667258 99186 667494
rect 99422 667258 106186 667494
rect 106422 667258 113186 667494
rect 113422 667258 120186 667494
rect 120422 667258 127186 667494
rect 127422 667258 134186 667494
rect 134422 667258 141186 667494
rect 141422 667258 148186 667494
rect 148422 667258 155186 667494
rect 155422 667258 162186 667494
rect 162422 667258 169186 667494
rect 169422 667258 176186 667494
rect 176422 667258 183186 667494
rect 183422 667258 190186 667494
rect 190422 667258 197186 667494
rect 197422 667258 204186 667494
rect 204422 667258 211186 667494
rect 211422 667258 218186 667494
rect 218422 667258 225186 667494
rect 225422 667258 232186 667494
rect 232422 667258 239186 667494
rect 239422 667258 246186 667494
rect 246422 667258 253186 667494
rect 253422 667258 260186 667494
rect 260422 667258 267186 667494
rect 267422 667258 274186 667494
rect 274422 667258 281186 667494
rect 281422 667258 288186 667494
rect 288422 667258 295186 667494
rect 295422 667258 302186 667494
rect 302422 667258 309186 667494
rect 309422 667258 316186 667494
rect 316422 667258 323186 667494
rect 323422 667258 330186 667494
rect 330422 667258 337186 667494
rect 337422 667258 344186 667494
rect 344422 667258 351186 667494
rect 351422 667258 358186 667494
rect 358422 667258 365186 667494
rect 365422 667258 372186 667494
rect 372422 667258 379186 667494
rect 379422 667258 386186 667494
rect 386422 667258 393186 667494
rect 393422 667258 400186 667494
rect 400422 667258 407186 667494
rect 407422 667258 414186 667494
rect 414422 667258 421186 667494
rect 421422 667258 428186 667494
rect 428422 667258 435186 667494
rect 435422 667258 442186 667494
rect 442422 667258 449186 667494
rect 449422 667258 456186 667494
rect 456422 667258 463186 667494
rect 463422 667258 470186 667494
rect 470422 667258 477186 667494
rect 477422 667258 484186 667494
rect 484422 667258 491186 667494
rect 491422 667258 498186 667494
rect 498422 667258 505186 667494
rect 505422 667258 512186 667494
rect 512422 667258 519186 667494
rect 519422 667258 526186 667494
rect 526422 667258 533186 667494
rect 533422 667258 540186 667494
rect 540422 667258 547186 667494
rect 547422 667258 554186 667494
rect 554422 667258 561186 667494
rect 561422 667258 568186 667494
rect 568422 667258 575186 667494
rect 575422 667258 582186 667494
rect 582422 667258 585818 667494
rect 586054 667258 586138 667494
rect 586374 667258 586458 667494
rect 586694 667258 586778 667494
rect 587014 667258 588874 667494
rect -4950 667216 588874 667258
rect -4950 661434 588874 661476
rect -4950 661198 -4842 661434
rect -4606 661198 -4522 661434
rect -4286 661198 -4202 661434
rect -3966 661198 -3882 661434
rect -3646 661198 2918 661434
rect 3154 661198 9918 661434
rect 10154 661198 16918 661434
rect 17154 661198 23918 661434
rect 24154 661198 30918 661434
rect 31154 661198 37918 661434
rect 38154 661198 44918 661434
rect 45154 661198 51918 661434
rect 52154 661198 58918 661434
rect 59154 661198 65918 661434
rect 66154 661198 72918 661434
rect 73154 661198 79918 661434
rect 80154 661198 86918 661434
rect 87154 661198 93918 661434
rect 94154 661198 100918 661434
rect 101154 661198 107918 661434
rect 108154 661198 114918 661434
rect 115154 661198 121918 661434
rect 122154 661198 128918 661434
rect 129154 661198 135918 661434
rect 136154 661198 142918 661434
rect 143154 661198 149918 661434
rect 150154 661198 156918 661434
rect 157154 661198 163918 661434
rect 164154 661198 170918 661434
rect 171154 661198 177918 661434
rect 178154 661198 184918 661434
rect 185154 661198 191918 661434
rect 192154 661198 198918 661434
rect 199154 661198 205918 661434
rect 206154 661198 212918 661434
rect 213154 661198 219918 661434
rect 220154 661198 226918 661434
rect 227154 661198 233918 661434
rect 234154 661198 240918 661434
rect 241154 661198 247918 661434
rect 248154 661198 254918 661434
rect 255154 661198 261918 661434
rect 262154 661198 268918 661434
rect 269154 661198 275918 661434
rect 276154 661198 282918 661434
rect 283154 661198 289918 661434
rect 290154 661198 296918 661434
rect 297154 661198 303918 661434
rect 304154 661198 310918 661434
rect 311154 661198 317918 661434
rect 318154 661198 324918 661434
rect 325154 661198 331918 661434
rect 332154 661198 338918 661434
rect 339154 661198 345918 661434
rect 346154 661198 352918 661434
rect 353154 661198 359918 661434
rect 360154 661198 366918 661434
rect 367154 661198 373918 661434
rect 374154 661198 380918 661434
rect 381154 661198 387918 661434
rect 388154 661198 394918 661434
rect 395154 661198 401918 661434
rect 402154 661198 408918 661434
rect 409154 661198 415918 661434
rect 416154 661198 422918 661434
rect 423154 661198 429918 661434
rect 430154 661198 436918 661434
rect 437154 661198 443918 661434
rect 444154 661198 450918 661434
rect 451154 661198 457918 661434
rect 458154 661198 464918 661434
rect 465154 661198 471918 661434
rect 472154 661198 478918 661434
rect 479154 661198 485918 661434
rect 486154 661198 492918 661434
rect 493154 661198 499918 661434
rect 500154 661198 506918 661434
rect 507154 661198 513918 661434
rect 514154 661198 520918 661434
rect 521154 661198 527918 661434
rect 528154 661198 534918 661434
rect 535154 661198 541918 661434
rect 542154 661198 548918 661434
rect 549154 661198 555918 661434
rect 556154 661198 562918 661434
rect 563154 661198 569918 661434
rect 570154 661198 576918 661434
rect 577154 661198 587570 661434
rect 587806 661198 587890 661434
rect 588126 661198 588210 661434
rect 588446 661198 588530 661434
rect 588766 661198 588874 661434
rect -4950 661156 588874 661198
rect -4950 660494 588874 660536
rect -4950 660258 -3090 660494
rect -2854 660258 -2770 660494
rect -2534 660258 -2450 660494
rect -2214 660258 -2130 660494
rect -1894 660258 1186 660494
rect 1422 660258 8186 660494
rect 8422 660258 15186 660494
rect 15422 660258 22186 660494
rect 22422 660258 29186 660494
rect 29422 660258 36186 660494
rect 36422 660258 43186 660494
rect 43422 660258 50186 660494
rect 50422 660258 57186 660494
rect 57422 660258 64186 660494
rect 64422 660258 71186 660494
rect 71422 660258 78186 660494
rect 78422 660258 85186 660494
rect 85422 660258 92186 660494
rect 92422 660258 99186 660494
rect 99422 660258 106186 660494
rect 106422 660258 113186 660494
rect 113422 660258 120186 660494
rect 120422 660258 127186 660494
rect 127422 660258 134186 660494
rect 134422 660258 141186 660494
rect 141422 660258 148186 660494
rect 148422 660258 155186 660494
rect 155422 660258 162186 660494
rect 162422 660258 169186 660494
rect 169422 660258 176186 660494
rect 176422 660258 183186 660494
rect 183422 660258 190186 660494
rect 190422 660258 197186 660494
rect 197422 660258 204186 660494
rect 204422 660258 211186 660494
rect 211422 660258 218186 660494
rect 218422 660258 225186 660494
rect 225422 660258 232186 660494
rect 232422 660258 239186 660494
rect 239422 660258 246186 660494
rect 246422 660258 253186 660494
rect 253422 660258 260186 660494
rect 260422 660258 267186 660494
rect 267422 660258 274186 660494
rect 274422 660258 281186 660494
rect 281422 660258 288186 660494
rect 288422 660258 295186 660494
rect 295422 660258 302186 660494
rect 302422 660258 309186 660494
rect 309422 660258 316186 660494
rect 316422 660258 323186 660494
rect 323422 660258 330186 660494
rect 330422 660258 337186 660494
rect 337422 660258 344186 660494
rect 344422 660258 351186 660494
rect 351422 660258 358186 660494
rect 358422 660258 365186 660494
rect 365422 660258 372186 660494
rect 372422 660258 379186 660494
rect 379422 660258 386186 660494
rect 386422 660258 393186 660494
rect 393422 660258 400186 660494
rect 400422 660258 407186 660494
rect 407422 660258 414186 660494
rect 414422 660258 421186 660494
rect 421422 660258 428186 660494
rect 428422 660258 435186 660494
rect 435422 660258 442186 660494
rect 442422 660258 449186 660494
rect 449422 660258 456186 660494
rect 456422 660258 463186 660494
rect 463422 660258 470186 660494
rect 470422 660258 477186 660494
rect 477422 660258 484186 660494
rect 484422 660258 491186 660494
rect 491422 660258 498186 660494
rect 498422 660258 505186 660494
rect 505422 660258 512186 660494
rect 512422 660258 519186 660494
rect 519422 660258 526186 660494
rect 526422 660258 533186 660494
rect 533422 660258 540186 660494
rect 540422 660258 547186 660494
rect 547422 660258 554186 660494
rect 554422 660258 561186 660494
rect 561422 660258 568186 660494
rect 568422 660258 575186 660494
rect 575422 660258 582186 660494
rect 582422 660258 585818 660494
rect 586054 660258 586138 660494
rect 586374 660258 586458 660494
rect 586694 660258 586778 660494
rect 587014 660258 588874 660494
rect -4950 660216 588874 660258
rect -4950 654434 588874 654476
rect -4950 654198 -4842 654434
rect -4606 654198 -4522 654434
rect -4286 654198 -4202 654434
rect -3966 654198 -3882 654434
rect -3646 654198 2918 654434
rect 3154 654198 9918 654434
rect 10154 654198 16918 654434
rect 17154 654198 23918 654434
rect 24154 654198 30918 654434
rect 31154 654198 37918 654434
rect 38154 654198 44918 654434
rect 45154 654198 51918 654434
rect 52154 654198 58918 654434
rect 59154 654198 65918 654434
rect 66154 654198 72918 654434
rect 73154 654198 79918 654434
rect 80154 654198 86918 654434
rect 87154 654198 93918 654434
rect 94154 654198 100918 654434
rect 101154 654198 107918 654434
rect 108154 654198 114918 654434
rect 115154 654198 121918 654434
rect 122154 654198 128918 654434
rect 129154 654198 135918 654434
rect 136154 654198 142918 654434
rect 143154 654198 149918 654434
rect 150154 654198 156918 654434
rect 157154 654198 163918 654434
rect 164154 654198 170918 654434
rect 171154 654198 177918 654434
rect 178154 654198 184918 654434
rect 185154 654198 191918 654434
rect 192154 654198 198918 654434
rect 199154 654198 205918 654434
rect 206154 654198 212918 654434
rect 213154 654198 219918 654434
rect 220154 654198 226918 654434
rect 227154 654198 233918 654434
rect 234154 654198 240918 654434
rect 241154 654198 247918 654434
rect 248154 654198 254918 654434
rect 255154 654198 261918 654434
rect 262154 654198 268918 654434
rect 269154 654198 275918 654434
rect 276154 654198 282918 654434
rect 283154 654198 289918 654434
rect 290154 654198 296918 654434
rect 297154 654198 303918 654434
rect 304154 654198 310918 654434
rect 311154 654198 317918 654434
rect 318154 654198 324918 654434
rect 325154 654198 331918 654434
rect 332154 654198 338918 654434
rect 339154 654198 345918 654434
rect 346154 654198 352918 654434
rect 353154 654198 359918 654434
rect 360154 654198 366918 654434
rect 367154 654198 373918 654434
rect 374154 654198 380918 654434
rect 381154 654198 387918 654434
rect 388154 654198 394918 654434
rect 395154 654198 401918 654434
rect 402154 654198 408918 654434
rect 409154 654198 415918 654434
rect 416154 654198 422918 654434
rect 423154 654198 429918 654434
rect 430154 654198 436918 654434
rect 437154 654198 443918 654434
rect 444154 654198 450918 654434
rect 451154 654198 457918 654434
rect 458154 654198 464918 654434
rect 465154 654198 471918 654434
rect 472154 654198 478918 654434
rect 479154 654198 485918 654434
rect 486154 654198 492918 654434
rect 493154 654198 499918 654434
rect 500154 654198 506918 654434
rect 507154 654198 513918 654434
rect 514154 654198 520918 654434
rect 521154 654198 527918 654434
rect 528154 654198 534918 654434
rect 535154 654198 541918 654434
rect 542154 654198 548918 654434
rect 549154 654198 555918 654434
rect 556154 654198 562918 654434
rect 563154 654198 569918 654434
rect 570154 654198 576918 654434
rect 577154 654198 587570 654434
rect 587806 654198 587890 654434
rect 588126 654198 588210 654434
rect 588446 654198 588530 654434
rect 588766 654198 588874 654434
rect -4950 654156 588874 654198
rect -4950 653494 588874 653536
rect -4950 653258 -3090 653494
rect -2854 653258 -2770 653494
rect -2534 653258 -2450 653494
rect -2214 653258 -2130 653494
rect -1894 653258 1186 653494
rect 1422 653258 8186 653494
rect 8422 653258 15186 653494
rect 15422 653258 22186 653494
rect 22422 653258 29186 653494
rect 29422 653258 36186 653494
rect 36422 653258 43186 653494
rect 43422 653258 50186 653494
rect 50422 653258 57186 653494
rect 57422 653258 64186 653494
rect 64422 653258 71186 653494
rect 71422 653258 78186 653494
rect 78422 653258 85186 653494
rect 85422 653258 92186 653494
rect 92422 653258 99186 653494
rect 99422 653258 106186 653494
rect 106422 653258 113186 653494
rect 113422 653258 120186 653494
rect 120422 653258 127186 653494
rect 127422 653258 134186 653494
rect 134422 653258 141186 653494
rect 141422 653258 148186 653494
rect 148422 653258 155186 653494
rect 155422 653258 162186 653494
rect 162422 653258 169186 653494
rect 169422 653258 176186 653494
rect 176422 653258 183186 653494
rect 183422 653258 190186 653494
rect 190422 653258 197186 653494
rect 197422 653258 204186 653494
rect 204422 653258 211186 653494
rect 211422 653258 218186 653494
rect 218422 653258 225186 653494
rect 225422 653258 232186 653494
rect 232422 653258 239186 653494
rect 239422 653258 246186 653494
rect 246422 653258 253186 653494
rect 253422 653258 260186 653494
rect 260422 653258 267186 653494
rect 267422 653258 274186 653494
rect 274422 653258 281186 653494
rect 281422 653258 288186 653494
rect 288422 653258 295186 653494
rect 295422 653258 302186 653494
rect 302422 653258 309186 653494
rect 309422 653258 316186 653494
rect 316422 653258 323186 653494
rect 323422 653258 330186 653494
rect 330422 653258 337186 653494
rect 337422 653258 344186 653494
rect 344422 653258 351186 653494
rect 351422 653258 358186 653494
rect 358422 653258 365186 653494
rect 365422 653258 372186 653494
rect 372422 653258 379186 653494
rect 379422 653258 386186 653494
rect 386422 653258 393186 653494
rect 393422 653258 400186 653494
rect 400422 653258 407186 653494
rect 407422 653258 414186 653494
rect 414422 653258 421186 653494
rect 421422 653258 428186 653494
rect 428422 653258 435186 653494
rect 435422 653258 442186 653494
rect 442422 653258 449186 653494
rect 449422 653258 456186 653494
rect 456422 653258 463186 653494
rect 463422 653258 470186 653494
rect 470422 653258 477186 653494
rect 477422 653258 484186 653494
rect 484422 653258 491186 653494
rect 491422 653258 498186 653494
rect 498422 653258 505186 653494
rect 505422 653258 512186 653494
rect 512422 653258 519186 653494
rect 519422 653258 526186 653494
rect 526422 653258 533186 653494
rect 533422 653258 540186 653494
rect 540422 653258 547186 653494
rect 547422 653258 554186 653494
rect 554422 653258 561186 653494
rect 561422 653258 568186 653494
rect 568422 653258 575186 653494
rect 575422 653258 582186 653494
rect 582422 653258 585818 653494
rect 586054 653258 586138 653494
rect 586374 653258 586458 653494
rect 586694 653258 586778 653494
rect 587014 653258 588874 653494
rect -4950 653216 588874 653258
rect -4950 647434 588874 647476
rect -4950 647198 -4842 647434
rect -4606 647198 -4522 647434
rect -4286 647198 -4202 647434
rect -3966 647198 -3882 647434
rect -3646 647198 2918 647434
rect 3154 647198 9918 647434
rect 10154 647198 16918 647434
rect 17154 647198 23918 647434
rect 24154 647198 30918 647434
rect 31154 647198 37918 647434
rect 38154 647198 44918 647434
rect 45154 647198 51918 647434
rect 52154 647198 58918 647434
rect 59154 647198 65918 647434
rect 66154 647198 72918 647434
rect 73154 647198 79918 647434
rect 80154 647198 86918 647434
rect 87154 647198 93918 647434
rect 94154 647198 100918 647434
rect 101154 647198 107918 647434
rect 108154 647198 114918 647434
rect 115154 647198 121918 647434
rect 122154 647198 128918 647434
rect 129154 647198 135918 647434
rect 136154 647198 142918 647434
rect 143154 647198 149918 647434
rect 150154 647198 156918 647434
rect 157154 647198 163918 647434
rect 164154 647198 170918 647434
rect 171154 647198 177918 647434
rect 178154 647198 184918 647434
rect 185154 647198 191918 647434
rect 192154 647198 198918 647434
rect 199154 647198 205918 647434
rect 206154 647198 212918 647434
rect 213154 647198 219918 647434
rect 220154 647198 226918 647434
rect 227154 647198 233918 647434
rect 234154 647198 240918 647434
rect 241154 647198 247918 647434
rect 248154 647198 254918 647434
rect 255154 647198 261918 647434
rect 262154 647198 268918 647434
rect 269154 647198 275918 647434
rect 276154 647198 282918 647434
rect 283154 647198 289918 647434
rect 290154 647198 296918 647434
rect 297154 647198 303918 647434
rect 304154 647198 310918 647434
rect 311154 647198 317918 647434
rect 318154 647198 324918 647434
rect 325154 647198 331918 647434
rect 332154 647198 338918 647434
rect 339154 647198 345918 647434
rect 346154 647198 352918 647434
rect 353154 647198 359918 647434
rect 360154 647198 366918 647434
rect 367154 647198 373918 647434
rect 374154 647198 380918 647434
rect 381154 647198 387918 647434
rect 388154 647198 394918 647434
rect 395154 647198 401918 647434
rect 402154 647198 408918 647434
rect 409154 647198 415918 647434
rect 416154 647198 422918 647434
rect 423154 647198 429918 647434
rect 430154 647198 436918 647434
rect 437154 647198 443918 647434
rect 444154 647198 450918 647434
rect 451154 647198 457918 647434
rect 458154 647198 464918 647434
rect 465154 647198 471918 647434
rect 472154 647198 478918 647434
rect 479154 647198 485918 647434
rect 486154 647198 492918 647434
rect 493154 647198 499918 647434
rect 500154 647198 506918 647434
rect 507154 647198 513918 647434
rect 514154 647198 520918 647434
rect 521154 647198 527918 647434
rect 528154 647198 534918 647434
rect 535154 647198 541918 647434
rect 542154 647198 548918 647434
rect 549154 647198 555918 647434
rect 556154 647198 562918 647434
rect 563154 647198 569918 647434
rect 570154 647198 576918 647434
rect 577154 647198 587570 647434
rect 587806 647198 587890 647434
rect 588126 647198 588210 647434
rect 588446 647198 588530 647434
rect 588766 647198 588874 647434
rect -4950 647156 588874 647198
rect -4950 646494 588874 646536
rect -4950 646258 -3090 646494
rect -2854 646258 -2770 646494
rect -2534 646258 -2450 646494
rect -2214 646258 -2130 646494
rect -1894 646258 1186 646494
rect 1422 646258 8186 646494
rect 8422 646258 15186 646494
rect 15422 646258 22186 646494
rect 22422 646258 29186 646494
rect 29422 646258 36186 646494
rect 36422 646258 43186 646494
rect 43422 646258 50186 646494
rect 50422 646258 57186 646494
rect 57422 646258 64186 646494
rect 64422 646258 71186 646494
rect 71422 646258 78186 646494
rect 78422 646258 85186 646494
rect 85422 646258 92186 646494
rect 92422 646258 99186 646494
rect 99422 646258 106186 646494
rect 106422 646258 113186 646494
rect 113422 646258 120186 646494
rect 120422 646258 127186 646494
rect 127422 646258 134186 646494
rect 134422 646258 141186 646494
rect 141422 646258 148186 646494
rect 148422 646258 155186 646494
rect 155422 646258 162186 646494
rect 162422 646258 169186 646494
rect 169422 646258 176186 646494
rect 176422 646258 183186 646494
rect 183422 646258 190186 646494
rect 190422 646258 197186 646494
rect 197422 646258 204186 646494
rect 204422 646258 211186 646494
rect 211422 646258 218186 646494
rect 218422 646258 225186 646494
rect 225422 646258 232186 646494
rect 232422 646258 239186 646494
rect 239422 646258 246186 646494
rect 246422 646258 253186 646494
rect 253422 646258 260186 646494
rect 260422 646258 267186 646494
rect 267422 646258 274186 646494
rect 274422 646258 281186 646494
rect 281422 646258 288186 646494
rect 288422 646258 295186 646494
rect 295422 646258 302186 646494
rect 302422 646258 309186 646494
rect 309422 646258 316186 646494
rect 316422 646258 323186 646494
rect 323422 646258 330186 646494
rect 330422 646258 337186 646494
rect 337422 646258 344186 646494
rect 344422 646258 351186 646494
rect 351422 646258 358186 646494
rect 358422 646258 365186 646494
rect 365422 646258 372186 646494
rect 372422 646258 379186 646494
rect 379422 646258 386186 646494
rect 386422 646258 393186 646494
rect 393422 646258 400186 646494
rect 400422 646258 407186 646494
rect 407422 646258 414186 646494
rect 414422 646258 421186 646494
rect 421422 646258 428186 646494
rect 428422 646258 435186 646494
rect 435422 646258 442186 646494
rect 442422 646258 449186 646494
rect 449422 646258 456186 646494
rect 456422 646258 463186 646494
rect 463422 646258 470186 646494
rect 470422 646258 477186 646494
rect 477422 646258 484186 646494
rect 484422 646258 491186 646494
rect 491422 646258 498186 646494
rect 498422 646258 505186 646494
rect 505422 646258 512186 646494
rect 512422 646258 519186 646494
rect 519422 646258 526186 646494
rect 526422 646258 533186 646494
rect 533422 646258 540186 646494
rect 540422 646258 547186 646494
rect 547422 646258 554186 646494
rect 554422 646258 561186 646494
rect 561422 646258 568186 646494
rect 568422 646258 575186 646494
rect 575422 646258 582186 646494
rect 582422 646258 585818 646494
rect 586054 646258 586138 646494
rect 586374 646258 586458 646494
rect 586694 646258 586778 646494
rect 587014 646258 588874 646494
rect -4950 646216 588874 646258
rect -4950 640434 588874 640476
rect -4950 640198 -4842 640434
rect -4606 640198 -4522 640434
rect -4286 640198 -4202 640434
rect -3966 640198 -3882 640434
rect -3646 640198 2918 640434
rect 3154 640198 9918 640434
rect 10154 640198 16918 640434
rect 17154 640198 23918 640434
rect 24154 640198 30918 640434
rect 31154 640198 37918 640434
rect 38154 640198 44918 640434
rect 45154 640198 51918 640434
rect 52154 640198 58918 640434
rect 59154 640198 65918 640434
rect 66154 640198 72918 640434
rect 73154 640198 79918 640434
rect 80154 640198 86918 640434
rect 87154 640198 93918 640434
rect 94154 640198 100918 640434
rect 101154 640198 107918 640434
rect 108154 640198 114918 640434
rect 115154 640198 121918 640434
rect 122154 640198 128918 640434
rect 129154 640198 135918 640434
rect 136154 640198 142918 640434
rect 143154 640198 149918 640434
rect 150154 640198 156918 640434
rect 157154 640198 163918 640434
rect 164154 640198 170918 640434
rect 171154 640198 177918 640434
rect 178154 640198 184918 640434
rect 185154 640198 191918 640434
rect 192154 640198 198918 640434
rect 199154 640198 205918 640434
rect 206154 640198 212918 640434
rect 213154 640198 219918 640434
rect 220154 640198 226918 640434
rect 227154 640198 233918 640434
rect 234154 640198 240918 640434
rect 241154 640198 247918 640434
rect 248154 640198 254918 640434
rect 255154 640198 261918 640434
rect 262154 640198 268918 640434
rect 269154 640198 275918 640434
rect 276154 640198 282918 640434
rect 283154 640198 289918 640434
rect 290154 640198 296918 640434
rect 297154 640198 303918 640434
rect 304154 640198 310918 640434
rect 311154 640198 317918 640434
rect 318154 640198 324918 640434
rect 325154 640198 331918 640434
rect 332154 640198 338918 640434
rect 339154 640198 345918 640434
rect 346154 640198 352918 640434
rect 353154 640198 359918 640434
rect 360154 640198 366918 640434
rect 367154 640198 373918 640434
rect 374154 640198 380918 640434
rect 381154 640198 387918 640434
rect 388154 640198 394918 640434
rect 395154 640198 401918 640434
rect 402154 640198 408918 640434
rect 409154 640198 415918 640434
rect 416154 640198 422918 640434
rect 423154 640198 429918 640434
rect 430154 640198 436918 640434
rect 437154 640198 443918 640434
rect 444154 640198 450918 640434
rect 451154 640198 457918 640434
rect 458154 640198 464918 640434
rect 465154 640198 471918 640434
rect 472154 640198 478918 640434
rect 479154 640198 485918 640434
rect 486154 640198 492918 640434
rect 493154 640198 499918 640434
rect 500154 640198 506918 640434
rect 507154 640198 513918 640434
rect 514154 640198 520918 640434
rect 521154 640198 527918 640434
rect 528154 640198 534918 640434
rect 535154 640198 541918 640434
rect 542154 640198 548918 640434
rect 549154 640198 555918 640434
rect 556154 640198 562918 640434
rect 563154 640198 569918 640434
rect 570154 640198 576918 640434
rect 577154 640198 587570 640434
rect 587806 640198 587890 640434
rect 588126 640198 588210 640434
rect 588446 640198 588530 640434
rect 588766 640198 588874 640434
rect -4950 640156 588874 640198
rect -4950 639494 588874 639536
rect -4950 639258 -3090 639494
rect -2854 639258 -2770 639494
rect -2534 639258 -2450 639494
rect -2214 639258 -2130 639494
rect -1894 639258 1186 639494
rect 1422 639258 8186 639494
rect 8422 639258 15186 639494
rect 15422 639258 22186 639494
rect 22422 639258 29186 639494
rect 29422 639258 36186 639494
rect 36422 639258 43186 639494
rect 43422 639258 50186 639494
rect 50422 639258 57186 639494
rect 57422 639258 64186 639494
rect 64422 639258 71186 639494
rect 71422 639258 78186 639494
rect 78422 639258 85186 639494
rect 85422 639258 92186 639494
rect 92422 639258 99186 639494
rect 99422 639258 106186 639494
rect 106422 639258 113186 639494
rect 113422 639258 120186 639494
rect 120422 639258 127186 639494
rect 127422 639258 134186 639494
rect 134422 639258 141186 639494
rect 141422 639258 148186 639494
rect 148422 639258 155186 639494
rect 155422 639258 162186 639494
rect 162422 639258 169186 639494
rect 169422 639258 176186 639494
rect 176422 639258 183186 639494
rect 183422 639258 190186 639494
rect 190422 639258 197186 639494
rect 197422 639258 204186 639494
rect 204422 639258 211186 639494
rect 211422 639258 218186 639494
rect 218422 639258 225186 639494
rect 225422 639258 232186 639494
rect 232422 639258 239186 639494
rect 239422 639258 246186 639494
rect 246422 639258 253186 639494
rect 253422 639258 260186 639494
rect 260422 639258 267186 639494
rect 267422 639258 274186 639494
rect 274422 639258 281186 639494
rect 281422 639258 288186 639494
rect 288422 639258 295186 639494
rect 295422 639258 302186 639494
rect 302422 639258 309186 639494
rect 309422 639258 316186 639494
rect 316422 639258 323186 639494
rect 323422 639258 330186 639494
rect 330422 639258 337186 639494
rect 337422 639258 344186 639494
rect 344422 639258 351186 639494
rect 351422 639258 358186 639494
rect 358422 639258 365186 639494
rect 365422 639258 372186 639494
rect 372422 639258 379186 639494
rect 379422 639258 386186 639494
rect 386422 639258 393186 639494
rect 393422 639258 400186 639494
rect 400422 639258 407186 639494
rect 407422 639258 414186 639494
rect 414422 639258 421186 639494
rect 421422 639258 428186 639494
rect 428422 639258 435186 639494
rect 435422 639258 442186 639494
rect 442422 639258 449186 639494
rect 449422 639258 456186 639494
rect 456422 639258 463186 639494
rect 463422 639258 470186 639494
rect 470422 639258 477186 639494
rect 477422 639258 484186 639494
rect 484422 639258 491186 639494
rect 491422 639258 498186 639494
rect 498422 639258 505186 639494
rect 505422 639258 512186 639494
rect 512422 639258 519186 639494
rect 519422 639258 526186 639494
rect 526422 639258 533186 639494
rect 533422 639258 540186 639494
rect 540422 639258 547186 639494
rect 547422 639258 554186 639494
rect 554422 639258 561186 639494
rect 561422 639258 568186 639494
rect 568422 639258 575186 639494
rect 575422 639258 582186 639494
rect 582422 639258 585818 639494
rect 586054 639258 586138 639494
rect 586374 639258 586458 639494
rect 586694 639258 586778 639494
rect 587014 639258 588874 639494
rect -4950 639216 588874 639258
rect -4950 633434 588874 633476
rect -4950 633198 -4842 633434
rect -4606 633198 -4522 633434
rect -4286 633198 -4202 633434
rect -3966 633198 -3882 633434
rect -3646 633198 2918 633434
rect 3154 633198 9918 633434
rect 10154 633198 16918 633434
rect 17154 633198 23918 633434
rect 24154 633198 30918 633434
rect 31154 633198 37918 633434
rect 38154 633198 44918 633434
rect 45154 633198 51918 633434
rect 52154 633198 58918 633434
rect 59154 633198 65918 633434
rect 66154 633198 72918 633434
rect 73154 633198 79918 633434
rect 80154 633198 86918 633434
rect 87154 633198 93918 633434
rect 94154 633198 100918 633434
rect 101154 633198 107918 633434
rect 108154 633198 114918 633434
rect 115154 633198 121918 633434
rect 122154 633198 128918 633434
rect 129154 633198 135918 633434
rect 136154 633198 142918 633434
rect 143154 633198 149918 633434
rect 150154 633198 156918 633434
rect 157154 633198 163918 633434
rect 164154 633198 170918 633434
rect 171154 633198 177918 633434
rect 178154 633198 184918 633434
rect 185154 633198 191918 633434
rect 192154 633198 198918 633434
rect 199154 633198 205918 633434
rect 206154 633198 212918 633434
rect 213154 633198 219918 633434
rect 220154 633198 226918 633434
rect 227154 633198 233918 633434
rect 234154 633198 240918 633434
rect 241154 633198 247918 633434
rect 248154 633198 254918 633434
rect 255154 633198 261918 633434
rect 262154 633198 268918 633434
rect 269154 633198 275918 633434
rect 276154 633198 282918 633434
rect 283154 633198 289918 633434
rect 290154 633198 296918 633434
rect 297154 633198 303918 633434
rect 304154 633198 310918 633434
rect 311154 633198 317918 633434
rect 318154 633198 324918 633434
rect 325154 633198 331918 633434
rect 332154 633198 338918 633434
rect 339154 633198 345918 633434
rect 346154 633198 352918 633434
rect 353154 633198 359918 633434
rect 360154 633198 366918 633434
rect 367154 633198 373918 633434
rect 374154 633198 380918 633434
rect 381154 633198 387918 633434
rect 388154 633198 394918 633434
rect 395154 633198 401918 633434
rect 402154 633198 408918 633434
rect 409154 633198 415918 633434
rect 416154 633198 422918 633434
rect 423154 633198 429918 633434
rect 430154 633198 436918 633434
rect 437154 633198 443918 633434
rect 444154 633198 450918 633434
rect 451154 633198 457918 633434
rect 458154 633198 464918 633434
rect 465154 633198 471918 633434
rect 472154 633198 478918 633434
rect 479154 633198 485918 633434
rect 486154 633198 492918 633434
rect 493154 633198 499918 633434
rect 500154 633198 506918 633434
rect 507154 633198 513918 633434
rect 514154 633198 520918 633434
rect 521154 633198 527918 633434
rect 528154 633198 534918 633434
rect 535154 633198 541918 633434
rect 542154 633198 548918 633434
rect 549154 633198 555918 633434
rect 556154 633198 562918 633434
rect 563154 633198 569918 633434
rect 570154 633198 576918 633434
rect 577154 633198 587570 633434
rect 587806 633198 587890 633434
rect 588126 633198 588210 633434
rect 588446 633198 588530 633434
rect 588766 633198 588874 633434
rect -4950 633156 588874 633198
rect -4950 632494 588874 632536
rect -4950 632258 -3090 632494
rect -2854 632258 -2770 632494
rect -2534 632258 -2450 632494
rect -2214 632258 -2130 632494
rect -1894 632258 1186 632494
rect 1422 632258 8186 632494
rect 8422 632258 15186 632494
rect 15422 632258 22186 632494
rect 22422 632258 29186 632494
rect 29422 632258 36186 632494
rect 36422 632258 43186 632494
rect 43422 632258 50186 632494
rect 50422 632258 57186 632494
rect 57422 632258 64186 632494
rect 64422 632258 71186 632494
rect 71422 632258 78186 632494
rect 78422 632258 85186 632494
rect 85422 632258 92186 632494
rect 92422 632258 99186 632494
rect 99422 632258 106186 632494
rect 106422 632258 113186 632494
rect 113422 632258 120186 632494
rect 120422 632258 127186 632494
rect 127422 632258 134186 632494
rect 134422 632258 141186 632494
rect 141422 632258 148186 632494
rect 148422 632258 155186 632494
rect 155422 632258 162186 632494
rect 162422 632258 169186 632494
rect 169422 632258 176186 632494
rect 176422 632258 183186 632494
rect 183422 632258 190186 632494
rect 190422 632258 197186 632494
rect 197422 632258 204186 632494
rect 204422 632258 211186 632494
rect 211422 632258 218186 632494
rect 218422 632258 225186 632494
rect 225422 632258 232186 632494
rect 232422 632258 239186 632494
rect 239422 632258 246186 632494
rect 246422 632258 253186 632494
rect 253422 632258 260186 632494
rect 260422 632258 267186 632494
rect 267422 632258 274186 632494
rect 274422 632258 281186 632494
rect 281422 632258 288186 632494
rect 288422 632258 295186 632494
rect 295422 632258 302186 632494
rect 302422 632258 309186 632494
rect 309422 632258 316186 632494
rect 316422 632258 323186 632494
rect 323422 632258 330186 632494
rect 330422 632258 337186 632494
rect 337422 632258 344186 632494
rect 344422 632258 351186 632494
rect 351422 632258 358186 632494
rect 358422 632258 365186 632494
rect 365422 632258 372186 632494
rect 372422 632258 379186 632494
rect 379422 632258 386186 632494
rect 386422 632258 393186 632494
rect 393422 632258 400186 632494
rect 400422 632258 407186 632494
rect 407422 632258 414186 632494
rect 414422 632258 421186 632494
rect 421422 632258 428186 632494
rect 428422 632258 435186 632494
rect 435422 632258 442186 632494
rect 442422 632258 449186 632494
rect 449422 632258 456186 632494
rect 456422 632258 463186 632494
rect 463422 632258 470186 632494
rect 470422 632258 477186 632494
rect 477422 632258 484186 632494
rect 484422 632258 491186 632494
rect 491422 632258 498186 632494
rect 498422 632258 505186 632494
rect 505422 632258 512186 632494
rect 512422 632258 519186 632494
rect 519422 632258 526186 632494
rect 526422 632258 533186 632494
rect 533422 632258 540186 632494
rect 540422 632258 547186 632494
rect 547422 632258 554186 632494
rect 554422 632258 561186 632494
rect 561422 632258 568186 632494
rect 568422 632258 575186 632494
rect 575422 632258 582186 632494
rect 582422 632258 585818 632494
rect 586054 632258 586138 632494
rect 586374 632258 586458 632494
rect 586694 632258 586778 632494
rect 587014 632258 588874 632494
rect -4950 632216 588874 632258
rect -4950 626434 588874 626476
rect -4950 626198 -4842 626434
rect -4606 626198 -4522 626434
rect -4286 626198 -4202 626434
rect -3966 626198 -3882 626434
rect -3646 626198 2918 626434
rect 3154 626198 9918 626434
rect 10154 626198 16918 626434
rect 17154 626198 23918 626434
rect 24154 626198 30918 626434
rect 31154 626198 37918 626434
rect 38154 626198 44918 626434
rect 45154 626198 51918 626434
rect 52154 626198 58918 626434
rect 59154 626198 65918 626434
rect 66154 626198 72918 626434
rect 73154 626198 79918 626434
rect 80154 626198 86918 626434
rect 87154 626198 93918 626434
rect 94154 626198 100918 626434
rect 101154 626198 107918 626434
rect 108154 626198 114918 626434
rect 115154 626198 121918 626434
rect 122154 626198 128918 626434
rect 129154 626198 135918 626434
rect 136154 626198 142918 626434
rect 143154 626198 149918 626434
rect 150154 626198 156918 626434
rect 157154 626198 163918 626434
rect 164154 626198 170918 626434
rect 171154 626198 177918 626434
rect 178154 626198 184918 626434
rect 185154 626198 191918 626434
rect 192154 626198 198918 626434
rect 199154 626198 205918 626434
rect 206154 626198 212918 626434
rect 213154 626198 219918 626434
rect 220154 626198 226918 626434
rect 227154 626198 233918 626434
rect 234154 626198 240918 626434
rect 241154 626198 247918 626434
rect 248154 626198 254918 626434
rect 255154 626198 261918 626434
rect 262154 626198 268918 626434
rect 269154 626198 275918 626434
rect 276154 626198 282918 626434
rect 283154 626198 289918 626434
rect 290154 626198 296918 626434
rect 297154 626198 303918 626434
rect 304154 626198 310918 626434
rect 311154 626198 317918 626434
rect 318154 626198 324918 626434
rect 325154 626198 331918 626434
rect 332154 626198 338918 626434
rect 339154 626198 345918 626434
rect 346154 626198 352918 626434
rect 353154 626198 359918 626434
rect 360154 626198 366918 626434
rect 367154 626198 373918 626434
rect 374154 626198 380918 626434
rect 381154 626198 387918 626434
rect 388154 626198 394918 626434
rect 395154 626198 401918 626434
rect 402154 626198 408918 626434
rect 409154 626198 415918 626434
rect 416154 626198 422918 626434
rect 423154 626198 429918 626434
rect 430154 626198 436918 626434
rect 437154 626198 443918 626434
rect 444154 626198 450918 626434
rect 451154 626198 457918 626434
rect 458154 626198 464918 626434
rect 465154 626198 471918 626434
rect 472154 626198 478918 626434
rect 479154 626198 485918 626434
rect 486154 626198 492918 626434
rect 493154 626198 499918 626434
rect 500154 626198 506918 626434
rect 507154 626198 513918 626434
rect 514154 626198 520918 626434
rect 521154 626198 527918 626434
rect 528154 626198 534918 626434
rect 535154 626198 541918 626434
rect 542154 626198 548918 626434
rect 549154 626198 555918 626434
rect 556154 626198 562918 626434
rect 563154 626198 569918 626434
rect 570154 626198 576918 626434
rect 577154 626198 587570 626434
rect 587806 626198 587890 626434
rect 588126 626198 588210 626434
rect 588446 626198 588530 626434
rect 588766 626198 588874 626434
rect -4950 626156 588874 626198
rect -4950 625494 588874 625536
rect -4950 625258 -3090 625494
rect -2854 625258 -2770 625494
rect -2534 625258 -2450 625494
rect -2214 625258 -2130 625494
rect -1894 625258 1186 625494
rect 1422 625258 8186 625494
rect 8422 625258 15186 625494
rect 15422 625258 22186 625494
rect 22422 625258 29186 625494
rect 29422 625258 36186 625494
rect 36422 625258 43186 625494
rect 43422 625258 50186 625494
rect 50422 625258 57186 625494
rect 57422 625258 64186 625494
rect 64422 625258 71186 625494
rect 71422 625258 78186 625494
rect 78422 625258 85186 625494
rect 85422 625258 92186 625494
rect 92422 625258 99186 625494
rect 99422 625258 106186 625494
rect 106422 625258 113186 625494
rect 113422 625258 120186 625494
rect 120422 625258 127186 625494
rect 127422 625258 134186 625494
rect 134422 625258 141186 625494
rect 141422 625258 148186 625494
rect 148422 625258 155186 625494
rect 155422 625258 162186 625494
rect 162422 625258 169186 625494
rect 169422 625258 176186 625494
rect 176422 625258 183186 625494
rect 183422 625258 190186 625494
rect 190422 625258 197186 625494
rect 197422 625258 204186 625494
rect 204422 625258 211186 625494
rect 211422 625258 218186 625494
rect 218422 625258 225186 625494
rect 225422 625258 232186 625494
rect 232422 625258 239186 625494
rect 239422 625258 246186 625494
rect 246422 625258 253186 625494
rect 253422 625258 260186 625494
rect 260422 625258 267186 625494
rect 267422 625258 274186 625494
rect 274422 625258 281186 625494
rect 281422 625258 288186 625494
rect 288422 625258 295186 625494
rect 295422 625258 302186 625494
rect 302422 625258 309186 625494
rect 309422 625258 316186 625494
rect 316422 625258 323186 625494
rect 323422 625258 330186 625494
rect 330422 625258 337186 625494
rect 337422 625258 344186 625494
rect 344422 625258 351186 625494
rect 351422 625258 358186 625494
rect 358422 625258 365186 625494
rect 365422 625258 372186 625494
rect 372422 625258 379186 625494
rect 379422 625258 386186 625494
rect 386422 625258 393186 625494
rect 393422 625258 400186 625494
rect 400422 625258 407186 625494
rect 407422 625258 414186 625494
rect 414422 625258 421186 625494
rect 421422 625258 428186 625494
rect 428422 625258 435186 625494
rect 435422 625258 442186 625494
rect 442422 625258 449186 625494
rect 449422 625258 456186 625494
rect 456422 625258 463186 625494
rect 463422 625258 470186 625494
rect 470422 625258 477186 625494
rect 477422 625258 484186 625494
rect 484422 625258 491186 625494
rect 491422 625258 498186 625494
rect 498422 625258 505186 625494
rect 505422 625258 512186 625494
rect 512422 625258 519186 625494
rect 519422 625258 526186 625494
rect 526422 625258 533186 625494
rect 533422 625258 540186 625494
rect 540422 625258 547186 625494
rect 547422 625258 554186 625494
rect 554422 625258 561186 625494
rect 561422 625258 568186 625494
rect 568422 625258 575186 625494
rect 575422 625258 582186 625494
rect 582422 625258 585818 625494
rect 586054 625258 586138 625494
rect 586374 625258 586458 625494
rect 586694 625258 586778 625494
rect 587014 625258 588874 625494
rect -4950 625216 588874 625258
rect -4950 619434 588874 619476
rect -4950 619198 -4842 619434
rect -4606 619198 -4522 619434
rect -4286 619198 -4202 619434
rect -3966 619198 -3882 619434
rect -3646 619198 2918 619434
rect 3154 619198 9918 619434
rect 10154 619198 16918 619434
rect 17154 619198 23918 619434
rect 24154 619198 30918 619434
rect 31154 619198 37918 619434
rect 38154 619198 44918 619434
rect 45154 619198 51918 619434
rect 52154 619198 58918 619434
rect 59154 619198 65918 619434
rect 66154 619198 72918 619434
rect 73154 619198 79918 619434
rect 80154 619198 86918 619434
rect 87154 619198 93918 619434
rect 94154 619198 100918 619434
rect 101154 619198 107918 619434
rect 108154 619198 114918 619434
rect 115154 619198 121918 619434
rect 122154 619198 128918 619434
rect 129154 619198 135918 619434
rect 136154 619198 142918 619434
rect 143154 619198 149918 619434
rect 150154 619198 156918 619434
rect 157154 619198 163918 619434
rect 164154 619198 170918 619434
rect 171154 619198 177918 619434
rect 178154 619198 184918 619434
rect 185154 619198 191918 619434
rect 192154 619198 198918 619434
rect 199154 619198 205918 619434
rect 206154 619198 212918 619434
rect 213154 619198 219918 619434
rect 220154 619198 226918 619434
rect 227154 619198 233918 619434
rect 234154 619198 240918 619434
rect 241154 619198 247918 619434
rect 248154 619198 254918 619434
rect 255154 619198 261918 619434
rect 262154 619198 268918 619434
rect 269154 619198 275918 619434
rect 276154 619198 282918 619434
rect 283154 619198 289918 619434
rect 290154 619198 296918 619434
rect 297154 619198 303918 619434
rect 304154 619198 310918 619434
rect 311154 619198 317918 619434
rect 318154 619198 324918 619434
rect 325154 619198 331918 619434
rect 332154 619198 338918 619434
rect 339154 619198 345918 619434
rect 346154 619198 352918 619434
rect 353154 619198 359918 619434
rect 360154 619198 366918 619434
rect 367154 619198 373918 619434
rect 374154 619198 380918 619434
rect 381154 619198 387918 619434
rect 388154 619198 394918 619434
rect 395154 619198 401918 619434
rect 402154 619198 408918 619434
rect 409154 619198 415918 619434
rect 416154 619198 422918 619434
rect 423154 619198 429918 619434
rect 430154 619198 436918 619434
rect 437154 619198 443918 619434
rect 444154 619198 450918 619434
rect 451154 619198 457918 619434
rect 458154 619198 464918 619434
rect 465154 619198 471918 619434
rect 472154 619198 478918 619434
rect 479154 619198 485918 619434
rect 486154 619198 492918 619434
rect 493154 619198 499918 619434
rect 500154 619198 506918 619434
rect 507154 619198 513918 619434
rect 514154 619198 520918 619434
rect 521154 619198 527918 619434
rect 528154 619198 534918 619434
rect 535154 619198 541918 619434
rect 542154 619198 548918 619434
rect 549154 619198 555918 619434
rect 556154 619198 562918 619434
rect 563154 619198 569918 619434
rect 570154 619198 576918 619434
rect 577154 619198 587570 619434
rect 587806 619198 587890 619434
rect 588126 619198 588210 619434
rect 588446 619198 588530 619434
rect 588766 619198 588874 619434
rect -4950 619156 588874 619198
rect -4950 618494 588874 618536
rect -4950 618258 -3090 618494
rect -2854 618258 -2770 618494
rect -2534 618258 -2450 618494
rect -2214 618258 -2130 618494
rect -1894 618258 1186 618494
rect 1422 618258 8186 618494
rect 8422 618258 15186 618494
rect 15422 618258 22186 618494
rect 22422 618258 29186 618494
rect 29422 618258 36186 618494
rect 36422 618258 43186 618494
rect 43422 618258 50186 618494
rect 50422 618258 57186 618494
rect 57422 618258 64186 618494
rect 64422 618258 71186 618494
rect 71422 618258 78186 618494
rect 78422 618258 85186 618494
rect 85422 618258 92186 618494
rect 92422 618258 99186 618494
rect 99422 618258 106186 618494
rect 106422 618258 113186 618494
rect 113422 618258 120186 618494
rect 120422 618258 127186 618494
rect 127422 618258 134186 618494
rect 134422 618258 141186 618494
rect 141422 618258 148186 618494
rect 148422 618258 155186 618494
rect 155422 618258 162186 618494
rect 162422 618258 169186 618494
rect 169422 618258 176186 618494
rect 176422 618258 183186 618494
rect 183422 618258 190186 618494
rect 190422 618258 197186 618494
rect 197422 618258 204186 618494
rect 204422 618258 211186 618494
rect 211422 618258 218186 618494
rect 218422 618258 225186 618494
rect 225422 618258 232186 618494
rect 232422 618258 239186 618494
rect 239422 618258 246186 618494
rect 246422 618258 253186 618494
rect 253422 618258 260186 618494
rect 260422 618258 267186 618494
rect 267422 618258 274186 618494
rect 274422 618258 281186 618494
rect 281422 618258 288186 618494
rect 288422 618258 295186 618494
rect 295422 618258 302186 618494
rect 302422 618258 309186 618494
rect 309422 618258 316186 618494
rect 316422 618258 323186 618494
rect 323422 618258 330186 618494
rect 330422 618258 337186 618494
rect 337422 618258 344186 618494
rect 344422 618258 351186 618494
rect 351422 618258 358186 618494
rect 358422 618258 365186 618494
rect 365422 618258 372186 618494
rect 372422 618258 379186 618494
rect 379422 618258 386186 618494
rect 386422 618258 393186 618494
rect 393422 618258 400186 618494
rect 400422 618258 407186 618494
rect 407422 618258 414186 618494
rect 414422 618258 421186 618494
rect 421422 618258 428186 618494
rect 428422 618258 435186 618494
rect 435422 618258 442186 618494
rect 442422 618258 449186 618494
rect 449422 618258 456186 618494
rect 456422 618258 463186 618494
rect 463422 618258 470186 618494
rect 470422 618258 477186 618494
rect 477422 618258 484186 618494
rect 484422 618258 491186 618494
rect 491422 618258 498186 618494
rect 498422 618258 505186 618494
rect 505422 618258 512186 618494
rect 512422 618258 519186 618494
rect 519422 618258 526186 618494
rect 526422 618258 533186 618494
rect 533422 618258 540186 618494
rect 540422 618258 547186 618494
rect 547422 618258 554186 618494
rect 554422 618258 561186 618494
rect 561422 618258 568186 618494
rect 568422 618258 575186 618494
rect 575422 618258 582186 618494
rect 582422 618258 585818 618494
rect 586054 618258 586138 618494
rect 586374 618258 586458 618494
rect 586694 618258 586778 618494
rect 587014 618258 588874 618494
rect -4950 618216 588874 618258
rect -4950 612434 588874 612476
rect -4950 612198 -4842 612434
rect -4606 612198 -4522 612434
rect -4286 612198 -4202 612434
rect -3966 612198 -3882 612434
rect -3646 612198 2918 612434
rect 3154 612198 9918 612434
rect 10154 612198 16918 612434
rect 17154 612198 23918 612434
rect 24154 612198 30918 612434
rect 31154 612198 37918 612434
rect 38154 612198 44918 612434
rect 45154 612198 51918 612434
rect 52154 612198 58918 612434
rect 59154 612198 65918 612434
rect 66154 612198 72918 612434
rect 73154 612198 79918 612434
rect 80154 612198 86918 612434
rect 87154 612198 93918 612434
rect 94154 612198 100918 612434
rect 101154 612198 107918 612434
rect 108154 612198 114918 612434
rect 115154 612198 121918 612434
rect 122154 612198 128918 612434
rect 129154 612198 135918 612434
rect 136154 612198 142918 612434
rect 143154 612198 149918 612434
rect 150154 612198 156918 612434
rect 157154 612198 163918 612434
rect 164154 612198 170918 612434
rect 171154 612198 177918 612434
rect 178154 612198 184918 612434
rect 185154 612198 191918 612434
rect 192154 612198 198918 612434
rect 199154 612198 205918 612434
rect 206154 612198 212918 612434
rect 213154 612198 219918 612434
rect 220154 612198 226918 612434
rect 227154 612198 233918 612434
rect 234154 612198 240918 612434
rect 241154 612198 247918 612434
rect 248154 612198 254918 612434
rect 255154 612198 261918 612434
rect 262154 612198 268918 612434
rect 269154 612198 275918 612434
rect 276154 612198 282918 612434
rect 283154 612198 289918 612434
rect 290154 612198 296918 612434
rect 297154 612198 303918 612434
rect 304154 612198 310918 612434
rect 311154 612198 317918 612434
rect 318154 612198 324918 612434
rect 325154 612198 331918 612434
rect 332154 612198 338918 612434
rect 339154 612198 345918 612434
rect 346154 612198 352918 612434
rect 353154 612198 359918 612434
rect 360154 612198 366918 612434
rect 367154 612198 373918 612434
rect 374154 612198 380918 612434
rect 381154 612198 387918 612434
rect 388154 612198 394918 612434
rect 395154 612198 401918 612434
rect 402154 612198 408918 612434
rect 409154 612198 415918 612434
rect 416154 612198 422918 612434
rect 423154 612198 429918 612434
rect 430154 612198 436918 612434
rect 437154 612198 443918 612434
rect 444154 612198 450918 612434
rect 451154 612198 457918 612434
rect 458154 612198 464918 612434
rect 465154 612198 471918 612434
rect 472154 612198 478918 612434
rect 479154 612198 485918 612434
rect 486154 612198 492918 612434
rect 493154 612198 499918 612434
rect 500154 612198 506918 612434
rect 507154 612198 513918 612434
rect 514154 612198 520918 612434
rect 521154 612198 527918 612434
rect 528154 612198 534918 612434
rect 535154 612198 541918 612434
rect 542154 612198 548918 612434
rect 549154 612198 555918 612434
rect 556154 612198 562918 612434
rect 563154 612198 569918 612434
rect 570154 612198 576918 612434
rect 577154 612198 587570 612434
rect 587806 612198 587890 612434
rect 588126 612198 588210 612434
rect 588446 612198 588530 612434
rect 588766 612198 588874 612434
rect -4950 612156 588874 612198
rect -4950 611494 588874 611536
rect -4950 611258 -3090 611494
rect -2854 611258 -2770 611494
rect -2534 611258 -2450 611494
rect -2214 611258 -2130 611494
rect -1894 611258 1186 611494
rect 1422 611258 8186 611494
rect 8422 611258 15186 611494
rect 15422 611258 22186 611494
rect 22422 611258 29186 611494
rect 29422 611258 36186 611494
rect 36422 611258 43186 611494
rect 43422 611258 50186 611494
rect 50422 611258 57186 611494
rect 57422 611258 64186 611494
rect 64422 611258 71186 611494
rect 71422 611258 78186 611494
rect 78422 611258 85186 611494
rect 85422 611258 92186 611494
rect 92422 611258 99186 611494
rect 99422 611258 106186 611494
rect 106422 611258 113186 611494
rect 113422 611258 120186 611494
rect 120422 611258 127186 611494
rect 127422 611258 134186 611494
rect 134422 611258 141186 611494
rect 141422 611258 148186 611494
rect 148422 611258 155186 611494
rect 155422 611258 162186 611494
rect 162422 611258 169186 611494
rect 169422 611258 176186 611494
rect 176422 611258 183186 611494
rect 183422 611258 190186 611494
rect 190422 611258 197186 611494
rect 197422 611258 204186 611494
rect 204422 611258 211186 611494
rect 211422 611258 218186 611494
rect 218422 611258 225186 611494
rect 225422 611258 232186 611494
rect 232422 611258 239186 611494
rect 239422 611258 246186 611494
rect 246422 611258 253186 611494
rect 253422 611258 260186 611494
rect 260422 611258 267186 611494
rect 267422 611258 274186 611494
rect 274422 611258 281186 611494
rect 281422 611258 288186 611494
rect 288422 611258 295186 611494
rect 295422 611258 302186 611494
rect 302422 611258 309186 611494
rect 309422 611258 316186 611494
rect 316422 611258 323186 611494
rect 323422 611258 330186 611494
rect 330422 611258 337186 611494
rect 337422 611258 344186 611494
rect 344422 611258 351186 611494
rect 351422 611258 358186 611494
rect 358422 611258 365186 611494
rect 365422 611258 372186 611494
rect 372422 611258 379186 611494
rect 379422 611258 386186 611494
rect 386422 611258 393186 611494
rect 393422 611258 400186 611494
rect 400422 611258 407186 611494
rect 407422 611258 414186 611494
rect 414422 611258 421186 611494
rect 421422 611258 428186 611494
rect 428422 611258 435186 611494
rect 435422 611258 442186 611494
rect 442422 611258 449186 611494
rect 449422 611258 456186 611494
rect 456422 611258 463186 611494
rect 463422 611258 470186 611494
rect 470422 611258 477186 611494
rect 477422 611258 484186 611494
rect 484422 611258 491186 611494
rect 491422 611258 498186 611494
rect 498422 611258 505186 611494
rect 505422 611258 512186 611494
rect 512422 611258 519186 611494
rect 519422 611258 526186 611494
rect 526422 611258 533186 611494
rect 533422 611258 540186 611494
rect 540422 611258 547186 611494
rect 547422 611258 554186 611494
rect 554422 611258 561186 611494
rect 561422 611258 568186 611494
rect 568422 611258 575186 611494
rect 575422 611258 582186 611494
rect 582422 611258 585818 611494
rect 586054 611258 586138 611494
rect 586374 611258 586458 611494
rect 586694 611258 586778 611494
rect 587014 611258 588874 611494
rect -4950 611216 588874 611258
rect -4950 605434 588874 605476
rect -4950 605198 -4842 605434
rect -4606 605198 -4522 605434
rect -4286 605198 -4202 605434
rect -3966 605198 -3882 605434
rect -3646 605198 2918 605434
rect 3154 605198 9918 605434
rect 10154 605198 16918 605434
rect 17154 605198 23918 605434
rect 24154 605198 30918 605434
rect 31154 605198 37918 605434
rect 38154 605198 44918 605434
rect 45154 605198 51918 605434
rect 52154 605198 58918 605434
rect 59154 605198 65918 605434
rect 66154 605198 72918 605434
rect 73154 605198 79918 605434
rect 80154 605198 86918 605434
rect 87154 605198 93918 605434
rect 94154 605198 100918 605434
rect 101154 605198 107918 605434
rect 108154 605198 114918 605434
rect 115154 605198 121918 605434
rect 122154 605198 128918 605434
rect 129154 605198 135918 605434
rect 136154 605198 142918 605434
rect 143154 605198 149918 605434
rect 150154 605198 156918 605434
rect 157154 605198 163918 605434
rect 164154 605198 170918 605434
rect 171154 605198 177918 605434
rect 178154 605198 184918 605434
rect 185154 605198 191918 605434
rect 192154 605198 198918 605434
rect 199154 605198 205918 605434
rect 206154 605198 212918 605434
rect 213154 605198 219918 605434
rect 220154 605198 226918 605434
rect 227154 605198 233918 605434
rect 234154 605198 240918 605434
rect 241154 605198 247918 605434
rect 248154 605198 254918 605434
rect 255154 605198 261918 605434
rect 262154 605198 268918 605434
rect 269154 605198 275918 605434
rect 276154 605198 282918 605434
rect 283154 605198 289918 605434
rect 290154 605198 296918 605434
rect 297154 605198 303918 605434
rect 304154 605198 310918 605434
rect 311154 605198 317918 605434
rect 318154 605198 324918 605434
rect 325154 605198 331918 605434
rect 332154 605198 338918 605434
rect 339154 605198 345918 605434
rect 346154 605198 352918 605434
rect 353154 605198 359918 605434
rect 360154 605198 366918 605434
rect 367154 605198 373918 605434
rect 374154 605198 380918 605434
rect 381154 605198 387918 605434
rect 388154 605198 394918 605434
rect 395154 605198 401918 605434
rect 402154 605198 408918 605434
rect 409154 605198 415918 605434
rect 416154 605198 422918 605434
rect 423154 605198 429918 605434
rect 430154 605198 436918 605434
rect 437154 605198 443918 605434
rect 444154 605198 450918 605434
rect 451154 605198 457918 605434
rect 458154 605198 464918 605434
rect 465154 605198 471918 605434
rect 472154 605198 478918 605434
rect 479154 605198 485918 605434
rect 486154 605198 492918 605434
rect 493154 605198 499918 605434
rect 500154 605198 506918 605434
rect 507154 605198 513918 605434
rect 514154 605198 520918 605434
rect 521154 605198 527918 605434
rect 528154 605198 534918 605434
rect 535154 605198 541918 605434
rect 542154 605198 548918 605434
rect 549154 605198 555918 605434
rect 556154 605198 562918 605434
rect 563154 605198 569918 605434
rect 570154 605198 576918 605434
rect 577154 605198 587570 605434
rect 587806 605198 587890 605434
rect 588126 605198 588210 605434
rect 588446 605198 588530 605434
rect 588766 605198 588874 605434
rect -4950 605156 588874 605198
rect -4950 604494 588874 604536
rect -4950 604258 -3090 604494
rect -2854 604258 -2770 604494
rect -2534 604258 -2450 604494
rect -2214 604258 -2130 604494
rect -1894 604258 1186 604494
rect 1422 604258 8186 604494
rect 8422 604258 15186 604494
rect 15422 604258 22186 604494
rect 22422 604258 29186 604494
rect 29422 604258 36186 604494
rect 36422 604258 43186 604494
rect 43422 604258 50186 604494
rect 50422 604258 57186 604494
rect 57422 604258 64186 604494
rect 64422 604258 71186 604494
rect 71422 604258 78186 604494
rect 78422 604258 85186 604494
rect 85422 604258 92186 604494
rect 92422 604258 99186 604494
rect 99422 604258 106186 604494
rect 106422 604258 113186 604494
rect 113422 604258 120186 604494
rect 120422 604258 127186 604494
rect 127422 604258 134186 604494
rect 134422 604258 141186 604494
rect 141422 604258 148186 604494
rect 148422 604258 155186 604494
rect 155422 604258 162186 604494
rect 162422 604258 169186 604494
rect 169422 604258 176186 604494
rect 176422 604258 183186 604494
rect 183422 604258 190186 604494
rect 190422 604258 197186 604494
rect 197422 604258 204186 604494
rect 204422 604258 211186 604494
rect 211422 604258 218186 604494
rect 218422 604258 225186 604494
rect 225422 604258 232186 604494
rect 232422 604258 239186 604494
rect 239422 604258 246186 604494
rect 246422 604258 253186 604494
rect 253422 604258 260186 604494
rect 260422 604258 267186 604494
rect 267422 604258 274186 604494
rect 274422 604258 281186 604494
rect 281422 604258 288186 604494
rect 288422 604258 295186 604494
rect 295422 604258 302186 604494
rect 302422 604258 309186 604494
rect 309422 604258 316186 604494
rect 316422 604258 323186 604494
rect 323422 604258 330186 604494
rect 330422 604258 337186 604494
rect 337422 604258 344186 604494
rect 344422 604258 351186 604494
rect 351422 604258 358186 604494
rect 358422 604258 365186 604494
rect 365422 604258 372186 604494
rect 372422 604258 379186 604494
rect 379422 604258 386186 604494
rect 386422 604258 393186 604494
rect 393422 604258 400186 604494
rect 400422 604258 407186 604494
rect 407422 604258 414186 604494
rect 414422 604258 421186 604494
rect 421422 604258 428186 604494
rect 428422 604258 435186 604494
rect 435422 604258 442186 604494
rect 442422 604258 449186 604494
rect 449422 604258 456186 604494
rect 456422 604258 463186 604494
rect 463422 604258 470186 604494
rect 470422 604258 477186 604494
rect 477422 604258 484186 604494
rect 484422 604258 491186 604494
rect 491422 604258 498186 604494
rect 498422 604258 505186 604494
rect 505422 604258 512186 604494
rect 512422 604258 519186 604494
rect 519422 604258 526186 604494
rect 526422 604258 533186 604494
rect 533422 604258 540186 604494
rect 540422 604258 547186 604494
rect 547422 604258 554186 604494
rect 554422 604258 561186 604494
rect 561422 604258 568186 604494
rect 568422 604258 575186 604494
rect 575422 604258 582186 604494
rect 582422 604258 585818 604494
rect 586054 604258 586138 604494
rect 586374 604258 586458 604494
rect 586694 604258 586778 604494
rect 587014 604258 588874 604494
rect -4950 604216 588874 604258
rect -4950 598434 588874 598476
rect -4950 598198 -4842 598434
rect -4606 598198 -4522 598434
rect -4286 598198 -4202 598434
rect -3966 598198 -3882 598434
rect -3646 598198 2918 598434
rect 3154 598198 9918 598434
rect 10154 598198 16918 598434
rect 17154 598198 23918 598434
rect 24154 598198 30918 598434
rect 31154 598198 37918 598434
rect 38154 598198 44918 598434
rect 45154 598198 51918 598434
rect 52154 598198 58918 598434
rect 59154 598198 65918 598434
rect 66154 598198 72918 598434
rect 73154 598198 79918 598434
rect 80154 598198 86918 598434
rect 87154 598198 93918 598434
rect 94154 598198 100918 598434
rect 101154 598198 107918 598434
rect 108154 598198 114918 598434
rect 115154 598198 121918 598434
rect 122154 598198 128918 598434
rect 129154 598198 135918 598434
rect 136154 598198 142918 598434
rect 143154 598198 149918 598434
rect 150154 598198 156918 598434
rect 157154 598198 163918 598434
rect 164154 598198 170918 598434
rect 171154 598198 177918 598434
rect 178154 598198 184918 598434
rect 185154 598198 191918 598434
rect 192154 598198 198918 598434
rect 199154 598198 205918 598434
rect 206154 598198 212918 598434
rect 213154 598198 219918 598434
rect 220154 598198 226918 598434
rect 227154 598198 233918 598434
rect 234154 598198 240918 598434
rect 241154 598198 247918 598434
rect 248154 598198 254918 598434
rect 255154 598198 261918 598434
rect 262154 598198 268918 598434
rect 269154 598198 275918 598434
rect 276154 598198 282918 598434
rect 283154 598198 289918 598434
rect 290154 598198 296918 598434
rect 297154 598198 303918 598434
rect 304154 598198 310918 598434
rect 311154 598198 317918 598434
rect 318154 598198 324918 598434
rect 325154 598198 331918 598434
rect 332154 598198 338918 598434
rect 339154 598198 345918 598434
rect 346154 598198 352918 598434
rect 353154 598198 359918 598434
rect 360154 598198 366918 598434
rect 367154 598198 373918 598434
rect 374154 598198 380918 598434
rect 381154 598198 387918 598434
rect 388154 598198 394918 598434
rect 395154 598198 401918 598434
rect 402154 598198 408918 598434
rect 409154 598198 415918 598434
rect 416154 598198 422918 598434
rect 423154 598198 429918 598434
rect 430154 598198 436918 598434
rect 437154 598198 443918 598434
rect 444154 598198 450918 598434
rect 451154 598198 457918 598434
rect 458154 598198 464918 598434
rect 465154 598198 471918 598434
rect 472154 598198 478918 598434
rect 479154 598198 485918 598434
rect 486154 598198 492918 598434
rect 493154 598198 499918 598434
rect 500154 598198 506918 598434
rect 507154 598198 513918 598434
rect 514154 598198 520918 598434
rect 521154 598198 527918 598434
rect 528154 598198 534918 598434
rect 535154 598198 541918 598434
rect 542154 598198 548918 598434
rect 549154 598198 555918 598434
rect 556154 598198 562918 598434
rect 563154 598198 569918 598434
rect 570154 598198 576918 598434
rect 577154 598198 587570 598434
rect 587806 598198 587890 598434
rect 588126 598198 588210 598434
rect 588446 598198 588530 598434
rect 588766 598198 588874 598434
rect -4950 598156 588874 598198
rect -4950 597494 588874 597536
rect -4950 597258 -3090 597494
rect -2854 597258 -2770 597494
rect -2534 597258 -2450 597494
rect -2214 597258 -2130 597494
rect -1894 597258 1186 597494
rect 1422 597258 8186 597494
rect 8422 597258 15186 597494
rect 15422 597258 22186 597494
rect 22422 597258 29186 597494
rect 29422 597258 36186 597494
rect 36422 597258 43186 597494
rect 43422 597258 50186 597494
rect 50422 597258 57186 597494
rect 57422 597258 64186 597494
rect 64422 597258 71186 597494
rect 71422 597258 78186 597494
rect 78422 597258 85186 597494
rect 85422 597258 92186 597494
rect 92422 597258 99186 597494
rect 99422 597258 106186 597494
rect 106422 597258 113186 597494
rect 113422 597258 120186 597494
rect 120422 597258 127186 597494
rect 127422 597258 134186 597494
rect 134422 597258 141186 597494
rect 141422 597258 148186 597494
rect 148422 597258 155186 597494
rect 155422 597258 162186 597494
rect 162422 597258 169186 597494
rect 169422 597258 176186 597494
rect 176422 597258 183186 597494
rect 183422 597258 190186 597494
rect 190422 597258 197186 597494
rect 197422 597258 204186 597494
rect 204422 597258 211186 597494
rect 211422 597258 218186 597494
rect 218422 597258 225186 597494
rect 225422 597258 232186 597494
rect 232422 597258 239186 597494
rect 239422 597258 246186 597494
rect 246422 597258 253186 597494
rect 253422 597258 260186 597494
rect 260422 597258 267186 597494
rect 267422 597258 274186 597494
rect 274422 597258 281186 597494
rect 281422 597258 288186 597494
rect 288422 597258 295186 597494
rect 295422 597258 302186 597494
rect 302422 597258 309186 597494
rect 309422 597258 316186 597494
rect 316422 597258 323186 597494
rect 323422 597258 330186 597494
rect 330422 597258 337186 597494
rect 337422 597258 344186 597494
rect 344422 597258 351186 597494
rect 351422 597258 358186 597494
rect 358422 597258 365186 597494
rect 365422 597258 372186 597494
rect 372422 597258 379186 597494
rect 379422 597258 386186 597494
rect 386422 597258 393186 597494
rect 393422 597258 400186 597494
rect 400422 597258 407186 597494
rect 407422 597258 414186 597494
rect 414422 597258 421186 597494
rect 421422 597258 428186 597494
rect 428422 597258 435186 597494
rect 435422 597258 442186 597494
rect 442422 597258 449186 597494
rect 449422 597258 456186 597494
rect 456422 597258 463186 597494
rect 463422 597258 470186 597494
rect 470422 597258 477186 597494
rect 477422 597258 484186 597494
rect 484422 597258 491186 597494
rect 491422 597258 498186 597494
rect 498422 597258 505186 597494
rect 505422 597258 512186 597494
rect 512422 597258 519186 597494
rect 519422 597258 526186 597494
rect 526422 597258 533186 597494
rect 533422 597258 540186 597494
rect 540422 597258 547186 597494
rect 547422 597258 554186 597494
rect 554422 597258 561186 597494
rect 561422 597258 568186 597494
rect 568422 597258 575186 597494
rect 575422 597258 582186 597494
rect 582422 597258 585818 597494
rect 586054 597258 586138 597494
rect 586374 597258 586458 597494
rect 586694 597258 586778 597494
rect 587014 597258 588874 597494
rect -4950 597216 588874 597258
rect -4950 591434 588874 591476
rect -4950 591198 -4842 591434
rect -4606 591198 -4522 591434
rect -4286 591198 -4202 591434
rect -3966 591198 -3882 591434
rect -3646 591198 2918 591434
rect 3154 591198 9918 591434
rect 10154 591198 16918 591434
rect 17154 591198 23918 591434
rect 24154 591198 30918 591434
rect 31154 591198 37918 591434
rect 38154 591198 44918 591434
rect 45154 591198 51918 591434
rect 52154 591198 58918 591434
rect 59154 591198 65918 591434
rect 66154 591198 72918 591434
rect 73154 591198 79918 591434
rect 80154 591198 86918 591434
rect 87154 591198 93918 591434
rect 94154 591198 100918 591434
rect 101154 591198 107918 591434
rect 108154 591198 114918 591434
rect 115154 591198 121918 591434
rect 122154 591198 128918 591434
rect 129154 591198 135918 591434
rect 136154 591198 142918 591434
rect 143154 591198 149918 591434
rect 150154 591198 156918 591434
rect 157154 591198 163918 591434
rect 164154 591198 170918 591434
rect 171154 591198 177918 591434
rect 178154 591198 184918 591434
rect 185154 591198 191918 591434
rect 192154 591198 198918 591434
rect 199154 591198 205918 591434
rect 206154 591198 212918 591434
rect 213154 591198 219918 591434
rect 220154 591198 226918 591434
rect 227154 591198 233918 591434
rect 234154 591198 240918 591434
rect 241154 591198 247918 591434
rect 248154 591198 254918 591434
rect 255154 591198 261918 591434
rect 262154 591198 268918 591434
rect 269154 591198 275918 591434
rect 276154 591198 282918 591434
rect 283154 591198 289918 591434
rect 290154 591198 296918 591434
rect 297154 591198 303918 591434
rect 304154 591198 310918 591434
rect 311154 591198 317918 591434
rect 318154 591198 324918 591434
rect 325154 591198 331918 591434
rect 332154 591198 338918 591434
rect 339154 591198 345918 591434
rect 346154 591198 352918 591434
rect 353154 591198 359918 591434
rect 360154 591198 366918 591434
rect 367154 591198 373918 591434
rect 374154 591198 380918 591434
rect 381154 591198 387918 591434
rect 388154 591198 394918 591434
rect 395154 591198 401918 591434
rect 402154 591198 408918 591434
rect 409154 591198 415918 591434
rect 416154 591198 422918 591434
rect 423154 591198 429918 591434
rect 430154 591198 436918 591434
rect 437154 591198 443918 591434
rect 444154 591198 450918 591434
rect 451154 591198 457918 591434
rect 458154 591198 464918 591434
rect 465154 591198 471918 591434
rect 472154 591198 478918 591434
rect 479154 591198 485918 591434
rect 486154 591198 492918 591434
rect 493154 591198 499918 591434
rect 500154 591198 506918 591434
rect 507154 591198 513918 591434
rect 514154 591198 520918 591434
rect 521154 591198 527918 591434
rect 528154 591198 534918 591434
rect 535154 591198 541918 591434
rect 542154 591198 548918 591434
rect 549154 591198 555918 591434
rect 556154 591198 562918 591434
rect 563154 591198 569918 591434
rect 570154 591198 576918 591434
rect 577154 591198 587570 591434
rect 587806 591198 587890 591434
rect 588126 591198 588210 591434
rect 588446 591198 588530 591434
rect 588766 591198 588874 591434
rect -4950 591156 588874 591198
rect -4950 590494 588874 590536
rect -4950 590258 -3090 590494
rect -2854 590258 -2770 590494
rect -2534 590258 -2450 590494
rect -2214 590258 -2130 590494
rect -1894 590258 1186 590494
rect 1422 590258 8186 590494
rect 8422 590258 15186 590494
rect 15422 590258 22186 590494
rect 22422 590258 29186 590494
rect 29422 590258 36186 590494
rect 36422 590258 43186 590494
rect 43422 590258 50186 590494
rect 50422 590258 57186 590494
rect 57422 590258 64186 590494
rect 64422 590258 71186 590494
rect 71422 590258 78186 590494
rect 78422 590258 85186 590494
rect 85422 590258 92186 590494
rect 92422 590258 99186 590494
rect 99422 590258 106186 590494
rect 106422 590258 113186 590494
rect 113422 590258 120186 590494
rect 120422 590258 127186 590494
rect 127422 590258 134186 590494
rect 134422 590258 141186 590494
rect 141422 590258 148186 590494
rect 148422 590258 155186 590494
rect 155422 590258 162186 590494
rect 162422 590258 169186 590494
rect 169422 590258 176186 590494
rect 176422 590258 183186 590494
rect 183422 590258 190186 590494
rect 190422 590258 197186 590494
rect 197422 590258 204186 590494
rect 204422 590258 211186 590494
rect 211422 590258 218186 590494
rect 218422 590258 225186 590494
rect 225422 590258 232186 590494
rect 232422 590258 239186 590494
rect 239422 590258 246186 590494
rect 246422 590258 253186 590494
rect 253422 590258 260186 590494
rect 260422 590258 267186 590494
rect 267422 590258 274186 590494
rect 274422 590258 281186 590494
rect 281422 590258 288186 590494
rect 288422 590258 295186 590494
rect 295422 590258 302186 590494
rect 302422 590258 309186 590494
rect 309422 590258 316186 590494
rect 316422 590258 323186 590494
rect 323422 590258 330186 590494
rect 330422 590258 337186 590494
rect 337422 590258 344186 590494
rect 344422 590258 351186 590494
rect 351422 590258 358186 590494
rect 358422 590258 365186 590494
rect 365422 590258 372186 590494
rect 372422 590258 379186 590494
rect 379422 590258 386186 590494
rect 386422 590258 393186 590494
rect 393422 590258 400186 590494
rect 400422 590258 407186 590494
rect 407422 590258 414186 590494
rect 414422 590258 421186 590494
rect 421422 590258 428186 590494
rect 428422 590258 435186 590494
rect 435422 590258 442186 590494
rect 442422 590258 449186 590494
rect 449422 590258 456186 590494
rect 456422 590258 463186 590494
rect 463422 590258 470186 590494
rect 470422 590258 477186 590494
rect 477422 590258 484186 590494
rect 484422 590258 491186 590494
rect 491422 590258 498186 590494
rect 498422 590258 505186 590494
rect 505422 590258 512186 590494
rect 512422 590258 519186 590494
rect 519422 590258 526186 590494
rect 526422 590258 533186 590494
rect 533422 590258 540186 590494
rect 540422 590258 547186 590494
rect 547422 590258 554186 590494
rect 554422 590258 561186 590494
rect 561422 590258 568186 590494
rect 568422 590258 575186 590494
rect 575422 590258 582186 590494
rect 582422 590258 585818 590494
rect 586054 590258 586138 590494
rect 586374 590258 586458 590494
rect 586694 590258 586778 590494
rect 587014 590258 588874 590494
rect -4950 590216 588874 590258
rect -4950 584434 588874 584476
rect -4950 584198 -4842 584434
rect -4606 584198 -4522 584434
rect -4286 584198 -4202 584434
rect -3966 584198 -3882 584434
rect -3646 584198 2918 584434
rect 3154 584198 9918 584434
rect 10154 584198 16918 584434
rect 17154 584198 23918 584434
rect 24154 584198 30918 584434
rect 31154 584198 37918 584434
rect 38154 584198 44918 584434
rect 45154 584198 51918 584434
rect 52154 584198 58918 584434
rect 59154 584198 65918 584434
rect 66154 584198 72918 584434
rect 73154 584198 79918 584434
rect 80154 584198 86918 584434
rect 87154 584198 93918 584434
rect 94154 584198 100918 584434
rect 101154 584198 107918 584434
rect 108154 584198 114918 584434
rect 115154 584198 121918 584434
rect 122154 584198 128918 584434
rect 129154 584198 135918 584434
rect 136154 584198 142918 584434
rect 143154 584198 149918 584434
rect 150154 584198 156918 584434
rect 157154 584198 163918 584434
rect 164154 584198 170918 584434
rect 171154 584198 177918 584434
rect 178154 584198 184918 584434
rect 185154 584198 191918 584434
rect 192154 584198 198918 584434
rect 199154 584198 205918 584434
rect 206154 584198 212918 584434
rect 213154 584198 219918 584434
rect 220154 584198 226918 584434
rect 227154 584198 233918 584434
rect 234154 584198 240918 584434
rect 241154 584198 247918 584434
rect 248154 584198 254918 584434
rect 255154 584198 261918 584434
rect 262154 584198 268918 584434
rect 269154 584198 275918 584434
rect 276154 584198 282918 584434
rect 283154 584198 289918 584434
rect 290154 584198 296918 584434
rect 297154 584198 303918 584434
rect 304154 584198 310918 584434
rect 311154 584198 317918 584434
rect 318154 584198 324918 584434
rect 325154 584198 331918 584434
rect 332154 584198 338918 584434
rect 339154 584198 345918 584434
rect 346154 584198 352918 584434
rect 353154 584198 359918 584434
rect 360154 584198 366918 584434
rect 367154 584198 373918 584434
rect 374154 584198 380918 584434
rect 381154 584198 387918 584434
rect 388154 584198 394918 584434
rect 395154 584198 401918 584434
rect 402154 584198 408918 584434
rect 409154 584198 415918 584434
rect 416154 584198 422918 584434
rect 423154 584198 429918 584434
rect 430154 584198 436918 584434
rect 437154 584198 443918 584434
rect 444154 584198 450918 584434
rect 451154 584198 457918 584434
rect 458154 584198 464918 584434
rect 465154 584198 471918 584434
rect 472154 584198 478918 584434
rect 479154 584198 485918 584434
rect 486154 584198 492918 584434
rect 493154 584198 499918 584434
rect 500154 584198 506918 584434
rect 507154 584198 513918 584434
rect 514154 584198 520918 584434
rect 521154 584198 527918 584434
rect 528154 584198 534918 584434
rect 535154 584198 541918 584434
rect 542154 584198 548918 584434
rect 549154 584198 555918 584434
rect 556154 584198 562918 584434
rect 563154 584198 569918 584434
rect 570154 584198 576918 584434
rect 577154 584198 587570 584434
rect 587806 584198 587890 584434
rect 588126 584198 588210 584434
rect 588446 584198 588530 584434
rect 588766 584198 588874 584434
rect -4950 584156 588874 584198
rect -4950 583494 588874 583536
rect -4950 583258 -3090 583494
rect -2854 583258 -2770 583494
rect -2534 583258 -2450 583494
rect -2214 583258 -2130 583494
rect -1894 583258 1186 583494
rect 1422 583258 8186 583494
rect 8422 583258 15186 583494
rect 15422 583258 22186 583494
rect 22422 583258 29186 583494
rect 29422 583258 36186 583494
rect 36422 583258 43186 583494
rect 43422 583258 50186 583494
rect 50422 583258 57186 583494
rect 57422 583258 64186 583494
rect 64422 583258 71186 583494
rect 71422 583258 78186 583494
rect 78422 583258 85186 583494
rect 85422 583258 92186 583494
rect 92422 583258 99186 583494
rect 99422 583258 106186 583494
rect 106422 583258 113186 583494
rect 113422 583258 120186 583494
rect 120422 583258 127186 583494
rect 127422 583258 134186 583494
rect 134422 583258 141186 583494
rect 141422 583258 148186 583494
rect 148422 583258 155186 583494
rect 155422 583258 162186 583494
rect 162422 583258 169186 583494
rect 169422 583258 176186 583494
rect 176422 583258 183186 583494
rect 183422 583258 190186 583494
rect 190422 583258 197186 583494
rect 197422 583258 204186 583494
rect 204422 583258 211186 583494
rect 211422 583258 218186 583494
rect 218422 583258 225186 583494
rect 225422 583258 232186 583494
rect 232422 583258 239186 583494
rect 239422 583258 246186 583494
rect 246422 583258 253186 583494
rect 253422 583258 260186 583494
rect 260422 583258 267186 583494
rect 267422 583258 274186 583494
rect 274422 583258 281186 583494
rect 281422 583258 288186 583494
rect 288422 583258 295186 583494
rect 295422 583258 302186 583494
rect 302422 583258 309186 583494
rect 309422 583258 316186 583494
rect 316422 583258 323186 583494
rect 323422 583258 330186 583494
rect 330422 583258 337186 583494
rect 337422 583258 344186 583494
rect 344422 583258 351186 583494
rect 351422 583258 358186 583494
rect 358422 583258 365186 583494
rect 365422 583258 372186 583494
rect 372422 583258 379186 583494
rect 379422 583258 386186 583494
rect 386422 583258 393186 583494
rect 393422 583258 400186 583494
rect 400422 583258 407186 583494
rect 407422 583258 414186 583494
rect 414422 583258 421186 583494
rect 421422 583258 428186 583494
rect 428422 583258 435186 583494
rect 435422 583258 442186 583494
rect 442422 583258 449186 583494
rect 449422 583258 456186 583494
rect 456422 583258 463186 583494
rect 463422 583258 470186 583494
rect 470422 583258 477186 583494
rect 477422 583258 484186 583494
rect 484422 583258 491186 583494
rect 491422 583258 498186 583494
rect 498422 583258 505186 583494
rect 505422 583258 512186 583494
rect 512422 583258 519186 583494
rect 519422 583258 526186 583494
rect 526422 583258 533186 583494
rect 533422 583258 540186 583494
rect 540422 583258 547186 583494
rect 547422 583258 554186 583494
rect 554422 583258 561186 583494
rect 561422 583258 568186 583494
rect 568422 583258 575186 583494
rect 575422 583258 582186 583494
rect 582422 583258 585818 583494
rect 586054 583258 586138 583494
rect 586374 583258 586458 583494
rect 586694 583258 586778 583494
rect 587014 583258 588874 583494
rect -4950 583216 588874 583258
rect -4950 577434 588874 577476
rect -4950 577198 -4842 577434
rect -4606 577198 -4522 577434
rect -4286 577198 -4202 577434
rect -3966 577198 -3882 577434
rect -3646 577198 2918 577434
rect 3154 577198 9918 577434
rect 10154 577198 16918 577434
rect 17154 577198 23918 577434
rect 24154 577198 30918 577434
rect 31154 577198 37918 577434
rect 38154 577198 44918 577434
rect 45154 577198 51918 577434
rect 52154 577198 58918 577434
rect 59154 577198 65918 577434
rect 66154 577198 72918 577434
rect 73154 577198 79918 577434
rect 80154 577198 86918 577434
rect 87154 577198 93918 577434
rect 94154 577198 100918 577434
rect 101154 577198 107918 577434
rect 108154 577198 114918 577434
rect 115154 577198 121918 577434
rect 122154 577198 128918 577434
rect 129154 577198 135918 577434
rect 136154 577198 142918 577434
rect 143154 577198 149918 577434
rect 150154 577198 156918 577434
rect 157154 577198 163918 577434
rect 164154 577198 170918 577434
rect 171154 577198 177918 577434
rect 178154 577198 184918 577434
rect 185154 577198 191918 577434
rect 192154 577198 198918 577434
rect 199154 577198 205918 577434
rect 206154 577198 212918 577434
rect 213154 577198 219918 577434
rect 220154 577198 226918 577434
rect 227154 577198 233918 577434
rect 234154 577198 240918 577434
rect 241154 577198 247918 577434
rect 248154 577198 254918 577434
rect 255154 577198 261918 577434
rect 262154 577198 268918 577434
rect 269154 577198 275918 577434
rect 276154 577198 282918 577434
rect 283154 577198 289918 577434
rect 290154 577198 296918 577434
rect 297154 577198 303918 577434
rect 304154 577198 310918 577434
rect 311154 577198 317918 577434
rect 318154 577198 324918 577434
rect 325154 577198 331918 577434
rect 332154 577198 338918 577434
rect 339154 577198 345918 577434
rect 346154 577198 352918 577434
rect 353154 577198 359918 577434
rect 360154 577198 366918 577434
rect 367154 577198 373918 577434
rect 374154 577198 380918 577434
rect 381154 577198 387918 577434
rect 388154 577198 394918 577434
rect 395154 577198 401918 577434
rect 402154 577198 408918 577434
rect 409154 577198 415918 577434
rect 416154 577198 422918 577434
rect 423154 577198 429918 577434
rect 430154 577198 436918 577434
rect 437154 577198 443918 577434
rect 444154 577198 450918 577434
rect 451154 577198 457918 577434
rect 458154 577198 464918 577434
rect 465154 577198 471918 577434
rect 472154 577198 478918 577434
rect 479154 577198 485918 577434
rect 486154 577198 492918 577434
rect 493154 577198 499918 577434
rect 500154 577198 506918 577434
rect 507154 577198 513918 577434
rect 514154 577198 520918 577434
rect 521154 577198 527918 577434
rect 528154 577198 534918 577434
rect 535154 577198 541918 577434
rect 542154 577198 548918 577434
rect 549154 577198 555918 577434
rect 556154 577198 562918 577434
rect 563154 577198 569918 577434
rect 570154 577198 576918 577434
rect 577154 577198 587570 577434
rect 587806 577198 587890 577434
rect 588126 577198 588210 577434
rect 588446 577198 588530 577434
rect 588766 577198 588874 577434
rect -4950 577156 588874 577198
rect -4950 576494 588874 576536
rect -4950 576258 -3090 576494
rect -2854 576258 -2770 576494
rect -2534 576258 -2450 576494
rect -2214 576258 -2130 576494
rect -1894 576258 1186 576494
rect 1422 576258 8186 576494
rect 8422 576258 15186 576494
rect 15422 576258 22186 576494
rect 22422 576258 29186 576494
rect 29422 576258 36186 576494
rect 36422 576258 43186 576494
rect 43422 576258 50186 576494
rect 50422 576258 57186 576494
rect 57422 576258 64186 576494
rect 64422 576258 71186 576494
rect 71422 576258 78186 576494
rect 78422 576258 85186 576494
rect 85422 576258 92186 576494
rect 92422 576258 99186 576494
rect 99422 576258 106186 576494
rect 106422 576258 113186 576494
rect 113422 576258 120186 576494
rect 120422 576258 127186 576494
rect 127422 576258 134186 576494
rect 134422 576258 141186 576494
rect 141422 576258 148186 576494
rect 148422 576258 155186 576494
rect 155422 576258 162186 576494
rect 162422 576258 169186 576494
rect 169422 576258 176186 576494
rect 176422 576258 183186 576494
rect 183422 576258 190186 576494
rect 190422 576258 197186 576494
rect 197422 576258 204186 576494
rect 204422 576258 211186 576494
rect 211422 576258 218186 576494
rect 218422 576258 225186 576494
rect 225422 576258 232186 576494
rect 232422 576258 239186 576494
rect 239422 576258 246186 576494
rect 246422 576258 253186 576494
rect 253422 576258 260186 576494
rect 260422 576258 267186 576494
rect 267422 576258 274186 576494
rect 274422 576258 281186 576494
rect 281422 576258 288186 576494
rect 288422 576258 295186 576494
rect 295422 576258 302186 576494
rect 302422 576258 309186 576494
rect 309422 576258 316186 576494
rect 316422 576258 323186 576494
rect 323422 576258 330186 576494
rect 330422 576258 337186 576494
rect 337422 576258 344186 576494
rect 344422 576258 351186 576494
rect 351422 576258 358186 576494
rect 358422 576258 365186 576494
rect 365422 576258 372186 576494
rect 372422 576258 379186 576494
rect 379422 576258 386186 576494
rect 386422 576258 393186 576494
rect 393422 576258 400186 576494
rect 400422 576258 407186 576494
rect 407422 576258 414186 576494
rect 414422 576258 421186 576494
rect 421422 576258 428186 576494
rect 428422 576258 435186 576494
rect 435422 576258 442186 576494
rect 442422 576258 449186 576494
rect 449422 576258 456186 576494
rect 456422 576258 463186 576494
rect 463422 576258 470186 576494
rect 470422 576258 477186 576494
rect 477422 576258 484186 576494
rect 484422 576258 491186 576494
rect 491422 576258 498186 576494
rect 498422 576258 505186 576494
rect 505422 576258 512186 576494
rect 512422 576258 519186 576494
rect 519422 576258 526186 576494
rect 526422 576258 533186 576494
rect 533422 576258 540186 576494
rect 540422 576258 547186 576494
rect 547422 576258 554186 576494
rect 554422 576258 561186 576494
rect 561422 576258 568186 576494
rect 568422 576258 575186 576494
rect 575422 576258 582186 576494
rect 582422 576258 585818 576494
rect 586054 576258 586138 576494
rect 586374 576258 586458 576494
rect 586694 576258 586778 576494
rect 587014 576258 588874 576494
rect -4950 576216 588874 576258
rect -4950 570434 588874 570476
rect -4950 570198 -4842 570434
rect -4606 570198 -4522 570434
rect -4286 570198 -4202 570434
rect -3966 570198 -3882 570434
rect -3646 570198 2918 570434
rect 3154 570198 9918 570434
rect 10154 570198 16918 570434
rect 17154 570198 23918 570434
rect 24154 570198 30918 570434
rect 31154 570198 37918 570434
rect 38154 570198 44918 570434
rect 45154 570198 51918 570434
rect 52154 570198 58918 570434
rect 59154 570198 65918 570434
rect 66154 570198 72918 570434
rect 73154 570198 79918 570434
rect 80154 570198 86918 570434
rect 87154 570198 93918 570434
rect 94154 570198 100918 570434
rect 101154 570198 107918 570434
rect 108154 570198 114918 570434
rect 115154 570198 121918 570434
rect 122154 570198 128918 570434
rect 129154 570198 135918 570434
rect 136154 570198 142918 570434
rect 143154 570198 149918 570434
rect 150154 570198 156918 570434
rect 157154 570198 163918 570434
rect 164154 570198 170918 570434
rect 171154 570198 177918 570434
rect 178154 570198 184918 570434
rect 185154 570198 191918 570434
rect 192154 570198 198918 570434
rect 199154 570198 205918 570434
rect 206154 570198 212918 570434
rect 213154 570198 219918 570434
rect 220154 570198 226918 570434
rect 227154 570198 233918 570434
rect 234154 570198 240918 570434
rect 241154 570198 247918 570434
rect 248154 570198 254918 570434
rect 255154 570198 261918 570434
rect 262154 570198 268918 570434
rect 269154 570198 275918 570434
rect 276154 570198 282918 570434
rect 283154 570198 289918 570434
rect 290154 570198 296918 570434
rect 297154 570198 303918 570434
rect 304154 570198 310918 570434
rect 311154 570198 317918 570434
rect 318154 570198 324918 570434
rect 325154 570198 331918 570434
rect 332154 570198 338918 570434
rect 339154 570198 345918 570434
rect 346154 570198 352918 570434
rect 353154 570198 359918 570434
rect 360154 570198 366918 570434
rect 367154 570198 373918 570434
rect 374154 570198 380918 570434
rect 381154 570198 387918 570434
rect 388154 570198 394918 570434
rect 395154 570198 401918 570434
rect 402154 570198 408918 570434
rect 409154 570198 415918 570434
rect 416154 570198 422918 570434
rect 423154 570198 429918 570434
rect 430154 570198 436918 570434
rect 437154 570198 443918 570434
rect 444154 570198 450918 570434
rect 451154 570198 457918 570434
rect 458154 570198 464918 570434
rect 465154 570198 471918 570434
rect 472154 570198 478918 570434
rect 479154 570198 485918 570434
rect 486154 570198 492918 570434
rect 493154 570198 499918 570434
rect 500154 570198 506918 570434
rect 507154 570198 513918 570434
rect 514154 570198 520918 570434
rect 521154 570198 527918 570434
rect 528154 570198 534918 570434
rect 535154 570198 541918 570434
rect 542154 570198 548918 570434
rect 549154 570198 555918 570434
rect 556154 570198 562918 570434
rect 563154 570198 569918 570434
rect 570154 570198 576918 570434
rect 577154 570198 587570 570434
rect 587806 570198 587890 570434
rect 588126 570198 588210 570434
rect 588446 570198 588530 570434
rect 588766 570198 588874 570434
rect -4950 570156 588874 570198
rect -4950 569494 588874 569536
rect -4950 569258 -3090 569494
rect -2854 569258 -2770 569494
rect -2534 569258 -2450 569494
rect -2214 569258 -2130 569494
rect -1894 569258 1186 569494
rect 1422 569258 8186 569494
rect 8422 569258 15186 569494
rect 15422 569258 22186 569494
rect 22422 569258 29186 569494
rect 29422 569258 36186 569494
rect 36422 569258 43186 569494
rect 43422 569258 50186 569494
rect 50422 569258 57186 569494
rect 57422 569258 64186 569494
rect 64422 569258 71186 569494
rect 71422 569258 78186 569494
rect 78422 569258 85186 569494
rect 85422 569258 92186 569494
rect 92422 569258 99186 569494
rect 99422 569258 106186 569494
rect 106422 569258 113186 569494
rect 113422 569258 120186 569494
rect 120422 569258 127186 569494
rect 127422 569258 134186 569494
rect 134422 569258 141186 569494
rect 141422 569258 148186 569494
rect 148422 569258 155186 569494
rect 155422 569258 162186 569494
rect 162422 569258 169186 569494
rect 169422 569258 176186 569494
rect 176422 569258 183186 569494
rect 183422 569258 190186 569494
rect 190422 569258 197186 569494
rect 197422 569258 204186 569494
rect 204422 569258 211186 569494
rect 211422 569258 218186 569494
rect 218422 569258 225186 569494
rect 225422 569258 232186 569494
rect 232422 569258 239186 569494
rect 239422 569258 246186 569494
rect 246422 569258 253186 569494
rect 253422 569258 260186 569494
rect 260422 569258 267186 569494
rect 267422 569258 274186 569494
rect 274422 569258 281186 569494
rect 281422 569258 288186 569494
rect 288422 569258 295186 569494
rect 295422 569258 302186 569494
rect 302422 569258 309186 569494
rect 309422 569258 316186 569494
rect 316422 569258 323186 569494
rect 323422 569258 330186 569494
rect 330422 569258 337186 569494
rect 337422 569258 344186 569494
rect 344422 569258 351186 569494
rect 351422 569258 358186 569494
rect 358422 569258 365186 569494
rect 365422 569258 372186 569494
rect 372422 569258 379186 569494
rect 379422 569258 386186 569494
rect 386422 569258 393186 569494
rect 393422 569258 400186 569494
rect 400422 569258 407186 569494
rect 407422 569258 414186 569494
rect 414422 569258 421186 569494
rect 421422 569258 428186 569494
rect 428422 569258 435186 569494
rect 435422 569258 442186 569494
rect 442422 569258 449186 569494
rect 449422 569258 456186 569494
rect 456422 569258 463186 569494
rect 463422 569258 470186 569494
rect 470422 569258 477186 569494
rect 477422 569258 484186 569494
rect 484422 569258 491186 569494
rect 491422 569258 498186 569494
rect 498422 569258 505186 569494
rect 505422 569258 512186 569494
rect 512422 569258 519186 569494
rect 519422 569258 526186 569494
rect 526422 569258 533186 569494
rect 533422 569258 540186 569494
rect 540422 569258 547186 569494
rect 547422 569258 554186 569494
rect 554422 569258 561186 569494
rect 561422 569258 568186 569494
rect 568422 569258 575186 569494
rect 575422 569258 582186 569494
rect 582422 569258 585818 569494
rect 586054 569258 586138 569494
rect 586374 569258 586458 569494
rect 586694 569258 586778 569494
rect 587014 569258 588874 569494
rect -4950 569216 588874 569258
rect -4950 563434 588874 563476
rect -4950 563198 -4842 563434
rect -4606 563198 -4522 563434
rect -4286 563198 -4202 563434
rect -3966 563198 -3882 563434
rect -3646 563198 2918 563434
rect 3154 563198 9918 563434
rect 10154 563198 16918 563434
rect 17154 563198 23918 563434
rect 24154 563198 30918 563434
rect 31154 563198 37918 563434
rect 38154 563198 44918 563434
rect 45154 563198 51918 563434
rect 52154 563198 58918 563434
rect 59154 563198 65918 563434
rect 66154 563198 72918 563434
rect 73154 563198 79918 563434
rect 80154 563198 86918 563434
rect 87154 563198 93918 563434
rect 94154 563198 100918 563434
rect 101154 563198 107918 563434
rect 108154 563198 114918 563434
rect 115154 563198 121918 563434
rect 122154 563198 128918 563434
rect 129154 563198 135918 563434
rect 136154 563198 142918 563434
rect 143154 563198 149918 563434
rect 150154 563198 156918 563434
rect 157154 563198 163918 563434
rect 164154 563198 170918 563434
rect 171154 563198 177918 563434
rect 178154 563198 184918 563434
rect 185154 563198 191918 563434
rect 192154 563198 198918 563434
rect 199154 563198 205918 563434
rect 206154 563198 212918 563434
rect 213154 563198 219918 563434
rect 220154 563198 226918 563434
rect 227154 563198 233918 563434
rect 234154 563198 240918 563434
rect 241154 563198 247918 563434
rect 248154 563198 254918 563434
rect 255154 563198 261918 563434
rect 262154 563198 268918 563434
rect 269154 563198 275918 563434
rect 276154 563198 282918 563434
rect 283154 563198 289918 563434
rect 290154 563198 296918 563434
rect 297154 563198 303918 563434
rect 304154 563198 310918 563434
rect 311154 563198 317918 563434
rect 318154 563198 324918 563434
rect 325154 563198 331918 563434
rect 332154 563198 338918 563434
rect 339154 563198 345918 563434
rect 346154 563198 352918 563434
rect 353154 563198 359918 563434
rect 360154 563198 366918 563434
rect 367154 563198 373918 563434
rect 374154 563198 380918 563434
rect 381154 563198 387918 563434
rect 388154 563198 394918 563434
rect 395154 563198 401918 563434
rect 402154 563198 408918 563434
rect 409154 563198 415918 563434
rect 416154 563198 422918 563434
rect 423154 563198 429918 563434
rect 430154 563198 436918 563434
rect 437154 563198 443918 563434
rect 444154 563198 450918 563434
rect 451154 563198 457918 563434
rect 458154 563198 464918 563434
rect 465154 563198 471918 563434
rect 472154 563198 478918 563434
rect 479154 563198 485918 563434
rect 486154 563198 492918 563434
rect 493154 563198 499918 563434
rect 500154 563198 506918 563434
rect 507154 563198 513918 563434
rect 514154 563198 520918 563434
rect 521154 563198 527918 563434
rect 528154 563198 534918 563434
rect 535154 563198 541918 563434
rect 542154 563198 548918 563434
rect 549154 563198 555918 563434
rect 556154 563198 562918 563434
rect 563154 563198 569918 563434
rect 570154 563198 576918 563434
rect 577154 563198 587570 563434
rect 587806 563198 587890 563434
rect 588126 563198 588210 563434
rect 588446 563198 588530 563434
rect 588766 563198 588874 563434
rect -4950 563156 588874 563198
rect -4950 562494 588874 562536
rect -4950 562258 -3090 562494
rect -2854 562258 -2770 562494
rect -2534 562258 -2450 562494
rect -2214 562258 -2130 562494
rect -1894 562258 1186 562494
rect 1422 562258 8186 562494
rect 8422 562258 15186 562494
rect 15422 562258 22186 562494
rect 22422 562258 29186 562494
rect 29422 562258 36186 562494
rect 36422 562258 43186 562494
rect 43422 562258 50186 562494
rect 50422 562258 57186 562494
rect 57422 562258 64186 562494
rect 64422 562258 71186 562494
rect 71422 562258 78186 562494
rect 78422 562258 85186 562494
rect 85422 562258 92186 562494
rect 92422 562258 99186 562494
rect 99422 562258 106186 562494
rect 106422 562258 113186 562494
rect 113422 562258 120186 562494
rect 120422 562258 127186 562494
rect 127422 562258 134186 562494
rect 134422 562258 141186 562494
rect 141422 562258 148186 562494
rect 148422 562258 155186 562494
rect 155422 562258 162186 562494
rect 162422 562258 169186 562494
rect 169422 562258 176186 562494
rect 176422 562258 183186 562494
rect 183422 562258 190186 562494
rect 190422 562258 197186 562494
rect 197422 562258 204186 562494
rect 204422 562258 211186 562494
rect 211422 562258 218186 562494
rect 218422 562258 225186 562494
rect 225422 562258 232186 562494
rect 232422 562258 239186 562494
rect 239422 562258 246186 562494
rect 246422 562258 253186 562494
rect 253422 562258 260186 562494
rect 260422 562258 267186 562494
rect 267422 562258 274186 562494
rect 274422 562258 281186 562494
rect 281422 562258 288186 562494
rect 288422 562258 295186 562494
rect 295422 562258 302186 562494
rect 302422 562258 309186 562494
rect 309422 562258 316186 562494
rect 316422 562258 323186 562494
rect 323422 562258 330186 562494
rect 330422 562258 337186 562494
rect 337422 562258 344186 562494
rect 344422 562258 351186 562494
rect 351422 562258 358186 562494
rect 358422 562258 365186 562494
rect 365422 562258 372186 562494
rect 372422 562258 379186 562494
rect 379422 562258 386186 562494
rect 386422 562258 393186 562494
rect 393422 562258 400186 562494
rect 400422 562258 407186 562494
rect 407422 562258 414186 562494
rect 414422 562258 421186 562494
rect 421422 562258 428186 562494
rect 428422 562258 435186 562494
rect 435422 562258 442186 562494
rect 442422 562258 449186 562494
rect 449422 562258 456186 562494
rect 456422 562258 463186 562494
rect 463422 562258 470186 562494
rect 470422 562258 477186 562494
rect 477422 562258 484186 562494
rect 484422 562258 491186 562494
rect 491422 562258 498186 562494
rect 498422 562258 505186 562494
rect 505422 562258 512186 562494
rect 512422 562258 519186 562494
rect 519422 562258 526186 562494
rect 526422 562258 533186 562494
rect 533422 562258 540186 562494
rect 540422 562258 547186 562494
rect 547422 562258 554186 562494
rect 554422 562258 561186 562494
rect 561422 562258 568186 562494
rect 568422 562258 575186 562494
rect 575422 562258 582186 562494
rect 582422 562258 585818 562494
rect 586054 562258 586138 562494
rect 586374 562258 586458 562494
rect 586694 562258 586778 562494
rect 587014 562258 588874 562494
rect -4950 562216 588874 562258
rect -4950 556434 588874 556476
rect -4950 556198 -4842 556434
rect -4606 556198 -4522 556434
rect -4286 556198 -4202 556434
rect -3966 556198 -3882 556434
rect -3646 556198 2918 556434
rect 3154 556198 9918 556434
rect 10154 556198 16918 556434
rect 17154 556198 23918 556434
rect 24154 556198 30918 556434
rect 31154 556198 37918 556434
rect 38154 556198 44918 556434
rect 45154 556198 51918 556434
rect 52154 556198 58918 556434
rect 59154 556198 65918 556434
rect 66154 556198 72918 556434
rect 73154 556198 79918 556434
rect 80154 556198 86918 556434
rect 87154 556198 93918 556434
rect 94154 556198 100918 556434
rect 101154 556198 107918 556434
rect 108154 556198 114918 556434
rect 115154 556198 121918 556434
rect 122154 556198 128918 556434
rect 129154 556198 135918 556434
rect 136154 556198 142918 556434
rect 143154 556198 149918 556434
rect 150154 556198 156918 556434
rect 157154 556198 163918 556434
rect 164154 556198 170918 556434
rect 171154 556198 177918 556434
rect 178154 556198 184918 556434
rect 185154 556198 191918 556434
rect 192154 556198 198918 556434
rect 199154 556198 205918 556434
rect 206154 556198 212918 556434
rect 213154 556198 219918 556434
rect 220154 556198 226918 556434
rect 227154 556198 233918 556434
rect 234154 556198 240918 556434
rect 241154 556198 247918 556434
rect 248154 556198 254918 556434
rect 255154 556198 261918 556434
rect 262154 556198 268918 556434
rect 269154 556198 275918 556434
rect 276154 556198 282918 556434
rect 283154 556198 289918 556434
rect 290154 556198 296918 556434
rect 297154 556198 303918 556434
rect 304154 556198 310918 556434
rect 311154 556198 317918 556434
rect 318154 556198 324918 556434
rect 325154 556198 331918 556434
rect 332154 556198 338918 556434
rect 339154 556198 345918 556434
rect 346154 556198 352918 556434
rect 353154 556198 359918 556434
rect 360154 556198 366918 556434
rect 367154 556198 373918 556434
rect 374154 556198 380918 556434
rect 381154 556198 387918 556434
rect 388154 556198 394918 556434
rect 395154 556198 401918 556434
rect 402154 556198 408918 556434
rect 409154 556198 415918 556434
rect 416154 556198 422918 556434
rect 423154 556198 429918 556434
rect 430154 556198 436918 556434
rect 437154 556198 443918 556434
rect 444154 556198 450918 556434
rect 451154 556198 457918 556434
rect 458154 556198 464918 556434
rect 465154 556198 471918 556434
rect 472154 556198 478918 556434
rect 479154 556198 485918 556434
rect 486154 556198 492918 556434
rect 493154 556198 499918 556434
rect 500154 556198 506918 556434
rect 507154 556198 513918 556434
rect 514154 556198 520918 556434
rect 521154 556198 527918 556434
rect 528154 556198 534918 556434
rect 535154 556198 541918 556434
rect 542154 556198 548918 556434
rect 549154 556198 555918 556434
rect 556154 556198 562918 556434
rect 563154 556198 569918 556434
rect 570154 556198 576918 556434
rect 577154 556198 587570 556434
rect 587806 556198 587890 556434
rect 588126 556198 588210 556434
rect 588446 556198 588530 556434
rect 588766 556198 588874 556434
rect -4950 556156 588874 556198
rect -4950 555494 588874 555536
rect -4950 555258 -3090 555494
rect -2854 555258 -2770 555494
rect -2534 555258 -2450 555494
rect -2214 555258 -2130 555494
rect -1894 555258 1186 555494
rect 1422 555258 8186 555494
rect 8422 555258 15186 555494
rect 15422 555258 22186 555494
rect 22422 555258 29186 555494
rect 29422 555258 36186 555494
rect 36422 555258 43186 555494
rect 43422 555258 50186 555494
rect 50422 555258 57186 555494
rect 57422 555258 64186 555494
rect 64422 555258 71186 555494
rect 71422 555258 78186 555494
rect 78422 555258 85186 555494
rect 85422 555258 92186 555494
rect 92422 555258 99186 555494
rect 99422 555258 106186 555494
rect 106422 555258 113186 555494
rect 113422 555258 120186 555494
rect 120422 555258 127186 555494
rect 127422 555258 134186 555494
rect 134422 555258 141186 555494
rect 141422 555258 148186 555494
rect 148422 555258 155186 555494
rect 155422 555258 162186 555494
rect 162422 555258 169186 555494
rect 169422 555258 176186 555494
rect 176422 555258 183186 555494
rect 183422 555258 190186 555494
rect 190422 555258 197186 555494
rect 197422 555258 204186 555494
rect 204422 555258 211186 555494
rect 211422 555258 218186 555494
rect 218422 555258 225186 555494
rect 225422 555258 232186 555494
rect 232422 555258 239186 555494
rect 239422 555258 246186 555494
rect 246422 555258 253186 555494
rect 253422 555258 260186 555494
rect 260422 555258 267186 555494
rect 267422 555258 274186 555494
rect 274422 555258 281186 555494
rect 281422 555258 288186 555494
rect 288422 555258 295186 555494
rect 295422 555258 302186 555494
rect 302422 555258 309186 555494
rect 309422 555258 316186 555494
rect 316422 555258 323186 555494
rect 323422 555258 330186 555494
rect 330422 555258 337186 555494
rect 337422 555258 344186 555494
rect 344422 555258 351186 555494
rect 351422 555258 358186 555494
rect 358422 555258 365186 555494
rect 365422 555258 372186 555494
rect 372422 555258 379186 555494
rect 379422 555258 386186 555494
rect 386422 555258 393186 555494
rect 393422 555258 400186 555494
rect 400422 555258 407186 555494
rect 407422 555258 414186 555494
rect 414422 555258 421186 555494
rect 421422 555258 428186 555494
rect 428422 555258 435186 555494
rect 435422 555258 442186 555494
rect 442422 555258 449186 555494
rect 449422 555258 456186 555494
rect 456422 555258 463186 555494
rect 463422 555258 470186 555494
rect 470422 555258 477186 555494
rect 477422 555258 484186 555494
rect 484422 555258 491186 555494
rect 491422 555258 498186 555494
rect 498422 555258 505186 555494
rect 505422 555258 512186 555494
rect 512422 555258 519186 555494
rect 519422 555258 526186 555494
rect 526422 555258 533186 555494
rect 533422 555258 540186 555494
rect 540422 555258 547186 555494
rect 547422 555258 554186 555494
rect 554422 555258 561186 555494
rect 561422 555258 568186 555494
rect 568422 555258 575186 555494
rect 575422 555258 582186 555494
rect 582422 555258 585818 555494
rect 586054 555258 586138 555494
rect 586374 555258 586458 555494
rect 586694 555258 586778 555494
rect 587014 555258 588874 555494
rect -4950 555216 588874 555258
rect -4950 549434 588874 549476
rect -4950 549198 -4842 549434
rect -4606 549198 -4522 549434
rect -4286 549198 -4202 549434
rect -3966 549198 -3882 549434
rect -3646 549198 2918 549434
rect 3154 549198 9918 549434
rect 10154 549198 16918 549434
rect 17154 549198 23918 549434
rect 24154 549198 30918 549434
rect 31154 549198 37918 549434
rect 38154 549198 44918 549434
rect 45154 549198 51918 549434
rect 52154 549198 58918 549434
rect 59154 549198 65918 549434
rect 66154 549198 72918 549434
rect 73154 549198 79918 549434
rect 80154 549198 86918 549434
rect 87154 549198 93918 549434
rect 94154 549198 100918 549434
rect 101154 549198 107918 549434
rect 108154 549198 114918 549434
rect 115154 549198 121918 549434
rect 122154 549198 128918 549434
rect 129154 549198 135918 549434
rect 136154 549198 142918 549434
rect 143154 549198 149918 549434
rect 150154 549198 156918 549434
rect 157154 549198 163918 549434
rect 164154 549198 170918 549434
rect 171154 549198 177918 549434
rect 178154 549198 184918 549434
rect 185154 549198 191918 549434
rect 192154 549198 198918 549434
rect 199154 549198 205918 549434
rect 206154 549198 212918 549434
rect 213154 549198 219918 549434
rect 220154 549198 226918 549434
rect 227154 549198 233918 549434
rect 234154 549198 240918 549434
rect 241154 549198 247918 549434
rect 248154 549198 254918 549434
rect 255154 549198 261918 549434
rect 262154 549198 268918 549434
rect 269154 549198 275918 549434
rect 276154 549198 282918 549434
rect 283154 549198 289918 549434
rect 290154 549198 296918 549434
rect 297154 549198 303918 549434
rect 304154 549198 310918 549434
rect 311154 549198 317918 549434
rect 318154 549198 324918 549434
rect 325154 549198 331918 549434
rect 332154 549198 338918 549434
rect 339154 549198 345918 549434
rect 346154 549198 352918 549434
rect 353154 549198 359918 549434
rect 360154 549198 366918 549434
rect 367154 549198 373918 549434
rect 374154 549198 380918 549434
rect 381154 549198 387918 549434
rect 388154 549198 394918 549434
rect 395154 549198 401918 549434
rect 402154 549198 408918 549434
rect 409154 549198 415918 549434
rect 416154 549198 422918 549434
rect 423154 549198 429918 549434
rect 430154 549198 436918 549434
rect 437154 549198 443918 549434
rect 444154 549198 450918 549434
rect 451154 549198 457918 549434
rect 458154 549198 464918 549434
rect 465154 549198 471918 549434
rect 472154 549198 478918 549434
rect 479154 549198 485918 549434
rect 486154 549198 492918 549434
rect 493154 549198 499918 549434
rect 500154 549198 506918 549434
rect 507154 549198 513918 549434
rect 514154 549198 520918 549434
rect 521154 549198 527918 549434
rect 528154 549198 534918 549434
rect 535154 549198 541918 549434
rect 542154 549198 548918 549434
rect 549154 549198 555918 549434
rect 556154 549198 562918 549434
rect 563154 549198 569918 549434
rect 570154 549198 576918 549434
rect 577154 549198 587570 549434
rect 587806 549198 587890 549434
rect 588126 549198 588210 549434
rect 588446 549198 588530 549434
rect 588766 549198 588874 549434
rect -4950 549156 588874 549198
rect -4950 548494 588874 548536
rect -4950 548258 -3090 548494
rect -2854 548258 -2770 548494
rect -2534 548258 -2450 548494
rect -2214 548258 -2130 548494
rect -1894 548258 1186 548494
rect 1422 548258 8186 548494
rect 8422 548258 15186 548494
rect 15422 548258 22186 548494
rect 22422 548258 29186 548494
rect 29422 548258 36186 548494
rect 36422 548258 43186 548494
rect 43422 548258 50186 548494
rect 50422 548258 57186 548494
rect 57422 548258 64186 548494
rect 64422 548258 71186 548494
rect 71422 548258 78186 548494
rect 78422 548258 85186 548494
rect 85422 548258 92186 548494
rect 92422 548258 99186 548494
rect 99422 548258 106186 548494
rect 106422 548258 113186 548494
rect 113422 548258 120186 548494
rect 120422 548258 127186 548494
rect 127422 548258 134186 548494
rect 134422 548258 141186 548494
rect 141422 548258 148186 548494
rect 148422 548258 155186 548494
rect 155422 548258 162186 548494
rect 162422 548258 169186 548494
rect 169422 548258 176186 548494
rect 176422 548258 183186 548494
rect 183422 548258 190186 548494
rect 190422 548258 197186 548494
rect 197422 548258 204186 548494
rect 204422 548258 211186 548494
rect 211422 548258 218186 548494
rect 218422 548258 225186 548494
rect 225422 548258 232186 548494
rect 232422 548258 239186 548494
rect 239422 548258 246186 548494
rect 246422 548258 253186 548494
rect 253422 548258 260186 548494
rect 260422 548258 267186 548494
rect 267422 548258 274186 548494
rect 274422 548258 281186 548494
rect 281422 548258 288186 548494
rect 288422 548258 295186 548494
rect 295422 548258 302186 548494
rect 302422 548258 309186 548494
rect 309422 548258 316186 548494
rect 316422 548258 323186 548494
rect 323422 548258 330186 548494
rect 330422 548258 337186 548494
rect 337422 548258 344186 548494
rect 344422 548258 351186 548494
rect 351422 548258 358186 548494
rect 358422 548258 365186 548494
rect 365422 548258 372186 548494
rect 372422 548258 379186 548494
rect 379422 548258 386186 548494
rect 386422 548258 393186 548494
rect 393422 548258 400186 548494
rect 400422 548258 407186 548494
rect 407422 548258 414186 548494
rect 414422 548258 421186 548494
rect 421422 548258 428186 548494
rect 428422 548258 435186 548494
rect 435422 548258 442186 548494
rect 442422 548258 449186 548494
rect 449422 548258 456186 548494
rect 456422 548258 463186 548494
rect 463422 548258 470186 548494
rect 470422 548258 477186 548494
rect 477422 548258 484186 548494
rect 484422 548258 491186 548494
rect 491422 548258 498186 548494
rect 498422 548258 505186 548494
rect 505422 548258 512186 548494
rect 512422 548258 519186 548494
rect 519422 548258 526186 548494
rect 526422 548258 533186 548494
rect 533422 548258 540186 548494
rect 540422 548258 547186 548494
rect 547422 548258 554186 548494
rect 554422 548258 561186 548494
rect 561422 548258 568186 548494
rect 568422 548258 575186 548494
rect 575422 548258 582186 548494
rect 582422 548258 585818 548494
rect 586054 548258 586138 548494
rect 586374 548258 586458 548494
rect 586694 548258 586778 548494
rect 587014 548258 588874 548494
rect -4950 548216 588874 548258
rect -4950 542434 588874 542476
rect -4950 542198 -4842 542434
rect -4606 542198 -4522 542434
rect -4286 542198 -4202 542434
rect -3966 542198 -3882 542434
rect -3646 542198 2918 542434
rect 3154 542198 9918 542434
rect 10154 542198 16918 542434
rect 17154 542198 23918 542434
rect 24154 542198 30918 542434
rect 31154 542198 37918 542434
rect 38154 542198 44918 542434
rect 45154 542198 51918 542434
rect 52154 542198 58918 542434
rect 59154 542198 65918 542434
rect 66154 542198 72918 542434
rect 73154 542198 79918 542434
rect 80154 542198 86918 542434
rect 87154 542198 93918 542434
rect 94154 542198 100918 542434
rect 101154 542198 107918 542434
rect 108154 542198 114918 542434
rect 115154 542198 121918 542434
rect 122154 542198 128918 542434
rect 129154 542198 135918 542434
rect 136154 542198 142918 542434
rect 143154 542198 149918 542434
rect 150154 542198 156918 542434
rect 157154 542198 163918 542434
rect 164154 542198 170918 542434
rect 171154 542198 177918 542434
rect 178154 542198 184918 542434
rect 185154 542198 191918 542434
rect 192154 542198 198918 542434
rect 199154 542198 205918 542434
rect 206154 542198 212918 542434
rect 213154 542198 219918 542434
rect 220154 542198 226918 542434
rect 227154 542198 233918 542434
rect 234154 542198 240918 542434
rect 241154 542198 247918 542434
rect 248154 542198 254918 542434
rect 255154 542198 261918 542434
rect 262154 542198 268918 542434
rect 269154 542198 275918 542434
rect 276154 542198 282918 542434
rect 283154 542198 289918 542434
rect 290154 542198 296918 542434
rect 297154 542198 303918 542434
rect 304154 542198 310918 542434
rect 311154 542198 317918 542434
rect 318154 542198 324918 542434
rect 325154 542198 331918 542434
rect 332154 542198 338918 542434
rect 339154 542198 345918 542434
rect 346154 542198 352918 542434
rect 353154 542198 359918 542434
rect 360154 542198 366918 542434
rect 367154 542198 373918 542434
rect 374154 542198 380918 542434
rect 381154 542198 387918 542434
rect 388154 542198 394918 542434
rect 395154 542198 401918 542434
rect 402154 542198 408918 542434
rect 409154 542198 415918 542434
rect 416154 542198 422918 542434
rect 423154 542198 429918 542434
rect 430154 542198 436918 542434
rect 437154 542198 443918 542434
rect 444154 542198 450918 542434
rect 451154 542198 457918 542434
rect 458154 542198 464918 542434
rect 465154 542198 471918 542434
rect 472154 542198 478918 542434
rect 479154 542198 485918 542434
rect 486154 542198 492918 542434
rect 493154 542198 499918 542434
rect 500154 542198 506918 542434
rect 507154 542198 513918 542434
rect 514154 542198 520918 542434
rect 521154 542198 527918 542434
rect 528154 542198 534918 542434
rect 535154 542198 541918 542434
rect 542154 542198 548918 542434
rect 549154 542198 555918 542434
rect 556154 542198 562918 542434
rect 563154 542198 569918 542434
rect 570154 542198 576918 542434
rect 577154 542198 587570 542434
rect 587806 542198 587890 542434
rect 588126 542198 588210 542434
rect 588446 542198 588530 542434
rect 588766 542198 588874 542434
rect -4950 542156 588874 542198
rect -4950 541494 588874 541536
rect -4950 541258 -3090 541494
rect -2854 541258 -2770 541494
rect -2534 541258 -2450 541494
rect -2214 541258 -2130 541494
rect -1894 541258 1186 541494
rect 1422 541258 8186 541494
rect 8422 541258 15186 541494
rect 15422 541258 22186 541494
rect 22422 541258 29186 541494
rect 29422 541258 36186 541494
rect 36422 541258 43186 541494
rect 43422 541258 50186 541494
rect 50422 541258 57186 541494
rect 57422 541258 64186 541494
rect 64422 541258 71186 541494
rect 71422 541258 78186 541494
rect 78422 541258 85186 541494
rect 85422 541258 92186 541494
rect 92422 541258 99186 541494
rect 99422 541258 106186 541494
rect 106422 541258 113186 541494
rect 113422 541258 120186 541494
rect 120422 541258 127186 541494
rect 127422 541258 134186 541494
rect 134422 541258 141186 541494
rect 141422 541258 148186 541494
rect 148422 541258 155186 541494
rect 155422 541258 162186 541494
rect 162422 541258 169186 541494
rect 169422 541258 176186 541494
rect 176422 541258 183186 541494
rect 183422 541258 190186 541494
rect 190422 541258 197186 541494
rect 197422 541258 204186 541494
rect 204422 541258 211186 541494
rect 211422 541258 218186 541494
rect 218422 541258 225186 541494
rect 225422 541258 232186 541494
rect 232422 541258 239186 541494
rect 239422 541258 246186 541494
rect 246422 541258 253186 541494
rect 253422 541258 260186 541494
rect 260422 541258 267186 541494
rect 267422 541258 274186 541494
rect 274422 541258 281186 541494
rect 281422 541258 288186 541494
rect 288422 541258 295186 541494
rect 295422 541258 302186 541494
rect 302422 541258 309186 541494
rect 309422 541258 316186 541494
rect 316422 541258 323186 541494
rect 323422 541258 330186 541494
rect 330422 541258 337186 541494
rect 337422 541258 344186 541494
rect 344422 541258 351186 541494
rect 351422 541258 358186 541494
rect 358422 541258 365186 541494
rect 365422 541258 372186 541494
rect 372422 541258 379186 541494
rect 379422 541258 386186 541494
rect 386422 541258 393186 541494
rect 393422 541258 400186 541494
rect 400422 541258 407186 541494
rect 407422 541258 414186 541494
rect 414422 541258 421186 541494
rect 421422 541258 428186 541494
rect 428422 541258 435186 541494
rect 435422 541258 442186 541494
rect 442422 541258 449186 541494
rect 449422 541258 456186 541494
rect 456422 541258 463186 541494
rect 463422 541258 470186 541494
rect 470422 541258 477186 541494
rect 477422 541258 484186 541494
rect 484422 541258 491186 541494
rect 491422 541258 498186 541494
rect 498422 541258 505186 541494
rect 505422 541258 512186 541494
rect 512422 541258 519186 541494
rect 519422 541258 526186 541494
rect 526422 541258 533186 541494
rect 533422 541258 540186 541494
rect 540422 541258 547186 541494
rect 547422 541258 554186 541494
rect 554422 541258 561186 541494
rect 561422 541258 568186 541494
rect 568422 541258 575186 541494
rect 575422 541258 582186 541494
rect 582422 541258 585818 541494
rect 586054 541258 586138 541494
rect 586374 541258 586458 541494
rect 586694 541258 586778 541494
rect 587014 541258 588874 541494
rect -4950 541216 588874 541258
rect -4950 535434 588874 535476
rect -4950 535198 -4842 535434
rect -4606 535198 -4522 535434
rect -4286 535198 -4202 535434
rect -3966 535198 -3882 535434
rect -3646 535198 2918 535434
rect 3154 535198 9918 535434
rect 10154 535198 16918 535434
rect 17154 535198 23918 535434
rect 24154 535198 30918 535434
rect 31154 535198 37918 535434
rect 38154 535198 44918 535434
rect 45154 535198 51918 535434
rect 52154 535198 58918 535434
rect 59154 535198 65918 535434
rect 66154 535198 72918 535434
rect 73154 535198 79918 535434
rect 80154 535198 86918 535434
rect 87154 535198 93918 535434
rect 94154 535198 100918 535434
rect 101154 535198 107918 535434
rect 108154 535198 114918 535434
rect 115154 535198 121918 535434
rect 122154 535198 128918 535434
rect 129154 535198 135918 535434
rect 136154 535198 142918 535434
rect 143154 535198 149918 535434
rect 150154 535198 156918 535434
rect 157154 535198 163918 535434
rect 164154 535198 170918 535434
rect 171154 535198 177918 535434
rect 178154 535198 184918 535434
rect 185154 535198 191918 535434
rect 192154 535198 198918 535434
rect 199154 535198 205918 535434
rect 206154 535198 212918 535434
rect 213154 535198 219918 535434
rect 220154 535198 226918 535434
rect 227154 535198 233918 535434
rect 234154 535198 240918 535434
rect 241154 535198 247918 535434
rect 248154 535198 254918 535434
rect 255154 535198 261918 535434
rect 262154 535198 268918 535434
rect 269154 535198 275918 535434
rect 276154 535198 282918 535434
rect 283154 535198 289918 535434
rect 290154 535198 296918 535434
rect 297154 535198 303918 535434
rect 304154 535198 310918 535434
rect 311154 535198 317918 535434
rect 318154 535198 324918 535434
rect 325154 535198 331918 535434
rect 332154 535198 338918 535434
rect 339154 535198 345918 535434
rect 346154 535198 352918 535434
rect 353154 535198 359918 535434
rect 360154 535198 366918 535434
rect 367154 535198 373918 535434
rect 374154 535198 380918 535434
rect 381154 535198 387918 535434
rect 388154 535198 394918 535434
rect 395154 535198 401918 535434
rect 402154 535198 408918 535434
rect 409154 535198 415918 535434
rect 416154 535198 422918 535434
rect 423154 535198 429918 535434
rect 430154 535198 436918 535434
rect 437154 535198 443918 535434
rect 444154 535198 450918 535434
rect 451154 535198 457918 535434
rect 458154 535198 464918 535434
rect 465154 535198 471918 535434
rect 472154 535198 478918 535434
rect 479154 535198 485918 535434
rect 486154 535198 492918 535434
rect 493154 535198 499918 535434
rect 500154 535198 506918 535434
rect 507154 535198 513918 535434
rect 514154 535198 520918 535434
rect 521154 535198 527918 535434
rect 528154 535198 534918 535434
rect 535154 535198 541918 535434
rect 542154 535198 548918 535434
rect 549154 535198 555918 535434
rect 556154 535198 562918 535434
rect 563154 535198 569918 535434
rect 570154 535198 576918 535434
rect 577154 535198 587570 535434
rect 587806 535198 587890 535434
rect 588126 535198 588210 535434
rect 588446 535198 588530 535434
rect 588766 535198 588874 535434
rect -4950 535156 588874 535198
rect -4950 534494 588874 534536
rect -4950 534258 -3090 534494
rect -2854 534258 -2770 534494
rect -2534 534258 -2450 534494
rect -2214 534258 -2130 534494
rect -1894 534258 1186 534494
rect 1422 534258 8186 534494
rect 8422 534258 15186 534494
rect 15422 534258 22186 534494
rect 22422 534258 29186 534494
rect 29422 534258 36186 534494
rect 36422 534258 43186 534494
rect 43422 534258 50186 534494
rect 50422 534258 57186 534494
rect 57422 534258 64186 534494
rect 64422 534258 71186 534494
rect 71422 534258 78186 534494
rect 78422 534258 85186 534494
rect 85422 534258 92186 534494
rect 92422 534258 99186 534494
rect 99422 534258 106186 534494
rect 106422 534258 113186 534494
rect 113422 534258 120186 534494
rect 120422 534258 127186 534494
rect 127422 534258 134186 534494
rect 134422 534258 141186 534494
rect 141422 534258 148186 534494
rect 148422 534258 155186 534494
rect 155422 534258 162186 534494
rect 162422 534258 169186 534494
rect 169422 534258 176186 534494
rect 176422 534258 183186 534494
rect 183422 534258 190186 534494
rect 190422 534258 197186 534494
rect 197422 534258 204186 534494
rect 204422 534258 211186 534494
rect 211422 534258 218186 534494
rect 218422 534258 225186 534494
rect 225422 534258 232186 534494
rect 232422 534258 239186 534494
rect 239422 534258 246186 534494
rect 246422 534258 253186 534494
rect 253422 534258 260186 534494
rect 260422 534258 267186 534494
rect 267422 534258 274186 534494
rect 274422 534258 281186 534494
rect 281422 534258 288186 534494
rect 288422 534258 295186 534494
rect 295422 534258 302186 534494
rect 302422 534258 309186 534494
rect 309422 534258 316186 534494
rect 316422 534258 323186 534494
rect 323422 534258 330186 534494
rect 330422 534258 337186 534494
rect 337422 534258 344186 534494
rect 344422 534258 351186 534494
rect 351422 534258 358186 534494
rect 358422 534258 365186 534494
rect 365422 534258 372186 534494
rect 372422 534258 379186 534494
rect 379422 534258 386186 534494
rect 386422 534258 393186 534494
rect 393422 534258 400186 534494
rect 400422 534258 407186 534494
rect 407422 534258 414186 534494
rect 414422 534258 421186 534494
rect 421422 534258 428186 534494
rect 428422 534258 435186 534494
rect 435422 534258 442186 534494
rect 442422 534258 449186 534494
rect 449422 534258 456186 534494
rect 456422 534258 463186 534494
rect 463422 534258 470186 534494
rect 470422 534258 477186 534494
rect 477422 534258 484186 534494
rect 484422 534258 491186 534494
rect 491422 534258 498186 534494
rect 498422 534258 505186 534494
rect 505422 534258 512186 534494
rect 512422 534258 519186 534494
rect 519422 534258 526186 534494
rect 526422 534258 533186 534494
rect 533422 534258 540186 534494
rect 540422 534258 547186 534494
rect 547422 534258 554186 534494
rect 554422 534258 561186 534494
rect 561422 534258 568186 534494
rect 568422 534258 575186 534494
rect 575422 534258 582186 534494
rect 582422 534258 585818 534494
rect 586054 534258 586138 534494
rect 586374 534258 586458 534494
rect 586694 534258 586778 534494
rect 587014 534258 588874 534494
rect -4950 534216 588874 534258
rect -4950 528434 588874 528476
rect -4950 528198 -4842 528434
rect -4606 528198 -4522 528434
rect -4286 528198 -4202 528434
rect -3966 528198 -3882 528434
rect -3646 528198 2918 528434
rect 3154 528198 9918 528434
rect 10154 528198 16918 528434
rect 17154 528198 23918 528434
rect 24154 528198 30918 528434
rect 31154 528198 37918 528434
rect 38154 528198 44918 528434
rect 45154 528198 51918 528434
rect 52154 528198 58918 528434
rect 59154 528198 65918 528434
rect 66154 528198 72918 528434
rect 73154 528198 79918 528434
rect 80154 528198 86918 528434
rect 87154 528198 93918 528434
rect 94154 528198 100918 528434
rect 101154 528198 107918 528434
rect 108154 528198 114918 528434
rect 115154 528198 121918 528434
rect 122154 528198 128918 528434
rect 129154 528198 135918 528434
rect 136154 528198 142918 528434
rect 143154 528198 149918 528434
rect 150154 528198 156918 528434
rect 157154 528198 163918 528434
rect 164154 528198 170918 528434
rect 171154 528198 177918 528434
rect 178154 528198 184918 528434
rect 185154 528198 191918 528434
rect 192154 528198 198918 528434
rect 199154 528198 205918 528434
rect 206154 528198 212918 528434
rect 213154 528198 219918 528434
rect 220154 528198 226918 528434
rect 227154 528198 233918 528434
rect 234154 528198 240918 528434
rect 241154 528198 247918 528434
rect 248154 528198 254918 528434
rect 255154 528198 261918 528434
rect 262154 528198 268918 528434
rect 269154 528198 275918 528434
rect 276154 528198 282918 528434
rect 283154 528198 289918 528434
rect 290154 528198 296918 528434
rect 297154 528198 303918 528434
rect 304154 528198 310918 528434
rect 311154 528198 317918 528434
rect 318154 528198 324918 528434
rect 325154 528198 331918 528434
rect 332154 528198 338918 528434
rect 339154 528198 345918 528434
rect 346154 528198 352918 528434
rect 353154 528198 359918 528434
rect 360154 528198 366918 528434
rect 367154 528198 373918 528434
rect 374154 528198 380918 528434
rect 381154 528198 387918 528434
rect 388154 528198 394918 528434
rect 395154 528198 401918 528434
rect 402154 528198 408918 528434
rect 409154 528198 415918 528434
rect 416154 528198 422918 528434
rect 423154 528198 429918 528434
rect 430154 528198 436918 528434
rect 437154 528198 443918 528434
rect 444154 528198 450918 528434
rect 451154 528198 457918 528434
rect 458154 528198 464918 528434
rect 465154 528198 471918 528434
rect 472154 528198 478918 528434
rect 479154 528198 485918 528434
rect 486154 528198 492918 528434
rect 493154 528198 499918 528434
rect 500154 528198 506918 528434
rect 507154 528198 513918 528434
rect 514154 528198 520918 528434
rect 521154 528198 527918 528434
rect 528154 528198 534918 528434
rect 535154 528198 541918 528434
rect 542154 528198 548918 528434
rect 549154 528198 555918 528434
rect 556154 528198 562918 528434
rect 563154 528198 569918 528434
rect 570154 528198 576918 528434
rect 577154 528198 587570 528434
rect 587806 528198 587890 528434
rect 588126 528198 588210 528434
rect 588446 528198 588530 528434
rect 588766 528198 588874 528434
rect -4950 528156 588874 528198
rect -4950 527494 588874 527536
rect -4950 527258 -3090 527494
rect -2854 527258 -2770 527494
rect -2534 527258 -2450 527494
rect -2214 527258 -2130 527494
rect -1894 527258 1186 527494
rect 1422 527258 8186 527494
rect 8422 527258 15186 527494
rect 15422 527258 22186 527494
rect 22422 527258 29186 527494
rect 29422 527258 36186 527494
rect 36422 527258 43186 527494
rect 43422 527258 50186 527494
rect 50422 527258 57186 527494
rect 57422 527258 64186 527494
rect 64422 527258 71186 527494
rect 71422 527258 78186 527494
rect 78422 527258 85186 527494
rect 85422 527258 92186 527494
rect 92422 527258 99186 527494
rect 99422 527258 106186 527494
rect 106422 527258 113186 527494
rect 113422 527258 120186 527494
rect 120422 527258 127186 527494
rect 127422 527258 134186 527494
rect 134422 527258 141186 527494
rect 141422 527258 148186 527494
rect 148422 527258 155186 527494
rect 155422 527258 162186 527494
rect 162422 527258 169186 527494
rect 169422 527258 176186 527494
rect 176422 527258 183186 527494
rect 183422 527258 190186 527494
rect 190422 527258 197186 527494
rect 197422 527258 204186 527494
rect 204422 527258 211186 527494
rect 211422 527258 218186 527494
rect 218422 527258 225186 527494
rect 225422 527258 232186 527494
rect 232422 527258 239186 527494
rect 239422 527258 246186 527494
rect 246422 527258 253186 527494
rect 253422 527258 260186 527494
rect 260422 527258 267186 527494
rect 267422 527258 274186 527494
rect 274422 527258 281186 527494
rect 281422 527258 288186 527494
rect 288422 527258 295186 527494
rect 295422 527258 302186 527494
rect 302422 527258 309186 527494
rect 309422 527258 316186 527494
rect 316422 527258 323186 527494
rect 323422 527258 330186 527494
rect 330422 527258 337186 527494
rect 337422 527258 344186 527494
rect 344422 527258 351186 527494
rect 351422 527258 358186 527494
rect 358422 527258 365186 527494
rect 365422 527258 372186 527494
rect 372422 527258 379186 527494
rect 379422 527258 386186 527494
rect 386422 527258 393186 527494
rect 393422 527258 400186 527494
rect 400422 527258 407186 527494
rect 407422 527258 414186 527494
rect 414422 527258 421186 527494
rect 421422 527258 428186 527494
rect 428422 527258 435186 527494
rect 435422 527258 442186 527494
rect 442422 527258 449186 527494
rect 449422 527258 456186 527494
rect 456422 527258 463186 527494
rect 463422 527258 470186 527494
rect 470422 527258 477186 527494
rect 477422 527258 484186 527494
rect 484422 527258 491186 527494
rect 491422 527258 498186 527494
rect 498422 527258 505186 527494
rect 505422 527258 512186 527494
rect 512422 527258 519186 527494
rect 519422 527258 526186 527494
rect 526422 527258 533186 527494
rect 533422 527258 540186 527494
rect 540422 527258 547186 527494
rect 547422 527258 554186 527494
rect 554422 527258 561186 527494
rect 561422 527258 568186 527494
rect 568422 527258 575186 527494
rect 575422 527258 582186 527494
rect 582422 527258 585818 527494
rect 586054 527258 586138 527494
rect 586374 527258 586458 527494
rect 586694 527258 586778 527494
rect 587014 527258 588874 527494
rect -4950 527216 588874 527258
rect -4950 521434 588874 521476
rect -4950 521198 -4842 521434
rect -4606 521198 -4522 521434
rect -4286 521198 -4202 521434
rect -3966 521198 -3882 521434
rect -3646 521198 2918 521434
rect 3154 521198 9918 521434
rect 10154 521198 16918 521434
rect 17154 521198 23918 521434
rect 24154 521198 30918 521434
rect 31154 521198 37918 521434
rect 38154 521198 44918 521434
rect 45154 521198 51918 521434
rect 52154 521198 58918 521434
rect 59154 521198 65918 521434
rect 66154 521198 72918 521434
rect 73154 521198 79918 521434
rect 80154 521198 86918 521434
rect 87154 521198 93918 521434
rect 94154 521198 100918 521434
rect 101154 521198 107918 521434
rect 108154 521198 114918 521434
rect 115154 521198 121918 521434
rect 122154 521198 128918 521434
rect 129154 521198 135918 521434
rect 136154 521198 142918 521434
rect 143154 521198 149918 521434
rect 150154 521198 156918 521434
rect 157154 521198 163918 521434
rect 164154 521198 170918 521434
rect 171154 521198 177918 521434
rect 178154 521198 184918 521434
rect 185154 521198 191918 521434
rect 192154 521198 198918 521434
rect 199154 521198 205918 521434
rect 206154 521198 212918 521434
rect 213154 521198 219918 521434
rect 220154 521198 226918 521434
rect 227154 521198 233918 521434
rect 234154 521198 240918 521434
rect 241154 521198 247918 521434
rect 248154 521198 254918 521434
rect 255154 521198 261918 521434
rect 262154 521198 268918 521434
rect 269154 521198 275918 521434
rect 276154 521198 282918 521434
rect 283154 521198 289918 521434
rect 290154 521198 296918 521434
rect 297154 521198 303918 521434
rect 304154 521198 310918 521434
rect 311154 521198 317918 521434
rect 318154 521198 324918 521434
rect 325154 521198 331918 521434
rect 332154 521198 338918 521434
rect 339154 521198 345918 521434
rect 346154 521198 352918 521434
rect 353154 521198 359918 521434
rect 360154 521198 366918 521434
rect 367154 521198 373918 521434
rect 374154 521198 380918 521434
rect 381154 521198 387918 521434
rect 388154 521198 394918 521434
rect 395154 521198 401918 521434
rect 402154 521198 408918 521434
rect 409154 521198 415918 521434
rect 416154 521198 422918 521434
rect 423154 521198 429918 521434
rect 430154 521198 436918 521434
rect 437154 521198 443918 521434
rect 444154 521198 450918 521434
rect 451154 521198 457918 521434
rect 458154 521198 464918 521434
rect 465154 521198 471918 521434
rect 472154 521198 478918 521434
rect 479154 521198 485918 521434
rect 486154 521198 492918 521434
rect 493154 521198 499918 521434
rect 500154 521198 506918 521434
rect 507154 521198 513918 521434
rect 514154 521198 520918 521434
rect 521154 521198 527918 521434
rect 528154 521198 534918 521434
rect 535154 521198 541918 521434
rect 542154 521198 548918 521434
rect 549154 521198 555918 521434
rect 556154 521198 562918 521434
rect 563154 521198 569918 521434
rect 570154 521198 576918 521434
rect 577154 521198 587570 521434
rect 587806 521198 587890 521434
rect 588126 521198 588210 521434
rect 588446 521198 588530 521434
rect 588766 521198 588874 521434
rect -4950 521156 588874 521198
rect -4950 520494 588874 520536
rect -4950 520258 -3090 520494
rect -2854 520258 -2770 520494
rect -2534 520258 -2450 520494
rect -2214 520258 -2130 520494
rect -1894 520258 1186 520494
rect 1422 520258 8186 520494
rect 8422 520258 15186 520494
rect 15422 520258 22186 520494
rect 22422 520258 29186 520494
rect 29422 520258 36186 520494
rect 36422 520258 43186 520494
rect 43422 520258 50186 520494
rect 50422 520258 57186 520494
rect 57422 520258 64186 520494
rect 64422 520258 71186 520494
rect 71422 520258 78186 520494
rect 78422 520258 85186 520494
rect 85422 520258 92186 520494
rect 92422 520258 99186 520494
rect 99422 520258 106186 520494
rect 106422 520258 113186 520494
rect 113422 520258 120186 520494
rect 120422 520258 127186 520494
rect 127422 520258 134186 520494
rect 134422 520258 141186 520494
rect 141422 520258 148186 520494
rect 148422 520258 155186 520494
rect 155422 520258 162186 520494
rect 162422 520258 169186 520494
rect 169422 520258 176186 520494
rect 176422 520258 183186 520494
rect 183422 520258 190186 520494
rect 190422 520258 197186 520494
rect 197422 520258 204186 520494
rect 204422 520258 211186 520494
rect 211422 520258 218186 520494
rect 218422 520258 225186 520494
rect 225422 520258 232186 520494
rect 232422 520258 239186 520494
rect 239422 520258 246186 520494
rect 246422 520258 253186 520494
rect 253422 520258 260186 520494
rect 260422 520258 267186 520494
rect 267422 520258 274186 520494
rect 274422 520258 281186 520494
rect 281422 520258 288186 520494
rect 288422 520258 295186 520494
rect 295422 520258 302186 520494
rect 302422 520258 309186 520494
rect 309422 520258 316186 520494
rect 316422 520258 323186 520494
rect 323422 520258 330186 520494
rect 330422 520258 337186 520494
rect 337422 520258 344186 520494
rect 344422 520258 351186 520494
rect 351422 520258 358186 520494
rect 358422 520258 365186 520494
rect 365422 520258 372186 520494
rect 372422 520258 379186 520494
rect 379422 520258 386186 520494
rect 386422 520258 393186 520494
rect 393422 520258 400186 520494
rect 400422 520258 407186 520494
rect 407422 520258 414186 520494
rect 414422 520258 421186 520494
rect 421422 520258 428186 520494
rect 428422 520258 435186 520494
rect 435422 520258 442186 520494
rect 442422 520258 449186 520494
rect 449422 520258 456186 520494
rect 456422 520258 463186 520494
rect 463422 520258 470186 520494
rect 470422 520258 477186 520494
rect 477422 520258 484186 520494
rect 484422 520258 491186 520494
rect 491422 520258 498186 520494
rect 498422 520258 505186 520494
rect 505422 520258 512186 520494
rect 512422 520258 519186 520494
rect 519422 520258 526186 520494
rect 526422 520258 533186 520494
rect 533422 520258 540186 520494
rect 540422 520258 547186 520494
rect 547422 520258 554186 520494
rect 554422 520258 561186 520494
rect 561422 520258 568186 520494
rect 568422 520258 575186 520494
rect 575422 520258 582186 520494
rect 582422 520258 585818 520494
rect 586054 520258 586138 520494
rect 586374 520258 586458 520494
rect 586694 520258 586778 520494
rect 587014 520258 588874 520494
rect -4950 520216 588874 520258
rect -4950 514434 588874 514476
rect -4950 514198 -4842 514434
rect -4606 514198 -4522 514434
rect -4286 514198 -4202 514434
rect -3966 514198 -3882 514434
rect -3646 514198 2918 514434
rect 3154 514198 9918 514434
rect 10154 514198 16918 514434
rect 17154 514198 23918 514434
rect 24154 514198 30918 514434
rect 31154 514198 37918 514434
rect 38154 514198 44918 514434
rect 45154 514198 51918 514434
rect 52154 514198 58918 514434
rect 59154 514198 65918 514434
rect 66154 514198 72918 514434
rect 73154 514198 79918 514434
rect 80154 514198 86918 514434
rect 87154 514198 93918 514434
rect 94154 514198 100918 514434
rect 101154 514198 107918 514434
rect 108154 514198 114918 514434
rect 115154 514198 121918 514434
rect 122154 514198 128918 514434
rect 129154 514198 135918 514434
rect 136154 514198 142918 514434
rect 143154 514198 149918 514434
rect 150154 514198 156918 514434
rect 157154 514198 163918 514434
rect 164154 514198 170918 514434
rect 171154 514198 177918 514434
rect 178154 514198 184918 514434
rect 185154 514198 191918 514434
rect 192154 514198 198918 514434
rect 199154 514198 205918 514434
rect 206154 514198 212918 514434
rect 213154 514198 219918 514434
rect 220154 514198 226918 514434
rect 227154 514198 233918 514434
rect 234154 514198 240918 514434
rect 241154 514198 247918 514434
rect 248154 514198 254918 514434
rect 255154 514198 261918 514434
rect 262154 514198 268918 514434
rect 269154 514198 275918 514434
rect 276154 514198 282918 514434
rect 283154 514198 289918 514434
rect 290154 514198 296918 514434
rect 297154 514198 303918 514434
rect 304154 514198 310918 514434
rect 311154 514198 317918 514434
rect 318154 514198 324918 514434
rect 325154 514198 331918 514434
rect 332154 514198 338918 514434
rect 339154 514198 345918 514434
rect 346154 514198 352918 514434
rect 353154 514198 359918 514434
rect 360154 514198 366918 514434
rect 367154 514198 373918 514434
rect 374154 514198 380918 514434
rect 381154 514198 387918 514434
rect 388154 514198 394918 514434
rect 395154 514198 401918 514434
rect 402154 514198 408918 514434
rect 409154 514198 415918 514434
rect 416154 514198 422918 514434
rect 423154 514198 429918 514434
rect 430154 514198 436918 514434
rect 437154 514198 443918 514434
rect 444154 514198 450918 514434
rect 451154 514198 457918 514434
rect 458154 514198 464918 514434
rect 465154 514198 471918 514434
rect 472154 514198 478918 514434
rect 479154 514198 485918 514434
rect 486154 514198 492918 514434
rect 493154 514198 499918 514434
rect 500154 514198 506918 514434
rect 507154 514198 513918 514434
rect 514154 514198 520918 514434
rect 521154 514198 527918 514434
rect 528154 514198 534918 514434
rect 535154 514198 541918 514434
rect 542154 514198 548918 514434
rect 549154 514198 555918 514434
rect 556154 514198 562918 514434
rect 563154 514198 569918 514434
rect 570154 514198 576918 514434
rect 577154 514198 587570 514434
rect 587806 514198 587890 514434
rect 588126 514198 588210 514434
rect 588446 514198 588530 514434
rect 588766 514198 588874 514434
rect -4950 514156 588874 514198
rect -4950 513494 588874 513536
rect -4950 513258 -3090 513494
rect -2854 513258 -2770 513494
rect -2534 513258 -2450 513494
rect -2214 513258 -2130 513494
rect -1894 513258 1186 513494
rect 1422 513258 8186 513494
rect 8422 513258 15186 513494
rect 15422 513258 22186 513494
rect 22422 513258 29186 513494
rect 29422 513258 36186 513494
rect 36422 513258 43186 513494
rect 43422 513258 50186 513494
rect 50422 513258 57186 513494
rect 57422 513258 64186 513494
rect 64422 513258 71186 513494
rect 71422 513258 78186 513494
rect 78422 513258 85186 513494
rect 85422 513258 92186 513494
rect 92422 513258 99186 513494
rect 99422 513258 106186 513494
rect 106422 513258 113186 513494
rect 113422 513258 120186 513494
rect 120422 513258 127186 513494
rect 127422 513258 134186 513494
rect 134422 513258 141186 513494
rect 141422 513258 148186 513494
rect 148422 513258 155186 513494
rect 155422 513258 162186 513494
rect 162422 513258 169186 513494
rect 169422 513258 176186 513494
rect 176422 513258 183186 513494
rect 183422 513258 190186 513494
rect 190422 513258 197186 513494
rect 197422 513258 204186 513494
rect 204422 513258 211186 513494
rect 211422 513258 218186 513494
rect 218422 513258 225186 513494
rect 225422 513258 232186 513494
rect 232422 513258 239186 513494
rect 239422 513258 246186 513494
rect 246422 513258 253186 513494
rect 253422 513258 260186 513494
rect 260422 513258 267186 513494
rect 267422 513258 274186 513494
rect 274422 513258 281186 513494
rect 281422 513258 288186 513494
rect 288422 513258 295186 513494
rect 295422 513258 302186 513494
rect 302422 513258 309186 513494
rect 309422 513258 316186 513494
rect 316422 513258 323186 513494
rect 323422 513258 330186 513494
rect 330422 513258 337186 513494
rect 337422 513258 344186 513494
rect 344422 513258 351186 513494
rect 351422 513258 358186 513494
rect 358422 513258 365186 513494
rect 365422 513258 372186 513494
rect 372422 513258 379186 513494
rect 379422 513258 386186 513494
rect 386422 513258 393186 513494
rect 393422 513258 400186 513494
rect 400422 513258 407186 513494
rect 407422 513258 414186 513494
rect 414422 513258 421186 513494
rect 421422 513258 428186 513494
rect 428422 513258 435186 513494
rect 435422 513258 442186 513494
rect 442422 513258 449186 513494
rect 449422 513258 456186 513494
rect 456422 513258 463186 513494
rect 463422 513258 470186 513494
rect 470422 513258 477186 513494
rect 477422 513258 484186 513494
rect 484422 513258 491186 513494
rect 491422 513258 498186 513494
rect 498422 513258 505186 513494
rect 505422 513258 512186 513494
rect 512422 513258 519186 513494
rect 519422 513258 526186 513494
rect 526422 513258 533186 513494
rect 533422 513258 540186 513494
rect 540422 513258 547186 513494
rect 547422 513258 554186 513494
rect 554422 513258 561186 513494
rect 561422 513258 568186 513494
rect 568422 513258 575186 513494
rect 575422 513258 582186 513494
rect 582422 513258 585818 513494
rect 586054 513258 586138 513494
rect 586374 513258 586458 513494
rect 586694 513258 586778 513494
rect 587014 513258 588874 513494
rect -4950 513216 588874 513258
rect -4950 507434 588874 507476
rect -4950 507198 -4842 507434
rect -4606 507198 -4522 507434
rect -4286 507198 -4202 507434
rect -3966 507198 -3882 507434
rect -3646 507198 2918 507434
rect 3154 507198 9918 507434
rect 10154 507198 16918 507434
rect 17154 507198 23918 507434
rect 24154 507198 30918 507434
rect 31154 507198 37918 507434
rect 38154 507198 44918 507434
rect 45154 507198 51918 507434
rect 52154 507198 58918 507434
rect 59154 507198 65918 507434
rect 66154 507198 72918 507434
rect 73154 507198 79918 507434
rect 80154 507198 86918 507434
rect 87154 507198 93918 507434
rect 94154 507198 100918 507434
rect 101154 507198 107918 507434
rect 108154 507198 114918 507434
rect 115154 507198 121918 507434
rect 122154 507198 128918 507434
rect 129154 507198 135918 507434
rect 136154 507198 142918 507434
rect 143154 507198 149918 507434
rect 150154 507198 156918 507434
rect 157154 507198 163918 507434
rect 164154 507198 170918 507434
rect 171154 507198 177918 507434
rect 178154 507198 184918 507434
rect 185154 507198 191918 507434
rect 192154 507198 198918 507434
rect 199154 507198 205918 507434
rect 206154 507198 212918 507434
rect 213154 507198 219918 507434
rect 220154 507198 226918 507434
rect 227154 507198 233918 507434
rect 234154 507198 240918 507434
rect 241154 507198 247918 507434
rect 248154 507198 254918 507434
rect 255154 507198 261918 507434
rect 262154 507198 268918 507434
rect 269154 507198 275918 507434
rect 276154 507198 282918 507434
rect 283154 507198 289918 507434
rect 290154 507198 296918 507434
rect 297154 507198 303918 507434
rect 304154 507198 310918 507434
rect 311154 507198 317918 507434
rect 318154 507198 324918 507434
rect 325154 507198 331918 507434
rect 332154 507198 338918 507434
rect 339154 507198 345918 507434
rect 346154 507198 352918 507434
rect 353154 507198 359918 507434
rect 360154 507198 366918 507434
rect 367154 507198 373918 507434
rect 374154 507198 380918 507434
rect 381154 507198 387918 507434
rect 388154 507198 394918 507434
rect 395154 507198 401918 507434
rect 402154 507198 408918 507434
rect 409154 507198 415918 507434
rect 416154 507198 422918 507434
rect 423154 507198 429918 507434
rect 430154 507198 436918 507434
rect 437154 507198 443918 507434
rect 444154 507198 450918 507434
rect 451154 507198 457918 507434
rect 458154 507198 464918 507434
rect 465154 507198 471918 507434
rect 472154 507198 478918 507434
rect 479154 507198 485918 507434
rect 486154 507198 492918 507434
rect 493154 507198 499918 507434
rect 500154 507198 506918 507434
rect 507154 507198 513918 507434
rect 514154 507198 520918 507434
rect 521154 507198 527918 507434
rect 528154 507198 534918 507434
rect 535154 507198 541918 507434
rect 542154 507198 548918 507434
rect 549154 507198 555918 507434
rect 556154 507198 562918 507434
rect 563154 507198 569918 507434
rect 570154 507198 576918 507434
rect 577154 507198 587570 507434
rect 587806 507198 587890 507434
rect 588126 507198 588210 507434
rect 588446 507198 588530 507434
rect 588766 507198 588874 507434
rect -4950 507156 588874 507198
rect -4950 506494 588874 506536
rect -4950 506258 -3090 506494
rect -2854 506258 -2770 506494
rect -2534 506258 -2450 506494
rect -2214 506258 -2130 506494
rect -1894 506258 1186 506494
rect 1422 506258 8186 506494
rect 8422 506258 15186 506494
rect 15422 506258 22186 506494
rect 22422 506258 29186 506494
rect 29422 506258 36186 506494
rect 36422 506258 43186 506494
rect 43422 506258 50186 506494
rect 50422 506258 57186 506494
rect 57422 506258 64186 506494
rect 64422 506258 71186 506494
rect 71422 506258 78186 506494
rect 78422 506258 85186 506494
rect 85422 506258 92186 506494
rect 92422 506258 99186 506494
rect 99422 506258 106186 506494
rect 106422 506258 113186 506494
rect 113422 506258 120186 506494
rect 120422 506258 127186 506494
rect 127422 506258 134186 506494
rect 134422 506258 141186 506494
rect 141422 506258 148186 506494
rect 148422 506258 155186 506494
rect 155422 506258 162186 506494
rect 162422 506258 169186 506494
rect 169422 506258 176186 506494
rect 176422 506258 183186 506494
rect 183422 506258 190186 506494
rect 190422 506258 197186 506494
rect 197422 506258 204186 506494
rect 204422 506258 211186 506494
rect 211422 506258 218186 506494
rect 218422 506258 225186 506494
rect 225422 506258 232186 506494
rect 232422 506258 239186 506494
rect 239422 506258 246186 506494
rect 246422 506258 253186 506494
rect 253422 506258 260186 506494
rect 260422 506258 267186 506494
rect 267422 506258 274186 506494
rect 274422 506258 281186 506494
rect 281422 506258 288186 506494
rect 288422 506258 295186 506494
rect 295422 506258 302186 506494
rect 302422 506258 309186 506494
rect 309422 506258 316186 506494
rect 316422 506258 323186 506494
rect 323422 506258 330186 506494
rect 330422 506258 337186 506494
rect 337422 506258 344186 506494
rect 344422 506258 351186 506494
rect 351422 506258 358186 506494
rect 358422 506258 365186 506494
rect 365422 506258 372186 506494
rect 372422 506258 379186 506494
rect 379422 506258 386186 506494
rect 386422 506258 393186 506494
rect 393422 506258 400186 506494
rect 400422 506258 407186 506494
rect 407422 506258 414186 506494
rect 414422 506258 421186 506494
rect 421422 506258 428186 506494
rect 428422 506258 435186 506494
rect 435422 506258 442186 506494
rect 442422 506258 449186 506494
rect 449422 506258 456186 506494
rect 456422 506258 463186 506494
rect 463422 506258 470186 506494
rect 470422 506258 477186 506494
rect 477422 506258 484186 506494
rect 484422 506258 491186 506494
rect 491422 506258 498186 506494
rect 498422 506258 505186 506494
rect 505422 506258 512186 506494
rect 512422 506258 519186 506494
rect 519422 506258 526186 506494
rect 526422 506258 533186 506494
rect 533422 506258 540186 506494
rect 540422 506258 547186 506494
rect 547422 506258 554186 506494
rect 554422 506258 561186 506494
rect 561422 506258 568186 506494
rect 568422 506258 575186 506494
rect 575422 506258 582186 506494
rect 582422 506258 585818 506494
rect 586054 506258 586138 506494
rect 586374 506258 586458 506494
rect 586694 506258 586778 506494
rect 587014 506258 588874 506494
rect -4950 506216 588874 506258
rect -4950 500434 588874 500476
rect -4950 500198 -4842 500434
rect -4606 500198 -4522 500434
rect -4286 500198 -4202 500434
rect -3966 500198 -3882 500434
rect -3646 500198 2918 500434
rect 3154 500198 9918 500434
rect 10154 500198 16918 500434
rect 17154 500198 23918 500434
rect 24154 500198 30918 500434
rect 31154 500198 37918 500434
rect 38154 500198 44918 500434
rect 45154 500198 51918 500434
rect 52154 500198 58918 500434
rect 59154 500198 65918 500434
rect 66154 500198 72918 500434
rect 73154 500198 79918 500434
rect 80154 500198 86918 500434
rect 87154 500198 93918 500434
rect 94154 500198 100918 500434
rect 101154 500198 107918 500434
rect 108154 500198 114918 500434
rect 115154 500198 121918 500434
rect 122154 500198 128918 500434
rect 129154 500198 135918 500434
rect 136154 500198 142918 500434
rect 143154 500198 149918 500434
rect 150154 500198 156918 500434
rect 157154 500198 163918 500434
rect 164154 500198 170918 500434
rect 171154 500198 177918 500434
rect 178154 500198 184918 500434
rect 185154 500198 191918 500434
rect 192154 500198 198918 500434
rect 199154 500198 205918 500434
rect 206154 500198 212918 500434
rect 213154 500198 219918 500434
rect 220154 500198 226918 500434
rect 227154 500198 233918 500434
rect 234154 500198 240918 500434
rect 241154 500198 247918 500434
rect 248154 500198 254918 500434
rect 255154 500198 261918 500434
rect 262154 500198 268918 500434
rect 269154 500198 275918 500434
rect 276154 500198 282918 500434
rect 283154 500198 289918 500434
rect 290154 500198 296918 500434
rect 297154 500198 303918 500434
rect 304154 500198 310918 500434
rect 311154 500198 317918 500434
rect 318154 500198 324918 500434
rect 325154 500198 331918 500434
rect 332154 500198 338918 500434
rect 339154 500198 345918 500434
rect 346154 500198 352918 500434
rect 353154 500198 359918 500434
rect 360154 500198 366918 500434
rect 367154 500198 373918 500434
rect 374154 500198 380918 500434
rect 381154 500198 387918 500434
rect 388154 500198 394918 500434
rect 395154 500198 401918 500434
rect 402154 500198 408918 500434
rect 409154 500198 415918 500434
rect 416154 500198 422918 500434
rect 423154 500198 429918 500434
rect 430154 500198 436918 500434
rect 437154 500198 443918 500434
rect 444154 500198 450918 500434
rect 451154 500198 457918 500434
rect 458154 500198 464918 500434
rect 465154 500198 471918 500434
rect 472154 500198 478918 500434
rect 479154 500198 485918 500434
rect 486154 500198 492918 500434
rect 493154 500198 499918 500434
rect 500154 500198 506918 500434
rect 507154 500198 513918 500434
rect 514154 500198 520918 500434
rect 521154 500198 527918 500434
rect 528154 500198 534918 500434
rect 535154 500198 541918 500434
rect 542154 500198 548918 500434
rect 549154 500198 555918 500434
rect 556154 500198 562918 500434
rect 563154 500198 569918 500434
rect 570154 500198 576918 500434
rect 577154 500198 587570 500434
rect 587806 500198 587890 500434
rect 588126 500198 588210 500434
rect 588446 500198 588530 500434
rect 588766 500198 588874 500434
rect -4950 500156 588874 500198
rect -4950 499494 588874 499536
rect -4950 499258 -3090 499494
rect -2854 499258 -2770 499494
rect -2534 499258 -2450 499494
rect -2214 499258 -2130 499494
rect -1894 499258 1186 499494
rect 1422 499258 8186 499494
rect 8422 499258 15186 499494
rect 15422 499258 22186 499494
rect 22422 499258 29186 499494
rect 29422 499258 36186 499494
rect 36422 499258 43186 499494
rect 43422 499258 50186 499494
rect 50422 499258 57186 499494
rect 57422 499258 64186 499494
rect 64422 499258 71186 499494
rect 71422 499258 78186 499494
rect 78422 499258 85186 499494
rect 85422 499258 92186 499494
rect 92422 499258 99186 499494
rect 99422 499258 106186 499494
rect 106422 499258 113186 499494
rect 113422 499258 120186 499494
rect 120422 499258 127186 499494
rect 127422 499258 134186 499494
rect 134422 499258 141186 499494
rect 141422 499258 148186 499494
rect 148422 499258 155186 499494
rect 155422 499258 162186 499494
rect 162422 499258 169186 499494
rect 169422 499258 176186 499494
rect 176422 499258 183186 499494
rect 183422 499258 190186 499494
rect 190422 499258 197186 499494
rect 197422 499258 204186 499494
rect 204422 499258 211186 499494
rect 211422 499258 218186 499494
rect 218422 499258 225186 499494
rect 225422 499258 232186 499494
rect 232422 499258 239186 499494
rect 239422 499258 246186 499494
rect 246422 499258 253186 499494
rect 253422 499258 260186 499494
rect 260422 499258 267186 499494
rect 267422 499258 274186 499494
rect 274422 499258 281186 499494
rect 281422 499258 288186 499494
rect 288422 499258 295186 499494
rect 295422 499258 302186 499494
rect 302422 499258 309186 499494
rect 309422 499258 316186 499494
rect 316422 499258 323186 499494
rect 323422 499258 330186 499494
rect 330422 499258 337186 499494
rect 337422 499258 344186 499494
rect 344422 499258 351186 499494
rect 351422 499258 358186 499494
rect 358422 499258 365186 499494
rect 365422 499258 372186 499494
rect 372422 499258 379186 499494
rect 379422 499258 386186 499494
rect 386422 499258 393186 499494
rect 393422 499258 400186 499494
rect 400422 499258 407186 499494
rect 407422 499258 414186 499494
rect 414422 499258 421186 499494
rect 421422 499258 428186 499494
rect 428422 499258 435186 499494
rect 435422 499258 442186 499494
rect 442422 499258 449186 499494
rect 449422 499258 456186 499494
rect 456422 499258 463186 499494
rect 463422 499258 470186 499494
rect 470422 499258 477186 499494
rect 477422 499258 484186 499494
rect 484422 499258 491186 499494
rect 491422 499258 498186 499494
rect 498422 499258 505186 499494
rect 505422 499258 512186 499494
rect 512422 499258 519186 499494
rect 519422 499258 526186 499494
rect 526422 499258 533186 499494
rect 533422 499258 540186 499494
rect 540422 499258 547186 499494
rect 547422 499258 554186 499494
rect 554422 499258 561186 499494
rect 561422 499258 568186 499494
rect 568422 499258 575186 499494
rect 575422 499258 582186 499494
rect 582422 499258 585818 499494
rect 586054 499258 586138 499494
rect 586374 499258 586458 499494
rect 586694 499258 586778 499494
rect 587014 499258 588874 499494
rect -4950 499216 588874 499258
rect -4950 493434 588874 493476
rect -4950 493198 -4842 493434
rect -4606 493198 -4522 493434
rect -4286 493198 -4202 493434
rect -3966 493198 -3882 493434
rect -3646 493198 2918 493434
rect 3154 493198 9918 493434
rect 10154 493198 16918 493434
rect 17154 493198 23918 493434
rect 24154 493198 30918 493434
rect 31154 493198 37918 493434
rect 38154 493198 44918 493434
rect 45154 493198 51918 493434
rect 52154 493198 58918 493434
rect 59154 493198 65918 493434
rect 66154 493198 72918 493434
rect 73154 493198 79918 493434
rect 80154 493198 86918 493434
rect 87154 493198 93918 493434
rect 94154 493198 100918 493434
rect 101154 493198 107918 493434
rect 108154 493198 114918 493434
rect 115154 493198 121918 493434
rect 122154 493198 128918 493434
rect 129154 493198 135918 493434
rect 136154 493198 142918 493434
rect 143154 493198 149918 493434
rect 150154 493198 156918 493434
rect 157154 493198 163918 493434
rect 164154 493198 170918 493434
rect 171154 493198 177918 493434
rect 178154 493198 184918 493434
rect 185154 493198 191918 493434
rect 192154 493198 198918 493434
rect 199154 493198 205918 493434
rect 206154 493198 212918 493434
rect 213154 493198 219918 493434
rect 220154 493198 226918 493434
rect 227154 493198 233918 493434
rect 234154 493198 240918 493434
rect 241154 493198 247918 493434
rect 248154 493198 254918 493434
rect 255154 493198 261918 493434
rect 262154 493198 268918 493434
rect 269154 493198 275918 493434
rect 276154 493198 282918 493434
rect 283154 493198 289918 493434
rect 290154 493198 296918 493434
rect 297154 493198 303918 493434
rect 304154 493198 310918 493434
rect 311154 493198 317918 493434
rect 318154 493198 324918 493434
rect 325154 493198 331918 493434
rect 332154 493198 338918 493434
rect 339154 493198 345918 493434
rect 346154 493198 352918 493434
rect 353154 493198 359918 493434
rect 360154 493198 366918 493434
rect 367154 493198 373918 493434
rect 374154 493198 380918 493434
rect 381154 493198 387918 493434
rect 388154 493198 394918 493434
rect 395154 493198 401918 493434
rect 402154 493198 408918 493434
rect 409154 493198 415918 493434
rect 416154 493198 422918 493434
rect 423154 493198 429918 493434
rect 430154 493198 436918 493434
rect 437154 493198 443918 493434
rect 444154 493198 450918 493434
rect 451154 493198 457918 493434
rect 458154 493198 464918 493434
rect 465154 493198 471918 493434
rect 472154 493198 478918 493434
rect 479154 493198 485918 493434
rect 486154 493198 492918 493434
rect 493154 493198 499918 493434
rect 500154 493198 506918 493434
rect 507154 493198 513918 493434
rect 514154 493198 520918 493434
rect 521154 493198 527918 493434
rect 528154 493198 534918 493434
rect 535154 493198 541918 493434
rect 542154 493198 548918 493434
rect 549154 493198 555918 493434
rect 556154 493198 562918 493434
rect 563154 493198 569918 493434
rect 570154 493198 576918 493434
rect 577154 493198 587570 493434
rect 587806 493198 587890 493434
rect 588126 493198 588210 493434
rect 588446 493198 588530 493434
rect 588766 493198 588874 493434
rect -4950 493156 588874 493198
rect -4950 492494 588874 492536
rect -4950 492258 -3090 492494
rect -2854 492258 -2770 492494
rect -2534 492258 -2450 492494
rect -2214 492258 -2130 492494
rect -1894 492258 1186 492494
rect 1422 492258 8186 492494
rect 8422 492258 15186 492494
rect 15422 492258 22186 492494
rect 22422 492258 29186 492494
rect 29422 492258 36186 492494
rect 36422 492258 43186 492494
rect 43422 492258 50186 492494
rect 50422 492258 57186 492494
rect 57422 492258 64186 492494
rect 64422 492258 71186 492494
rect 71422 492258 78186 492494
rect 78422 492258 85186 492494
rect 85422 492258 92186 492494
rect 92422 492258 99186 492494
rect 99422 492258 106186 492494
rect 106422 492258 113186 492494
rect 113422 492258 120186 492494
rect 120422 492258 127186 492494
rect 127422 492258 134186 492494
rect 134422 492258 141186 492494
rect 141422 492258 148186 492494
rect 148422 492258 155186 492494
rect 155422 492258 162186 492494
rect 162422 492258 169186 492494
rect 169422 492258 176186 492494
rect 176422 492258 183186 492494
rect 183422 492258 190186 492494
rect 190422 492258 197186 492494
rect 197422 492258 204186 492494
rect 204422 492258 211186 492494
rect 211422 492258 218186 492494
rect 218422 492258 225186 492494
rect 225422 492258 232186 492494
rect 232422 492258 239186 492494
rect 239422 492258 246186 492494
rect 246422 492258 253186 492494
rect 253422 492258 260186 492494
rect 260422 492258 267186 492494
rect 267422 492258 274186 492494
rect 274422 492258 281186 492494
rect 281422 492258 288186 492494
rect 288422 492258 295186 492494
rect 295422 492258 302186 492494
rect 302422 492258 309186 492494
rect 309422 492258 316186 492494
rect 316422 492258 323186 492494
rect 323422 492258 330186 492494
rect 330422 492258 337186 492494
rect 337422 492258 344186 492494
rect 344422 492258 351186 492494
rect 351422 492258 358186 492494
rect 358422 492258 365186 492494
rect 365422 492258 372186 492494
rect 372422 492258 379186 492494
rect 379422 492258 386186 492494
rect 386422 492258 393186 492494
rect 393422 492258 400186 492494
rect 400422 492258 407186 492494
rect 407422 492258 414186 492494
rect 414422 492258 421186 492494
rect 421422 492258 428186 492494
rect 428422 492258 435186 492494
rect 435422 492258 442186 492494
rect 442422 492258 449186 492494
rect 449422 492258 456186 492494
rect 456422 492258 463186 492494
rect 463422 492258 470186 492494
rect 470422 492258 477186 492494
rect 477422 492258 484186 492494
rect 484422 492258 491186 492494
rect 491422 492258 498186 492494
rect 498422 492258 505186 492494
rect 505422 492258 512186 492494
rect 512422 492258 519186 492494
rect 519422 492258 526186 492494
rect 526422 492258 533186 492494
rect 533422 492258 540186 492494
rect 540422 492258 547186 492494
rect 547422 492258 554186 492494
rect 554422 492258 561186 492494
rect 561422 492258 568186 492494
rect 568422 492258 575186 492494
rect 575422 492258 582186 492494
rect 582422 492258 585818 492494
rect 586054 492258 586138 492494
rect 586374 492258 586458 492494
rect 586694 492258 586778 492494
rect 587014 492258 588874 492494
rect -4950 492216 588874 492258
rect -4950 486434 588874 486476
rect -4950 486198 -4842 486434
rect -4606 486198 -4522 486434
rect -4286 486198 -4202 486434
rect -3966 486198 -3882 486434
rect -3646 486198 2918 486434
rect 3154 486198 9918 486434
rect 10154 486198 16918 486434
rect 17154 486198 23918 486434
rect 24154 486198 30918 486434
rect 31154 486198 37918 486434
rect 38154 486198 44918 486434
rect 45154 486198 51918 486434
rect 52154 486198 58918 486434
rect 59154 486198 65918 486434
rect 66154 486198 72918 486434
rect 73154 486198 79918 486434
rect 80154 486198 86918 486434
rect 87154 486198 93918 486434
rect 94154 486198 100918 486434
rect 101154 486198 107918 486434
rect 108154 486198 114918 486434
rect 115154 486198 121918 486434
rect 122154 486198 128918 486434
rect 129154 486198 135918 486434
rect 136154 486198 142918 486434
rect 143154 486198 149918 486434
rect 150154 486198 156918 486434
rect 157154 486198 163918 486434
rect 164154 486198 170918 486434
rect 171154 486198 177918 486434
rect 178154 486198 184918 486434
rect 185154 486198 191918 486434
rect 192154 486198 198918 486434
rect 199154 486198 205918 486434
rect 206154 486198 212918 486434
rect 213154 486198 219918 486434
rect 220154 486198 226918 486434
rect 227154 486198 233918 486434
rect 234154 486198 240918 486434
rect 241154 486198 247918 486434
rect 248154 486198 254918 486434
rect 255154 486198 261918 486434
rect 262154 486198 268918 486434
rect 269154 486198 275918 486434
rect 276154 486198 282918 486434
rect 283154 486198 289918 486434
rect 290154 486198 296918 486434
rect 297154 486198 303918 486434
rect 304154 486198 310918 486434
rect 311154 486198 317918 486434
rect 318154 486198 324918 486434
rect 325154 486198 331918 486434
rect 332154 486198 338918 486434
rect 339154 486198 345918 486434
rect 346154 486198 352918 486434
rect 353154 486198 359918 486434
rect 360154 486198 366918 486434
rect 367154 486198 373918 486434
rect 374154 486198 380918 486434
rect 381154 486198 387918 486434
rect 388154 486198 394918 486434
rect 395154 486198 401918 486434
rect 402154 486198 408918 486434
rect 409154 486198 415918 486434
rect 416154 486198 422918 486434
rect 423154 486198 429918 486434
rect 430154 486198 436918 486434
rect 437154 486198 443918 486434
rect 444154 486198 450918 486434
rect 451154 486198 457918 486434
rect 458154 486198 464918 486434
rect 465154 486198 471918 486434
rect 472154 486198 478918 486434
rect 479154 486198 485918 486434
rect 486154 486198 492918 486434
rect 493154 486198 499918 486434
rect 500154 486198 506918 486434
rect 507154 486198 513918 486434
rect 514154 486198 520918 486434
rect 521154 486198 527918 486434
rect 528154 486198 534918 486434
rect 535154 486198 541918 486434
rect 542154 486198 548918 486434
rect 549154 486198 555918 486434
rect 556154 486198 562918 486434
rect 563154 486198 569918 486434
rect 570154 486198 576918 486434
rect 577154 486198 587570 486434
rect 587806 486198 587890 486434
rect 588126 486198 588210 486434
rect 588446 486198 588530 486434
rect 588766 486198 588874 486434
rect -4950 486156 588874 486198
rect -4950 485494 588874 485536
rect -4950 485258 -3090 485494
rect -2854 485258 -2770 485494
rect -2534 485258 -2450 485494
rect -2214 485258 -2130 485494
rect -1894 485258 1186 485494
rect 1422 485258 8186 485494
rect 8422 485258 15186 485494
rect 15422 485258 22186 485494
rect 22422 485258 29186 485494
rect 29422 485258 36186 485494
rect 36422 485258 43186 485494
rect 43422 485258 50186 485494
rect 50422 485258 57186 485494
rect 57422 485258 64186 485494
rect 64422 485258 71186 485494
rect 71422 485258 78186 485494
rect 78422 485258 85186 485494
rect 85422 485258 92186 485494
rect 92422 485258 99186 485494
rect 99422 485258 106186 485494
rect 106422 485258 113186 485494
rect 113422 485258 120186 485494
rect 120422 485258 127186 485494
rect 127422 485258 134186 485494
rect 134422 485258 141186 485494
rect 141422 485258 148186 485494
rect 148422 485258 155186 485494
rect 155422 485258 162186 485494
rect 162422 485258 169186 485494
rect 169422 485258 176186 485494
rect 176422 485258 183186 485494
rect 183422 485258 190186 485494
rect 190422 485258 197186 485494
rect 197422 485258 204186 485494
rect 204422 485258 211186 485494
rect 211422 485258 218186 485494
rect 218422 485258 225186 485494
rect 225422 485258 232186 485494
rect 232422 485258 239186 485494
rect 239422 485258 246186 485494
rect 246422 485258 253186 485494
rect 253422 485258 260186 485494
rect 260422 485258 267186 485494
rect 267422 485258 274186 485494
rect 274422 485258 281186 485494
rect 281422 485258 288186 485494
rect 288422 485258 295186 485494
rect 295422 485258 302186 485494
rect 302422 485258 309186 485494
rect 309422 485258 316186 485494
rect 316422 485258 323186 485494
rect 323422 485258 330186 485494
rect 330422 485258 337186 485494
rect 337422 485258 344186 485494
rect 344422 485258 351186 485494
rect 351422 485258 358186 485494
rect 358422 485258 365186 485494
rect 365422 485258 372186 485494
rect 372422 485258 379186 485494
rect 379422 485258 386186 485494
rect 386422 485258 393186 485494
rect 393422 485258 400186 485494
rect 400422 485258 407186 485494
rect 407422 485258 414186 485494
rect 414422 485258 421186 485494
rect 421422 485258 428186 485494
rect 428422 485258 435186 485494
rect 435422 485258 442186 485494
rect 442422 485258 449186 485494
rect 449422 485258 456186 485494
rect 456422 485258 463186 485494
rect 463422 485258 470186 485494
rect 470422 485258 477186 485494
rect 477422 485258 484186 485494
rect 484422 485258 491186 485494
rect 491422 485258 498186 485494
rect 498422 485258 505186 485494
rect 505422 485258 512186 485494
rect 512422 485258 519186 485494
rect 519422 485258 526186 485494
rect 526422 485258 533186 485494
rect 533422 485258 540186 485494
rect 540422 485258 547186 485494
rect 547422 485258 554186 485494
rect 554422 485258 561186 485494
rect 561422 485258 568186 485494
rect 568422 485258 575186 485494
rect 575422 485258 582186 485494
rect 582422 485258 585818 485494
rect 586054 485258 586138 485494
rect 586374 485258 586458 485494
rect 586694 485258 586778 485494
rect 587014 485258 588874 485494
rect -4950 485216 588874 485258
rect -4950 479434 588874 479476
rect -4950 479198 -4842 479434
rect -4606 479198 -4522 479434
rect -4286 479198 -4202 479434
rect -3966 479198 -3882 479434
rect -3646 479198 2918 479434
rect 3154 479198 9918 479434
rect 10154 479198 16918 479434
rect 17154 479198 23918 479434
rect 24154 479198 30918 479434
rect 31154 479198 37918 479434
rect 38154 479198 44918 479434
rect 45154 479198 51918 479434
rect 52154 479198 58918 479434
rect 59154 479198 65918 479434
rect 66154 479198 72918 479434
rect 73154 479198 79918 479434
rect 80154 479198 86918 479434
rect 87154 479198 93918 479434
rect 94154 479198 100918 479434
rect 101154 479198 107918 479434
rect 108154 479198 114918 479434
rect 115154 479198 121918 479434
rect 122154 479198 128918 479434
rect 129154 479198 135918 479434
rect 136154 479198 142918 479434
rect 143154 479198 149918 479434
rect 150154 479198 156918 479434
rect 157154 479198 163918 479434
rect 164154 479198 170918 479434
rect 171154 479198 177918 479434
rect 178154 479198 184918 479434
rect 185154 479198 191918 479434
rect 192154 479198 198918 479434
rect 199154 479198 205918 479434
rect 206154 479198 212918 479434
rect 213154 479198 219918 479434
rect 220154 479198 226918 479434
rect 227154 479198 233918 479434
rect 234154 479198 240918 479434
rect 241154 479198 247918 479434
rect 248154 479198 254918 479434
rect 255154 479198 261918 479434
rect 262154 479198 268918 479434
rect 269154 479198 275918 479434
rect 276154 479198 282918 479434
rect 283154 479198 289918 479434
rect 290154 479198 296918 479434
rect 297154 479198 303918 479434
rect 304154 479198 310918 479434
rect 311154 479198 317918 479434
rect 318154 479198 324918 479434
rect 325154 479198 331918 479434
rect 332154 479198 338918 479434
rect 339154 479198 345918 479434
rect 346154 479198 352918 479434
rect 353154 479198 359918 479434
rect 360154 479198 366918 479434
rect 367154 479198 373918 479434
rect 374154 479198 380918 479434
rect 381154 479198 387918 479434
rect 388154 479198 394918 479434
rect 395154 479198 401918 479434
rect 402154 479198 408918 479434
rect 409154 479198 415918 479434
rect 416154 479198 422918 479434
rect 423154 479198 429918 479434
rect 430154 479198 436918 479434
rect 437154 479198 443918 479434
rect 444154 479198 450918 479434
rect 451154 479198 457918 479434
rect 458154 479198 464918 479434
rect 465154 479198 471918 479434
rect 472154 479198 478918 479434
rect 479154 479198 485918 479434
rect 486154 479198 492918 479434
rect 493154 479198 499918 479434
rect 500154 479198 506918 479434
rect 507154 479198 513918 479434
rect 514154 479198 520918 479434
rect 521154 479198 527918 479434
rect 528154 479198 534918 479434
rect 535154 479198 541918 479434
rect 542154 479198 548918 479434
rect 549154 479198 555918 479434
rect 556154 479198 562918 479434
rect 563154 479198 569918 479434
rect 570154 479198 576918 479434
rect 577154 479198 587570 479434
rect 587806 479198 587890 479434
rect 588126 479198 588210 479434
rect 588446 479198 588530 479434
rect 588766 479198 588874 479434
rect -4950 479156 588874 479198
rect -4950 478494 588874 478536
rect -4950 478258 -3090 478494
rect -2854 478258 -2770 478494
rect -2534 478258 -2450 478494
rect -2214 478258 -2130 478494
rect -1894 478258 1186 478494
rect 1422 478258 8186 478494
rect 8422 478258 15186 478494
rect 15422 478258 22186 478494
rect 22422 478258 29186 478494
rect 29422 478258 36186 478494
rect 36422 478258 43186 478494
rect 43422 478258 50186 478494
rect 50422 478258 57186 478494
rect 57422 478258 64186 478494
rect 64422 478258 71186 478494
rect 71422 478258 78186 478494
rect 78422 478258 85186 478494
rect 85422 478258 92186 478494
rect 92422 478258 99186 478494
rect 99422 478258 106186 478494
rect 106422 478258 113186 478494
rect 113422 478258 120186 478494
rect 120422 478258 127186 478494
rect 127422 478258 134186 478494
rect 134422 478258 141186 478494
rect 141422 478258 148186 478494
rect 148422 478258 155186 478494
rect 155422 478258 162186 478494
rect 162422 478258 169186 478494
rect 169422 478258 176186 478494
rect 176422 478258 183186 478494
rect 183422 478258 190186 478494
rect 190422 478258 197186 478494
rect 197422 478258 204186 478494
rect 204422 478258 211186 478494
rect 211422 478258 218186 478494
rect 218422 478258 225186 478494
rect 225422 478258 232186 478494
rect 232422 478258 239186 478494
rect 239422 478258 246186 478494
rect 246422 478258 253186 478494
rect 253422 478258 260186 478494
rect 260422 478258 267186 478494
rect 267422 478258 274186 478494
rect 274422 478258 281186 478494
rect 281422 478258 288186 478494
rect 288422 478258 295186 478494
rect 295422 478258 302186 478494
rect 302422 478258 309186 478494
rect 309422 478258 316186 478494
rect 316422 478258 323186 478494
rect 323422 478258 330186 478494
rect 330422 478258 337186 478494
rect 337422 478258 344186 478494
rect 344422 478258 351186 478494
rect 351422 478258 358186 478494
rect 358422 478258 365186 478494
rect 365422 478258 372186 478494
rect 372422 478258 379186 478494
rect 379422 478258 386186 478494
rect 386422 478258 393186 478494
rect 393422 478258 400186 478494
rect 400422 478258 407186 478494
rect 407422 478258 414186 478494
rect 414422 478258 421186 478494
rect 421422 478258 428186 478494
rect 428422 478258 435186 478494
rect 435422 478258 442186 478494
rect 442422 478258 449186 478494
rect 449422 478258 456186 478494
rect 456422 478258 463186 478494
rect 463422 478258 470186 478494
rect 470422 478258 477186 478494
rect 477422 478258 484186 478494
rect 484422 478258 491186 478494
rect 491422 478258 498186 478494
rect 498422 478258 505186 478494
rect 505422 478258 512186 478494
rect 512422 478258 519186 478494
rect 519422 478258 526186 478494
rect 526422 478258 533186 478494
rect 533422 478258 540186 478494
rect 540422 478258 547186 478494
rect 547422 478258 554186 478494
rect 554422 478258 561186 478494
rect 561422 478258 568186 478494
rect 568422 478258 575186 478494
rect 575422 478258 582186 478494
rect 582422 478258 585818 478494
rect 586054 478258 586138 478494
rect 586374 478258 586458 478494
rect 586694 478258 586778 478494
rect 587014 478258 588874 478494
rect -4950 478216 588874 478258
rect -4950 472434 588874 472476
rect -4950 472198 -4842 472434
rect -4606 472198 -4522 472434
rect -4286 472198 -4202 472434
rect -3966 472198 -3882 472434
rect -3646 472198 2918 472434
rect 3154 472198 9918 472434
rect 10154 472198 16918 472434
rect 17154 472198 23918 472434
rect 24154 472198 30918 472434
rect 31154 472198 37918 472434
rect 38154 472198 44918 472434
rect 45154 472198 51918 472434
rect 52154 472198 58918 472434
rect 59154 472198 65918 472434
rect 66154 472198 72918 472434
rect 73154 472198 79918 472434
rect 80154 472198 86918 472434
rect 87154 472198 93918 472434
rect 94154 472198 100918 472434
rect 101154 472198 107918 472434
rect 108154 472198 114918 472434
rect 115154 472198 121918 472434
rect 122154 472198 128918 472434
rect 129154 472198 135918 472434
rect 136154 472198 142918 472434
rect 143154 472198 149918 472434
rect 150154 472198 156918 472434
rect 157154 472198 163918 472434
rect 164154 472198 170918 472434
rect 171154 472198 177918 472434
rect 178154 472198 184918 472434
rect 185154 472198 191918 472434
rect 192154 472198 198918 472434
rect 199154 472198 205918 472434
rect 206154 472198 212918 472434
rect 213154 472198 219918 472434
rect 220154 472198 226918 472434
rect 227154 472198 233918 472434
rect 234154 472198 240918 472434
rect 241154 472198 247918 472434
rect 248154 472198 254918 472434
rect 255154 472198 261918 472434
rect 262154 472198 268918 472434
rect 269154 472198 275918 472434
rect 276154 472198 282918 472434
rect 283154 472198 289918 472434
rect 290154 472198 296918 472434
rect 297154 472198 303918 472434
rect 304154 472198 310918 472434
rect 311154 472198 317918 472434
rect 318154 472198 324918 472434
rect 325154 472198 331918 472434
rect 332154 472198 338918 472434
rect 339154 472198 345918 472434
rect 346154 472198 352918 472434
rect 353154 472198 359918 472434
rect 360154 472198 366918 472434
rect 367154 472198 373918 472434
rect 374154 472198 380918 472434
rect 381154 472198 387918 472434
rect 388154 472198 394918 472434
rect 395154 472198 401918 472434
rect 402154 472198 408918 472434
rect 409154 472198 415918 472434
rect 416154 472198 422918 472434
rect 423154 472198 429918 472434
rect 430154 472198 436918 472434
rect 437154 472198 443918 472434
rect 444154 472198 450918 472434
rect 451154 472198 457918 472434
rect 458154 472198 464918 472434
rect 465154 472198 471918 472434
rect 472154 472198 478918 472434
rect 479154 472198 485918 472434
rect 486154 472198 492918 472434
rect 493154 472198 499918 472434
rect 500154 472198 506918 472434
rect 507154 472198 513918 472434
rect 514154 472198 520918 472434
rect 521154 472198 527918 472434
rect 528154 472198 534918 472434
rect 535154 472198 541918 472434
rect 542154 472198 548918 472434
rect 549154 472198 555918 472434
rect 556154 472198 562918 472434
rect 563154 472198 569918 472434
rect 570154 472198 576918 472434
rect 577154 472198 587570 472434
rect 587806 472198 587890 472434
rect 588126 472198 588210 472434
rect 588446 472198 588530 472434
rect 588766 472198 588874 472434
rect -4950 472156 588874 472198
rect -4950 471494 588874 471536
rect -4950 471258 -3090 471494
rect -2854 471258 -2770 471494
rect -2534 471258 -2450 471494
rect -2214 471258 -2130 471494
rect -1894 471258 1186 471494
rect 1422 471258 8186 471494
rect 8422 471258 15186 471494
rect 15422 471258 22186 471494
rect 22422 471258 29186 471494
rect 29422 471258 36186 471494
rect 36422 471258 43186 471494
rect 43422 471258 50186 471494
rect 50422 471258 57186 471494
rect 57422 471258 64186 471494
rect 64422 471258 71186 471494
rect 71422 471258 78186 471494
rect 78422 471258 85186 471494
rect 85422 471258 92186 471494
rect 92422 471258 99186 471494
rect 99422 471258 106186 471494
rect 106422 471258 113186 471494
rect 113422 471258 120186 471494
rect 120422 471258 127186 471494
rect 127422 471258 134186 471494
rect 134422 471258 141186 471494
rect 141422 471258 148186 471494
rect 148422 471258 155186 471494
rect 155422 471258 162186 471494
rect 162422 471258 169186 471494
rect 169422 471258 176186 471494
rect 176422 471258 183186 471494
rect 183422 471258 190186 471494
rect 190422 471258 197186 471494
rect 197422 471258 204186 471494
rect 204422 471258 211186 471494
rect 211422 471258 218186 471494
rect 218422 471258 225186 471494
rect 225422 471258 232186 471494
rect 232422 471258 239186 471494
rect 239422 471258 246186 471494
rect 246422 471258 253186 471494
rect 253422 471258 260186 471494
rect 260422 471258 267186 471494
rect 267422 471258 274186 471494
rect 274422 471258 281186 471494
rect 281422 471258 288186 471494
rect 288422 471258 295186 471494
rect 295422 471258 302186 471494
rect 302422 471258 309186 471494
rect 309422 471258 316186 471494
rect 316422 471258 323186 471494
rect 323422 471258 330186 471494
rect 330422 471258 337186 471494
rect 337422 471258 344186 471494
rect 344422 471258 351186 471494
rect 351422 471258 358186 471494
rect 358422 471258 365186 471494
rect 365422 471258 372186 471494
rect 372422 471258 379186 471494
rect 379422 471258 386186 471494
rect 386422 471258 393186 471494
rect 393422 471258 400186 471494
rect 400422 471258 407186 471494
rect 407422 471258 414186 471494
rect 414422 471258 421186 471494
rect 421422 471258 428186 471494
rect 428422 471258 435186 471494
rect 435422 471258 442186 471494
rect 442422 471258 449186 471494
rect 449422 471258 456186 471494
rect 456422 471258 463186 471494
rect 463422 471258 470186 471494
rect 470422 471258 477186 471494
rect 477422 471258 484186 471494
rect 484422 471258 491186 471494
rect 491422 471258 498186 471494
rect 498422 471258 505186 471494
rect 505422 471258 512186 471494
rect 512422 471258 519186 471494
rect 519422 471258 526186 471494
rect 526422 471258 533186 471494
rect 533422 471258 540186 471494
rect 540422 471258 547186 471494
rect 547422 471258 554186 471494
rect 554422 471258 561186 471494
rect 561422 471258 568186 471494
rect 568422 471258 575186 471494
rect 575422 471258 582186 471494
rect 582422 471258 585818 471494
rect 586054 471258 586138 471494
rect 586374 471258 586458 471494
rect 586694 471258 586778 471494
rect 587014 471258 588874 471494
rect -4950 471216 588874 471258
rect -4950 465434 588874 465476
rect -4950 465198 -4842 465434
rect -4606 465198 -4522 465434
rect -4286 465198 -4202 465434
rect -3966 465198 -3882 465434
rect -3646 465198 2918 465434
rect 3154 465198 9918 465434
rect 10154 465198 16918 465434
rect 17154 465198 23918 465434
rect 24154 465198 30918 465434
rect 31154 465198 37918 465434
rect 38154 465198 44918 465434
rect 45154 465198 51918 465434
rect 52154 465198 58918 465434
rect 59154 465198 65918 465434
rect 66154 465198 72918 465434
rect 73154 465198 79918 465434
rect 80154 465198 86918 465434
rect 87154 465198 93918 465434
rect 94154 465198 100918 465434
rect 101154 465198 107918 465434
rect 108154 465198 114918 465434
rect 115154 465198 121918 465434
rect 122154 465198 128918 465434
rect 129154 465198 135918 465434
rect 136154 465198 142918 465434
rect 143154 465198 149918 465434
rect 150154 465198 156918 465434
rect 157154 465198 163918 465434
rect 164154 465198 170918 465434
rect 171154 465198 177918 465434
rect 178154 465198 184918 465434
rect 185154 465198 191918 465434
rect 192154 465198 198918 465434
rect 199154 465198 205918 465434
rect 206154 465198 212918 465434
rect 213154 465198 219918 465434
rect 220154 465198 226918 465434
rect 227154 465198 233918 465434
rect 234154 465198 240918 465434
rect 241154 465198 247918 465434
rect 248154 465198 254918 465434
rect 255154 465198 261918 465434
rect 262154 465198 268918 465434
rect 269154 465198 275918 465434
rect 276154 465198 282918 465434
rect 283154 465198 289918 465434
rect 290154 465198 296918 465434
rect 297154 465198 303918 465434
rect 304154 465198 310918 465434
rect 311154 465198 317918 465434
rect 318154 465198 324918 465434
rect 325154 465198 331918 465434
rect 332154 465198 338918 465434
rect 339154 465198 345918 465434
rect 346154 465198 352918 465434
rect 353154 465198 359918 465434
rect 360154 465198 366918 465434
rect 367154 465198 373918 465434
rect 374154 465198 380918 465434
rect 381154 465198 387918 465434
rect 388154 465198 394918 465434
rect 395154 465198 401918 465434
rect 402154 465198 408918 465434
rect 409154 465198 415918 465434
rect 416154 465198 422918 465434
rect 423154 465198 429918 465434
rect 430154 465198 436918 465434
rect 437154 465198 443918 465434
rect 444154 465198 450918 465434
rect 451154 465198 457918 465434
rect 458154 465198 464918 465434
rect 465154 465198 471918 465434
rect 472154 465198 478918 465434
rect 479154 465198 485918 465434
rect 486154 465198 492918 465434
rect 493154 465198 499918 465434
rect 500154 465198 506918 465434
rect 507154 465198 513918 465434
rect 514154 465198 520918 465434
rect 521154 465198 527918 465434
rect 528154 465198 534918 465434
rect 535154 465198 541918 465434
rect 542154 465198 548918 465434
rect 549154 465198 555918 465434
rect 556154 465198 562918 465434
rect 563154 465198 569918 465434
rect 570154 465198 576918 465434
rect 577154 465198 587570 465434
rect 587806 465198 587890 465434
rect 588126 465198 588210 465434
rect 588446 465198 588530 465434
rect 588766 465198 588874 465434
rect -4950 465156 588874 465198
rect -4950 464494 588874 464536
rect -4950 464258 -3090 464494
rect -2854 464258 -2770 464494
rect -2534 464258 -2450 464494
rect -2214 464258 -2130 464494
rect -1894 464258 1186 464494
rect 1422 464258 8186 464494
rect 8422 464258 15186 464494
rect 15422 464258 22186 464494
rect 22422 464258 29186 464494
rect 29422 464258 36186 464494
rect 36422 464258 43186 464494
rect 43422 464258 50186 464494
rect 50422 464258 57186 464494
rect 57422 464258 64186 464494
rect 64422 464258 71186 464494
rect 71422 464258 78186 464494
rect 78422 464258 85186 464494
rect 85422 464258 92186 464494
rect 92422 464258 99186 464494
rect 99422 464258 106186 464494
rect 106422 464258 113186 464494
rect 113422 464258 120186 464494
rect 120422 464258 127186 464494
rect 127422 464258 134186 464494
rect 134422 464258 141186 464494
rect 141422 464258 148186 464494
rect 148422 464258 155186 464494
rect 155422 464258 162186 464494
rect 162422 464258 169186 464494
rect 169422 464258 176186 464494
rect 176422 464258 183186 464494
rect 183422 464258 190186 464494
rect 190422 464258 197186 464494
rect 197422 464258 204186 464494
rect 204422 464258 211186 464494
rect 211422 464258 218186 464494
rect 218422 464258 225186 464494
rect 225422 464258 232186 464494
rect 232422 464258 239186 464494
rect 239422 464258 246186 464494
rect 246422 464258 253186 464494
rect 253422 464258 260186 464494
rect 260422 464258 267186 464494
rect 267422 464258 274186 464494
rect 274422 464258 281186 464494
rect 281422 464258 288186 464494
rect 288422 464258 295186 464494
rect 295422 464258 302186 464494
rect 302422 464258 309186 464494
rect 309422 464258 316186 464494
rect 316422 464258 323186 464494
rect 323422 464258 330186 464494
rect 330422 464258 337186 464494
rect 337422 464258 344186 464494
rect 344422 464258 351186 464494
rect 351422 464258 358186 464494
rect 358422 464258 365186 464494
rect 365422 464258 372186 464494
rect 372422 464258 379186 464494
rect 379422 464258 386186 464494
rect 386422 464258 393186 464494
rect 393422 464258 400186 464494
rect 400422 464258 407186 464494
rect 407422 464258 414186 464494
rect 414422 464258 421186 464494
rect 421422 464258 428186 464494
rect 428422 464258 435186 464494
rect 435422 464258 442186 464494
rect 442422 464258 449186 464494
rect 449422 464258 456186 464494
rect 456422 464258 463186 464494
rect 463422 464258 470186 464494
rect 470422 464258 477186 464494
rect 477422 464258 484186 464494
rect 484422 464258 491186 464494
rect 491422 464258 498186 464494
rect 498422 464258 505186 464494
rect 505422 464258 512186 464494
rect 512422 464258 519186 464494
rect 519422 464258 526186 464494
rect 526422 464258 533186 464494
rect 533422 464258 540186 464494
rect 540422 464258 547186 464494
rect 547422 464258 554186 464494
rect 554422 464258 561186 464494
rect 561422 464258 568186 464494
rect 568422 464258 575186 464494
rect 575422 464258 582186 464494
rect 582422 464258 585818 464494
rect 586054 464258 586138 464494
rect 586374 464258 586458 464494
rect 586694 464258 586778 464494
rect 587014 464258 588874 464494
rect -4950 464216 588874 464258
rect -4950 458434 588874 458476
rect -4950 458198 -4842 458434
rect -4606 458198 -4522 458434
rect -4286 458198 -4202 458434
rect -3966 458198 -3882 458434
rect -3646 458198 2918 458434
rect 3154 458198 9918 458434
rect 10154 458198 16918 458434
rect 17154 458198 23918 458434
rect 24154 458198 30918 458434
rect 31154 458198 37918 458434
rect 38154 458198 44918 458434
rect 45154 458198 51918 458434
rect 52154 458198 58918 458434
rect 59154 458198 65918 458434
rect 66154 458198 72918 458434
rect 73154 458198 79918 458434
rect 80154 458198 86918 458434
rect 87154 458198 93918 458434
rect 94154 458198 100918 458434
rect 101154 458198 107918 458434
rect 108154 458198 114918 458434
rect 115154 458198 121918 458434
rect 122154 458198 128918 458434
rect 129154 458198 135918 458434
rect 136154 458198 142918 458434
rect 143154 458198 149918 458434
rect 150154 458198 156918 458434
rect 157154 458198 163918 458434
rect 164154 458198 170918 458434
rect 171154 458198 177918 458434
rect 178154 458198 184918 458434
rect 185154 458198 191918 458434
rect 192154 458198 198918 458434
rect 199154 458198 205918 458434
rect 206154 458198 212918 458434
rect 213154 458198 219918 458434
rect 220154 458198 226918 458434
rect 227154 458198 233918 458434
rect 234154 458198 240918 458434
rect 241154 458198 247918 458434
rect 248154 458198 254918 458434
rect 255154 458198 261918 458434
rect 262154 458198 268918 458434
rect 269154 458198 275918 458434
rect 276154 458198 282918 458434
rect 283154 458198 289918 458434
rect 290154 458198 296918 458434
rect 297154 458198 303918 458434
rect 304154 458198 310918 458434
rect 311154 458198 317918 458434
rect 318154 458198 324918 458434
rect 325154 458198 331918 458434
rect 332154 458198 338918 458434
rect 339154 458198 345918 458434
rect 346154 458198 352918 458434
rect 353154 458198 359918 458434
rect 360154 458198 366918 458434
rect 367154 458198 373918 458434
rect 374154 458198 380918 458434
rect 381154 458198 387918 458434
rect 388154 458198 394918 458434
rect 395154 458198 401918 458434
rect 402154 458198 408918 458434
rect 409154 458198 415918 458434
rect 416154 458198 422918 458434
rect 423154 458198 429918 458434
rect 430154 458198 436918 458434
rect 437154 458198 443918 458434
rect 444154 458198 450918 458434
rect 451154 458198 457918 458434
rect 458154 458198 464918 458434
rect 465154 458198 471918 458434
rect 472154 458198 478918 458434
rect 479154 458198 485918 458434
rect 486154 458198 492918 458434
rect 493154 458198 499918 458434
rect 500154 458198 506918 458434
rect 507154 458198 513918 458434
rect 514154 458198 520918 458434
rect 521154 458198 527918 458434
rect 528154 458198 534918 458434
rect 535154 458198 541918 458434
rect 542154 458198 548918 458434
rect 549154 458198 555918 458434
rect 556154 458198 562918 458434
rect 563154 458198 569918 458434
rect 570154 458198 576918 458434
rect 577154 458198 587570 458434
rect 587806 458198 587890 458434
rect 588126 458198 588210 458434
rect 588446 458198 588530 458434
rect 588766 458198 588874 458434
rect -4950 458156 588874 458198
rect -4950 457494 588874 457536
rect -4950 457258 -3090 457494
rect -2854 457258 -2770 457494
rect -2534 457258 -2450 457494
rect -2214 457258 -2130 457494
rect -1894 457258 1186 457494
rect 1422 457258 8186 457494
rect 8422 457258 15186 457494
rect 15422 457258 22186 457494
rect 22422 457258 29186 457494
rect 29422 457258 36186 457494
rect 36422 457258 43186 457494
rect 43422 457258 50186 457494
rect 50422 457258 57186 457494
rect 57422 457258 64186 457494
rect 64422 457258 71186 457494
rect 71422 457258 78186 457494
rect 78422 457258 85186 457494
rect 85422 457258 92186 457494
rect 92422 457258 99186 457494
rect 99422 457258 106186 457494
rect 106422 457258 113186 457494
rect 113422 457258 120186 457494
rect 120422 457258 127186 457494
rect 127422 457258 134186 457494
rect 134422 457258 141186 457494
rect 141422 457258 148186 457494
rect 148422 457258 155186 457494
rect 155422 457258 162186 457494
rect 162422 457258 169186 457494
rect 169422 457258 176186 457494
rect 176422 457258 183186 457494
rect 183422 457258 190186 457494
rect 190422 457258 197186 457494
rect 197422 457258 204186 457494
rect 204422 457258 211186 457494
rect 211422 457258 218186 457494
rect 218422 457258 225186 457494
rect 225422 457258 232186 457494
rect 232422 457258 239186 457494
rect 239422 457258 246186 457494
rect 246422 457258 253186 457494
rect 253422 457258 260186 457494
rect 260422 457258 267186 457494
rect 267422 457258 274186 457494
rect 274422 457258 281186 457494
rect 281422 457258 288186 457494
rect 288422 457258 295186 457494
rect 295422 457258 302186 457494
rect 302422 457258 309186 457494
rect 309422 457258 316186 457494
rect 316422 457258 323186 457494
rect 323422 457258 330186 457494
rect 330422 457258 337186 457494
rect 337422 457258 344186 457494
rect 344422 457258 351186 457494
rect 351422 457258 358186 457494
rect 358422 457258 365186 457494
rect 365422 457258 372186 457494
rect 372422 457258 379186 457494
rect 379422 457258 386186 457494
rect 386422 457258 393186 457494
rect 393422 457258 400186 457494
rect 400422 457258 407186 457494
rect 407422 457258 414186 457494
rect 414422 457258 421186 457494
rect 421422 457258 428186 457494
rect 428422 457258 435186 457494
rect 435422 457258 442186 457494
rect 442422 457258 449186 457494
rect 449422 457258 456186 457494
rect 456422 457258 463186 457494
rect 463422 457258 470186 457494
rect 470422 457258 477186 457494
rect 477422 457258 484186 457494
rect 484422 457258 491186 457494
rect 491422 457258 498186 457494
rect 498422 457258 505186 457494
rect 505422 457258 512186 457494
rect 512422 457258 519186 457494
rect 519422 457258 526186 457494
rect 526422 457258 533186 457494
rect 533422 457258 540186 457494
rect 540422 457258 547186 457494
rect 547422 457258 554186 457494
rect 554422 457258 561186 457494
rect 561422 457258 568186 457494
rect 568422 457258 575186 457494
rect 575422 457258 582186 457494
rect 582422 457258 585818 457494
rect 586054 457258 586138 457494
rect 586374 457258 586458 457494
rect 586694 457258 586778 457494
rect 587014 457258 588874 457494
rect -4950 457216 588874 457258
rect -4950 451434 588874 451476
rect -4950 451198 -4842 451434
rect -4606 451198 -4522 451434
rect -4286 451198 -4202 451434
rect -3966 451198 -3882 451434
rect -3646 451198 2918 451434
rect 3154 451198 9918 451434
rect 10154 451198 16918 451434
rect 17154 451198 23918 451434
rect 24154 451198 30918 451434
rect 31154 451198 37918 451434
rect 38154 451198 44918 451434
rect 45154 451198 51918 451434
rect 52154 451198 58918 451434
rect 59154 451198 65918 451434
rect 66154 451198 72918 451434
rect 73154 451198 79918 451434
rect 80154 451198 86918 451434
rect 87154 451198 93918 451434
rect 94154 451198 100918 451434
rect 101154 451198 107918 451434
rect 108154 451198 114918 451434
rect 115154 451198 121918 451434
rect 122154 451198 128918 451434
rect 129154 451198 135918 451434
rect 136154 451198 142918 451434
rect 143154 451198 149918 451434
rect 150154 451198 156918 451434
rect 157154 451198 163918 451434
rect 164154 451198 170918 451434
rect 171154 451198 177918 451434
rect 178154 451198 184918 451434
rect 185154 451198 191918 451434
rect 192154 451198 198918 451434
rect 199154 451198 205918 451434
rect 206154 451198 212918 451434
rect 213154 451198 219918 451434
rect 220154 451198 226918 451434
rect 227154 451198 233918 451434
rect 234154 451198 240918 451434
rect 241154 451198 247918 451434
rect 248154 451198 254918 451434
rect 255154 451198 261918 451434
rect 262154 451198 268918 451434
rect 269154 451198 275918 451434
rect 276154 451198 282918 451434
rect 283154 451198 289918 451434
rect 290154 451198 296918 451434
rect 297154 451198 303918 451434
rect 304154 451198 310918 451434
rect 311154 451198 317918 451434
rect 318154 451198 324918 451434
rect 325154 451198 331918 451434
rect 332154 451198 338918 451434
rect 339154 451198 345918 451434
rect 346154 451198 352918 451434
rect 353154 451198 359918 451434
rect 360154 451198 366918 451434
rect 367154 451198 373918 451434
rect 374154 451198 380918 451434
rect 381154 451198 387918 451434
rect 388154 451198 394918 451434
rect 395154 451198 401918 451434
rect 402154 451198 408918 451434
rect 409154 451198 415918 451434
rect 416154 451198 422918 451434
rect 423154 451198 429918 451434
rect 430154 451198 436918 451434
rect 437154 451198 443918 451434
rect 444154 451198 450918 451434
rect 451154 451198 457918 451434
rect 458154 451198 464918 451434
rect 465154 451198 471918 451434
rect 472154 451198 478918 451434
rect 479154 451198 485918 451434
rect 486154 451198 492918 451434
rect 493154 451198 499918 451434
rect 500154 451198 506918 451434
rect 507154 451198 513918 451434
rect 514154 451198 520918 451434
rect 521154 451198 527918 451434
rect 528154 451198 534918 451434
rect 535154 451198 541918 451434
rect 542154 451198 548918 451434
rect 549154 451198 555918 451434
rect 556154 451198 562918 451434
rect 563154 451198 569918 451434
rect 570154 451198 576918 451434
rect 577154 451198 587570 451434
rect 587806 451198 587890 451434
rect 588126 451198 588210 451434
rect 588446 451198 588530 451434
rect 588766 451198 588874 451434
rect -4950 451156 588874 451198
rect -4950 450494 588874 450536
rect -4950 450258 -3090 450494
rect -2854 450258 -2770 450494
rect -2534 450258 -2450 450494
rect -2214 450258 -2130 450494
rect -1894 450258 1186 450494
rect 1422 450258 8186 450494
rect 8422 450258 15186 450494
rect 15422 450258 22186 450494
rect 22422 450258 29186 450494
rect 29422 450258 36186 450494
rect 36422 450258 43186 450494
rect 43422 450258 50186 450494
rect 50422 450258 57186 450494
rect 57422 450258 64186 450494
rect 64422 450258 71186 450494
rect 71422 450258 78186 450494
rect 78422 450258 85186 450494
rect 85422 450258 92186 450494
rect 92422 450258 99186 450494
rect 99422 450258 106186 450494
rect 106422 450258 113186 450494
rect 113422 450258 120186 450494
rect 120422 450258 127186 450494
rect 127422 450258 134186 450494
rect 134422 450258 141186 450494
rect 141422 450258 148186 450494
rect 148422 450258 155186 450494
rect 155422 450258 162186 450494
rect 162422 450258 169186 450494
rect 169422 450258 176186 450494
rect 176422 450258 183186 450494
rect 183422 450258 190186 450494
rect 190422 450258 197186 450494
rect 197422 450258 204186 450494
rect 204422 450258 211186 450494
rect 211422 450258 218186 450494
rect 218422 450258 225186 450494
rect 225422 450258 232186 450494
rect 232422 450258 239186 450494
rect 239422 450258 246186 450494
rect 246422 450258 253186 450494
rect 253422 450258 260186 450494
rect 260422 450258 267186 450494
rect 267422 450258 274186 450494
rect 274422 450258 281186 450494
rect 281422 450258 288186 450494
rect 288422 450258 295186 450494
rect 295422 450258 302186 450494
rect 302422 450258 309186 450494
rect 309422 450258 316186 450494
rect 316422 450258 323186 450494
rect 323422 450258 330186 450494
rect 330422 450258 337186 450494
rect 337422 450258 344186 450494
rect 344422 450258 351186 450494
rect 351422 450258 358186 450494
rect 358422 450258 365186 450494
rect 365422 450258 372186 450494
rect 372422 450258 379186 450494
rect 379422 450258 386186 450494
rect 386422 450258 393186 450494
rect 393422 450258 400186 450494
rect 400422 450258 407186 450494
rect 407422 450258 414186 450494
rect 414422 450258 421186 450494
rect 421422 450258 428186 450494
rect 428422 450258 435186 450494
rect 435422 450258 442186 450494
rect 442422 450258 449186 450494
rect 449422 450258 456186 450494
rect 456422 450258 463186 450494
rect 463422 450258 470186 450494
rect 470422 450258 477186 450494
rect 477422 450258 484186 450494
rect 484422 450258 491186 450494
rect 491422 450258 498186 450494
rect 498422 450258 505186 450494
rect 505422 450258 512186 450494
rect 512422 450258 519186 450494
rect 519422 450258 526186 450494
rect 526422 450258 533186 450494
rect 533422 450258 540186 450494
rect 540422 450258 547186 450494
rect 547422 450258 554186 450494
rect 554422 450258 561186 450494
rect 561422 450258 568186 450494
rect 568422 450258 575186 450494
rect 575422 450258 582186 450494
rect 582422 450258 585818 450494
rect 586054 450258 586138 450494
rect 586374 450258 586458 450494
rect 586694 450258 586778 450494
rect 587014 450258 588874 450494
rect -4950 450216 588874 450258
rect -4950 444434 588874 444476
rect -4950 444198 -4842 444434
rect -4606 444198 -4522 444434
rect -4286 444198 -4202 444434
rect -3966 444198 -3882 444434
rect -3646 444198 2918 444434
rect 3154 444198 9918 444434
rect 10154 444198 16918 444434
rect 17154 444198 23918 444434
rect 24154 444198 30918 444434
rect 31154 444198 37918 444434
rect 38154 444198 44918 444434
rect 45154 444198 51918 444434
rect 52154 444198 58918 444434
rect 59154 444198 65918 444434
rect 66154 444198 72918 444434
rect 73154 444198 79918 444434
rect 80154 444198 86918 444434
rect 87154 444198 93918 444434
rect 94154 444198 100918 444434
rect 101154 444198 107918 444434
rect 108154 444198 114918 444434
rect 115154 444198 121918 444434
rect 122154 444198 128918 444434
rect 129154 444198 135918 444434
rect 136154 444198 142918 444434
rect 143154 444198 149918 444434
rect 150154 444198 156918 444434
rect 157154 444198 163918 444434
rect 164154 444198 170918 444434
rect 171154 444198 177918 444434
rect 178154 444198 184918 444434
rect 185154 444198 191918 444434
rect 192154 444198 198918 444434
rect 199154 444198 205918 444434
rect 206154 444198 212918 444434
rect 213154 444198 219918 444434
rect 220154 444198 226918 444434
rect 227154 444198 233918 444434
rect 234154 444198 240918 444434
rect 241154 444198 247918 444434
rect 248154 444198 254918 444434
rect 255154 444198 261918 444434
rect 262154 444198 268918 444434
rect 269154 444198 275918 444434
rect 276154 444198 282918 444434
rect 283154 444198 289918 444434
rect 290154 444198 296918 444434
rect 297154 444198 303918 444434
rect 304154 444198 310918 444434
rect 311154 444198 317918 444434
rect 318154 444198 324918 444434
rect 325154 444198 331918 444434
rect 332154 444198 338918 444434
rect 339154 444198 345918 444434
rect 346154 444198 352918 444434
rect 353154 444198 359918 444434
rect 360154 444198 366918 444434
rect 367154 444198 373918 444434
rect 374154 444198 380918 444434
rect 381154 444198 387918 444434
rect 388154 444198 394918 444434
rect 395154 444198 401918 444434
rect 402154 444198 408918 444434
rect 409154 444198 415918 444434
rect 416154 444198 422918 444434
rect 423154 444198 429918 444434
rect 430154 444198 436918 444434
rect 437154 444198 443918 444434
rect 444154 444198 450918 444434
rect 451154 444198 457918 444434
rect 458154 444198 464918 444434
rect 465154 444198 471918 444434
rect 472154 444198 478918 444434
rect 479154 444198 485918 444434
rect 486154 444198 492918 444434
rect 493154 444198 499918 444434
rect 500154 444198 506918 444434
rect 507154 444198 513918 444434
rect 514154 444198 520918 444434
rect 521154 444198 527918 444434
rect 528154 444198 534918 444434
rect 535154 444198 541918 444434
rect 542154 444198 548918 444434
rect 549154 444198 555918 444434
rect 556154 444198 562918 444434
rect 563154 444198 569918 444434
rect 570154 444198 576918 444434
rect 577154 444198 587570 444434
rect 587806 444198 587890 444434
rect 588126 444198 588210 444434
rect 588446 444198 588530 444434
rect 588766 444198 588874 444434
rect -4950 444156 588874 444198
rect -4950 443494 588874 443536
rect -4950 443258 -3090 443494
rect -2854 443258 -2770 443494
rect -2534 443258 -2450 443494
rect -2214 443258 -2130 443494
rect -1894 443258 1186 443494
rect 1422 443258 8186 443494
rect 8422 443258 15186 443494
rect 15422 443258 22186 443494
rect 22422 443258 29186 443494
rect 29422 443258 36186 443494
rect 36422 443258 43186 443494
rect 43422 443258 50186 443494
rect 50422 443258 57186 443494
rect 57422 443258 64186 443494
rect 64422 443258 71186 443494
rect 71422 443258 78186 443494
rect 78422 443258 85186 443494
rect 85422 443258 92186 443494
rect 92422 443258 99186 443494
rect 99422 443258 106186 443494
rect 106422 443258 113186 443494
rect 113422 443258 120186 443494
rect 120422 443258 127186 443494
rect 127422 443258 134186 443494
rect 134422 443258 141186 443494
rect 141422 443258 148186 443494
rect 148422 443258 155186 443494
rect 155422 443258 162186 443494
rect 162422 443258 169186 443494
rect 169422 443258 176186 443494
rect 176422 443258 183186 443494
rect 183422 443258 190186 443494
rect 190422 443258 197186 443494
rect 197422 443258 204186 443494
rect 204422 443258 211186 443494
rect 211422 443258 218186 443494
rect 218422 443258 225186 443494
rect 225422 443258 232186 443494
rect 232422 443258 239186 443494
rect 239422 443258 246186 443494
rect 246422 443258 253186 443494
rect 253422 443258 260186 443494
rect 260422 443258 267186 443494
rect 267422 443258 274186 443494
rect 274422 443258 281186 443494
rect 281422 443258 288186 443494
rect 288422 443258 295186 443494
rect 295422 443258 302186 443494
rect 302422 443258 309186 443494
rect 309422 443258 316186 443494
rect 316422 443258 323186 443494
rect 323422 443258 330186 443494
rect 330422 443258 337186 443494
rect 337422 443258 344186 443494
rect 344422 443258 351186 443494
rect 351422 443258 358186 443494
rect 358422 443258 365186 443494
rect 365422 443258 372186 443494
rect 372422 443258 379186 443494
rect 379422 443258 386186 443494
rect 386422 443258 393186 443494
rect 393422 443258 400186 443494
rect 400422 443258 407186 443494
rect 407422 443258 414186 443494
rect 414422 443258 421186 443494
rect 421422 443258 428186 443494
rect 428422 443258 435186 443494
rect 435422 443258 442186 443494
rect 442422 443258 449186 443494
rect 449422 443258 456186 443494
rect 456422 443258 463186 443494
rect 463422 443258 470186 443494
rect 470422 443258 477186 443494
rect 477422 443258 484186 443494
rect 484422 443258 491186 443494
rect 491422 443258 498186 443494
rect 498422 443258 505186 443494
rect 505422 443258 512186 443494
rect 512422 443258 519186 443494
rect 519422 443258 526186 443494
rect 526422 443258 533186 443494
rect 533422 443258 540186 443494
rect 540422 443258 547186 443494
rect 547422 443258 554186 443494
rect 554422 443258 561186 443494
rect 561422 443258 568186 443494
rect 568422 443258 575186 443494
rect 575422 443258 582186 443494
rect 582422 443258 585818 443494
rect 586054 443258 586138 443494
rect 586374 443258 586458 443494
rect 586694 443258 586778 443494
rect 587014 443258 588874 443494
rect -4950 443216 588874 443258
rect -4950 437434 588874 437476
rect -4950 437198 -4842 437434
rect -4606 437198 -4522 437434
rect -4286 437198 -4202 437434
rect -3966 437198 -3882 437434
rect -3646 437198 2918 437434
rect 3154 437198 9918 437434
rect 10154 437198 16918 437434
rect 17154 437198 23918 437434
rect 24154 437198 30918 437434
rect 31154 437198 37918 437434
rect 38154 437198 44918 437434
rect 45154 437198 51918 437434
rect 52154 437198 58918 437434
rect 59154 437198 65918 437434
rect 66154 437198 72918 437434
rect 73154 437198 79918 437434
rect 80154 437198 86918 437434
rect 87154 437198 93918 437434
rect 94154 437198 100918 437434
rect 101154 437198 107918 437434
rect 108154 437198 114918 437434
rect 115154 437198 121918 437434
rect 122154 437198 128918 437434
rect 129154 437198 135918 437434
rect 136154 437198 142918 437434
rect 143154 437198 149918 437434
rect 150154 437198 156918 437434
rect 157154 437198 163918 437434
rect 164154 437198 170918 437434
rect 171154 437198 177918 437434
rect 178154 437198 184918 437434
rect 185154 437198 191918 437434
rect 192154 437198 198918 437434
rect 199154 437198 205918 437434
rect 206154 437198 212918 437434
rect 213154 437198 219918 437434
rect 220154 437198 226918 437434
rect 227154 437198 233918 437434
rect 234154 437198 240918 437434
rect 241154 437198 247918 437434
rect 248154 437198 254918 437434
rect 255154 437198 261918 437434
rect 262154 437198 268918 437434
rect 269154 437198 275918 437434
rect 276154 437198 282918 437434
rect 283154 437198 289918 437434
rect 290154 437198 296918 437434
rect 297154 437198 303918 437434
rect 304154 437198 310918 437434
rect 311154 437198 317918 437434
rect 318154 437198 324918 437434
rect 325154 437198 331918 437434
rect 332154 437198 338918 437434
rect 339154 437198 345918 437434
rect 346154 437198 352918 437434
rect 353154 437198 359918 437434
rect 360154 437198 366918 437434
rect 367154 437198 373918 437434
rect 374154 437198 380918 437434
rect 381154 437198 387918 437434
rect 388154 437198 394918 437434
rect 395154 437198 401918 437434
rect 402154 437198 408918 437434
rect 409154 437198 415918 437434
rect 416154 437198 422918 437434
rect 423154 437198 429918 437434
rect 430154 437198 436918 437434
rect 437154 437198 443918 437434
rect 444154 437198 450918 437434
rect 451154 437198 457918 437434
rect 458154 437198 464918 437434
rect 465154 437198 471918 437434
rect 472154 437198 478918 437434
rect 479154 437198 485918 437434
rect 486154 437198 492918 437434
rect 493154 437198 499918 437434
rect 500154 437198 506918 437434
rect 507154 437198 513918 437434
rect 514154 437198 520918 437434
rect 521154 437198 527918 437434
rect 528154 437198 534918 437434
rect 535154 437198 541918 437434
rect 542154 437198 548918 437434
rect 549154 437198 555918 437434
rect 556154 437198 562918 437434
rect 563154 437198 569918 437434
rect 570154 437198 576918 437434
rect 577154 437198 587570 437434
rect 587806 437198 587890 437434
rect 588126 437198 588210 437434
rect 588446 437198 588530 437434
rect 588766 437198 588874 437434
rect -4950 437156 588874 437198
rect -4950 436494 588874 436536
rect -4950 436258 -3090 436494
rect -2854 436258 -2770 436494
rect -2534 436258 -2450 436494
rect -2214 436258 -2130 436494
rect -1894 436258 1186 436494
rect 1422 436258 8186 436494
rect 8422 436258 15186 436494
rect 15422 436258 22186 436494
rect 22422 436258 29186 436494
rect 29422 436258 36186 436494
rect 36422 436258 43186 436494
rect 43422 436258 50186 436494
rect 50422 436258 57186 436494
rect 57422 436258 64186 436494
rect 64422 436258 71186 436494
rect 71422 436258 78186 436494
rect 78422 436258 85186 436494
rect 85422 436258 92186 436494
rect 92422 436258 99186 436494
rect 99422 436258 106186 436494
rect 106422 436258 113186 436494
rect 113422 436258 120186 436494
rect 120422 436258 127186 436494
rect 127422 436258 134186 436494
rect 134422 436258 141186 436494
rect 141422 436258 148186 436494
rect 148422 436258 155186 436494
rect 155422 436258 162186 436494
rect 162422 436258 169186 436494
rect 169422 436258 176186 436494
rect 176422 436258 183186 436494
rect 183422 436258 190186 436494
rect 190422 436258 197186 436494
rect 197422 436258 204186 436494
rect 204422 436258 211186 436494
rect 211422 436258 218186 436494
rect 218422 436258 225186 436494
rect 225422 436258 232186 436494
rect 232422 436258 239186 436494
rect 239422 436258 246186 436494
rect 246422 436258 253186 436494
rect 253422 436258 260186 436494
rect 260422 436258 267186 436494
rect 267422 436258 274186 436494
rect 274422 436258 281186 436494
rect 281422 436258 288186 436494
rect 288422 436258 295186 436494
rect 295422 436258 302186 436494
rect 302422 436258 309186 436494
rect 309422 436258 316186 436494
rect 316422 436258 323186 436494
rect 323422 436258 330186 436494
rect 330422 436258 337186 436494
rect 337422 436258 344186 436494
rect 344422 436258 351186 436494
rect 351422 436258 358186 436494
rect 358422 436258 365186 436494
rect 365422 436258 372186 436494
rect 372422 436258 379186 436494
rect 379422 436258 386186 436494
rect 386422 436258 393186 436494
rect 393422 436258 400186 436494
rect 400422 436258 407186 436494
rect 407422 436258 414186 436494
rect 414422 436258 421186 436494
rect 421422 436258 428186 436494
rect 428422 436258 435186 436494
rect 435422 436258 442186 436494
rect 442422 436258 449186 436494
rect 449422 436258 456186 436494
rect 456422 436258 463186 436494
rect 463422 436258 470186 436494
rect 470422 436258 477186 436494
rect 477422 436258 484186 436494
rect 484422 436258 491186 436494
rect 491422 436258 498186 436494
rect 498422 436258 505186 436494
rect 505422 436258 512186 436494
rect 512422 436258 519186 436494
rect 519422 436258 526186 436494
rect 526422 436258 533186 436494
rect 533422 436258 540186 436494
rect 540422 436258 547186 436494
rect 547422 436258 554186 436494
rect 554422 436258 561186 436494
rect 561422 436258 568186 436494
rect 568422 436258 575186 436494
rect 575422 436258 582186 436494
rect 582422 436258 585818 436494
rect 586054 436258 586138 436494
rect 586374 436258 586458 436494
rect 586694 436258 586778 436494
rect 587014 436258 588874 436494
rect -4950 436216 588874 436258
rect -4950 430434 588874 430476
rect -4950 430198 -4842 430434
rect -4606 430198 -4522 430434
rect -4286 430198 -4202 430434
rect -3966 430198 -3882 430434
rect -3646 430198 2918 430434
rect 3154 430198 9918 430434
rect 10154 430198 16918 430434
rect 17154 430198 23918 430434
rect 24154 430198 30918 430434
rect 31154 430198 37918 430434
rect 38154 430198 44918 430434
rect 45154 430198 51918 430434
rect 52154 430198 58918 430434
rect 59154 430198 65918 430434
rect 66154 430198 72918 430434
rect 73154 430198 79918 430434
rect 80154 430198 86918 430434
rect 87154 430198 93918 430434
rect 94154 430198 100918 430434
rect 101154 430198 107918 430434
rect 108154 430198 114918 430434
rect 115154 430198 121918 430434
rect 122154 430198 128918 430434
rect 129154 430198 135918 430434
rect 136154 430198 142918 430434
rect 143154 430198 149918 430434
rect 150154 430198 156918 430434
rect 157154 430198 163918 430434
rect 164154 430198 170918 430434
rect 171154 430198 177918 430434
rect 178154 430198 184918 430434
rect 185154 430198 191918 430434
rect 192154 430198 198918 430434
rect 199154 430198 205918 430434
rect 206154 430198 212918 430434
rect 213154 430198 219918 430434
rect 220154 430198 226918 430434
rect 227154 430198 233918 430434
rect 234154 430198 240918 430434
rect 241154 430198 247918 430434
rect 248154 430198 254918 430434
rect 255154 430198 261918 430434
rect 262154 430198 268918 430434
rect 269154 430198 275918 430434
rect 276154 430198 282918 430434
rect 283154 430198 289918 430434
rect 290154 430198 296918 430434
rect 297154 430198 303918 430434
rect 304154 430198 310918 430434
rect 311154 430198 317918 430434
rect 318154 430198 324918 430434
rect 325154 430198 331918 430434
rect 332154 430198 338918 430434
rect 339154 430198 345918 430434
rect 346154 430198 352918 430434
rect 353154 430198 359918 430434
rect 360154 430198 366918 430434
rect 367154 430198 373918 430434
rect 374154 430198 380918 430434
rect 381154 430198 387918 430434
rect 388154 430198 394918 430434
rect 395154 430198 401918 430434
rect 402154 430198 408918 430434
rect 409154 430198 415918 430434
rect 416154 430198 422918 430434
rect 423154 430198 429918 430434
rect 430154 430198 436918 430434
rect 437154 430198 443918 430434
rect 444154 430198 450918 430434
rect 451154 430198 457918 430434
rect 458154 430198 464918 430434
rect 465154 430198 471918 430434
rect 472154 430198 478918 430434
rect 479154 430198 485918 430434
rect 486154 430198 492918 430434
rect 493154 430198 499918 430434
rect 500154 430198 506918 430434
rect 507154 430198 513918 430434
rect 514154 430198 520918 430434
rect 521154 430198 527918 430434
rect 528154 430198 534918 430434
rect 535154 430198 541918 430434
rect 542154 430198 548918 430434
rect 549154 430198 555918 430434
rect 556154 430198 562918 430434
rect 563154 430198 569918 430434
rect 570154 430198 576918 430434
rect 577154 430198 587570 430434
rect 587806 430198 587890 430434
rect 588126 430198 588210 430434
rect 588446 430198 588530 430434
rect 588766 430198 588874 430434
rect -4950 430156 588874 430198
rect -4950 429494 588874 429536
rect -4950 429258 -3090 429494
rect -2854 429258 -2770 429494
rect -2534 429258 -2450 429494
rect -2214 429258 -2130 429494
rect -1894 429258 1186 429494
rect 1422 429258 8186 429494
rect 8422 429258 15186 429494
rect 15422 429258 22186 429494
rect 22422 429258 29186 429494
rect 29422 429258 36186 429494
rect 36422 429258 43186 429494
rect 43422 429258 50186 429494
rect 50422 429258 57186 429494
rect 57422 429258 64186 429494
rect 64422 429258 71186 429494
rect 71422 429258 78186 429494
rect 78422 429258 85186 429494
rect 85422 429258 92186 429494
rect 92422 429258 99186 429494
rect 99422 429258 106186 429494
rect 106422 429258 113186 429494
rect 113422 429258 120186 429494
rect 120422 429258 127186 429494
rect 127422 429258 134186 429494
rect 134422 429258 141186 429494
rect 141422 429258 148186 429494
rect 148422 429258 155186 429494
rect 155422 429258 162186 429494
rect 162422 429258 169186 429494
rect 169422 429258 176186 429494
rect 176422 429258 183186 429494
rect 183422 429258 190186 429494
rect 190422 429258 197186 429494
rect 197422 429258 204186 429494
rect 204422 429258 211186 429494
rect 211422 429258 218186 429494
rect 218422 429258 225186 429494
rect 225422 429258 232186 429494
rect 232422 429258 239186 429494
rect 239422 429258 246186 429494
rect 246422 429258 253186 429494
rect 253422 429258 260186 429494
rect 260422 429258 267186 429494
rect 267422 429258 274186 429494
rect 274422 429258 281186 429494
rect 281422 429258 288186 429494
rect 288422 429258 295186 429494
rect 295422 429258 302186 429494
rect 302422 429258 309186 429494
rect 309422 429258 316186 429494
rect 316422 429258 323186 429494
rect 323422 429258 330186 429494
rect 330422 429258 337186 429494
rect 337422 429258 344186 429494
rect 344422 429258 351186 429494
rect 351422 429258 358186 429494
rect 358422 429258 365186 429494
rect 365422 429258 372186 429494
rect 372422 429258 379186 429494
rect 379422 429258 386186 429494
rect 386422 429258 393186 429494
rect 393422 429258 400186 429494
rect 400422 429258 407186 429494
rect 407422 429258 414186 429494
rect 414422 429258 421186 429494
rect 421422 429258 428186 429494
rect 428422 429258 435186 429494
rect 435422 429258 442186 429494
rect 442422 429258 449186 429494
rect 449422 429258 456186 429494
rect 456422 429258 463186 429494
rect 463422 429258 470186 429494
rect 470422 429258 477186 429494
rect 477422 429258 484186 429494
rect 484422 429258 491186 429494
rect 491422 429258 498186 429494
rect 498422 429258 505186 429494
rect 505422 429258 512186 429494
rect 512422 429258 519186 429494
rect 519422 429258 526186 429494
rect 526422 429258 533186 429494
rect 533422 429258 540186 429494
rect 540422 429258 547186 429494
rect 547422 429258 554186 429494
rect 554422 429258 561186 429494
rect 561422 429258 568186 429494
rect 568422 429258 575186 429494
rect 575422 429258 582186 429494
rect 582422 429258 585818 429494
rect 586054 429258 586138 429494
rect 586374 429258 586458 429494
rect 586694 429258 586778 429494
rect 587014 429258 588874 429494
rect -4950 429216 588874 429258
rect -4950 423434 588874 423476
rect -4950 423198 -4842 423434
rect -4606 423198 -4522 423434
rect -4286 423198 -4202 423434
rect -3966 423198 -3882 423434
rect -3646 423198 2918 423434
rect 3154 423198 9918 423434
rect 10154 423198 16918 423434
rect 17154 423198 23918 423434
rect 24154 423198 30918 423434
rect 31154 423198 37918 423434
rect 38154 423198 44918 423434
rect 45154 423198 51918 423434
rect 52154 423198 58918 423434
rect 59154 423198 65918 423434
rect 66154 423198 72918 423434
rect 73154 423198 79918 423434
rect 80154 423198 86918 423434
rect 87154 423198 93918 423434
rect 94154 423198 100918 423434
rect 101154 423198 107918 423434
rect 108154 423198 114918 423434
rect 115154 423198 121918 423434
rect 122154 423198 128918 423434
rect 129154 423198 135918 423434
rect 136154 423198 142918 423434
rect 143154 423198 149918 423434
rect 150154 423198 156918 423434
rect 157154 423198 163918 423434
rect 164154 423198 170918 423434
rect 171154 423198 177918 423434
rect 178154 423198 184918 423434
rect 185154 423198 191918 423434
rect 192154 423198 198918 423434
rect 199154 423198 205918 423434
rect 206154 423198 212918 423434
rect 213154 423198 219918 423434
rect 220154 423198 226918 423434
rect 227154 423198 233918 423434
rect 234154 423198 240918 423434
rect 241154 423198 247918 423434
rect 248154 423198 254918 423434
rect 255154 423198 261918 423434
rect 262154 423198 268918 423434
rect 269154 423198 275918 423434
rect 276154 423198 282918 423434
rect 283154 423198 289918 423434
rect 290154 423198 296918 423434
rect 297154 423198 303918 423434
rect 304154 423198 310918 423434
rect 311154 423198 317918 423434
rect 318154 423198 324918 423434
rect 325154 423198 331918 423434
rect 332154 423198 338918 423434
rect 339154 423198 345918 423434
rect 346154 423198 352918 423434
rect 353154 423198 359918 423434
rect 360154 423198 366918 423434
rect 367154 423198 373918 423434
rect 374154 423198 380918 423434
rect 381154 423198 387918 423434
rect 388154 423198 394918 423434
rect 395154 423198 401918 423434
rect 402154 423198 408918 423434
rect 409154 423198 415918 423434
rect 416154 423198 422918 423434
rect 423154 423198 429918 423434
rect 430154 423198 436918 423434
rect 437154 423198 443918 423434
rect 444154 423198 450918 423434
rect 451154 423198 457918 423434
rect 458154 423198 464918 423434
rect 465154 423198 471918 423434
rect 472154 423198 478918 423434
rect 479154 423198 485918 423434
rect 486154 423198 492918 423434
rect 493154 423198 499918 423434
rect 500154 423198 506918 423434
rect 507154 423198 513918 423434
rect 514154 423198 520918 423434
rect 521154 423198 527918 423434
rect 528154 423198 534918 423434
rect 535154 423198 541918 423434
rect 542154 423198 548918 423434
rect 549154 423198 555918 423434
rect 556154 423198 562918 423434
rect 563154 423198 569918 423434
rect 570154 423198 576918 423434
rect 577154 423198 587570 423434
rect 587806 423198 587890 423434
rect 588126 423198 588210 423434
rect 588446 423198 588530 423434
rect 588766 423198 588874 423434
rect -4950 423156 588874 423198
rect -4950 422494 588874 422536
rect -4950 422258 -3090 422494
rect -2854 422258 -2770 422494
rect -2534 422258 -2450 422494
rect -2214 422258 -2130 422494
rect -1894 422258 1186 422494
rect 1422 422258 8186 422494
rect 8422 422258 15186 422494
rect 15422 422258 22186 422494
rect 22422 422258 29186 422494
rect 29422 422258 36186 422494
rect 36422 422258 43186 422494
rect 43422 422258 50186 422494
rect 50422 422258 57186 422494
rect 57422 422258 64186 422494
rect 64422 422258 71186 422494
rect 71422 422258 78186 422494
rect 78422 422258 85186 422494
rect 85422 422258 92186 422494
rect 92422 422258 99186 422494
rect 99422 422258 106186 422494
rect 106422 422258 113186 422494
rect 113422 422258 120186 422494
rect 120422 422258 127186 422494
rect 127422 422258 134186 422494
rect 134422 422258 141186 422494
rect 141422 422258 148186 422494
rect 148422 422258 155186 422494
rect 155422 422258 162186 422494
rect 162422 422258 169186 422494
rect 169422 422258 176186 422494
rect 176422 422258 183186 422494
rect 183422 422258 190186 422494
rect 190422 422258 197186 422494
rect 197422 422258 204186 422494
rect 204422 422258 211186 422494
rect 211422 422258 218186 422494
rect 218422 422258 225186 422494
rect 225422 422258 232186 422494
rect 232422 422258 239186 422494
rect 239422 422258 246186 422494
rect 246422 422258 253186 422494
rect 253422 422258 260186 422494
rect 260422 422258 267186 422494
rect 267422 422258 274186 422494
rect 274422 422258 281186 422494
rect 281422 422258 288186 422494
rect 288422 422258 295186 422494
rect 295422 422258 302186 422494
rect 302422 422258 309186 422494
rect 309422 422258 316186 422494
rect 316422 422258 323186 422494
rect 323422 422258 330186 422494
rect 330422 422258 337186 422494
rect 337422 422258 344186 422494
rect 344422 422258 351186 422494
rect 351422 422258 358186 422494
rect 358422 422258 365186 422494
rect 365422 422258 372186 422494
rect 372422 422258 379186 422494
rect 379422 422258 386186 422494
rect 386422 422258 393186 422494
rect 393422 422258 400186 422494
rect 400422 422258 407186 422494
rect 407422 422258 414186 422494
rect 414422 422258 421186 422494
rect 421422 422258 428186 422494
rect 428422 422258 435186 422494
rect 435422 422258 442186 422494
rect 442422 422258 449186 422494
rect 449422 422258 456186 422494
rect 456422 422258 463186 422494
rect 463422 422258 470186 422494
rect 470422 422258 477186 422494
rect 477422 422258 484186 422494
rect 484422 422258 491186 422494
rect 491422 422258 498186 422494
rect 498422 422258 505186 422494
rect 505422 422258 512186 422494
rect 512422 422258 519186 422494
rect 519422 422258 526186 422494
rect 526422 422258 533186 422494
rect 533422 422258 540186 422494
rect 540422 422258 547186 422494
rect 547422 422258 554186 422494
rect 554422 422258 561186 422494
rect 561422 422258 568186 422494
rect 568422 422258 575186 422494
rect 575422 422258 582186 422494
rect 582422 422258 585818 422494
rect 586054 422258 586138 422494
rect 586374 422258 586458 422494
rect 586694 422258 586778 422494
rect 587014 422258 588874 422494
rect -4950 422216 588874 422258
rect -4950 416434 588874 416476
rect -4950 416198 -4842 416434
rect -4606 416198 -4522 416434
rect -4286 416198 -4202 416434
rect -3966 416198 -3882 416434
rect -3646 416198 2918 416434
rect 3154 416198 9918 416434
rect 10154 416198 16918 416434
rect 17154 416198 23918 416434
rect 24154 416198 30918 416434
rect 31154 416198 37918 416434
rect 38154 416198 44918 416434
rect 45154 416198 51918 416434
rect 52154 416198 58918 416434
rect 59154 416198 65918 416434
rect 66154 416198 72918 416434
rect 73154 416198 79918 416434
rect 80154 416198 86918 416434
rect 87154 416198 93918 416434
rect 94154 416198 100918 416434
rect 101154 416198 107918 416434
rect 108154 416198 114918 416434
rect 115154 416198 121918 416434
rect 122154 416198 128918 416434
rect 129154 416198 135918 416434
rect 136154 416198 142918 416434
rect 143154 416198 149918 416434
rect 150154 416198 156918 416434
rect 157154 416198 163918 416434
rect 164154 416198 170918 416434
rect 171154 416198 177918 416434
rect 178154 416198 184918 416434
rect 185154 416198 191918 416434
rect 192154 416198 198918 416434
rect 199154 416198 205918 416434
rect 206154 416198 212918 416434
rect 213154 416198 219918 416434
rect 220154 416198 226918 416434
rect 227154 416198 233918 416434
rect 234154 416198 240918 416434
rect 241154 416198 247918 416434
rect 248154 416198 254918 416434
rect 255154 416198 261918 416434
rect 262154 416198 268918 416434
rect 269154 416198 275918 416434
rect 276154 416198 282918 416434
rect 283154 416198 289918 416434
rect 290154 416198 296918 416434
rect 297154 416198 303918 416434
rect 304154 416198 310918 416434
rect 311154 416198 317918 416434
rect 318154 416198 324918 416434
rect 325154 416198 331918 416434
rect 332154 416198 338918 416434
rect 339154 416198 345918 416434
rect 346154 416198 352918 416434
rect 353154 416198 359918 416434
rect 360154 416198 366918 416434
rect 367154 416198 373918 416434
rect 374154 416198 380918 416434
rect 381154 416198 387918 416434
rect 388154 416198 394918 416434
rect 395154 416198 401918 416434
rect 402154 416198 408918 416434
rect 409154 416198 415918 416434
rect 416154 416198 422918 416434
rect 423154 416198 429918 416434
rect 430154 416198 436918 416434
rect 437154 416198 443918 416434
rect 444154 416198 450918 416434
rect 451154 416198 457918 416434
rect 458154 416198 464918 416434
rect 465154 416198 471918 416434
rect 472154 416198 478918 416434
rect 479154 416198 485918 416434
rect 486154 416198 492918 416434
rect 493154 416198 499918 416434
rect 500154 416198 506918 416434
rect 507154 416198 513918 416434
rect 514154 416198 520918 416434
rect 521154 416198 522850 416434
rect 523086 416198 524782 416434
rect 525018 416198 526714 416434
rect 526950 416198 527918 416434
rect 528154 416198 534918 416434
rect 535154 416198 541918 416434
rect 542154 416198 548918 416434
rect 549154 416198 555918 416434
rect 556154 416198 562918 416434
rect 563154 416198 569918 416434
rect 570154 416198 576918 416434
rect 577154 416198 587570 416434
rect 587806 416198 587890 416434
rect 588126 416198 588210 416434
rect 588446 416198 588530 416434
rect 588766 416198 588874 416434
rect -4950 416156 588874 416198
rect -4950 415494 588874 415536
rect -4950 415258 -3090 415494
rect -2854 415258 -2770 415494
rect -2534 415258 -2450 415494
rect -2214 415258 -2130 415494
rect -1894 415258 1186 415494
rect 1422 415258 8186 415494
rect 8422 415258 15186 415494
rect 15422 415258 22186 415494
rect 22422 415258 29186 415494
rect 29422 415258 36186 415494
rect 36422 415258 43186 415494
rect 43422 415258 50186 415494
rect 50422 415258 57186 415494
rect 57422 415258 64186 415494
rect 64422 415258 71186 415494
rect 71422 415258 78186 415494
rect 78422 415258 85186 415494
rect 85422 415258 92186 415494
rect 92422 415258 99186 415494
rect 99422 415258 106186 415494
rect 106422 415258 113186 415494
rect 113422 415258 120186 415494
rect 120422 415258 127186 415494
rect 127422 415258 134186 415494
rect 134422 415258 141186 415494
rect 141422 415258 148186 415494
rect 148422 415258 155186 415494
rect 155422 415258 162186 415494
rect 162422 415258 169186 415494
rect 169422 415258 176186 415494
rect 176422 415258 183186 415494
rect 183422 415258 190186 415494
rect 190422 415258 197186 415494
rect 197422 415258 204186 415494
rect 204422 415258 211186 415494
rect 211422 415258 218186 415494
rect 218422 415258 225186 415494
rect 225422 415258 232186 415494
rect 232422 415258 239186 415494
rect 239422 415258 246186 415494
rect 246422 415258 253186 415494
rect 253422 415258 260186 415494
rect 260422 415258 267186 415494
rect 267422 415258 274186 415494
rect 274422 415258 281186 415494
rect 281422 415258 288186 415494
rect 288422 415258 295186 415494
rect 295422 415258 302186 415494
rect 302422 415258 309186 415494
rect 309422 415258 316186 415494
rect 316422 415258 323186 415494
rect 323422 415258 330186 415494
rect 330422 415258 337186 415494
rect 337422 415258 344186 415494
rect 344422 415258 351186 415494
rect 351422 415258 358186 415494
rect 358422 415258 365186 415494
rect 365422 415258 372186 415494
rect 372422 415258 379186 415494
rect 379422 415258 386186 415494
rect 386422 415258 393186 415494
rect 393422 415258 400186 415494
rect 400422 415258 407186 415494
rect 407422 415258 414186 415494
rect 414422 415258 421186 415494
rect 421422 415258 428186 415494
rect 428422 415258 435186 415494
rect 435422 415258 442186 415494
rect 442422 415258 449186 415494
rect 449422 415258 456186 415494
rect 456422 415258 463186 415494
rect 463422 415258 470186 415494
rect 470422 415258 477186 415494
rect 477422 415258 484186 415494
rect 484422 415258 491186 415494
rect 491422 415258 498186 415494
rect 498422 415258 505186 415494
rect 505422 415258 512186 415494
rect 512422 415258 519186 415494
rect 519422 415258 519952 415494
rect 520188 415258 521884 415494
rect 522120 415258 523816 415494
rect 524052 415258 525748 415494
rect 525984 415258 533186 415494
rect 533422 415258 540186 415494
rect 540422 415258 547186 415494
rect 547422 415258 554186 415494
rect 554422 415258 561186 415494
rect 561422 415258 568186 415494
rect 568422 415258 575186 415494
rect 575422 415258 582186 415494
rect 582422 415258 585818 415494
rect 586054 415258 586138 415494
rect 586374 415258 586458 415494
rect 586694 415258 586778 415494
rect 587014 415258 588874 415494
rect -4950 415216 588874 415258
rect -4950 409434 588874 409476
rect -4950 409198 -4842 409434
rect -4606 409198 -4522 409434
rect -4286 409198 -4202 409434
rect -3966 409198 -3882 409434
rect -3646 409198 2918 409434
rect 3154 409198 9918 409434
rect 10154 409198 16918 409434
rect 17154 409198 23918 409434
rect 24154 409198 30918 409434
rect 31154 409198 37918 409434
rect 38154 409198 44918 409434
rect 45154 409198 51918 409434
rect 52154 409198 58918 409434
rect 59154 409198 65918 409434
rect 66154 409198 72918 409434
rect 73154 409198 79918 409434
rect 80154 409198 86918 409434
rect 87154 409198 93918 409434
rect 94154 409198 100918 409434
rect 101154 409198 107918 409434
rect 108154 409198 114918 409434
rect 115154 409198 121918 409434
rect 122154 409198 128918 409434
rect 129154 409198 135918 409434
rect 136154 409198 142918 409434
rect 143154 409198 149918 409434
rect 150154 409198 156918 409434
rect 157154 409198 163918 409434
rect 164154 409198 170918 409434
rect 171154 409198 177918 409434
rect 178154 409198 184918 409434
rect 185154 409198 191918 409434
rect 192154 409198 198918 409434
rect 199154 409198 205918 409434
rect 206154 409198 212918 409434
rect 213154 409198 219918 409434
rect 220154 409198 226918 409434
rect 227154 409198 233918 409434
rect 234154 409198 240918 409434
rect 241154 409198 247918 409434
rect 248154 409198 254918 409434
rect 255154 409198 261918 409434
rect 262154 409198 268918 409434
rect 269154 409198 275918 409434
rect 276154 409198 282918 409434
rect 283154 409198 289918 409434
rect 290154 409198 296918 409434
rect 297154 409198 303918 409434
rect 304154 409198 310918 409434
rect 311154 409198 317918 409434
rect 318154 409198 324918 409434
rect 325154 409198 331918 409434
rect 332154 409198 338918 409434
rect 339154 409198 345918 409434
rect 346154 409198 352918 409434
rect 353154 409198 359918 409434
rect 360154 409198 366918 409434
rect 367154 409198 373918 409434
rect 374154 409198 380918 409434
rect 381154 409198 387918 409434
rect 388154 409198 394918 409434
rect 395154 409198 401918 409434
rect 402154 409198 408918 409434
rect 409154 409198 415918 409434
rect 416154 409198 422918 409434
rect 423154 409198 429918 409434
rect 430154 409198 436918 409434
rect 437154 409198 443918 409434
rect 444154 409198 450918 409434
rect 451154 409198 457918 409434
rect 458154 409198 464918 409434
rect 465154 409198 471918 409434
rect 472154 409198 478918 409434
rect 479154 409198 485918 409434
rect 486154 409198 492918 409434
rect 493154 409198 499918 409434
rect 500154 409198 506918 409434
rect 507154 409198 513918 409434
rect 514154 409198 520918 409434
rect 521154 409198 522850 409434
rect 523086 409198 524782 409434
rect 525018 409198 526714 409434
rect 526950 409198 527918 409434
rect 528154 409198 534918 409434
rect 535154 409198 541918 409434
rect 542154 409198 548918 409434
rect 549154 409198 555918 409434
rect 556154 409198 562918 409434
rect 563154 409198 569918 409434
rect 570154 409198 576918 409434
rect 577154 409198 587570 409434
rect 587806 409198 587890 409434
rect 588126 409198 588210 409434
rect 588446 409198 588530 409434
rect 588766 409198 588874 409434
rect -4950 409156 588874 409198
rect -4950 408494 588874 408536
rect -4950 408258 -3090 408494
rect -2854 408258 -2770 408494
rect -2534 408258 -2450 408494
rect -2214 408258 -2130 408494
rect -1894 408258 1186 408494
rect 1422 408258 8186 408494
rect 8422 408258 15186 408494
rect 15422 408258 22186 408494
rect 22422 408258 29186 408494
rect 29422 408258 36186 408494
rect 36422 408258 43186 408494
rect 43422 408258 50186 408494
rect 50422 408258 57186 408494
rect 57422 408258 64186 408494
rect 64422 408258 71186 408494
rect 71422 408258 78186 408494
rect 78422 408258 85186 408494
rect 85422 408258 92186 408494
rect 92422 408258 99186 408494
rect 99422 408258 106186 408494
rect 106422 408258 113186 408494
rect 113422 408258 120186 408494
rect 120422 408258 127186 408494
rect 127422 408258 134186 408494
rect 134422 408258 141186 408494
rect 141422 408258 148186 408494
rect 148422 408258 155186 408494
rect 155422 408258 162186 408494
rect 162422 408258 169186 408494
rect 169422 408258 176186 408494
rect 176422 408258 183186 408494
rect 183422 408258 190186 408494
rect 190422 408258 197186 408494
rect 197422 408258 204186 408494
rect 204422 408258 211186 408494
rect 211422 408258 218186 408494
rect 218422 408258 225186 408494
rect 225422 408258 232186 408494
rect 232422 408258 239186 408494
rect 239422 408258 246186 408494
rect 246422 408258 253186 408494
rect 253422 408258 260186 408494
rect 260422 408258 267186 408494
rect 267422 408258 274186 408494
rect 274422 408258 281186 408494
rect 281422 408258 288186 408494
rect 288422 408258 295186 408494
rect 295422 408258 302186 408494
rect 302422 408258 309186 408494
rect 309422 408258 316186 408494
rect 316422 408258 323186 408494
rect 323422 408258 330186 408494
rect 330422 408258 337186 408494
rect 337422 408258 344186 408494
rect 344422 408258 351186 408494
rect 351422 408258 358186 408494
rect 358422 408258 365186 408494
rect 365422 408258 372186 408494
rect 372422 408258 379186 408494
rect 379422 408258 386186 408494
rect 386422 408258 393186 408494
rect 393422 408258 400186 408494
rect 400422 408258 407186 408494
rect 407422 408258 414186 408494
rect 414422 408258 421186 408494
rect 421422 408258 428186 408494
rect 428422 408258 435186 408494
rect 435422 408258 442186 408494
rect 442422 408258 449186 408494
rect 449422 408258 456186 408494
rect 456422 408258 463186 408494
rect 463422 408258 470186 408494
rect 470422 408258 477186 408494
rect 477422 408258 484186 408494
rect 484422 408258 491186 408494
rect 491422 408258 498186 408494
rect 498422 408258 505186 408494
rect 505422 408258 512186 408494
rect 512422 408258 519186 408494
rect 519422 408258 519952 408494
rect 520188 408258 521884 408494
rect 522120 408258 523816 408494
rect 524052 408258 525748 408494
rect 525984 408258 533186 408494
rect 533422 408258 540186 408494
rect 540422 408258 547186 408494
rect 547422 408258 554186 408494
rect 554422 408258 561186 408494
rect 561422 408258 568186 408494
rect 568422 408258 575186 408494
rect 575422 408258 582186 408494
rect 582422 408258 585818 408494
rect 586054 408258 586138 408494
rect 586374 408258 586458 408494
rect 586694 408258 586778 408494
rect 587014 408258 588874 408494
rect -4950 408216 588874 408258
rect -4950 402434 588874 402476
rect -4950 402198 -4842 402434
rect -4606 402198 -4522 402434
rect -4286 402198 -4202 402434
rect -3966 402198 -3882 402434
rect -3646 402198 2918 402434
rect 3154 402198 9918 402434
rect 10154 402198 16918 402434
rect 17154 402198 23918 402434
rect 24154 402198 30918 402434
rect 31154 402198 37918 402434
rect 38154 402198 44918 402434
rect 45154 402198 51918 402434
rect 52154 402198 58918 402434
rect 59154 402198 65918 402434
rect 66154 402198 72918 402434
rect 73154 402198 79918 402434
rect 80154 402198 86918 402434
rect 87154 402198 93918 402434
rect 94154 402198 100918 402434
rect 101154 402198 107918 402434
rect 108154 402198 114918 402434
rect 115154 402198 121918 402434
rect 122154 402198 128918 402434
rect 129154 402198 135918 402434
rect 136154 402198 142918 402434
rect 143154 402198 149918 402434
rect 150154 402198 156918 402434
rect 157154 402198 163918 402434
rect 164154 402198 170918 402434
rect 171154 402198 177918 402434
rect 178154 402198 184918 402434
rect 185154 402198 191918 402434
rect 192154 402198 198918 402434
rect 199154 402198 205918 402434
rect 206154 402198 212918 402434
rect 213154 402198 219918 402434
rect 220154 402198 226918 402434
rect 227154 402198 233918 402434
rect 234154 402198 240918 402434
rect 241154 402198 247918 402434
rect 248154 402198 254918 402434
rect 255154 402198 261918 402434
rect 262154 402198 268918 402434
rect 269154 402198 275918 402434
rect 276154 402198 282918 402434
rect 283154 402198 289918 402434
rect 290154 402198 296918 402434
rect 297154 402198 303918 402434
rect 304154 402198 310918 402434
rect 311154 402198 317918 402434
rect 318154 402198 324918 402434
rect 325154 402198 331918 402434
rect 332154 402198 338918 402434
rect 339154 402198 345918 402434
rect 346154 402198 352918 402434
rect 353154 402198 359918 402434
rect 360154 402198 366918 402434
rect 367154 402198 373918 402434
rect 374154 402198 380918 402434
rect 381154 402198 387918 402434
rect 388154 402198 394918 402434
rect 395154 402198 401918 402434
rect 402154 402198 408918 402434
rect 409154 402198 415918 402434
rect 416154 402198 422918 402434
rect 423154 402198 429918 402434
rect 430154 402198 436918 402434
rect 437154 402198 443918 402434
rect 444154 402198 450918 402434
rect 451154 402198 457918 402434
rect 458154 402198 464918 402434
rect 465154 402198 471918 402434
rect 472154 402198 478918 402434
rect 479154 402198 485918 402434
rect 486154 402198 492918 402434
rect 493154 402198 499918 402434
rect 500154 402198 506918 402434
rect 507154 402198 513918 402434
rect 514154 402198 520918 402434
rect 521154 402198 522850 402434
rect 523086 402198 524782 402434
rect 525018 402198 526714 402434
rect 526950 402198 527918 402434
rect 528154 402198 534918 402434
rect 535154 402198 541918 402434
rect 542154 402198 548918 402434
rect 549154 402198 555918 402434
rect 556154 402198 562918 402434
rect 563154 402198 569918 402434
rect 570154 402198 576918 402434
rect 577154 402198 587570 402434
rect 587806 402198 587890 402434
rect 588126 402198 588210 402434
rect 588446 402198 588530 402434
rect 588766 402198 588874 402434
rect -4950 402156 588874 402198
rect -4950 401494 588874 401536
rect -4950 401258 -3090 401494
rect -2854 401258 -2770 401494
rect -2534 401258 -2450 401494
rect -2214 401258 -2130 401494
rect -1894 401258 1186 401494
rect 1422 401258 8186 401494
rect 8422 401258 15186 401494
rect 15422 401258 22186 401494
rect 22422 401258 29186 401494
rect 29422 401258 36186 401494
rect 36422 401258 43186 401494
rect 43422 401258 50186 401494
rect 50422 401258 57186 401494
rect 57422 401258 64186 401494
rect 64422 401258 71186 401494
rect 71422 401258 78186 401494
rect 78422 401258 85186 401494
rect 85422 401258 92186 401494
rect 92422 401258 99186 401494
rect 99422 401258 106186 401494
rect 106422 401258 113186 401494
rect 113422 401258 120186 401494
rect 120422 401258 127186 401494
rect 127422 401258 134186 401494
rect 134422 401258 141186 401494
rect 141422 401258 148186 401494
rect 148422 401258 155186 401494
rect 155422 401258 162186 401494
rect 162422 401258 169186 401494
rect 169422 401258 176186 401494
rect 176422 401258 183186 401494
rect 183422 401258 190186 401494
rect 190422 401258 197186 401494
rect 197422 401258 204186 401494
rect 204422 401258 211186 401494
rect 211422 401258 218186 401494
rect 218422 401258 225186 401494
rect 225422 401258 232186 401494
rect 232422 401258 239186 401494
rect 239422 401258 246186 401494
rect 246422 401258 253186 401494
rect 253422 401258 260186 401494
rect 260422 401258 267186 401494
rect 267422 401258 274186 401494
rect 274422 401258 281186 401494
rect 281422 401258 288186 401494
rect 288422 401258 295186 401494
rect 295422 401258 302186 401494
rect 302422 401258 309186 401494
rect 309422 401258 316186 401494
rect 316422 401258 323186 401494
rect 323422 401258 330186 401494
rect 330422 401258 337186 401494
rect 337422 401258 344186 401494
rect 344422 401258 351186 401494
rect 351422 401258 358186 401494
rect 358422 401258 365186 401494
rect 365422 401258 372186 401494
rect 372422 401258 379186 401494
rect 379422 401258 386186 401494
rect 386422 401258 393186 401494
rect 393422 401258 400186 401494
rect 400422 401258 407186 401494
rect 407422 401258 414186 401494
rect 414422 401258 421186 401494
rect 421422 401258 428186 401494
rect 428422 401258 435186 401494
rect 435422 401258 442186 401494
rect 442422 401258 449186 401494
rect 449422 401258 456186 401494
rect 456422 401258 463186 401494
rect 463422 401258 470186 401494
rect 470422 401258 477186 401494
rect 477422 401258 484186 401494
rect 484422 401258 491186 401494
rect 491422 401258 498186 401494
rect 498422 401258 505186 401494
rect 505422 401258 512186 401494
rect 512422 401258 519186 401494
rect 519422 401258 533186 401494
rect 533422 401258 540186 401494
rect 540422 401258 547186 401494
rect 547422 401258 554186 401494
rect 554422 401258 561186 401494
rect 561422 401258 568186 401494
rect 568422 401258 575186 401494
rect 575422 401258 582186 401494
rect 582422 401258 585818 401494
rect 586054 401258 586138 401494
rect 586374 401258 586458 401494
rect 586694 401258 586778 401494
rect 587014 401258 588874 401494
rect -4950 401216 588874 401258
rect -4950 395434 588874 395476
rect -4950 395198 -4842 395434
rect -4606 395198 -4522 395434
rect -4286 395198 -4202 395434
rect -3966 395198 -3882 395434
rect -3646 395198 2918 395434
rect 3154 395198 9918 395434
rect 10154 395198 16918 395434
rect 17154 395198 23918 395434
rect 24154 395198 30918 395434
rect 31154 395198 37918 395434
rect 38154 395198 44918 395434
rect 45154 395198 51918 395434
rect 52154 395198 58918 395434
rect 59154 395198 65918 395434
rect 66154 395198 72918 395434
rect 73154 395198 79918 395434
rect 80154 395198 86918 395434
rect 87154 395198 93918 395434
rect 94154 395198 100918 395434
rect 101154 395198 107918 395434
rect 108154 395198 114918 395434
rect 115154 395198 121918 395434
rect 122154 395198 128918 395434
rect 129154 395198 135918 395434
rect 136154 395198 142918 395434
rect 143154 395198 149918 395434
rect 150154 395198 156918 395434
rect 157154 395198 163918 395434
rect 164154 395198 170918 395434
rect 171154 395198 177918 395434
rect 178154 395198 184918 395434
rect 185154 395198 191918 395434
rect 192154 395198 198918 395434
rect 199154 395198 205918 395434
rect 206154 395198 212918 395434
rect 213154 395198 219918 395434
rect 220154 395198 226918 395434
rect 227154 395198 233918 395434
rect 234154 395198 240918 395434
rect 241154 395198 247918 395434
rect 248154 395198 254918 395434
rect 255154 395198 261918 395434
rect 262154 395198 268918 395434
rect 269154 395198 275918 395434
rect 276154 395198 282918 395434
rect 283154 395198 289918 395434
rect 290154 395198 296918 395434
rect 297154 395198 303918 395434
rect 304154 395198 310918 395434
rect 311154 395198 317918 395434
rect 318154 395198 324918 395434
rect 325154 395198 331918 395434
rect 332154 395198 338918 395434
rect 339154 395198 345918 395434
rect 346154 395198 352918 395434
rect 353154 395198 359918 395434
rect 360154 395198 366918 395434
rect 367154 395198 373918 395434
rect 374154 395198 380918 395434
rect 381154 395198 387918 395434
rect 388154 395198 394918 395434
rect 395154 395198 401918 395434
rect 402154 395198 408918 395434
rect 409154 395198 415918 395434
rect 416154 395198 422918 395434
rect 423154 395198 429918 395434
rect 430154 395198 436918 395434
rect 437154 395198 443918 395434
rect 444154 395198 450918 395434
rect 451154 395198 457918 395434
rect 458154 395198 464918 395434
rect 465154 395198 471918 395434
rect 472154 395198 478918 395434
rect 479154 395198 485918 395434
rect 486154 395198 492918 395434
rect 493154 395198 499918 395434
rect 500154 395198 506918 395434
rect 507154 395198 513918 395434
rect 514154 395198 520918 395434
rect 521154 395198 527918 395434
rect 528154 395198 534918 395434
rect 535154 395198 541918 395434
rect 542154 395198 548918 395434
rect 549154 395198 555918 395434
rect 556154 395198 562918 395434
rect 563154 395198 569918 395434
rect 570154 395198 576918 395434
rect 577154 395198 587570 395434
rect 587806 395198 587890 395434
rect 588126 395198 588210 395434
rect 588446 395198 588530 395434
rect 588766 395198 588874 395434
rect -4950 395156 588874 395198
rect -4950 394494 588874 394536
rect -4950 394258 -3090 394494
rect -2854 394258 -2770 394494
rect -2534 394258 -2450 394494
rect -2214 394258 -2130 394494
rect -1894 394258 1186 394494
rect 1422 394258 8186 394494
rect 8422 394258 15186 394494
rect 15422 394258 22186 394494
rect 22422 394258 29186 394494
rect 29422 394258 36186 394494
rect 36422 394258 43186 394494
rect 43422 394258 50186 394494
rect 50422 394258 57186 394494
rect 57422 394258 64186 394494
rect 64422 394258 71186 394494
rect 71422 394258 78186 394494
rect 78422 394258 85186 394494
rect 85422 394258 92186 394494
rect 92422 394258 99186 394494
rect 99422 394258 106186 394494
rect 106422 394258 113186 394494
rect 113422 394258 120186 394494
rect 120422 394258 127186 394494
rect 127422 394258 134186 394494
rect 134422 394258 141186 394494
rect 141422 394258 148186 394494
rect 148422 394258 155186 394494
rect 155422 394258 162186 394494
rect 162422 394258 169186 394494
rect 169422 394258 176186 394494
rect 176422 394258 183186 394494
rect 183422 394258 190186 394494
rect 190422 394258 197186 394494
rect 197422 394258 204186 394494
rect 204422 394258 211186 394494
rect 211422 394258 218186 394494
rect 218422 394258 225186 394494
rect 225422 394258 232186 394494
rect 232422 394258 239186 394494
rect 239422 394258 246186 394494
rect 246422 394258 253186 394494
rect 253422 394258 260186 394494
rect 260422 394258 267186 394494
rect 267422 394258 274186 394494
rect 274422 394258 281186 394494
rect 281422 394258 288186 394494
rect 288422 394258 295186 394494
rect 295422 394258 302186 394494
rect 302422 394258 309186 394494
rect 309422 394258 316186 394494
rect 316422 394258 323186 394494
rect 323422 394258 330186 394494
rect 330422 394258 337186 394494
rect 337422 394258 344186 394494
rect 344422 394258 351186 394494
rect 351422 394258 358186 394494
rect 358422 394258 365186 394494
rect 365422 394258 372186 394494
rect 372422 394258 379186 394494
rect 379422 394258 386186 394494
rect 386422 394258 393186 394494
rect 393422 394258 400186 394494
rect 400422 394258 407186 394494
rect 407422 394258 414186 394494
rect 414422 394258 421186 394494
rect 421422 394258 428186 394494
rect 428422 394258 435186 394494
rect 435422 394258 442186 394494
rect 442422 394258 449186 394494
rect 449422 394258 456186 394494
rect 456422 394258 463186 394494
rect 463422 394258 470186 394494
rect 470422 394258 477186 394494
rect 477422 394258 484186 394494
rect 484422 394258 491186 394494
rect 491422 394258 498186 394494
rect 498422 394258 505186 394494
rect 505422 394258 512186 394494
rect 512422 394258 519186 394494
rect 519422 394258 526186 394494
rect 526422 394258 533186 394494
rect 533422 394258 540186 394494
rect 540422 394258 547186 394494
rect 547422 394258 554186 394494
rect 554422 394258 561186 394494
rect 561422 394258 568186 394494
rect 568422 394258 575186 394494
rect 575422 394258 582186 394494
rect 582422 394258 585818 394494
rect 586054 394258 586138 394494
rect 586374 394258 586458 394494
rect 586694 394258 586778 394494
rect 587014 394258 588874 394494
rect -4950 394216 588874 394258
rect -4950 388434 588874 388476
rect -4950 388198 -4842 388434
rect -4606 388198 -4522 388434
rect -4286 388198 -4202 388434
rect -3966 388198 -3882 388434
rect -3646 388198 2918 388434
rect 3154 388198 9918 388434
rect 10154 388198 16918 388434
rect 17154 388198 23918 388434
rect 24154 388198 30918 388434
rect 31154 388198 37918 388434
rect 38154 388198 44918 388434
rect 45154 388198 51918 388434
rect 52154 388198 58918 388434
rect 59154 388198 65918 388434
rect 66154 388198 72918 388434
rect 73154 388198 79918 388434
rect 80154 388198 86918 388434
rect 87154 388198 93918 388434
rect 94154 388198 100918 388434
rect 101154 388198 107918 388434
rect 108154 388198 114918 388434
rect 115154 388198 121918 388434
rect 122154 388198 128918 388434
rect 129154 388198 135918 388434
rect 136154 388198 142918 388434
rect 143154 388198 149918 388434
rect 150154 388198 156918 388434
rect 157154 388198 163918 388434
rect 164154 388198 170918 388434
rect 171154 388198 177918 388434
rect 178154 388198 184918 388434
rect 185154 388198 191918 388434
rect 192154 388198 198918 388434
rect 199154 388198 205918 388434
rect 206154 388198 212918 388434
rect 213154 388198 219918 388434
rect 220154 388198 226918 388434
rect 227154 388198 233918 388434
rect 234154 388198 240918 388434
rect 241154 388198 247918 388434
rect 248154 388198 254918 388434
rect 255154 388198 261918 388434
rect 262154 388198 268918 388434
rect 269154 388198 275918 388434
rect 276154 388198 282918 388434
rect 283154 388198 289918 388434
rect 290154 388198 296918 388434
rect 297154 388198 303918 388434
rect 304154 388198 310918 388434
rect 311154 388198 317918 388434
rect 318154 388198 324918 388434
rect 325154 388198 331918 388434
rect 332154 388198 338918 388434
rect 339154 388198 345918 388434
rect 346154 388198 352918 388434
rect 353154 388198 359918 388434
rect 360154 388198 366918 388434
rect 367154 388198 373918 388434
rect 374154 388198 380918 388434
rect 381154 388198 387918 388434
rect 388154 388198 394918 388434
rect 395154 388198 401918 388434
rect 402154 388198 408918 388434
rect 409154 388198 415918 388434
rect 416154 388198 422918 388434
rect 423154 388198 429918 388434
rect 430154 388198 436918 388434
rect 437154 388198 443918 388434
rect 444154 388198 450918 388434
rect 451154 388198 457918 388434
rect 458154 388198 464918 388434
rect 465154 388198 471918 388434
rect 472154 388198 478918 388434
rect 479154 388198 485918 388434
rect 486154 388198 492918 388434
rect 493154 388198 499918 388434
rect 500154 388198 506918 388434
rect 507154 388198 513918 388434
rect 514154 388198 520918 388434
rect 521154 388198 527918 388434
rect 528154 388198 534918 388434
rect 535154 388198 541918 388434
rect 542154 388198 548918 388434
rect 549154 388198 555918 388434
rect 556154 388198 562918 388434
rect 563154 388198 569918 388434
rect 570154 388198 576918 388434
rect 577154 388198 587570 388434
rect 587806 388198 587890 388434
rect 588126 388198 588210 388434
rect 588446 388198 588530 388434
rect 588766 388198 588874 388434
rect -4950 388156 588874 388198
rect -4950 387494 588874 387536
rect -4950 387258 -3090 387494
rect -2854 387258 -2770 387494
rect -2534 387258 -2450 387494
rect -2214 387258 -2130 387494
rect -1894 387258 1186 387494
rect 1422 387258 8186 387494
rect 8422 387258 15186 387494
rect 15422 387258 22186 387494
rect 22422 387258 29186 387494
rect 29422 387258 36186 387494
rect 36422 387258 43186 387494
rect 43422 387258 50186 387494
rect 50422 387258 57186 387494
rect 57422 387258 64186 387494
rect 64422 387258 71186 387494
rect 71422 387258 78186 387494
rect 78422 387258 85186 387494
rect 85422 387258 92186 387494
rect 92422 387258 99186 387494
rect 99422 387258 106186 387494
rect 106422 387258 113186 387494
rect 113422 387258 120186 387494
rect 120422 387258 127186 387494
rect 127422 387258 134186 387494
rect 134422 387258 141186 387494
rect 141422 387258 148186 387494
rect 148422 387258 155186 387494
rect 155422 387258 162186 387494
rect 162422 387258 169186 387494
rect 169422 387258 176186 387494
rect 176422 387258 183186 387494
rect 183422 387258 190186 387494
rect 190422 387258 197186 387494
rect 197422 387258 204186 387494
rect 204422 387258 211186 387494
rect 211422 387258 218186 387494
rect 218422 387258 225186 387494
rect 225422 387258 232186 387494
rect 232422 387258 239186 387494
rect 239422 387258 246186 387494
rect 246422 387258 253186 387494
rect 253422 387258 260186 387494
rect 260422 387258 267186 387494
rect 267422 387258 274186 387494
rect 274422 387258 281186 387494
rect 281422 387258 288186 387494
rect 288422 387258 295186 387494
rect 295422 387258 302186 387494
rect 302422 387258 309186 387494
rect 309422 387258 316186 387494
rect 316422 387258 323186 387494
rect 323422 387258 330186 387494
rect 330422 387258 337186 387494
rect 337422 387258 344186 387494
rect 344422 387258 351186 387494
rect 351422 387258 358186 387494
rect 358422 387258 365186 387494
rect 365422 387258 372186 387494
rect 372422 387258 379186 387494
rect 379422 387258 386186 387494
rect 386422 387258 393186 387494
rect 393422 387258 400186 387494
rect 400422 387258 407186 387494
rect 407422 387258 414186 387494
rect 414422 387258 421186 387494
rect 421422 387258 428186 387494
rect 428422 387258 435186 387494
rect 435422 387258 442186 387494
rect 442422 387258 449186 387494
rect 449422 387258 456186 387494
rect 456422 387258 463186 387494
rect 463422 387258 470186 387494
rect 470422 387258 477186 387494
rect 477422 387258 484186 387494
rect 484422 387258 491186 387494
rect 491422 387258 498186 387494
rect 498422 387258 505186 387494
rect 505422 387258 512186 387494
rect 512422 387258 519186 387494
rect 519422 387258 526186 387494
rect 526422 387258 533186 387494
rect 533422 387258 540186 387494
rect 540422 387258 547186 387494
rect 547422 387258 554186 387494
rect 554422 387258 561186 387494
rect 561422 387258 568186 387494
rect 568422 387258 575186 387494
rect 575422 387258 582186 387494
rect 582422 387258 585818 387494
rect 586054 387258 586138 387494
rect 586374 387258 586458 387494
rect 586694 387258 586778 387494
rect 587014 387258 588874 387494
rect -4950 387216 588874 387258
rect -4950 381434 588874 381476
rect -4950 381198 -4842 381434
rect -4606 381198 -4522 381434
rect -4286 381198 -4202 381434
rect -3966 381198 -3882 381434
rect -3646 381198 2918 381434
rect 3154 381198 9918 381434
rect 10154 381198 16918 381434
rect 17154 381198 23918 381434
rect 24154 381198 30918 381434
rect 31154 381198 37918 381434
rect 38154 381198 44918 381434
rect 45154 381198 51918 381434
rect 52154 381198 58918 381434
rect 59154 381198 65918 381434
rect 66154 381198 72918 381434
rect 73154 381198 79918 381434
rect 80154 381198 86918 381434
rect 87154 381198 93918 381434
rect 94154 381198 100918 381434
rect 101154 381198 107918 381434
rect 108154 381198 114918 381434
rect 115154 381198 121918 381434
rect 122154 381198 128918 381434
rect 129154 381198 135918 381434
rect 136154 381198 142918 381434
rect 143154 381198 149918 381434
rect 150154 381198 156918 381434
rect 157154 381198 163918 381434
rect 164154 381198 170918 381434
rect 171154 381198 177918 381434
rect 178154 381198 184918 381434
rect 185154 381198 191918 381434
rect 192154 381198 198918 381434
rect 199154 381198 205918 381434
rect 206154 381198 212918 381434
rect 213154 381198 219918 381434
rect 220154 381198 226918 381434
rect 227154 381198 233918 381434
rect 234154 381198 240918 381434
rect 241154 381198 247918 381434
rect 248154 381198 254918 381434
rect 255154 381198 261918 381434
rect 262154 381198 268918 381434
rect 269154 381198 275918 381434
rect 276154 381198 282918 381434
rect 283154 381198 289918 381434
rect 290154 381198 296918 381434
rect 297154 381198 303918 381434
rect 304154 381198 310918 381434
rect 311154 381198 317918 381434
rect 318154 381198 324918 381434
rect 325154 381198 331918 381434
rect 332154 381198 338918 381434
rect 339154 381198 345918 381434
rect 346154 381198 352918 381434
rect 353154 381198 359918 381434
rect 360154 381198 366918 381434
rect 367154 381198 373918 381434
rect 374154 381198 380918 381434
rect 381154 381198 387918 381434
rect 388154 381198 394918 381434
rect 395154 381198 401918 381434
rect 402154 381198 408918 381434
rect 409154 381198 415918 381434
rect 416154 381198 422918 381434
rect 423154 381198 429918 381434
rect 430154 381198 436918 381434
rect 437154 381198 443918 381434
rect 444154 381198 450918 381434
rect 451154 381198 457918 381434
rect 458154 381198 464918 381434
rect 465154 381198 471918 381434
rect 472154 381198 478918 381434
rect 479154 381198 485918 381434
rect 486154 381198 492918 381434
rect 493154 381198 499918 381434
rect 500154 381198 506918 381434
rect 507154 381198 513918 381434
rect 514154 381198 527918 381434
rect 528154 381198 534918 381434
rect 535154 381198 541918 381434
rect 542154 381198 548918 381434
rect 549154 381198 555918 381434
rect 556154 381198 562918 381434
rect 563154 381198 569918 381434
rect 570154 381198 576918 381434
rect 577154 381198 587570 381434
rect 587806 381198 587890 381434
rect 588126 381198 588210 381434
rect 588446 381198 588530 381434
rect 588766 381198 588874 381434
rect -4950 381156 588874 381198
rect -4950 380494 588874 380536
rect -4950 380258 -3090 380494
rect -2854 380258 -2770 380494
rect -2534 380258 -2450 380494
rect -2214 380258 -2130 380494
rect -1894 380258 1186 380494
rect 1422 380258 8186 380494
rect 8422 380258 15186 380494
rect 15422 380258 22186 380494
rect 22422 380258 29186 380494
rect 29422 380258 36186 380494
rect 36422 380258 43186 380494
rect 43422 380258 50186 380494
rect 50422 380258 57186 380494
rect 57422 380258 64186 380494
rect 64422 380258 71186 380494
rect 71422 380258 78186 380494
rect 78422 380258 85186 380494
rect 85422 380258 92186 380494
rect 92422 380258 99186 380494
rect 99422 380258 106186 380494
rect 106422 380258 113186 380494
rect 113422 380258 120186 380494
rect 120422 380258 127186 380494
rect 127422 380258 134186 380494
rect 134422 380258 141186 380494
rect 141422 380258 148186 380494
rect 148422 380258 155186 380494
rect 155422 380258 162186 380494
rect 162422 380258 169186 380494
rect 169422 380258 176186 380494
rect 176422 380258 183186 380494
rect 183422 380258 190186 380494
rect 190422 380258 197186 380494
rect 197422 380258 204186 380494
rect 204422 380258 211186 380494
rect 211422 380258 218186 380494
rect 218422 380258 225186 380494
rect 225422 380258 232186 380494
rect 232422 380258 239186 380494
rect 239422 380258 246186 380494
rect 246422 380258 253186 380494
rect 253422 380258 260186 380494
rect 260422 380258 267186 380494
rect 267422 380258 274186 380494
rect 274422 380258 281186 380494
rect 281422 380258 288186 380494
rect 288422 380258 295186 380494
rect 295422 380258 302186 380494
rect 302422 380258 309186 380494
rect 309422 380258 316186 380494
rect 316422 380258 323186 380494
rect 323422 380258 330186 380494
rect 330422 380258 337186 380494
rect 337422 380258 344186 380494
rect 344422 380258 351186 380494
rect 351422 380258 358186 380494
rect 358422 380258 365186 380494
rect 365422 380258 372186 380494
rect 372422 380258 379186 380494
rect 379422 380258 386186 380494
rect 386422 380258 393186 380494
rect 393422 380258 400186 380494
rect 400422 380258 407186 380494
rect 407422 380258 414186 380494
rect 414422 380258 421186 380494
rect 421422 380258 428186 380494
rect 428422 380258 435186 380494
rect 435422 380258 442186 380494
rect 442422 380258 449186 380494
rect 449422 380258 456186 380494
rect 456422 380258 463186 380494
rect 463422 380258 470186 380494
rect 470422 380258 477186 380494
rect 477422 380258 484186 380494
rect 484422 380258 491186 380494
rect 491422 380258 498186 380494
rect 498422 380258 505186 380494
rect 505422 380258 512186 380494
rect 512422 380258 519186 380494
rect 519422 380258 533186 380494
rect 533422 380258 540186 380494
rect 540422 380258 547186 380494
rect 547422 380258 554186 380494
rect 554422 380258 561186 380494
rect 561422 380258 568186 380494
rect 568422 380258 575186 380494
rect 575422 380258 582186 380494
rect 582422 380258 585818 380494
rect 586054 380258 586138 380494
rect 586374 380258 586458 380494
rect 586694 380258 586778 380494
rect 587014 380258 588874 380494
rect -4950 380216 588874 380258
rect -4950 374434 588874 374476
rect -4950 374198 -4842 374434
rect -4606 374198 -4522 374434
rect -4286 374198 -4202 374434
rect -3966 374198 -3882 374434
rect -3646 374198 2918 374434
rect 3154 374198 9918 374434
rect 10154 374198 16918 374434
rect 17154 374198 23918 374434
rect 24154 374198 30918 374434
rect 31154 374198 37918 374434
rect 38154 374198 44918 374434
rect 45154 374198 51918 374434
rect 52154 374198 58918 374434
rect 59154 374198 65918 374434
rect 66154 374198 72918 374434
rect 73154 374198 79918 374434
rect 80154 374198 86918 374434
rect 87154 374198 93918 374434
rect 94154 374198 100918 374434
rect 101154 374198 107918 374434
rect 108154 374198 114918 374434
rect 115154 374198 121918 374434
rect 122154 374198 128918 374434
rect 129154 374198 135918 374434
rect 136154 374198 142918 374434
rect 143154 374198 149918 374434
rect 150154 374198 156918 374434
rect 157154 374198 163918 374434
rect 164154 374198 170918 374434
rect 171154 374198 177918 374434
rect 178154 374198 184918 374434
rect 185154 374198 191918 374434
rect 192154 374198 198918 374434
rect 199154 374198 205918 374434
rect 206154 374198 212918 374434
rect 213154 374198 219918 374434
rect 220154 374198 226918 374434
rect 227154 374198 233918 374434
rect 234154 374198 240918 374434
rect 241154 374198 247918 374434
rect 248154 374198 254918 374434
rect 255154 374198 261918 374434
rect 262154 374198 268918 374434
rect 269154 374198 275918 374434
rect 276154 374198 282918 374434
rect 283154 374198 289918 374434
rect 290154 374198 296918 374434
rect 297154 374198 303918 374434
rect 304154 374198 310918 374434
rect 311154 374198 317918 374434
rect 318154 374198 324918 374434
rect 325154 374198 331918 374434
rect 332154 374198 338918 374434
rect 339154 374198 345918 374434
rect 346154 374198 352918 374434
rect 353154 374198 359918 374434
rect 360154 374198 366918 374434
rect 367154 374198 373918 374434
rect 374154 374198 380918 374434
rect 381154 374198 387918 374434
rect 388154 374198 394918 374434
rect 395154 374198 401918 374434
rect 402154 374198 408918 374434
rect 409154 374198 415918 374434
rect 416154 374198 422918 374434
rect 423154 374198 429918 374434
rect 430154 374198 436918 374434
rect 437154 374198 443918 374434
rect 444154 374198 450918 374434
rect 451154 374198 457918 374434
rect 458154 374198 464918 374434
rect 465154 374198 471918 374434
rect 472154 374198 478918 374434
rect 479154 374198 485918 374434
rect 486154 374198 492918 374434
rect 493154 374198 499918 374434
rect 500154 374198 506918 374434
rect 507154 374198 513918 374434
rect 514154 374198 520918 374434
rect 521154 374198 522850 374434
rect 523086 374198 524782 374434
rect 525018 374198 526714 374434
rect 526950 374198 527918 374434
rect 528154 374198 534918 374434
rect 535154 374198 541918 374434
rect 542154 374198 548918 374434
rect 549154 374198 555918 374434
rect 556154 374198 562918 374434
rect 563154 374198 569918 374434
rect 570154 374198 576918 374434
rect 577154 374198 587570 374434
rect 587806 374198 587890 374434
rect 588126 374198 588210 374434
rect 588446 374198 588530 374434
rect 588766 374198 588874 374434
rect -4950 374156 588874 374198
rect -4950 373494 588874 373536
rect -4950 373258 -3090 373494
rect -2854 373258 -2770 373494
rect -2534 373258 -2450 373494
rect -2214 373258 -2130 373494
rect -1894 373258 1186 373494
rect 1422 373258 8186 373494
rect 8422 373258 15186 373494
rect 15422 373258 22186 373494
rect 22422 373258 29186 373494
rect 29422 373258 36186 373494
rect 36422 373258 43186 373494
rect 43422 373258 50186 373494
rect 50422 373258 57186 373494
rect 57422 373258 64186 373494
rect 64422 373258 71186 373494
rect 71422 373258 78186 373494
rect 78422 373258 85186 373494
rect 85422 373258 92186 373494
rect 92422 373258 99186 373494
rect 99422 373258 106186 373494
rect 106422 373258 113186 373494
rect 113422 373258 120186 373494
rect 120422 373258 127186 373494
rect 127422 373258 134186 373494
rect 134422 373258 141186 373494
rect 141422 373258 148186 373494
rect 148422 373258 155186 373494
rect 155422 373258 162186 373494
rect 162422 373258 169186 373494
rect 169422 373258 176186 373494
rect 176422 373258 183186 373494
rect 183422 373258 190186 373494
rect 190422 373258 197186 373494
rect 197422 373258 204186 373494
rect 204422 373258 211186 373494
rect 211422 373258 218186 373494
rect 218422 373258 225186 373494
rect 225422 373258 232186 373494
rect 232422 373258 239186 373494
rect 239422 373258 246186 373494
rect 246422 373258 253186 373494
rect 253422 373258 260186 373494
rect 260422 373258 267186 373494
rect 267422 373258 274186 373494
rect 274422 373258 281186 373494
rect 281422 373258 288186 373494
rect 288422 373258 295186 373494
rect 295422 373258 302186 373494
rect 302422 373258 309186 373494
rect 309422 373258 316186 373494
rect 316422 373258 323186 373494
rect 323422 373258 330186 373494
rect 330422 373258 337186 373494
rect 337422 373258 344186 373494
rect 344422 373258 351186 373494
rect 351422 373258 358186 373494
rect 358422 373258 365186 373494
rect 365422 373258 372186 373494
rect 372422 373258 379186 373494
rect 379422 373258 386186 373494
rect 386422 373258 393186 373494
rect 393422 373258 400186 373494
rect 400422 373258 407186 373494
rect 407422 373258 414186 373494
rect 414422 373258 421186 373494
rect 421422 373258 428186 373494
rect 428422 373258 435186 373494
rect 435422 373258 442186 373494
rect 442422 373258 449186 373494
rect 449422 373258 456186 373494
rect 456422 373258 463186 373494
rect 463422 373258 470186 373494
rect 470422 373258 477186 373494
rect 477422 373258 484186 373494
rect 484422 373258 491186 373494
rect 491422 373258 498186 373494
rect 498422 373258 505186 373494
rect 505422 373258 512186 373494
rect 512422 373258 519186 373494
rect 519422 373258 519952 373494
rect 520188 373258 521884 373494
rect 522120 373258 523816 373494
rect 524052 373258 525748 373494
rect 525984 373258 533186 373494
rect 533422 373258 540186 373494
rect 540422 373258 547186 373494
rect 547422 373258 554186 373494
rect 554422 373258 561186 373494
rect 561422 373258 568186 373494
rect 568422 373258 575186 373494
rect 575422 373258 582186 373494
rect 582422 373258 585818 373494
rect 586054 373258 586138 373494
rect 586374 373258 586458 373494
rect 586694 373258 586778 373494
rect 587014 373258 588874 373494
rect -4950 373216 588874 373258
rect -4950 367434 588874 367476
rect -4950 367198 -4842 367434
rect -4606 367198 -4522 367434
rect -4286 367198 -4202 367434
rect -3966 367198 -3882 367434
rect -3646 367198 2918 367434
rect 3154 367198 9918 367434
rect 10154 367198 16918 367434
rect 17154 367198 23918 367434
rect 24154 367198 30918 367434
rect 31154 367198 37918 367434
rect 38154 367198 44918 367434
rect 45154 367198 51918 367434
rect 52154 367198 58918 367434
rect 59154 367198 65918 367434
rect 66154 367198 72918 367434
rect 73154 367198 79918 367434
rect 80154 367198 86918 367434
rect 87154 367198 93918 367434
rect 94154 367198 100918 367434
rect 101154 367198 107918 367434
rect 108154 367198 114918 367434
rect 115154 367198 121918 367434
rect 122154 367198 128918 367434
rect 129154 367198 135918 367434
rect 136154 367198 142918 367434
rect 143154 367198 149918 367434
rect 150154 367198 156918 367434
rect 157154 367198 163918 367434
rect 164154 367198 170918 367434
rect 171154 367198 177918 367434
rect 178154 367198 184918 367434
rect 185154 367198 191918 367434
rect 192154 367198 198918 367434
rect 199154 367198 205918 367434
rect 206154 367198 212918 367434
rect 213154 367198 219918 367434
rect 220154 367198 226918 367434
rect 227154 367198 233918 367434
rect 234154 367198 240918 367434
rect 241154 367198 247918 367434
rect 248154 367198 254918 367434
rect 255154 367198 261918 367434
rect 262154 367198 268918 367434
rect 269154 367198 275918 367434
rect 276154 367198 282918 367434
rect 283154 367198 289918 367434
rect 290154 367198 310918 367434
rect 311154 367198 317918 367434
rect 318154 367198 324918 367434
rect 325154 367198 331918 367434
rect 332154 367198 338918 367434
rect 339154 367198 345918 367434
rect 346154 367198 352918 367434
rect 353154 367198 359918 367434
rect 360154 367198 366918 367434
rect 367154 367198 373918 367434
rect 374154 367198 380918 367434
rect 381154 367198 387918 367434
rect 388154 367198 394918 367434
rect 395154 367198 401918 367434
rect 402154 367198 408918 367434
rect 409154 367198 415918 367434
rect 416154 367198 422918 367434
rect 423154 367198 429918 367434
rect 430154 367198 436918 367434
rect 437154 367198 443918 367434
rect 444154 367198 450918 367434
rect 451154 367198 457918 367434
rect 458154 367198 464918 367434
rect 465154 367198 471918 367434
rect 472154 367198 478918 367434
rect 479154 367198 485918 367434
rect 486154 367198 492918 367434
rect 493154 367198 499918 367434
rect 500154 367198 506918 367434
rect 507154 367198 513918 367434
rect 514154 367198 520918 367434
rect 521154 367198 522850 367434
rect 523086 367198 524782 367434
rect 525018 367198 526714 367434
rect 526950 367198 527918 367434
rect 528154 367198 534918 367434
rect 535154 367198 541918 367434
rect 542154 367198 548918 367434
rect 549154 367198 555918 367434
rect 556154 367198 562918 367434
rect 563154 367198 569918 367434
rect 570154 367198 576918 367434
rect 577154 367198 587570 367434
rect 587806 367198 587890 367434
rect 588126 367198 588210 367434
rect 588446 367198 588530 367434
rect 588766 367198 588874 367434
rect -4950 367156 588874 367198
rect -4950 366494 588874 366536
rect -4950 366258 -3090 366494
rect -2854 366258 -2770 366494
rect -2534 366258 -2450 366494
rect -2214 366258 -2130 366494
rect -1894 366258 1186 366494
rect 1422 366258 8186 366494
rect 8422 366258 15186 366494
rect 15422 366258 22186 366494
rect 22422 366258 29186 366494
rect 29422 366258 36186 366494
rect 36422 366258 43186 366494
rect 43422 366258 50186 366494
rect 50422 366258 57186 366494
rect 57422 366258 64186 366494
rect 64422 366258 71186 366494
rect 71422 366258 78186 366494
rect 78422 366258 85186 366494
rect 85422 366258 92186 366494
rect 92422 366258 99186 366494
rect 99422 366258 106186 366494
rect 106422 366258 113186 366494
rect 113422 366258 120186 366494
rect 120422 366258 127186 366494
rect 127422 366258 134186 366494
rect 134422 366258 141186 366494
rect 141422 366258 148186 366494
rect 148422 366258 155186 366494
rect 155422 366258 162186 366494
rect 162422 366258 169186 366494
rect 169422 366258 176186 366494
rect 176422 366258 183186 366494
rect 183422 366258 190186 366494
rect 190422 366258 197186 366494
rect 197422 366258 204186 366494
rect 204422 366258 211186 366494
rect 211422 366258 218186 366494
rect 218422 366258 225186 366494
rect 225422 366258 232186 366494
rect 232422 366258 239186 366494
rect 239422 366258 246186 366494
rect 246422 366258 253186 366494
rect 253422 366258 260186 366494
rect 260422 366258 267186 366494
rect 267422 366258 274186 366494
rect 274422 366258 281186 366494
rect 281422 366258 288186 366494
rect 288422 366258 309186 366494
rect 309422 366258 316186 366494
rect 316422 366258 323186 366494
rect 323422 366258 330186 366494
rect 330422 366258 337186 366494
rect 337422 366258 344186 366494
rect 344422 366258 351186 366494
rect 351422 366258 358186 366494
rect 358422 366258 365186 366494
rect 365422 366258 372186 366494
rect 372422 366258 379186 366494
rect 379422 366258 386186 366494
rect 386422 366258 393186 366494
rect 393422 366258 400186 366494
rect 400422 366258 407186 366494
rect 407422 366258 414186 366494
rect 414422 366258 421186 366494
rect 421422 366258 428186 366494
rect 428422 366258 435186 366494
rect 435422 366258 442186 366494
rect 442422 366258 449186 366494
rect 449422 366258 456186 366494
rect 456422 366258 463186 366494
rect 463422 366258 470186 366494
rect 470422 366258 477186 366494
rect 477422 366258 484186 366494
rect 484422 366258 491186 366494
rect 491422 366258 498186 366494
rect 498422 366258 505186 366494
rect 505422 366258 512186 366494
rect 512422 366258 519186 366494
rect 519422 366258 519952 366494
rect 520188 366258 521884 366494
rect 522120 366258 523816 366494
rect 524052 366258 525748 366494
rect 525984 366258 533186 366494
rect 533422 366258 540186 366494
rect 540422 366258 547186 366494
rect 547422 366258 554186 366494
rect 554422 366258 561186 366494
rect 561422 366258 568186 366494
rect 568422 366258 575186 366494
rect 575422 366258 582186 366494
rect 582422 366258 585818 366494
rect 586054 366258 586138 366494
rect 586374 366258 586458 366494
rect 586694 366258 586778 366494
rect 587014 366258 588874 366494
rect -4950 366216 588874 366258
rect -4950 360434 588874 360476
rect -4950 360198 -4842 360434
rect -4606 360198 -4522 360434
rect -4286 360198 -4202 360434
rect -3966 360198 -3882 360434
rect -3646 360198 2918 360434
rect 3154 360198 9918 360434
rect 10154 360198 16918 360434
rect 17154 360198 23918 360434
rect 24154 360198 30918 360434
rect 31154 360198 37918 360434
rect 38154 360198 44918 360434
rect 45154 360198 51918 360434
rect 52154 360198 58918 360434
rect 59154 360198 65918 360434
rect 66154 360198 72918 360434
rect 73154 360198 79918 360434
rect 80154 360198 86918 360434
rect 87154 360198 93918 360434
rect 94154 360198 100918 360434
rect 101154 360198 107918 360434
rect 108154 360198 114918 360434
rect 115154 360198 121918 360434
rect 122154 360198 128918 360434
rect 129154 360198 135918 360434
rect 136154 360198 142918 360434
rect 143154 360198 149918 360434
rect 150154 360198 156918 360434
rect 157154 360198 163918 360434
rect 164154 360198 170918 360434
rect 171154 360198 177918 360434
rect 178154 360198 184918 360434
rect 185154 360198 191918 360434
rect 192154 360198 198918 360434
rect 199154 360198 205918 360434
rect 206154 360198 212918 360434
rect 213154 360198 219918 360434
rect 220154 360198 226918 360434
rect 227154 360198 233918 360434
rect 234154 360198 240918 360434
rect 241154 360198 247918 360434
rect 248154 360198 254918 360434
rect 255154 360198 261918 360434
rect 262154 360198 268918 360434
rect 269154 360198 275918 360434
rect 276154 360198 282918 360434
rect 283154 360198 289918 360434
rect 290154 360198 296918 360434
rect 297154 360198 303918 360434
rect 304154 360198 310918 360434
rect 311154 360198 317918 360434
rect 318154 360198 324918 360434
rect 325154 360198 331918 360434
rect 332154 360198 338918 360434
rect 339154 360198 345918 360434
rect 346154 360198 352918 360434
rect 353154 360198 359918 360434
rect 360154 360198 366918 360434
rect 367154 360198 373918 360434
rect 374154 360198 380918 360434
rect 381154 360198 387918 360434
rect 388154 360198 394918 360434
rect 395154 360198 401918 360434
rect 402154 360198 408918 360434
rect 409154 360198 415918 360434
rect 416154 360198 422918 360434
rect 423154 360198 429918 360434
rect 430154 360198 436918 360434
rect 437154 360198 443918 360434
rect 444154 360198 450918 360434
rect 451154 360198 457918 360434
rect 458154 360198 464918 360434
rect 465154 360198 471918 360434
rect 472154 360198 478918 360434
rect 479154 360198 485918 360434
rect 486154 360198 492918 360434
rect 493154 360198 499918 360434
rect 500154 360198 506918 360434
rect 507154 360198 513918 360434
rect 514154 360198 527918 360434
rect 528154 360198 534918 360434
rect 535154 360198 541918 360434
rect 542154 360198 548918 360434
rect 549154 360198 555918 360434
rect 556154 360198 562918 360434
rect 563154 360198 569918 360434
rect 570154 360198 576918 360434
rect 577154 360198 587570 360434
rect 587806 360198 587890 360434
rect 588126 360198 588210 360434
rect 588446 360198 588530 360434
rect 588766 360198 588874 360434
rect -4950 360156 588874 360198
rect -4950 359494 588874 359536
rect -4950 359258 -3090 359494
rect -2854 359258 -2770 359494
rect -2534 359258 -2450 359494
rect -2214 359258 -2130 359494
rect -1894 359258 1186 359494
rect 1422 359258 8186 359494
rect 8422 359258 15186 359494
rect 15422 359258 22186 359494
rect 22422 359258 29186 359494
rect 29422 359258 36186 359494
rect 36422 359258 43186 359494
rect 43422 359258 50186 359494
rect 50422 359258 57186 359494
rect 57422 359258 64186 359494
rect 64422 359258 71186 359494
rect 71422 359258 78186 359494
rect 78422 359258 85186 359494
rect 85422 359258 92186 359494
rect 92422 359258 99186 359494
rect 99422 359258 106186 359494
rect 106422 359258 113186 359494
rect 113422 359258 120186 359494
rect 120422 359258 127186 359494
rect 127422 359258 134186 359494
rect 134422 359258 141186 359494
rect 141422 359258 148186 359494
rect 148422 359258 155186 359494
rect 155422 359258 162186 359494
rect 162422 359258 169186 359494
rect 169422 359258 176186 359494
rect 176422 359258 183186 359494
rect 183422 359258 190186 359494
rect 190422 359258 197186 359494
rect 197422 359258 204186 359494
rect 204422 359258 211186 359494
rect 211422 359258 218186 359494
rect 218422 359258 225186 359494
rect 225422 359258 232186 359494
rect 232422 359258 239186 359494
rect 239422 359258 246186 359494
rect 246422 359258 253186 359494
rect 253422 359258 260186 359494
rect 260422 359258 267186 359494
rect 267422 359258 274186 359494
rect 274422 359258 281186 359494
rect 281422 359258 288186 359494
rect 288422 359258 295186 359494
rect 295422 359258 302186 359494
rect 302422 359258 309186 359494
rect 309422 359258 316186 359494
rect 316422 359258 323186 359494
rect 323422 359258 330186 359494
rect 330422 359258 337186 359494
rect 337422 359258 344186 359494
rect 344422 359258 351186 359494
rect 351422 359258 358186 359494
rect 358422 359258 365186 359494
rect 365422 359258 372186 359494
rect 372422 359258 379186 359494
rect 379422 359258 386186 359494
rect 386422 359258 393186 359494
rect 393422 359258 400186 359494
rect 400422 359258 407186 359494
rect 407422 359258 414186 359494
rect 414422 359258 421186 359494
rect 421422 359258 428186 359494
rect 428422 359258 435186 359494
rect 435422 359258 442186 359494
rect 442422 359258 449186 359494
rect 449422 359258 456186 359494
rect 456422 359258 463186 359494
rect 463422 359258 470186 359494
rect 470422 359258 477186 359494
rect 477422 359258 484186 359494
rect 484422 359258 491186 359494
rect 491422 359258 498186 359494
rect 498422 359258 505186 359494
rect 505422 359258 512186 359494
rect 512422 359258 519186 359494
rect 519422 359258 526186 359494
rect 526422 359258 533186 359494
rect 533422 359258 540186 359494
rect 540422 359258 547186 359494
rect 547422 359258 554186 359494
rect 554422 359258 561186 359494
rect 561422 359258 568186 359494
rect 568422 359258 575186 359494
rect 575422 359258 582186 359494
rect 582422 359258 585818 359494
rect 586054 359258 586138 359494
rect 586374 359258 586458 359494
rect 586694 359258 586778 359494
rect 587014 359258 588874 359494
rect -4950 359216 588874 359258
rect -4950 353434 588874 353476
rect -4950 353198 -4842 353434
rect -4606 353198 -4522 353434
rect -4286 353198 -4202 353434
rect -3966 353198 -3882 353434
rect -3646 353198 2918 353434
rect 3154 353198 9918 353434
rect 10154 353198 16918 353434
rect 17154 353198 23918 353434
rect 24154 353198 30918 353434
rect 31154 353198 37918 353434
rect 38154 353198 44918 353434
rect 45154 353198 51918 353434
rect 52154 353198 58918 353434
rect 59154 353198 65918 353434
rect 66154 353198 72918 353434
rect 73154 353198 79918 353434
rect 80154 353198 86918 353434
rect 87154 353198 93918 353434
rect 94154 353198 100918 353434
rect 101154 353198 107918 353434
rect 108154 353198 114918 353434
rect 115154 353198 121918 353434
rect 122154 353198 128918 353434
rect 129154 353198 135918 353434
rect 136154 353198 142918 353434
rect 143154 353198 149918 353434
rect 150154 353198 156918 353434
rect 157154 353198 163918 353434
rect 164154 353198 170918 353434
rect 171154 353198 177918 353434
rect 178154 353198 184918 353434
rect 185154 353198 191918 353434
rect 192154 353198 198918 353434
rect 199154 353198 205918 353434
rect 206154 353198 212918 353434
rect 213154 353198 219918 353434
rect 220154 353198 226918 353434
rect 227154 353198 233918 353434
rect 234154 353198 240918 353434
rect 241154 353198 247918 353434
rect 248154 353198 254918 353434
rect 255154 353198 261918 353434
rect 262154 353198 268918 353434
rect 269154 353198 275918 353434
rect 276154 353198 282918 353434
rect 283154 353198 289918 353434
rect 290154 353198 296918 353434
rect 297154 353198 303918 353434
rect 304154 353198 310918 353434
rect 311154 353198 317918 353434
rect 318154 353198 324918 353434
rect 325154 353198 331918 353434
rect 332154 353198 338918 353434
rect 339154 353198 345918 353434
rect 346154 353198 352918 353434
rect 353154 353198 359918 353434
rect 360154 353198 366918 353434
rect 367154 353198 373918 353434
rect 374154 353198 380918 353434
rect 381154 353198 387918 353434
rect 388154 353198 394918 353434
rect 395154 353198 401918 353434
rect 402154 353198 408918 353434
rect 409154 353198 415918 353434
rect 416154 353198 422918 353434
rect 423154 353198 429918 353434
rect 430154 353198 436918 353434
rect 437154 353198 443918 353434
rect 444154 353198 450918 353434
rect 451154 353198 457918 353434
rect 458154 353198 464918 353434
rect 465154 353198 471918 353434
rect 472154 353198 478918 353434
rect 479154 353198 485918 353434
rect 486154 353198 492918 353434
rect 493154 353198 499918 353434
rect 500154 353198 506918 353434
rect 507154 353198 513918 353434
rect 514154 353198 520918 353434
rect 521154 353198 527918 353434
rect 528154 353198 534918 353434
rect 535154 353198 541918 353434
rect 542154 353198 548918 353434
rect 549154 353198 555918 353434
rect 556154 353198 562918 353434
rect 563154 353198 569918 353434
rect 570154 353198 576918 353434
rect 577154 353198 587570 353434
rect 587806 353198 587890 353434
rect 588126 353198 588210 353434
rect 588446 353198 588530 353434
rect 588766 353198 588874 353434
rect -4950 353156 588874 353198
rect -4950 352494 588874 352536
rect -4950 352258 -3090 352494
rect -2854 352258 -2770 352494
rect -2534 352258 -2450 352494
rect -2214 352258 -2130 352494
rect -1894 352258 1186 352494
rect 1422 352258 8186 352494
rect 8422 352258 15186 352494
rect 15422 352258 22186 352494
rect 22422 352258 29186 352494
rect 29422 352258 36186 352494
rect 36422 352258 43186 352494
rect 43422 352258 50186 352494
rect 50422 352258 57186 352494
rect 57422 352258 64186 352494
rect 64422 352258 71186 352494
rect 71422 352258 78186 352494
rect 78422 352258 85186 352494
rect 85422 352258 92186 352494
rect 92422 352258 99186 352494
rect 99422 352258 106186 352494
rect 106422 352258 113186 352494
rect 113422 352258 120186 352494
rect 120422 352258 127186 352494
rect 127422 352258 134186 352494
rect 134422 352258 141186 352494
rect 141422 352258 148186 352494
rect 148422 352258 155186 352494
rect 155422 352258 162186 352494
rect 162422 352258 169186 352494
rect 169422 352258 176186 352494
rect 176422 352258 183186 352494
rect 183422 352258 190186 352494
rect 190422 352258 197186 352494
rect 197422 352258 204186 352494
rect 204422 352258 211186 352494
rect 211422 352258 218186 352494
rect 218422 352258 225186 352494
rect 225422 352258 232186 352494
rect 232422 352258 239186 352494
rect 239422 352258 246186 352494
rect 246422 352258 253186 352494
rect 253422 352258 260186 352494
rect 260422 352258 267186 352494
rect 267422 352258 274186 352494
rect 274422 352258 281186 352494
rect 281422 352258 288186 352494
rect 288422 352258 295186 352494
rect 295422 352258 302186 352494
rect 302422 352258 309186 352494
rect 309422 352258 316186 352494
rect 316422 352258 323186 352494
rect 323422 352258 330186 352494
rect 330422 352258 337186 352494
rect 337422 352258 344186 352494
rect 344422 352258 351186 352494
rect 351422 352258 358186 352494
rect 358422 352258 365186 352494
rect 365422 352258 372186 352494
rect 372422 352258 379186 352494
rect 379422 352258 386186 352494
rect 386422 352258 393186 352494
rect 393422 352258 400186 352494
rect 400422 352258 407186 352494
rect 407422 352258 414186 352494
rect 414422 352258 421186 352494
rect 421422 352258 428186 352494
rect 428422 352258 435186 352494
rect 435422 352258 442186 352494
rect 442422 352258 449186 352494
rect 449422 352258 456186 352494
rect 456422 352258 463186 352494
rect 463422 352258 470186 352494
rect 470422 352258 477186 352494
rect 477422 352258 484186 352494
rect 484422 352258 491186 352494
rect 491422 352258 498186 352494
rect 498422 352258 505186 352494
rect 505422 352258 512186 352494
rect 512422 352258 519186 352494
rect 519422 352258 526186 352494
rect 526422 352258 533186 352494
rect 533422 352258 540186 352494
rect 540422 352258 547186 352494
rect 547422 352258 554186 352494
rect 554422 352258 561186 352494
rect 561422 352258 568186 352494
rect 568422 352258 575186 352494
rect 575422 352258 582186 352494
rect 582422 352258 585818 352494
rect 586054 352258 586138 352494
rect 586374 352258 586458 352494
rect 586694 352258 586778 352494
rect 587014 352258 588874 352494
rect -4950 352216 588874 352258
rect -4950 346434 588874 346476
rect -4950 346198 -4842 346434
rect -4606 346198 -4522 346434
rect -4286 346198 -4202 346434
rect -3966 346198 -3882 346434
rect -3646 346198 2918 346434
rect 3154 346198 9918 346434
rect 10154 346198 16918 346434
rect 17154 346198 23918 346434
rect 24154 346198 30918 346434
rect 31154 346198 37918 346434
rect 38154 346198 44918 346434
rect 45154 346198 51918 346434
rect 52154 346198 58918 346434
rect 59154 346198 65918 346434
rect 66154 346198 72918 346434
rect 73154 346198 79918 346434
rect 80154 346198 86918 346434
rect 87154 346198 93918 346434
rect 94154 346198 100918 346434
rect 101154 346198 107918 346434
rect 108154 346198 114918 346434
rect 115154 346198 121918 346434
rect 122154 346198 128918 346434
rect 129154 346198 135918 346434
rect 136154 346198 142918 346434
rect 143154 346198 149918 346434
rect 150154 346198 156918 346434
rect 157154 346198 163918 346434
rect 164154 346198 170918 346434
rect 171154 346198 177918 346434
rect 178154 346198 184918 346434
rect 185154 346198 191918 346434
rect 192154 346198 198918 346434
rect 199154 346198 205918 346434
rect 206154 346198 212918 346434
rect 213154 346198 219918 346434
rect 220154 346198 226918 346434
rect 227154 346198 233918 346434
rect 234154 346198 240918 346434
rect 241154 346198 247918 346434
rect 248154 346198 254918 346434
rect 255154 346198 261918 346434
rect 262154 346198 268918 346434
rect 269154 346198 275918 346434
rect 276154 346198 282918 346434
rect 283154 346198 289918 346434
rect 290154 346198 296918 346434
rect 297154 346198 303918 346434
rect 304154 346198 310918 346434
rect 311154 346198 317918 346434
rect 318154 346198 324918 346434
rect 325154 346198 331918 346434
rect 332154 346198 338918 346434
rect 339154 346198 345918 346434
rect 346154 346198 352918 346434
rect 353154 346198 359918 346434
rect 360154 346198 366918 346434
rect 367154 346198 373918 346434
rect 374154 346198 380918 346434
rect 381154 346198 387918 346434
rect 388154 346198 394918 346434
rect 395154 346198 401918 346434
rect 402154 346198 408918 346434
rect 409154 346198 415918 346434
rect 416154 346198 422918 346434
rect 423154 346198 429918 346434
rect 430154 346198 436918 346434
rect 437154 346198 443918 346434
rect 444154 346198 450918 346434
rect 451154 346198 457918 346434
rect 458154 346198 464918 346434
rect 465154 346198 471918 346434
rect 472154 346198 478918 346434
rect 479154 346198 485918 346434
rect 486154 346198 492918 346434
rect 493154 346198 499918 346434
rect 500154 346198 506918 346434
rect 507154 346198 513918 346434
rect 514154 346198 520918 346434
rect 521154 346198 527918 346434
rect 528154 346198 534918 346434
rect 535154 346198 541918 346434
rect 542154 346198 548918 346434
rect 549154 346198 555918 346434
rect 556154 346198 562918 346434
rect 563154 346198 569918 346434
rect 570154 346198 576918 346434
rect 577154 346198 587570 346434
rect 587806 346198 587890 346434
rect 588126 346198 588210 346434
rect 588446 346198 588530 346434
rect 588766 346198 588874 346434
rect -4950 346156 588874 346198
rect -4950 345494 588874 345536
rect -4950 345258 -3090 345494
rect -2854 345258 -2770 345494
rect -2534 345258 -2450 345494
rect -2214 345258 -2130 345494
rect -1894 345258 1186 345494
rect 1422 345258 8186 345494
rect 8422 345258 15186 345494
rect 15422 345258 22186 345494
rect 22422 345258 29186 345494
rect 29422 345258 36186 345494
rect 36422 345258 43186 345494
rect 43422 345258 50186 345494
rect 50422 345258 57186 345494
rect 57422 345258 64186 345494
rect 64422 345258 71186 345494
rect 71422 345258 78186 345494
rect 78422 345258 85186 345494
rect 85422 345258 92186 345494
rect 92422 345258 99186 345494
rect 99422 345258 106186 345494
rect 106422 345258 113186 345494
rect 113422 345258 120186 345494
rect 120422 345258 127186 345494
rect 127422 345258 134186 345494
rect 134422 345258 141186 345494
rect 141422 345258 148186 345494
rect 148422 345258 155186 345494
rect 155422 345258 162186 345494
rect 162422 345258 169186 345494
rect 169422 345258 176186 345494
rect 176422 345258 183186 345494
rect 183422 345258 190186 345494
rect 190422 345258 197186 345494
rect 197422 345258 204186 345494
rect 204422 345258 211186 345494
rect 211422 345258 218186 345494
rect 218422 345258 225186 345494
rect 225422 345258 232186 345494
rect 232422 345258 239186 345494
rect 239422 345258 246186 345494
rect 246422 345258 253186 345494
rect 253422 345258 260186 345494
rect 260422 345258 267186 345494
rect 267422 345258 274186 345494
rect 274422 345258 281186 345494
rect 281422 345258 288186 345494
rect 288422 345258 295186 345494
rect 295422 345258 302186 345494
rect 302422 345258 309186 345494
rect 309422 345258 316186 345494
rect 316422 345258 323186 345494
rect 323422 345258 330186 345494
rect 330422 345258 337186 345494
rect 337422 345258 344186 345494
rect 344422 345258 351186 345494
rect 351422 345258 358186 345494
rect 358422 345258 365186 345494
rect 365422 345258 372186 345494
rect 372422 345258 379186 345494
rect 379422 345258 386186 345494
rect 386422 345258 393186 345494
rect 393422 345258 400186 345494
rect 400422 345258 407186 345494
rect 407422 345258 414186 345494
rect 414422 345258 421186 345494
rect 421422 345258 428186 345494
rect 428422 345258 435186 345494
rect 435422 345258 442186 345494
rect 442422 345258 449186 345494
rect 449422 345258 456186 345494
rect 456422 345258 463186 345494
rect 463422 345258 470186 345494
rect 470422 345258 477186 345494
rect 477422 345258 484186 345494
rect 484422 345258 491186 345494
rect 491422 345258 498186 345494
rect 498422 345258 505186 345494
rect 505422 345258 512186 345494
rect 512422 345258 519186 345494
rect 519422 345258 526186 345494
rect 526422 345258 533186 345494
rect 533422 345258 540186 345494
rect 540422 345258 547186 345494
rect 547422 345258 554186 345494
rect 554422 345258 561186 345494
rect 561422 345258 568186 345494
rect 568422 345258 575186 345494
rect 575422 345258 582186 345494
rect 582422 345258 585818 345494
rect 586054 345258 586138 345494
rect 586374 345258 586458 345494
rect 586694 345258 586778 345494
rect 587014 345258 588874 345494
rect -4950 345216 588874 345258
rect -4950 339434 588874 339476
rect -4950 339198 -4842 339434
rect -4606 339198 -4522 339434
rect -4286 339198 -4202 339434
rect -3966 339198 -3882 339434
rect -3646 339198 2918 339434
rect 3154 339198 9918 339434
rect 10154 339198 16918 339434
rect 17154 339198 23918 339434
rect 24154 339198 30918 339434
rect 31154 339198 37918 339434
rect 38154 339198 44918 339434
rect 45154 339198 51918 339434
rect 52154 339198 58918 339434
rect 59154 339198 65918 339434
rect 66154 339198 72918 339434
rect 73154 339198 79918 339434
rect 80154 339198 86918 339434
rect 87154 339198 93918 339434
rect 94154 339198 100918 339434
rect 101154 339198 107918 339434
rect 108154 339198 114918 339434
rect 115154 339198 121918 339434
rect 122154 339198 128918 339434
rect 129154 339198 135918 339434
rect 136154 339198 142918 339434
rect 143154 339198 149918 339434
rect 150154 339198 156918 339434
rect 157154 339198 163918 339434
rect 164154 339198 170918 339434
rect 171154 339198 177918 339434
rect 178154 339198 184918 339434
rect 185154 339198 191918 339434
rect 192154 339198 198918 339434
rect 199154 339198 205918 339434
rect 206154 339198 212918 339434
rect 213154 339198 219918 339434
rect 220154 339198 226918 339434
rect 227154 339198 233918 339434
rect 234154 339198 240918 339434
rect 241154 339198 247918 339434
rect 248154 339198 254918 339434
rect 255154 339198 261918 339434
rect 262154 339198 268918 339434
rect 269154 339198 275918 339434
rect 276154 339198 282918 339434
rect 283154 339198 289918 339434
rect 290154 339198 296918 339434
rect 297154 339198 303918 339434
rect 304154 339198 310918 339434
rect 311154 339198 317918 339434
rect 318154 339198 324918 339434
rect 325154 339198 331918 339434
rect 332154 339198 338918 339434
rect 339154 339198 345918 339434
rect 346154 339198 352918 339434
rect 353154 339198 359918 339434
rect 360154 339198 366918 339434
rect 367154 339198 373918 339434
rect 374154 339198 380918 339434
rect 381154 339198 387918 339434
rect 388154 339198 394918 339434
rect 395154 339198 401918 339434
rect 402154 339198 408918 339434
rect 409154 339198 415918 339434
rect 416154 339198 422918 339434
rect 423154 339198 429918 339434
rect 430154 339198 436918 339434
rect 437154 339198 443918 339434
rect 444154 339198 450918 339434
rect 451154 339198 457918 339434
rect 458154 339198 464918 339434
rect 465154 339198 471918 339434
rect 472154 339198 478918 339434
rect 479154 339198 485918 339434
rect 486154 339198 492918 339434
rect 493154 339198 499918 339434
rect 500154 339198 506918 339434
rect 507154 339198 513918 339434
rect 514154 339198 520918 339434
rect 521154 339198 522850 339434
rect 523086 339198 524782 339434
rect 525018 339198 526714 339434
rect 526950 339198 527918 339434
rect 528154 339198 534918 339434
rect 535154 339198 541918 339434
rect 542154 339198 548918 339434
rect 549154 339198 555918 339434
rect 556154 339198 562918 339434
rect 563154 339198 569918 339434
rect 570154 339198 576918 339434
rect 577154 339198 587570 339434
rect 587806 339198 587890 339434
rect 588126 339198 588210 339434
rect 588446 339198 588530 339434
rect 588766 339198 588874 339434
rect -4950 339156 588874 339198
rect -4950 338494 588874 338536
rect -4950 338258 -3090 338494
rect -2854 338258 -2770 338494
rect -2534 338258 -2450 338494
rect -2214 338258 -2130 338494
rect -1894 338258 1186 338494
rect 1422 338258 8186 338494
rect 8422 338258 15186 338494
rect 15422 338258 22186 338494
rect 22422 338258 29186 338494
rect 29422 338258 36186 338494
rect 36422 338258 43186 338494
rect 43422 338258 50186 338494
rect 50422 338258 57186 338494
rect 57422 338258 64186 338494
rect 64422 338258 71186 338494
rect 71422 338258 78186 338494
rect 78422 338258 85186 338494
rect 85422 338258 92186 338494
rect 92422 338258 99186 338494
rect 99422 338258 106186 338494
rect 106422 338258 113186 338494
rect 113422 338258 120186 338494
rect 120422 338258 127186 338494
rect 127422 338258 134186 338494
rect 134422 338258 141186 338494
rect 141422 338258 148186 338494
rect 148422 338258 155186 338494
rect 155422 338258 162186 338494
rect 162422 338258 169186 338494
rect 169422 338258 176186 338494
rect 176422 338258 183186 338494
rect 183422 338258 190186 338494
rect 190422 338258 197186 338494
rect 197422 338258 204186 338494
rect 204422 338258 211186 338494
rect 211422 338258 218186 338494
rect 218422 338258 225186 338494
rect 225422 338258 232186 338494
rect 232422 338258 239186 338494
rect 239422 338258 246186 338494
rect 246422 338258 253186 338494
rect 253422 338258 260186 338494
rect 260422 338258 267186 338494
rect 267422 338258 274186 338494
rect 274422 338258 281186 338494
rect 281422 338258 288186 338494
rect 288422 338258 295186 338494
rect 295422 338258 302186 338494
rect 302422 338258 309186 338494
rect 309422 338258 316186 338494
rect 316422 338258 323186 338494
rect 323422 338258 330186 338494
rect 330422 338258 337186 338494
rect 337422 338258 344186 338494
rect 344422 338258 351186 338494
rect 351422 338258 358186 338494
rect 358422 338258 365186 338494
rect 365422 338258 372186 338494
rect 372422 338258 379186 338494
rect 379422 338258 386186 338494
rect 386422 338258 393186 338494
rect 393422 338258 400186 338494
rect 400422 338258 407186 338494
rect 407422 338258 414186 338494
rect 414422 338258 421186 338494
rect 421422 338258 428186 338494
rect 428422 338258 435186 338494
rect 435422 338258 442186 338494
rect 442422 338258 449186 338494
rect 449422 338258 456186 338494
rect 456422 338258 463186 338494
rect 463422 338258 470186 338494
rect 470422 338258 477186 338494
rect 477422 338258 484186 338494
rect 484422 338258 491186 338494
rect 491422 338258 498186 338494
rect 498422 338258 505186 338494
rect 505422 338258 512186 338494
rect 512422 338258 519186 338494
rect 519422 338258 519952 338494
rect 520188 338258 521884 338494
rect 522120 338258 523816 338494
rect 524052 338258 525748 338494
rect 525984 338258 533186 338494
rect 533422 338258 540186 338494
rect 540422 338258 547186 338494
rect 547422 338258 554186 338494
rect 554422 338258 561186 338494
rect 561422 338258 568186 338494
rect 568422 338258 575186 338494
rect 575422 338258 582186 338494
rect 582422 338258 585818 338494
rect 586054 338258 586138 338494
rect 586374 338258 586458 338494
rect 586694 338258 586778 338494
rect 587014 338258 588874 338494
rect -4950 338216 588874 338258
rect -4950 332434 588874 332476
rect -4950 332198 -4842 332434
rect -4606 332198 -4522 332434
rect -4286 332198 -4202 332434
rect -3966 332198 -3882 332434
rect -3646 332198 2918 332434
rect 3154 332198 9918 332434
rect 10154 332198 16918 332434
rect 17154 332198 23918 332434
rect 24154 332198 30918 332434
rect 31154 332198 37918 332434
rect 38154 332198 44918 332434
rect 45154 332198 51918 332434
rect 52154 332198 58918 332434
rect 59154 332198 65918 332434
rect 66154 332198 72918 332434
rect 73154 332198 79918 332434
rect 80154 332198 86918 332434
rect 87154 332198 93918 332434
rect 94154 332198 100918 332434
rect 101154 332198 107918 332434
rect 108154 332198 114918 332434
rect 115154 332198 121918 332434
rect 122154 332198 128918 332434
rect 129154 332198 135918 332434
rect 136154 332198 142918 332434
rect 143154 332198 149918 332434
rect 150154 332198 156918 332434
rect 157154 332198 163918 332434
rect 164154 332198 170918 332434
rect 171154 332198 177918 332434
rect 178154 332198 184918 332434
rect 185154 332198 191918 332434
rect 192154 332198 198918 332434
rect 199154 332198 205918 332434
rect 206154 332198 212918 332434
rect 213154 332198 219918 332434
rect 220154 332198 226918 332434
rect 227154 332198 233918 332434
rect 234154 332198 240918 332434
rect 241154 332198 247918 332434
rect 248154 332198 254918 332434
rect 255154 332198 261918 332434
rect 262154 332198 268918 332434
rect 269154 332198 275918 332434
rect 276154 332198 282918 332434
rect 283154 332198 289918 332434
rect 290154 332198 296918 332434
rect 297154 332198 303918 332434
rect 304154 332198 310918 332434
rect 311154 332198 317918 332434
rect 318154 332198 324918 332434
rect 325154 332198 331918 332434
rect 332154 332198 338918 332434
rect 339154 332198 345918 332434
rect 346154 332198 352918 332434
rect 353154 332198 359918 332434
rect 360154 332198 366918 332434
rect 367154 332198 373918 332434
rect 374154 332198 380918 332434
rect 381154 332198 387918 332434
rect 388154 332198 394918 332434
rect 395154 332198 401918 332434
rect 402154 332198 408918 332434
rect 409154 332198 415918 332434
rect 416154 332198 422918 332434
rect 423154 332198 429918 332434
rect 430154 332198 436918 332434
rect 437154 332198 443918 332434
rect 444154 332198 450918 332434
rect 451154 332198 457918 332434
rect 458154 332198 464918 332434
rect 465154 332198 471918 332434
rect 472154 332198 478918 332434
rect 479154 332198 485918 332434
rect 486154 332198 492918 332434
rect 493154 332198 499918 332434
rect 500154 332198 506918 332434
rect 507154 332198 513918 332434
rect 514154 332198 520918 332434
rect 521154 332198 522850 332434
rect 523086 332198 524782 332434
rect 525018 332198 526714 332434
rect 526950 332198 527918 332434
rect 528154 332198 534918 332434
rect 535154 332198 541918 332434
rect 542154 332198 548918 332434
rect 549154 332198 555918 332434
rect 556154 332198 562918 332434
rect 563154 332198 569918 332434
rect 570154 332198 576918 332434
rect 577154 332198 587570 332434
rect 587806 332198 587890 332434
rect 588126 332198 588210 332434
rect 588446 332198 588530 332434
rect 588766 332198 588874 332434
rect -4950 332156 588874 332198
rect -4950 331494 588874 331536
rect -4950 331258 -3090 331494
rect -2854 331258 -2770 331494
rect -2534 331258 -2450 331494
rect -2214 331258 -2130 331494
rect -1894 331258 1186 331494
rect 1422 331258 8186 331494
rect 8422 331258 15186 331494
rect 15422 331258 22186 331494
rect 22422 331258 29186 331494
rect 29422 331258 36186 331494
rect 36422 331258 43186 331494
rect 43422 331258 50186 331494
rect 50422 331258 57186 331494
rect 57422 331258 64186 331494
rect 64422 331258 71186 331494
rect 71422 331258 78186 331494
rect 78422 331258 85186 331494
rect 85422 331258 92186 331494
rect 92422 331258 99186 331494
rect 99422 331258 106186 331494
rect 106422 331258 113186 331494
rect 113422 331258 120186 331494
rect 120422 331258 127186 331494
rect 127422 331258 134186 331494
rect 134422 331258 141186 331494
rect 141422 331258 148186 331494
rect 148422 331258 155186 331494
rect 155422 331258 162186 331494
rect 162422 331258 169186 331494
rect 169422 331258 176186 331494
rect 176422 331258 183186 331494
rect 183422 331258 190186 331494
rect 190422 331258 197186 331494
rect 197422 331258 204186 331494
rect 204422 331258 211186 331494
rect 211422 331258 218186 331494
rect 218422 331258 225186 331494
rect 225422 331258 232186 331494
rect 232422 331258 239186 331494
rect 239422 331258 246186 331494
rect 246422 331258 253186 331494
rect 253422 331258 260186 331494
rect 260422 331258 267186 331494
rect 267422 331258 274186 331494
rect 274422 331258 281186 331494
rect 281422 331258 288186 331494
rect 288422 331258 295186 331494
rect 295422 331258 302186 331494
rect 302422 331258 309186 331494
rect 309422 331258 316186 331494
rect 316422 331258 323186 331494
rect 323422 331258 330186 331494
rect 330422 331258 337186 331494
rect 337422 331258 344186 331494
rect 344422 331258 351186 331494
rect 351422 331258 358186 331494
rect 358422 331258 365186 331494
rect 365422 331258 372186 331494
rect 372422 331258 379186 331494
rect 379422 331258 386186 331494
rect 386422 331258 393186 331494
rect 393422 331258 400186 331494
rect 400422 331258 407186 331494
rect 407422 331258 414186 331494
rect 414422 331258 421186 331494
rect 421422 331258 428186 331494
rect 428422 331258 435186 331494
rect 435422 331258 442186 331494
rect 442422 331258 449186 331494
rect 449422 331258 456186 331494
rect 456422 331258 463186 331494
rect 463422 331258 470186 331494
rect 470422 331258 477186 331494
rect 477422 331258 484186 331494
rect 484422 331258 491186 331494
rect 491422 331258 498186 331494
rect 498422 331258 505186 331494
rect 505422 331258 512186 331494
rect 512422 331258 519186 331494
rect 519422 331258 519952 331494
rect 520188 331258 521884 331494
rect 522120 331258 523816 331494
rect 524052 331258 525748 331494
rect 525984 331258 533186 331494
rect 533422 331258 540186 331494
rect 540422 331258 547186 331494
rect 547422 331258 554186 331494
rect 554422 331258 561186 331494
rect 561422 331258 568186 331494
rect 568422 331258 575186 331494
rect 575422 331258 582186 331494
rect 582422 331258 585818 331494
rect 586054 331258 586138 331494
rect 586374 331258 586458 331494
rect 586694 331258 586778 331494
rect 587014 331258 588874 331494
rect -4950 331216 588874 331258
rect -4950 325434 588874 325476
rect -4950 325198 -4842 325434
rect -4606 325198 -4522 325434
rect -4286 325198 -4202 325434
rect -3966 325198 -3882 325434
rect -3646 325198 2918 325434
rect 3154 325198 9918 325434
rect 10154 325198 16918 325434
rect 17154 325198 23918 325434
rect 24154 325198 30918 325434
rect 31154 325198 37918 325434
rect 38154 325198 44918 325434
rect 45154 325198 51918 325434
rect 52154 325198 58918 325434
rect 59154 325198 65918 325434
rect 66154 325198 72918 325434
rect 73154 325198 79918 325434
rect 80154 325198 86918 325434
rect 87154 325198 93918 325434
rect 94154 325198 100918 325434
rect 101154 325198 107918 325434
rect 108154 325198 114918 325434
rect 115154 325198 121918 325434
rect 122154 325198 128918 325434
rect 129154 325198 135918 325434
rect 136154 325198 142918 325434
rect 143154 325198 149918 325434
rect 150154 325198 156918 325434
rect 157154 325198 163918 325434
rect 164154 325198 170918 325434
rect 171154 325198 177918 325434
rect 178154 325198 184918 325434
rect 185154 325198 191918 325434
rect 192154 325198 198918 325434
rect 199154 325198 205918 325434
rect 206154 325198 212918 325434
rect 213154 325198 219918 325434
rect 220154 325198 226918 325434
rect 227154 325198 233918 325434
rect 234154 325198 240918 325434
rect 241154 325198 247918 325434
rect 248154 325198 254918 325434
rect 255154 325198 261918 325434
rect 262154 325198 268918 325434
rect 269154 325198 275918 325434
rect 276154 325198 282918 325434
rect 283154 325198 289918 325434
rect 290154 325198 296918 325434
rect 297154 325198 303918 325434
rect 304154 325198 310918 325434
rect 311154 325198 317918 325434
rect 318154 325198 324918 325434
rect 325154 325198 331918 325434
rect 332154 325198 338918 325434
rect 339154 325198 345918 325434
rect 346154 325198 352918 325434
rect 353154 325198 359918 325434
rect 360154 325198 366918 325434
rect 367154 325198 373918 325434
rect 374154 325198 380918 325434
rect 381154 325198 387918 325434
rect 388154 325198 394918 325434
rect 395154 325198 401918 325434
rect 402154 325198 408918 325434
rect 409154 325198 415918 325434
rect 416154 325198 422918 325434
rect 423154 325198 429918 325434
rect 430154 325198 436918 325434
rect 437154 325198 443918 325434
rect 444154 325198 450918 325434
rect 451154 325198 457918 325434
rect 458154 325198 464918 325434
rect 465154 325198 471918 325434
rect 472154 325198 478918 325434
rect 479154 325198 485918 325434
rect 486154 325198 492918 325434
rect 493154 325198 499918 325434
rect 500154 325198 506918 325434
rect 507154 325198 513918 325434
rect 514154 325198 520918 325434
rect 521154 325198 522850 325434
rect 523086 325198 524782 325434
rect 525018 325198 526714 325434
rect 526950 325198 527918 325434
rect 528154 325198 534918 325434
rect 535154 325198 541918 325434
rect 542154 325198 548918 325434
rect 549154 325198 555918 325434
rect 556154 325198 562918 325434
rect 563154 325198 569918 325434
rect 570154 325198 576918 325434
rect 577154 325198 587570 325434
rect 587806 325198 587890 325434
rect 588126 325198 588210 325434
rect 588446 325198 588530 325434
rect 588766 325198 588874 325434
rect -4950 325156 588874 325198
rect -4950 324494 588874 324536
rect -4950 324258 -3090 324494
rect -2854 324258 -2770 324494
rect -2534 324258 -2450 324494
rect -2214 324258 -2130 324494
rect -1894 324258 1186 324494
rect 1422 324258 8186 324494
rect 8422 324258 15186 324494
rect 15422 324258 22186 324494
rect 22422 324258 29186 324494
rect 29422 324258 36186 324494
rect 36422 324258 43186 324494
rect 43422 324258 50186 324494
rect 50422 324258 57186 324494
rect 57422 324258 64186 324494
rect 64422 324258 71186 324494
rect 71422 324258 78186 324494
rect 78422 324258 85186 324494
rect 85422 324258 92186 324494
rect 92422 324258 99186 324494
rect 99422 324258 106186 324494
rect 106422 324258 113186 324494
rect 113422 324258 120186 324494
rect 120422 324258 127186 324494
rect 127422 324258 134186 324494
rect 134422 324258 141186 324494
rect 141422 324258 148186 324494
rect 148422 324258 155186 324494
rect 155422 324258 162186 324494
rect 162422 324258 169186 324494
rect 169422 324258 176186 324494
rect 176422 324258 183186 324494
rect 183422 324258 190186 324494
rect 190422 324258 197186 324494
rect 197422 324258 204186 324494
rect 204422 324258 211186 324494
rect 211422 324258 218186 324494
rect 218422 324258 225186 324494
rect 225422 324258 232186 324494
rect 232422 324258 239186 324494
rect 239422 324258 246186 324494
rect 246422 324258 253186 324494
rect 253422 324258 260186 324494
rect 260422 324258 267186 324494
rect 267422 324258 274186 324494
rect 274422 324258 281186 324494
rect 281422 324258 288186 324494
rect 288422 324258 295186 324494
rect 295422 324258 302186 324494
rect 302422 324258 309186 324494
rect 309422 324258 316186 324494
rect 316422 324258 323186 324494
rect 323422 324258 330186 324494
rect 330422 324258 337186 324494
rect 337422 324258 344186 324494
rect 344422 324258 351186 324494
rect 351422 324258 358186 324494
rect 358422 324258 365186 324494
rect 365422 324258 372186 324494
rect 372422 324258 379186 324494
rect 379422 324258 386186 324494
rect 386422 324258 393186 324494
rect 393422 324258 400186 324494
rect 400422 324258 407186 324494
rect 407422 324258 414186 324494
rect 414422 324258 421186 324494
rect 421422 324258 428186 324494
rect 428422 324258 435186 324494
rect 435422 324258 442186 324494
rect 442422 324258 449186 324494
rect 449422 324258 456186 324494
rect 456422 324258 463186 324494
rect 463422 324258 470186 324494
rect 470422 324258 477186 324494
rect 477422 324258 484186 324494
rect 484422 324258 491186 324494
rect 491422 324258 498186 324494
rect 498422 324258 505186 324494
rect 505422 324258 512186 324494
rect 512422 324258 519186 324494
rect 519422 324258 519952 324494
rect 520188 324258 521884 324494
rect 522120 324258 523816 324494
rect 524052 324258 525748 324494
rect 525984 324258 533186 324494
rect 533422 324258 540186 324494
rect 540422 324258 547186 324494
rect 547422 324258 554186 324494
rect 554422 324258 561186 324494
rect 561422 324258 568186 324494
rect 568422 324258 575186 324494
rect 575422 324258 582186 324494
rect 582422 324258 585818 324494
rect 586054 324258 586138 324494
rect 586374 324258 586458 324494
rect 586694 324258 586778 324494
rect 587014 324258 588874 324494
rect -4950 324216 588874 324258
rect -4950 318434 588874 318476
rect -4950 318198 -4842 318434
rect -4606 318198 -4522 318434
rect -4286 318198 -4202 318434
rect -3966 318198 -3882 318434
rect -3646 318198 2918 318434
rect 3154 318198 9918 318434
rect 10154 318198 16918 318434
rect 17154 318198 23918 318434
rect 24154 318198 30918 318434
rect 31154 318198 37918 318434
rect 38154 318198 44918 318434
rect 45154 318198 51918 318434
rect 52154 318198 58918 318434
rect 59154 318198 65918 318434
rect 66154 318198 72918 318434
rect 73154 318198 79918 318434
rect 80154 318198 86918 318434
rect 87154 318198 93918 318434
rect 94154 318198 100918 318434
rect 101154 318198 107918 318434
rect 108154 318198 114918 318434
rect 115154 318198 121918 318434
rect 122154 318198 128918 318434
rect 129154 318198 135918 318434
rect 136154 318198 142918 318434
rect 143154 318198 149918 318434
rect 150154 318198 156918 318434
rect 157154 318198 163918 318434
rect 164154 318198 170918 318434
rect 171154 318198 177918 318434
rect 178154 318198 184918 318434
rect 185154 318198 191918 318434
rect 192154 318198 198918 318434
rect 199154 318198 205918 318434
rect 206154 318198 212918 318434
rect 213154 318198 219918 318434
rect 220154 318198 226918 318434
rect 227154 318198 233918 318434
rect 234154 318198 240918 318434
rect 241154 318198 247918 318434
rect 248154 318198 254918 318434
rect 255154 318198 261918 318434
rect 262154 318198 268918 318434
rect 269154 318198 275918 318434
rect 276154 318198 282918 318434
rect 283154 318198 289918 318434
rect 290154 318198 296918 318434
rect 297154 318198 303918 318434
rect 304154 318198 310918 318434
rect 311154 318198 317918 318434
rect 318154 318198 324918 318434
rect 325154 318198 331918 318434
rect 332154 318198 338918 318434
rect 339154 318198 345918 318434
rect 346154 318198 352918 318434
rect 353154 318198 359918 318434
rect 360154 318198 366918 318434
rect 367154 318198 373918 318434
rect 374154 318198 380918 318434
rect 381154 318198 387918 318434
rect 388154 318198 394918 318434
rect 395154 318198 401918 318434
rect 402154 318198 408918 318434
rect 409154 318198 415918 318434
rect 416154 318198 422918 318434
rect 423154 318198 429918 318434
rect 430154 318198 436918 318434
rect 437154 318198 443918 318434
rect 444154 318198 450918 318434
rect 451154 318198 457918 318434
rect 458154 318198 464918 318434
rect 465154 318198 471918 318434
rect 472154 318198 478918 318434
rect 479154 318198 485918 318434
rect 486154 318198 492918 318434
rect 493154 318198 499918 318434
rect 500154 318198 506918 318434
rect 507154 318198 513918 318434
rect 514154 318198 520918 318434
rect 521154 318198 527918 318434
rect 528154 318198 534918 318434
rect 535154 318198 541918 318434
rect 542154 318198 548918 318434
rect 549154 318198 555918 318434
rect 556154 318198 562918 318434
rect 563154 318198 569918 318434
rect 570154 318198 576918 318434
rect 577154 318198 587570 318434
rect 587806 318198 587890 318434
rect 588126 318198 588210 318434
rect 588446 318198 588530 318434
rect 588766 318198 588874 318434
rect -4950 318156 588874 318198
rect -4950 317494 588874 317536
rect -4950 317258 -3090 317494
rect -2854 317258 -2770 317494
rect -2534 317258 -2450 317494
rect -2214 317258 -2130 317494
rect -1894 317258 1186 317494
rect 1422 317258 8186 317494
rect 8422 317258 15186 317494
rect 15422 317258 22186 317494
rect 22422 317258 29186 317494
rect 29422 317258 36186 317494
rect 36422 317258 43186 317494
rect 43422 317258 50186 317494
rect 50422 317258 57186 317494
rect 57422 317258 64186 317494
rect 64422 317258 71186 317494
rect 71422 317258 78186 317494
rect 78422 317258 85186 317494
rect 85422 317258 92186 317494
rect 92422 317258 99186 317494
rect 99422 317258 106186 317494
rect 106422 317258 113186 317494
rect 113422 317258 120186 317494
rect 120422 317258 127186 317494
rect 127422 317258 134186 317494
rect 134422 317258 141186 317494
rect 141422 317258 148186 317494
rect 148422 317258 155186 317494
rect 155422 317258 162186 317494
rect 162422 317258 169186 317494
rect 169422 317258 176186 317494
rect 176422 317258 183186 317494
rect 183422 317258 190186 317494
rect 190422 317258 197186 317494
rect 197422 317258 204186 317494
rect 204422 317258 211186 317494
rect 211422 317258 218186 317494
rect 218422 317258 225186 317494
rect 225422 317258 232186 317494
rect 232422 317258 239186 317494
rect 239422 317258 246186 317494
rect 246422 317258 253186 317494
rect 253422 317258 260186 317494
rect 260422 317258 267186 317494
rect 267422 317258 274186 317494
rect 274422 317258 281186 317494
rect 281422 317258 288186 317494
rect 288422 317258 295186 317494
rect 295422 317258 302186 317494
rect 302422 317258 309186 317494
rect 309422 317258 316186 317494
rect 316422 317258 323186 317494
rect 323422 317258 330186 317494
rect 330422 317258 337186 317494
rect 337422 317258 344186 317494
rect 344422 317258 351186 317494
rect 351422 317258 358186 317494
rect 358422 317258 365186 317494
rect 365422 317258 372186 317494
rect 372422 317258 379186 317494
rect 379422 317258 386186 317494
rect 386422 317258 393186 317494
rect 393422 317258 400186 317494
rect 400422 317258 407186 317494
rect 407422 317258 414186 317494
rect 414422 317258 421186 317494
rect 421422 317258 428186 317494
rect 428422 317258 435186 317494
rect 435422 317258 442186 317494
rect 442422 317258 449186 317494
rect 449422 317258 456186 317494
rect 456422 317258 463186 317494
rect 463422 317258 470186 317494
rect 470422 317258 477186 317494
rect 477422 317258 484186 317494
rect 484422 317258 491186 317494
rect 491422 317258 498186 317494
rect 498422 317258 505186 317494
rect 505422 317258 512186 317494
rect 512422 317258 519186 317494
rect 519422 317258 526186 317494
rect 526422 317258 533186 317494
rect 533422 317258 540186 317494
rect 540422 317258 547186 317494
rect 547422 317258 554186 317494
rect 554422 317258 561186 317494
rect 561422 317258 568186 317494
rect 568422 317258 575186 317494
rect 575422 317258 582186 317494
rect 582422 317258 585818 317494
rect 586054 317258 586138 317494
rect 586374 317258 586458 317494
rect 586694 317258 586778 317494
rect 587014 317258 588874 317494
rect -4950 317216 588874 317258
rect -4950 311434 588874 311476
rect -4950 311198 -4842 311434
rect -4606 311198 -4522 311434
rect -4286 311198 -4202 311434
rect -3966 311198 -3882 311434
rect -3646 311198 2918 311434
rect 3154 311198 9918 311434
rect 10154 311198 16918 311434
rect 17154 311198 23918 311434
rect 24154 311198 30918 311434
rect 31154 311198 37918 311434
rect 38154 311198 44918 311434
rect 45154 311198 51918 311434
rect 52154 311198 58918 311434
rect 59154 311198 65918 311434
rect 66154 311198 72918 311434
rect 73154 311198 79918 311434
rect 80154 311198 86918 311434
rect 87154 311198 93918 311434
rect 94154 311198 100918 311434
rect 101154 311198 107918 311434
rect 108154 311198 114918 311434
rect 115154 311198 121918 311434
rect 122154 311198 128918 311434
rect 129154 311198 135918 311434
rect 136154 311198 142918 311434
rect 143154 311198 149918 311434
rect 150154 311198 156918 311434
rect 157154 311198 163918 311434
rect 164154 311198 170918 311434
rect 171154 311198 177918 311434
rect 178154 311198 184918 311434
rect 185154 311198 191918 311434
rect 192154 311198 198918 311434
rect 199154 311198 205918 311434
rect 206154 311198 212918 311434
rect 213154 311198 219918 311434
rect 220154 311198 226918 311434
rect 227154 311198 233918 311434
rect 234154 311198 240918 311434
rect 241154 311198 247918 311434
rect 248154 311198 254918 311434
rect 255154 311198 261918 311434
rect 262154 311198 268918 311434
rect 269154 311198 275918 311434
rect 276154 311198 282918 311434
rect 283154 311198 289918 311434
rect 290154 311198 296918 311434
rect 297154 311198 303918 311434
rect 304154 311198 310918 311434
rect 311154 311198 317918 311434
rect 318154 311198 324918 311434
rect 325154 311198 331918 311434
rect 332154 311198 338918 311434
rect 339154 311198 345918 311434
rect 346154 311198 352918 311434
rect 353154 311198 359918 311434
rect 360154 311198 366918 311434
rect 367154 311198 373918 311434
rect 374154 311198 380918 311434
rect 381154 311198 387918 311434
rect 388154 311198 394918 311434
rect 395154 311198 401918 311434
rect 402154 311198 408918 311434
rect 409154 311198 415918 311434
rect 416154 311198 422918 311434
rect 423154 311198 429918 311434
rect 430154 311198 436918 311434
rect 437154 311198 443918 311434
rect 444154 311198 450918 311434
rect 451154 311198 457918 311434
rect 458154 311198 464918 311434
rect 465154 311198 471918 311434
rect 472154 311198 478918 311434
rect 479154 311198 485918 311434
rect 486154 311198 492918 311434
rect 493154 311198 499918 311434
rect 500154 311198 506918 311434
rect 507154 311198 513918 311434
rect 514154 311198 520918 311434
rect 521154 311198 527918 311434
rect 528154 311198 534918 311434
rect 535154 311198 541918 311434
rect 542154 311198 548918 311434
rect 549154 311198 555918 311434
rect 556154 311198 562918 311434
rect 563154 311198 569918 311434
rect 570154 311198 576918 311434
rect 577154 311198 587570 311434
rect 587806 311198 587890 311434
rect 588126 311198 588210 311434
rect 588446 311198 588530 311434
rect 588766 311198 588874 311434
rect -4950 311156 588874 311198
rect -4950 310494 588874 310536
rect -4950 310258 -3090 310494
rect -2854 310258 -2770 310494
rect -2534 310258 -2450 310494
rect -2214 310258 -2130 310494
rect -1894 310258 1186 310494
rect 1422 310258 8186 310494
rect 8422 310258 15186 310494
rect 15422 310258 22186 310494
rect 22422 310258 29186 310494
rect 29422 310258 36186 310494
rect 36422 310258 43186 310494
rect 43422 310258 50186 310494
rect 50422 310258 57186 310494
rect 57422 310258 64186 310494
rect 64422 310258 71186 310494
rect 71422 310258 78186 310494
rect 78422 310258 85186 310494
rect 85422 310258 92186 310494
rect 92422 310258 99186 310494
rect 99422 310258 106186 310494
rect 106422 310258 113186 310494
rect 113422 310258 120186 310494
rect 120422 310258 127186 310494
rect 127422 310258 134186 310494
rect 134422 310258 141186 310494
rect 141422 310258 148186 310494
rect 148422 310258 155186 310494
rect 155422 310258 162186 310494
rect 162422 310258 169186 310494
rect 169422 310258 176186 310494
rect 176422 310258 183186 310494
rect 183422 310258 190186 310494
rect 190422 310258 197186 310494
rect 197422 310258 204186 310494
rect 204422 310258 211186 310494
rect 211422 310258 218186 310494
rect 218422 310258 225186 310494
rect 225422 310258 232186 310494
rect 232422 310258 239186 310494
rect 239422 310258 246186 310494
rect 246422 310258 253186 310494
rect 253422 310258 260186 310494
rect 260422 310258 267186 310494
rect 267422 310258 274186 310494
rect 274422 310258 281186 310494
rect 281422 310258 288186 310494
rect 288422 310258 295186 310494
rect 295422 310258 302186 310494
rect 302422 310258 309186 310494
rect 309422 310258 316186 310494
rect 316422 310258 323186 310494
rect 323422 310258 330186 310494
rect 330422 310258 337186 310494
rect 337422 310258 344186 310494
rect 344422 310258 351186 310494
rect 351422 310258 358186 310494
rect 358422 310258 365186 310494
rect 365422 310258 372186 310494
rect 372422 310258 379186 310494
rect 379422 310258 386186 310494
rect 386422 310258 393186 310494
rect 393422 310258 400186 310494
rect 400422 310258 407186 310494
rect 407422 310258 414186 310494
rect 414422 310258 421186 310494
rect 421422 310258 428186 310494
rect 428422 310258 435186 310494
rect 435422 310258 442186 310494
rect 442422 310258 449186 310494
rect 449422 310258 456186 310494
rect 456422 310258 463186 310494
rect 463422 310258 470186 310494
rect 470422 310258 477186 310494
rect 477422 310258 484186 310494
rect 484422 310258 491186 310494
rect 491422 310258 498186 310494
rect 498422 310258 505186 310494
rect 505422 310258 512186 310494
rect 512422 310258 519186 310494
rect 519422 310258 526186 310494
rect 526422 310258 533186 310494
rect 533422 310258 540186 310494
rect 540422 310258 547186 310494
rect 547422 310258 554186 310494
rect 554422 310258 561186 310494
rect 561422 310258 568186 310494
rect 568422 310258 575186 310494
rect 575422 310258 582186 310494
rect 582422 310258 585818 310494
rect 586054 310258 586138 310494
rect 586374 310258 586458 310494
rect 586694 310258 586778 310494
rect 587014 310258 588874 310494
rect -4950 310216 588874 310258
rect -4950 304434 588874 304476
rect -4950 304198 -4842 304434
rect -4606 304198 -4522 304434
rect -4286 304198 -4202 304434
rect -3966 304198 -3882 304434
rect -3646 304198 2918 304434
rect 3154 304198 9918 304434
rect 10154 304198 16918 304434
rect 17154 304198 23918 304434
rect 24154 304198 30918 304434
rect 31154 304198 37918 304434
rect 38154 304198 44918 304434
rect 45154 304198 51918 304434
rect 52154 304198 58918 304434
rect 59154 304198 65918 304434
rect 66154 304198 72918 304434
rect 73154 304198 79918 304434
rect 80154 304198 86918 304434
rect 87154 304198 93918 304434
rect 94154 304198 100918 304434
rect 101154 304198 107918 304434
rect 108154 304198 114918 304434
rect 115154 304198 121918 304434
rect 122154 304198 128918 304434
rect 129154 304198 135918 304434
rect 136154 304198 142918 304434
rect 143154 304198 149918 304434
rect 150154 304198 156918 304434
rect 157154 304198 163918 304434
rect 164154 304198 170918 304434
rect 171154 304198 177918 304434
rect 178154 304198 184918 304434
rect 185154 304198 191918 304434
rect 192154 304198 198918 304434
rect 199154 304198 205918 304434
rect 206154 304198 212918 304434
rect 213154 304198 219918 304434
rect 220154 304198 226918 304434
rect 227154 304198 233918 304434
rect 234154 304198 240918 304434
rect 241154 304198 247918 304434
rect 248154 304198 254918 304434
rect 255154 304198 261918 304434
rect 262154 304198 268918 304434
rect 269154 304198 275918 304434
rect 276154 304198 282918 304434
rect 283154 304198 289918 304434
rect 290154 304198 296918 304434
rect 297154 304198 303918 304434
rect 304154 304198 310918 304434
rect 311154 304198 317918 304434
rect 318154 304198 324918 304434
rect 325154 304198 331918 304434
rect 332154 304198 338918 304434
rect 339154 304198 345918 304434
rect 346154 304198 352918 304434
rect 353154 304198 359918 304434
rect 360154 304198 366918 304434
rect 367154 304198 373918 304434
rect 374154 304198 380918 304434
rect 381154 304198 387918 304434
rect 388154 304198 394918 304434
rect 395154 304198 401918 304434
rect 402154 304198 408918 304434
rect 409154 304198 415918 304434
rect 416154 304198 422918 304434
rect 423154 304198 429918 304434
rect 430154 304198 436918 304434
rect 437154 304198 443918 304434
rect 444154 304198 450918 304434
rect 451154 304198 457918 304434
rect 458154 304198 464918 304434
rect 465154 304198 471918 304434
rect 472154 304198 478918 304434
rect 479154 304198 485918 304434
rect 486154 304198 492918 304434
rect 493154 304198 499918 304434
rect 500154 304198 506918 304434
rect 507154 304198 513918 304434
rect 514154 304198 520918 304434
rect 521154 304198 527918 304434
rect 528154 304198 534918 304434
rect 535154 304198 541918 304434
rect 542154 304198 548918 304434
rect 549154 304198 555918 304434
rect 556154 304198 562918 304434
rect 563154 304198 569918 304434
rect 570154 304198 576918 304434
rect 577154 304198 587570 304434
rect 587806 304198 587890 304434
rect 588126 304198 588210 304434
rect 588446 304198 588530 304434
rect 588766 304198 588874 304434
rect -4950 304156 588874 304198
rect -4950 303494 588874 303536
rect -4950 303258 -3090 303494
rect -2854 303258 -2770 303494
rect -2534 303258 -2450 303494
rect -2214 303258 -2130 303494
rect -1894 303258 1186 303494
rect 1422 303258 8186 303494
rect 8422 303258 15186 303494
rect 15422 303258 22186 303494
rect 22422 303258 29186 303494
rect 29422 303258 36186 303494
rect 36422 303258 43186 303494
rect 43422 303258 50186 303494
rect 50422 303258 57186 303494
rect 57422 303258 64186 303494
rect 64422 303258 71186 303494
rect 71422 303258 78186 303494
rect 78422 303258 85186 303494
rect 85422 303258 92186 303494
rect 92422 303258 99186 303494
rect 99422 303258 106186 303494
rect 106422 303258 113186 303494
rect 113422 303258 120186 303494
rect 120422 303258 127186 303494
rect 127422 303258 134186 303494
rect 134422 303258 141186 303494
rect 141422 303258 148186 303494
rect 148422 303258 155186 303494
rect 155422 303258 162186 303494
rect 162422 303258 169186 303494
rect 169422 303258 176186 303494
rect 176422 303258 183186 303494
rect 183422 303258 190186 303494
rect 190422 303258 197186 303494
rect 197422 303258 204186 303494
rect 204422 303258 211186 303494
rect 211422 303258 218186 303494
rect 218422 303258 225186 303494
rect 225422 303258 232186 303494
rect 232422 303258 239186 303494
rect 239422 303258 246186 303494
rect 246422 303258 253186 303494
rect 253422 303258 260186 303494
rect 260422 303258 267186 303494
rect 267422 303258 274186 303494
rect 274422 303258 281186 303494
rect 281422 303258 288186 303494
rect 288422 303258 295186 303494
rect 295422 303258 302186 303494
rect 302422 303258 309186 303494
rect 309422 303258 316186 303494
rect 316422 303258 323186 303494
rect 323422 303258 330186 303494
rect 330422 303258 337186 303494
rect 337422 303258 344186 303494
rect 344422 303258 351186 303494
rect 351422 303258 358186 303494
rect 358422 303258 365186 303494
rect 365422 303258 372186 303494
rect 372422 303258 379186 303494
rect 379422 303258 386186 303494
rect 386422 303258 393186 303494
rect 393422 303258 400186 303494
rect 400422 303258 407186 303494
rect 407422 303258 414186 303494
rect 414422 303258 421186 303494
rect 421422 303258 428186 303494
rect 428422 303258 435186 303494
rect 435422 303258 442186 303494
rect 442422 303258 449186 303494
rect 449422 303258 456186 303494
rect 456422 303258 463186 303494
rect 463422 303258 470186 303494
rect 470422 303258 477186 303494
rect 477422 303258 484186 303494
rect 484422 303258 491186 303494
rect 491422 303258 498186 303494
rect 498422 303258 505186 303494
rect 505422 303258 512186 303494
rect 512422 303258 519186 303494
rect 519422 303258 526186 303494
rect 526422 303258 533186 303494
rect 533422 303258 540186 303494
rect 540422 303258 547186 303494
rect 547422 303258 554186 303494
rect 554422 303258 561186 303494
rect 561422 303258 568186 303494
rect 568422 303258 575186 303494
rect 575422 303258 582186 303494
rect 582422 303258 585818 303494
rect 586054 303258 586138 303494
rect 586374 303258 586458 303494
rect 586694 303258 586778 303494
rect 587014 303258 588874 303494
rect -4950 303216 588874 303258
rect -4950 297434 588874 297476
rect -4950 297198 -4842 297434
rect -4606 297198 -4522 297434
rect -4286 297198 -4202 297434
rect -3966 297198 -3882 297434
rect -3646 297198 2918 297434
rect 3154 297198 9918 297434
rect 10154 297198 16918 297434
rect 17154 297198 23918 297434
rect 24154 297198 30918 297434
rect 31154 297198 37918 297434
rect 38154 297198 44918 297434
rect 45154 297198 51918 297434
rect 52154 297198 58918 297434
rect 59154 297198 65918 297434
rect 66154 297198 72918 297434
rect 73154 297198 79918 297434
rect 80154 297198 86918 297434
rect 87154 297198 93918 297434
rect 94154 297198 100918 297434
rect 101154 297198 107918 297434
rect 108154 297198 114918 297434
rect 115154 297198 121918 297434
rect 122154 297198 128918 297434
rect 129154 297198 135918 297434
rect 136154 297198 142918 297434
rect 143154 297198 149918 297434
rect 150154 297198 156918 297434
rect 157154 297198 163918 297434
rect 164154 297198 170918 297434
rect 171154 297198 177918 297434
rect 178154 297198 184918 297434
rect 185154 297198 191918 297434
rect 192154 297198 198918 297434
rect 199154 297198 205918 297434
rect 206154 297198 212918 297434
rect 213154 297198 219918 297434
rect 220154 297198 226918 297434
rect 227154 297198 233918 297434
rect 234154 297198 240918 297434
rect 241154 297198 247918 297434
rect 248154 297198 254918 297434
rect 255154 297198 261918 297434
rect 262154 297198 268918 297434
rect 269154 297198 275918 297434
rect 276154 297198 282918 297434
rect 283154 297198 289918 297434
rect 290154 297198 296918 297434
rect 297154 297198 303918 297434
rect 304154 297198 310918 297434
rect 311154 297198 317918 297434
rect 318154 297198 324918 297434
rect 325154 297198 331918 297434
rect 332154 297198 338918 297434
rect 339154 297198 345918 297434
rect 346154 297198 352918 297434
rect 353154 297198 359918 297434
rect 360154 297198 366918 297434
rect 367154 297198 373918 297434
rect 374154 297198 380918 297434
rect 381154 297198 387918 297434
rect 388154 297198 394918 297434
rect 395154 297198 401918 297434
rect 402154 297198 408918 297434
rect 409154 297198 415918 297434
rect 416154 297198 422918 297434
rect 423154 297198 429918 297434
rect 430154 297198 436918 297434
rect 437154 297198 443918 297434
rect 444154 297198 450918 297434
rect 451154 297198 457918 297434
rect 458154 297198 464918 297434
rect 465154 297198 471918 297434
rect 472154 297198 478918 297434
rect 479154 297198 485918 297434
rect 486154 297198 492918 297434
rect 493154 297198 499918 297434
rect 500154 297198 506918 297434
rect 507154 297198 513918 297434
rect 514154 297198 520918 297434
rect 521154 297198 522850 297434
rect 523086 297198 524782 297434
rect 525018 297198 526714 297434
rect 526950 297198 527918 297434
rect 528154 297198 534918 297434
rect 535154 297198 541918 297434
rect 542154 297198 548918 297434
rect 549154 297198 555918 297434
rect 556154 297198 562918 297434
rect 563154 297198 569918 297434
rect 570154 297198 576918 297434
rect 577154 297198 587570 297434
rect 587806 297198 587890 297434
rect 588126 297198 588210 297434
rect 588446 297198 588530 297434
rect 588766 297198 588874 297434
rect -4950 297156 588874 297198
rect -4950 296494 588874 296536
rect -4950 296258 -3090 296494
rect -2854 296258 -2770 296494
rect -2534 296258 -2450 296494
rect -2214 296258 -2130 296494
rect -1894 296258 1186 296494
rect 1422 296258 8186 296494
rect 8422 296258 15186 296494
rect 15422 296258 22186 296494
rect 22422 296258 29186 296494
rect 29422 296258 36186 296494
rect 36422 296258 43186 296494
rect 43422 296258 50186 296494
rect 50422 296258 57186 296494
rect 57422 296258 64186 296494
rect 64422 296258 71186 296494
rect 71422 296258 78186 296494
rect 78422 296258 85186 296494
rect 85422 296258 92186 296494
rect 92422 296258 99186 296494
rect 99422 296258 106186 296494
rect 106422 296258 113186 296494
rect 113422 296258 120186 296494
rect 120422 296258 127186 296494
rect 127422 296258 134186 296494
rect 134422 296258 141186 296494
rect 141422 296258 148186 296494
rect 148422 296258 155186 296494
rect 155422 296258 162186 296494
rect 162422 296258 169186 296494
rect 169422 296258 176186 296494
rect 176422 296258 183186 296494
rect 183422 296258 190186 296494
rect 190422 296258 197186 296494
rect 197422 296258 204186 296494
rect 204422 296258 211186 296494
rect 211422 296258 218186 296494
rect 218422 296258 225186 296494
rect 225422 296258 232186 296494
rect 232422 296258 239186 296494
rect 239422 296258 246186 296494
rect 246422 296258 253186 296494
rect 253422 296258 260186 296494
rect 260422 296258 267186 296494
rect 267422 296258 274186 296494
rect 274422 296258 281186 296494
rect 281422 296258 288186 296494
rect 288422 296258 295186 296494
rect 295422 296258 302186 296494
rect 302422 296258 309186 296494
rect 309422 296258 316186 296494
rect 316422 296258 323186 296494
rect 323422 296258 330186 296494
rect 330422 296258 337186 296494
rect 337422 296258 344186 296494
rect 344422 296258 351186 296494
rect 351422 296258 358186 296494
rect 358422 296258 365186 296494
rect 365422 296258 372186 296494
rect 372422 296258 379186 296494
rect 379422 296258 386186 296494
rect 386422 296258 393186 296494
rect 393422 296258 400186 296494
rect 400422 296258 407186 296494
rect 407422 296258 414186 296494
rect 414422 296258 421186 296494
rect 421422 296258 428186 296494
rect 428422 296258 435186 296494
rect 435422 296258 442186 296494
rect 442422 296258 449186 296494
rect 449422 296258 456186 296494
rect 456422 296258 463186 296494
rect 463422 296258 470186 296494
rect 470422 296258 477186 296494
rect 477422 296258 484186 296494
rect 484422 296258 491186 296494
rect 491422 296258 498186 296494
rect 498422 296258 505186 296494
rect 505422 296258 512186 296494
rect 512422 296258 519186 296494
rect 519422 296258 519952 296494
rect 520188 296258 521884 296494
rect 522120 296258 523816 296494
rect 524052 296258 525748 296494
rect 525984 296258 533186 296494
rect 533422 296258 540186 296494
rect 540422 296258 547186 296494
rect 547422 296258 554186 296494
rect 554422 296258 561186 296494
rect 561422 296258 568186 296494
rect 568422 296258 575186 296494
rect 575422 296258 582186 296494
rect 582422 296258 585818 296494
rect 586054 296258 586138 296494
rect 586374 296258 586458 296494
rect 586694 296258 586778 296494
rect 587014 296258 588874 296494
rect -4950 296216 588874 296258
rect -4950 290434 588874 290476
rect -4950 290198 -4842 290434
rect -4606 290198 -4522 290434
rect -4286 290198 -4202 290434
rect -3966 290198 -3882 290434
rect -3646 290198 2918 290434
rect 3154 290198 9918 290434
rect 10154 290198 16918 290434
rect 17154 290198 23918 290434
rect 24154 290198 30918 290434
rect 31154 290198 37918 290434
rect 38154 290198 44918 290434
rect 45154 290198 51918 290434
rect 52154 290198 58918 290434
rect 59154 290198 65918 290434
rect 66154 290198 72918 290434
rect 73154 290198 79918 290434
rect 80154 290198 86918 290434
rect 87154 290198 93918 290434
rect 94154 290198 100918 290434
rect 101154 290198 107918 290434
rect 108154 290198 114918 290434
rect 115154 290198 121918 290434
rect 122154 290198 128918 290434
rect 129154 290198 135918 290434
rect 136154 290198 142918 290434
rect 143154 290198 149918 290434
rect 150154 290198 156918 290434
rect 157154 290198 163918 290434
rect 164154 290198 170918 290434
rect 171154 290198 177918 290434
rect 178154 290198 184918 290434
rect 185154 290198 191918 290434
rect 192154 290198 198918 290434
rect 199154 290198 205918 290434
rect 206154 290198 212918 290434
rect 213154 290198 219918 290434
rect 220154 290198 226918 290434
rect 227154 290198 233918 290434
rect 234154 290198 240918 290434
rect 241154 290198 247918 290434
rect 248154 290198 254918 290434
rect 255154 290198 261918 290434
rect 262154 290198 268918 290434
rect 269154 290198 275918 290434
rect 276154 290198 282918 290434
rect 283154 290198 289918 290434
rect 290154 290198 296918 290434
rect 297154 290198 303918 290434
rect 304154 290198 310918 290434
rect 311154 290198 317918 290434
rect 318154 290198 324918 290434
rect 325154 290198 331918 290434
rect 332154 290198 338918 290434
rect 339154 290198 345918 290434
rect 346154 290198 352918 290434
rect 353154 290198 359918 290434
rect 360154 290198 366918 290434
rect 367154 290198 373918 290434
rect 374154 290198 380918 290434
rect 381154 290198 387918 290434
rect 388154 290198 394918 290434
rect 395154 290198 401918 290434
rect 402154 290198 408918 290434
rect 409154 290198 415918 290434
rect 416154 290198 422918 290434
rect 423154 290198 429918 290434
rect 430154 290198 436918 290434
rect 437154 290198 443918 290434
rect 444154 290198 450918 290434
rect 451154 290198 457918 290434
rect 458154 290198 464918 290434
rect 465154 290198 471918 290434
rect 472154 290198 478918 290434
rect 479154 290198 485918 290434
rect 486154 290198 492918 290434
rect 493154 290198 499918 290434
rect 500154 290198 506918 290434
rect 507154 290198 513918 290434
rect 514154 290198 520918 290434
rect 521154 290198 522850 290434
rect 523086 290198 524782 290434
rect 525018 290198 526714 290434
rect 526950 290198 527918 290434
rect 528154 290198 534918 290434
rect 535154 290198 541918 290434
rect 542154 290198 548918 290434
rect 549154 290198 555918 290434
rect 556154 290198 562918 290434
rect 563154 290198 569918 290434
rect 570154 290198 576918 290434
rect 577154 290198 587570 290434
rect 587806 290198 587890 290434
rect 588126 290198 588210 290434
rect 588446 290198 588530 290434
rect 588766 290198 588874 290434
rect -4950 290156 588874 290198
rect -4950 289494 588874 289536
rect -4950 289258 -3090 289494
rect -2854 289258 -2770 289494
rect -2534 289258 -2450 289494
rect -2214 289258 -2130 289494
rect -1894 289258 1186 289494
rect 1422 289258 8186 289494
rect 8422 289258 15186 289494
rect 15422 289258 22186 289494
rect 22422 289258 29186 289494
rect 29422 289258 36186 289494
rect 36422 289258 43186 289494
rect 43422 289258 50186 289494
rect 50422 289258 57186 289494
rect 57422 289258 64186 289494
rect 64422 289258 71186 289494
rect 71422 289258 78186 289494
rect 78422 289258 85186 289494
rect 85422 289258 92186 289494
rect 92422 289258 99186 289494
rect 99422 289258 106186 289494
rect 106422 289258 113186 289494
rect 113422 289258 120186 289494
rect 120422 289258 127186 289494
rect 127422 289258 134186 289494
rect 134422 289258 141186 289494
rect 141422 289258 148186 289494
rect 148422 289258 155186 289494
rect 155422 289258 162186 289494
rect 162422 289258 169186 289494
rect 169422 289258 176186 289494
rect 176422 289258 183186 289494
rect 183422 289258 190186 289494
rect 190422 289258 197186 289494
rect 197422 289258 204186 289494
rect 204422 289258 211186 289494
rect 211422 289258 218186 289494
rect 218422 289258 225186 289494
rect 225422 289258 232186 289494
rect 232422 289258 239186 289494
rect 239422 289258 246186 289494
rect 246422 289258 253186 289494
rect 253422 289258 260186 289494
rect 260422 289258 267186 289494
rect 267422 289258 274186 289494
rect 274422 289258 281186 289494
rect 281422 289258 288186 289494
rect 288422 289258 295186 289494
rect 295422 289258 302186 289494
rect 302422 289258 309186 289494
rect 309422 289258 316186 289494
rect 316422 289258 323186 289494
rect 323422 289258 330186 289494
rect 330422 289258 337186 289494
rect 337422 289258 344186 289494
rect 344422 289258 351186 289494
rect 351422 289258 358186 289494
rect 358422 289258 365186 289494
rect 365422 289258 372186 289494
rect 372422 289258 379186 289494
rect 379422 289258 386186 289494
rect 386422 289258 393186 289494
rect 393422 289258 400186 289494
rect 400422 289258 407186 289494
rect 407422 289258 414186 289494
rect 414422 289258 421186 289494
rect 421422 289258 428186 289494
rect 428422 289258 435186 289494
rect 435422 289258 442186 289494
rect 442422 289258 449186 289494
rect 449422 289258 456186 289494
rect 456422 289258 463186 289494
rect 463422 289258 470186 289494
rect 470422 289258 477186 289494
rect 477422 289258 484186 289494
rect 484422 289258 491186 289494
rect 491422 289258 498186 289494
rect 498422 289258 505186 289494
rect 505422 289258 512186 289494
rect 512422 289258 519186 289494
rect 519422 289258 519952 289494
rect 520188 289258 521884 289494
rect 522120 289258 523816 289494
rect 524052 289258 525748 289494
rect 525984 289258 533186 289494
rect 533422 289258 540186 289494
rect 540422 289258 547186 289494
rect 547422 289258 554186 289494
rect 554422 289258 561186 289494
rect 561422 289258 568186 289494
rect 568422 289258 575186 289494
rect 575422 289258 582186 289494
rect 582422 289258 585818 289494
rect 586054 289258 586138 289494
rect 586374 289258 586458 289494
rect 586694 289258 586778 289494
rect 587014 289258 588874 289494
rect -4950 289216 588874 289258
rect -4950 283434 588874 283476
rect -4950 283198 -4842 283434
rect -4606 283198 -4522 283434
rect -4286 283198 -4202 283434
rect -3966 283198 -3882 283434
rect -3646 283198 2918 283434
rect 3154 283198 9918 283434
rect 10154 283198 16918 283434
rect 17154 283198 23918 283434
rect 24154 283198 30918 283434
rect 31154 283198 37918 283434
rect 38154 283198 44918 283434
rect 45154 283198 51918 283434
rect 52154 283198 58918 283434
rect 59154 283198 65918 283434
rect 66154 283198 72918 283434
rect 73154 283198 79918 283434
rect 80154 283198 86918 283434
rect 87154 283198 93918 283434
rect 94154 283198 100918 283434
rect 101154 283198 107918 283434
rect 108154 283198 114918 283434
rect 115154 283198 121918 283434
rect 122154 283198 128918 283434
rect 129154 283198 135918 283434
rect 136154 283198 142918 283434
rect 143154 283198 149918 283434
rect 150154 283198 156918 283434
rect 157154 283198 163918 283434
rect 164154 283198 170918 283434
rect 171154 283198 177918 283434
rect 178154 283198 184918 283434
rect 185154 283198 191918 283434
rect 192154 283198 198918 283434
rect 199154 283198 205918 283434
rect 206154 283198 212918 283434
rect 213154 283198 219918 283434
rect 220154 283198 226918 283434
rect 227154 283198 233918 283434
rect 234154 283198 240918 283434
rect 241154 283198 247918 283434
rect 248154 283198 254918 283434
rect 255154 283198 261918 283434
rect 262154 283198 268918 283434
rect 269154 283198 275918 283434
rect 276154 283198 282918 283434
rect 283154 283198 289918 283434
rect 290154 283198 296918 283434
rect 297154 283198 303918 283434
rect 304154 283198 310918 283434
rect 311154 283198 317918 283434
rect 318154 283198 324918 283434
rect 325154 283198 331918 283434
rect 332154 283198 338918 283434
rect 339154 283198 345918 283434
rect 346154 283198 352918 283434
rect 353154 283198 359918 283434
rect 360154 283198 366918 283434
rect 367154 283198 373918 283434
rect 374154 283198 380918 283434
rect 381154 283198 387918 283434
rect 388154 283198 394918 283434
rect 395154 283198 401918 283434
rect 402154 283198 408918 283434
rect 409154 283198 415918 283434
rect 416154 283198 422918 283434
rect 423154 283198 429918 283434
rect 430154 283198 436918 283434
rect 437154 283198 443918 283434
rect 444154 283198 450918 283434
rect 451154 283198 457918 283434
rect 458154 283198 464918 283434
rect 465154 283198 471918 283434
rect 472154 283198 478918 283434
rect 479154 283198 485918 283434
rect 486154 283198 492918 283434
rect 493154 283198 499918 283434
rect 500154 283198 506918 283434
rect 507154 283198 513918 283434
rect 514154 283198 520918 283434
rect 521154 283198 522850 283434
rect 523086 283198 524782 283434
rect 525018 283198 526714 283434
rect 526950 283198 527918 283434
rect 528154 283198 534918 283434
rect 535154 283198 541918 283434
rect 542154 283198 548918 283434
rect 549154 283198 555918 283434
rect 556154 283198 562918 283434
rect 563154 283198 569918 283434
rect 570154 283198 576918 283434
rect 577154 283198 587570 283434
rect 587806 283198 587890 283434
rect 588126 283198 588210 283434
rect 588446 283198 588530 283434
rect 588766 283198 588874 283434
rect -4950 283156 588874 283198
rect -4950 282494 588874 282536
rect -4950 282258 -3090 282494
rect -2854 282258 -2770 282494
rect -2534 282258 -2450 282494
rect -2214 282258 -2130 282494
rect -1894 282258 1186 282494
rect 1422 282258 8186 282494
rect 8422 282258 15186 282494
rect 15422 282258 22186 282494
rect 22422 282258 29186 282494
rect 29422 282258 36186 282494
rect 36422 282258 43186 282494
rect 43422 282258 50186 282494
rect 50422 282258 57186 282494
rect 57422 282258 64186 282494
rect 64422 282258 71186 282494
rect 71422 282258 78186 282494
rect 78422 282258 85186 282494
rect 85422 282258 92186 282494
rect 92422 282258 99186 282494
rect 99422 282258 106186 282494
rect 106422 282258 113186 282494
rect 113422 282258 120186 282494
rect 120422 282258 127186 282494
rect 127422 282258 134186 282494
rect 134422 282258 141186 282494
rect 141422 282258 148186 282494
rect 148422 282258 155186 282494
rect 155422 282258 162186 282494
rect 162422 282258 169186 282494
rect 169422 282258 176186 282494
rect 176422 282258 183186 282494
rect 183422 282258 190186 282494
rect 190422 282258 197186 282494
rect 197422 282258 204186 282494
rect 204422 282258 211186 282494
rect 211422 282258 218186 282494
rect 218422 282258 225186 282494
rect 225422 282258 232186 282494
rect 232422 282258 239186 282494
rect 239422 282258 246186 282494
rect 246422 282258 253186 282494
rect 253422 282258 260186 282494
rect 260422 282258 267186 282494
rect 267422 282258 274186 282494
rect 274422 282258 281186 282494
rect 281422 282258 288186 282494
rect 288422 282258 295186 282494
rect 295422 282258 302186 282494
rect 302422 282258 309186 282494
rect 309422 282258 316186 282494
rect 316422 282258 323186 282494
rect 323422 282258 330186 282494
rect 330422 282258 337186 282494
rect 337422 282258 344186 282494
rect 344422 282258 351186 282494
rect 351422 282258 358186 282494
rect 358422 282258 365186 282494
rect 365422 282258 372186 282494
rect 372422 282258 379186 282494
rect 379422 282258 386186 282494
rect 386422 282258 393186 282494
rect 393422 282258 400186 282494
rect 400422 282258 407186 282494
rect 407422 282258 414186 282494
rect 414422 282258 421186 282494
rect 421422 282258 428186 282494
rect 428422 282258 435186 282494
rect 435422 282258 442186 282494
rect 442422 282258 449186 282494
rect 449422 282258 456186 282494
rect 456422 282258 463186 282494
rect 463422 282258 470186 282494
rect 470422 282258 477186 282494
rect 477422 282258 484186 282494
rect 484422 282258 491186 282494
rect 491422 282258 498186 282494
rect 498422 282258 505186 282494
rect 505422 282258 512186 282494
rect 512422 282258 519186 282494
rect 519422 282258 519952 282494
rect 520188 282258 521884 282494
rect 522120 282258 523816 282494
rect 524052 282258 525748 282494
rect 525984 282258 533186 282494
rect 533422 282258 540186 282494
rect 540422 282258 547186 282494
rect 547422 282258 554186 282494
rect 554422 282258 561186 282494
rect 561422 282258 568186 282494
rect 568422 282258 575186 282494
rect 575422 282258 582186 282494
rect 582422 282258 585818 282494
rect 586054 282258 586138 282494
rect 586374 282258 586458 282494
rect 586694 282258 586778 282494
rect 587014 282258 588874 282494
rect -4950 282216 588874 282258
rect -4950 276434 588874 276476
rect -4950 276198 -4842 276434
rect -4606 276198 -4522 276434
rect -4286 276198 -4202 276434
rect -3966 276198 -3882 276434
rect -3646 276198 2918 276434
rect 3154 276198 9918 276434
rect 10154 276198 16918 276434
rect 17154 276198 23918 276434
rect 24154 276198 30918 276434
rect 31154 276198 37918 276434
rect 38154 276198 44918 276434
rect 45154 276198 51918 276434
rect 52154 276198 58918 276434
rect 59154 276198 65918 276434
rect 66154 276198 72918 276434
rect 73154 276198 79918 276434
rect 80154 276198 86918 276434
rect 87154 276198 93918 276434
rect 94154 276198 100918 276434
rect 101154 276198 107918 276434
rect 108154 276198 114918 276434
rect 115154 276198 121918 276434
rect 122154 276198 128918 276434
rect 129154 276198 135918 276434
rect 136154 276198 142918 276434
rect 143154 276198 149918 276434
rect 150154 276198 156918 276434
rect 157154 276198 163918 276434
rect 164154 276198 170918 276434
rect 171154 276198 177918 276434
rect 178154 276198 184918 276434
rect 185154 276198 191918 276434
rect 192154 276198 198918 276434
rect 199154 276198 205918 276434
rect 206154 276198 212918 276434
rect 213154 276198 219918 276434
rect 220154 276198 226918 276434
rect 227154 276198 233918 276434
rect 234154 276198 240918 276434
rect 241154 276198 247918 276434
rect 248154 276198 254918 276434
rect 255154 276198 261918 276434
rect 262154 276198 268918 276434
rect 269154 276198 275918 276434
rect 276154 276198 282918 276434
rect 283154 276198 289918 276434
rect 290154 276198 296918 276434
rect 297154 276198 303918 276434
rect 304154 276198 310918 276434
rect 311154 276198 317918 276434
rect 318154 276198 324918 276434
rect 325154 276198 331918 276434
rect 332154 276198 338918 276434
rect 339154 276198 345918 276434
rect 346154 276198 352918 276434
rect 353154 276198 359918 276434
rect 360154 276198 366918 276434
rect 367154 276198 373918 276434
rect 374154 276198 380918 276434
rect 381154 276198 387918 276434
rect 388154 276198 394918 276434
rect 395154 276198 401918 276434
rect 402154 276198 408918 276434
rect 409154 276198 415918 276434
rect 416154 276198 422918 276434
rect 423154 276198 429918 276434
rect 430154 276198 436918 276434
rect 437154 276198 443918 276434
rect 444154 276198 450918 276434
rect 451154 276198 457918 276434
rect 458154 276198 464918 276434
rect 465154 276198 471918 276434
rect 472154 276198 478918 276434
rect 479154 276198 485918 276434
rect 486154 276198 492918 276434
rect 493154 276198 499918 276434
rect 500154 276198 506918 276434
rect 507154 276198 513918 276434
rect 514154 276198 520918 276434
rect 521154 276198 527918 276434
rect 528154 276198 534918 276434
rect 535154 276198 541918 276434
rect 542154 276198 548918 276434
rect 549154 276198 555918 276434
rect 556154 276198 562918 276434
rect 563154 276198 569918 276434
rect 570154 276198 576918 276434
rect 577154 276198 587570 276434
rect 587806 276198 587890 276434
rect 588126 276198 588210 276434
rect 588446 276198 588530 276434
rect 588766 276198 588874 276434
rect -4950 276156 588874 276198
rect -4950 275494 588874 275536
rect -4950 275258 -3090 275494
rect -2854 275258 -2770 275494
rect -2534 275258 -2450 275494
rect -2214 275258 -2130 275494
rect -1894 275258 1186 275494
rect 1422 275258 8186 275494
rect 8422 275258 15186 275494
rect 15422 275258 22186 275494
rect 22422 275258 29186 275494
rect 29422 275258 36186 275494
rect 36422 275258 43186 275494
rect 43422 275258 50186 275494
rect 50422 275258 57186 275494
rect 57422 275258 64186 275494
rect 64422 275258 71186 275494
rect 71422 275258 78186 275494
rect 78422 275258 85186 275494
rect 85422 275258 92186 275494
rect 92422 275258 99186 275494
rect 99422 275258 106186 275494
rect 106422 275258 113186 275494
rect 113422 275258 120186 275494
rect 120422 275258 127186 275494
rect 127422 275258 134186 275494
rect 134422 275258 141186 275494
rect 141422 275258 148186 275494
rect 148422 275258 155186 275494
rect 155422 275258 162186 275494
rect 162422 275258 169186 275494
rect 169422 275258 176186 275494
rect 176422 275258 183186 275494
rect 183422 275258 190186 275494
rect 190422 275258 197186 275494
rect 197422 275258 204186 275494
rect 204422 275258 211186 275494
rect 211422 275258 218186 275494
rect 218422 275258 225186 275494
rect 225422 275258 232186 275494
rect 232422 275258 239186 275494
rect 239422 275258 246186 275494
rect 246422 275258 253186 275494
rect 253422 275258 260186 275494
rect 260422 275258 267186 275494
rect 267422 275258 274186 275494
rect 274422 275258 281186 275494
rect 281422 275258 288186 275494
rect 288422 275258 295186 275494
rect 295422 275258 302186 275494
rect 302422 275258 309186 275494
rect 309422 275258 316186 275494
rect 316422 275258 323186 275494
rect 323422 275258 330186 275494
rect 330422 275258 337186 275494
rect 337422 275258 344186 275494
rect 344422 275258 351186 275494
rect 351422 275258 358186 275494
rect 358422 275258 365186 275494
rect 365422 275258 372186 275494
rect 372422 275258 379186 275494
rect 379422 275258 386186 275494
rect 386422 275258 393186 275494
rect 393422 275258 400186 275494
rect 400422 275258 407186 275494
rect 407422 275258 414186 275494
rect 414422 275258 421186 275494
rect 421422 275258 428186 275494
rect 428422 275258 435186 275494
rect 435422 275258 442186 275494
rect 442422 275258 449186 275494
rect 449422 275258 456186 275494
rect 456422 275258 463186 275494
rect 463422 275258 470186 275494
rect 470422 275258 477186 275494
rect 477422 275258 484186 275494
rect 484422 275258 491186 275494
rect 491422 275258 498186 275494
rect 498422 275258 505186 275494
rect 505422 275258 512186 275494
rect 512422 275258 519186 275494
rect 519422 275258 526186 275494
rect 526422 275258 533186 275494
rect 533422 275258 540186 275494
rect 540422 275258 547186 275494
rect 547422 275258 554186 275494
rect 554422 275258 561186 275494
rect 561422 275258 568186 275494
rect 568422 275258 575186 275494
rect 575422 275258 582186 275494
rect 582422 275258 585818 275494
rect 586054 275258 586138 275494
rect 586374 275258 586458 275494
rect 586694 275258 586778 275494
rect 587014 275258 588874 275494
rect -4950 275216 588874 275258
rect -4950 269434 588874 269476
rect -4950 269198 -4842 269434
rect -4606 269198 -4522 269434
rect -4286 269198 -4202 269434
rect -3966 269198 -3882 269434
rect -3646 269198 2918 269434
rect 3154 269198 9918 269434
rect 10154 269198 16918 269434
rect 17154 269198 23918 269434
rect 24154 269198 30918 269434
rect 31154 269198 37918 269434
rect 38154 269198 44918 269434
rect 45154 269198 51918 269434
rect 52154 269198 58918 269434
rect 59154 269198 65918 269434
rect 66154 269198 72918 269434
rect 73154 269198 79918 269434
rect 80154 269198 86918 269434
rect 87154 269198 93918 269434
rect 94154 269198 100918 269434
rect 101154 269198 107918 269434
rect 108154 269198 114918 269434
rect 115154 269198 121918 269434
rect 122154 269198 128918 269434
rect 129154 269198 135918 269434
rect 136154 269198 142918 269434
rect 143154 269198 149918 269434
rect 150154 269198 156918 269434
rect 157154 269198 163918 269434
rect 164154 269198 170918 269434
rect 171154 269198 177918 269434
rect 178154 269198 184918 269434
rect 185154 269198 191918 269434
rect 192154 269198 198918 269434
rect 199154 269198 205918 269434
rect 206154 269198 212918 269434
rect 213154 269198 219918 269434
rect 220154 269198 226918 269434
rect 227154 269198 233918 269434
rect 234154 269198 240918 269434
rect 241154 269198 247918 269434
rect 248154 269198 254918 269434
rect 255154 269198 261918 269434
rect 262154 269198 268918 269434
rect 269154 269198 275918 269434
rect 276154 269198 282918 269434
rect 283154 269198 289918 269434
rect 290154 269198 296918 269434
rect 297154 269198 303918 269434
rect 304154 269198 310918 269434
rect 311154 269198 317918 269434
rect 318154 269198 324918 269434
rect 325154 269198 331918 269434
rect 332154 269198 338918 269434
rect 339154 269198 345918 269434
rect 346154 269198 352918 269434
rect 353154 269198 359918 269434
rect 360154 269198 366918 269434
rect 367154 269198 373918 269434
rect 374154 269198 380918 269434
rect 381154 269198 387918 269434
rect 388154 269198 394918 269434
rect 395154 269198 401918 269434
rect 402154 269198 408918 269434
rect 409154 269198 415918 269434
rect 416154 269198 422918 269434
rect 423154 269198 429918 269434
rect 430154 269198 436918 269434
rect 437154 269198 443918 269434
rect 444154 269198 450918 269434
rect 451154 269198 457918 269434
rect 458154 269198 464918 269434
rect 465154 269198 471918 269434
rect 472154 269198 478918 269434
rect 479154 269198 485918 269434
rect 486154 269198 492918 269434
rect 493154 269198 499918 269434
rect 500154 269198 506918 269434
rect 507154 269198 513918 269434
rect 514154 269198 520918 269434
rect 521154 269198 527918 269434
rect 528154 269198 534918 269434
rect 535154 269198 541918 269434
rect 542154 269198 548918 269434
rect 549154 269198 555918 269434
rect 556154 269198 562918 269434
rect 563154 269198 569918 269434
rect 570154 269198 576918 269434
rect 577154 269198 587570 269434
rect 587806 269198 587890 269434
rect 588126 269198 588210 269434
rect 588446 269198 588530 269434
rect 588766 269198 588874 269434
rect -4950 269156 588874 269198
rect -4950 268494 588874 268536
rect -4950 268258 -3090 268494
rect -2854 268258 -2770 268494
rect -2534 268258 -2450 268494
rect -2214 268258 -2130 268494
rect -1894 268258 1186 268494
rect 1422 268258 8186 268494
rect 8422 268258 15186 268494
rect 15422 268258 22186 268494
rect 22422 268258 29186 268494
rect 29422 268258 36186 268494
rect 36422 268258 43186 268494
rect 43422 268258 50186 268494
rect 50422 268258 57186 268494
rect 57422 268258 64186 268494
rect 64422 268258 71186 268494
rect 71422 268258 78186 268494
rect 78422 268258 85186 268494
rect 85422 268258 92186 268494
rect 92422 268258 99186 268494
rect 99422 268258 106186 268494
rect 106422 268258 113186 268494
rect 113422 268258 120186 268494
rect 120422 268258 127186 268494
rect 127422 268258 134186 268494
rect 134422 268258 141186 268494
rect 141422 268258 148186 268494
rect 148422 268258 155186 268494
rect 155422 268258 162186 268494
rect 162422 268258 169186 268494
rect 169422 268258 176186 268494
rect 176422 268258 183186 268494
rect 183422 268258 190186 268494
rect 190422 268258 197186 268494
rect 197422 268258 204186 268494
rect 204422 268258 211186 268494
rect 211422 268258 218186 268494
rect 218422 268258 225186 268494
rect 225422 268258 232186 268494
rect 232422 268258 239186 268494
rect 239422 268258 246186 268494
rect 246422 268258 253186 268494
rect 253422 268258 260186 268494
rect 260422 268258 267186 268494
rect 267422 268258 274186 268494
rect 274422 268258 281186 268494
rect 281422 268258 288186 268494
rect 288422 268258 295186 268494
rect 295422 268258 302186 268494
rect 302422 268258 309186 268494
rect 309422 268258 316186 268494
rect 316422 268258 323186 268494
rect 323422 268258 330186 268494
rect 330422 268258 337186 268494
rect 337422 268258 344186 268494
rect 344422 268258 351186 268494
rect 351422 268258 358186 268494
rect 358422 268258 365186 268494
rect 365422 268258 372186 268494
rect 372422 268258 379186 268494
rect 379422 268258 386186 268494
rect 386422 268258 393186 268494
rect 393422 268258 400186 268494
rect 400422 268258 407186 268494
rect 407422 268258 414186 268494
rect 414422 268258 421186 268494
rect 421422 268258 428186 268494
rect 428422 268258 435186 268494
rect 435422 268258 442186 268494
rect 442422 268258 449186 268494
rect 449422 268258 456186 268494
rect 456422 268258 463186 268494
rect 463422 268258 470186 268494
rect 470422 268258 477186 268494
rect 477422 268258 484186 268494
rect 484422 268258 491186 268494
rect 491422 268258 498186 268494
rect 498422 268258 505186 268494
rect 505422 268258 512186 268494
rect 512422 268258 519186 268494
rect 519422 268258 526186 268494
rect 526422 268258 533186 268494
rect 533422 268258 540186 268494
rect 540422 268258 547186 268494
rect 547422 268258 554186 268494
rect 554422 268258 561186 268494
rect 561422 268258 568186 268494
rect 568422 268258 575186 268494
rect 575422 268258 582186 268494
rect 582422 268258 585818 268494
rect 586054 268258 586138 268494
rect 586374 268258 586458 268494
rect 586694 268258 586778 268494
rect 587014 268258 588874 268494
rect -4950 268216 588874 268258
rect -4950 262434 588874 262476
rect -4950 262198 -4842 262434
rect -4606 262198 -4522 262434
rect -4286 262198 -4202 262434
rect -3966 262198 -3882 262434
rect -3646 262198 2918 262434
rect 3154 262198 9918 262434
rect 10154 262198 16918 262434
rect 17154 262198 23918 262434
rect 24154 262198 30918 262434
rect 31154 262198 37918 262434
rect 38154 262198 44918 262434
rect 45154 262198 51918 262434
rect 52154 262198 58918 262434
rect 59154 262198 65918 262434
rect 66154 262198 72918 262434
rect 73154 262198 79918 262434
rect 80154 262198 86918 262434
rect 87154 262198 93918 262434
rect 94154 262198 100918 262434
rect 101154 262198 107918 262434
rect 108154 262198 114918 262434
rect 115154 262198 121918 262434
rect 122154 262198 128918 262434
rect 129154 262198 135918 262434
rect 136154 262198 142918 262434
rect 143154 262198 149918 262434
rect 150154 262198 156918 262434
rect 157154 262198 163918 262434
rect 164154 262198 170918 262434
rect 171154 262198 177918 262434
rect 178154 262198 184918 262434
rect 185154 262198 191918 262434
rect 192154 262198 198918 262434
rect 199154 262198 205918 262434
rect 206154 262198 212918 262434
rect 213154 262198 219918 262434
rect 220154 262198 226918 262434
rect 227154 262198 233918 262434
rect 234154 262198 240918 262434
rect 241154 262198 247918 262434
rect 248154 262198 254918 262434
rect 255154 262198 261918 262434
rect 262154 262198 268918 262434
rect 269154 262198 275918 262434
rect 276154 262198 282918 262434
rect 283154 262198 289918 262434
rect 290154 262198 296918 262434
rect 297154 262198 303918 262434
rect 304154 262198 310918 262434
rect 311154 262198 317918 262434
rect 318154 262198 324918 262434
rect 325154 262198 331918 262434
rect 332154 262198 338918 262434
rect 339154 262198 345918 262434
rect 346154 262198 352918 262434
rect 353154 262198 359918 262434
rect 360154 262198 366918 262434
rect 367154 262198 373918 262434
rect 374154 262198 380918 262434
rect 381154 262198 387918 262434
rect 388154 262198 394918 262434
rect 395154 262198 401918 262434
rect 402154 262198 408918 262434
rect 409154 262198 415918 262434
rect 416154 262198 422918 262434
rect 423154 262198 429918 262434
rect 430154 262198 436918 262434
rect 437154 262198 443918 262434
rect 444154 262198 450918 262434
rect 451154 262198 457918 262434
rect 458154 262198 464918 262434
rect 465154 262198 471918 262434
rect 472154 262198 478918 262434
rect 479154 262198 485918 262434
rect 486154 262198 492918 262434
rect 493154 262198 499918 262434
rect 500154 262198 506918 262434
rect 507154 262198 513918 262434
rect 514154 262198 520918 262434
rect 521154 262198 527918 262434
rect 528154 262198 534918 262434
rect 535154 262198 541918 262434
rect 542154 262198 548918 262434
rect 549154 262198 555918 262434
rect 556154 262198 562918 262434
rect 563154 262198 569918 262434
rect 570154 262198 576918 262434
rect 577154 262198 587570 262434
rect 587806 262198 587890 262434
rect 588126 262198 588210 262434
rect 588446 262198 588530 262434
rect 588766 262198 588874 262434
rect -4950 262156 588874 262198
rect -4950 261494 588874 261536
rect -4950 261258 -3090 261494
rect -2854 261258 -2770 261494
rect -2534 261258 -2450 261494
rect -2214 261258 -2130 261494
rect -1894 261258 1186 261494
rect 1422 261258 8186 261494
rect 8422 261258 15186 261494
rect 15422 261258 22186 261494
rect 22422 261258 29186 261494
rect 29422 261258 36186 261494
rect 36422 261258 43186 261494
rect 43422 261258 50186 261494
rect 50422 261258 57186 261494
rect 57422 261258 64186 261494
rect 64422 261258 71186 261494
rect 71422 261258 78186 261494
rect 78422 261258 85186 261494
rect 85422 261258 92186 261494
rect 92422 261258 99186 261494
rect 99422 261258 106186 261494
rect 106422 261258 113186 261494
rect 113422 261258 120186 261494
rect 120422 261258 127186 261494
rect 127422 261258 134186 261494
rect 134422 261258 141186 261494
rect 141422 261258 148186 261494
rect 148422 261258 155186 261494
rect 155422 261258 162186 261494
rect 162422 261258 169186 261494
rect 169422 261258 176186 261494
rect 176422 261258 183186 261494
rect 183422 261258 190186 261494
rect 190422 261258 197186 261494
rect 197422 261258 204186 261494
rect 204422 261258 211186 261494
rect 211422 261258 218186 261494
rect 218422 261258 225186 261494
rect 225422 261258 232186 261494
rect 232422 261258 239186 261494
rect 239422 261258 246186 261494
rect 246422 261258 253186 261494
rect 253422 261258 260186 261494
rect 260422 261258 267186 261494
rect 267422 261258 274186 261494
rect 274422 261258 281186 261494
rect 281422 261258 288186 261494
rect 288422 261258 295186 261494
rect 295422 261258 302186 261494
rect 302422 261258 309186 261494
rect 309422 261258 316186 261494
rect 316422 261258 323186 261494
rect 323422 261258 330186 261494
rect 330422 261258 337186 261494
rect 337422 261258 344186 261494
rect 344422 261258 351186 261494
rect 351422 261258 358186 261494
rect 358422 261258 365186 261494
rect 365422 261258 372186 261494
rect 372422 261258 379186 261494
rect 379422 261258 386186 261494
rect 386422 261258 393186 261494
rect 393422 261258 400186 261494
rect 400422 261258 407186 261494
rect 407422 261258 414186 261494
rect 414422 261258 421186 261494
rect 421422 261258 428186 261494
rect 428422 261258 435186 261494
rect 435422 261258 442186 261494
rect 442422 261258 449186 261494
rect 449422 261258 456186 261494
rect 456422 261258 463186 261494
rect 463422 261258 470186 261494
rect 470422 261258 477186 261494
rect 477422 261258 484186 261494
rect 484422 261258 491186 261494
rect 491422 261258 498186 261494
rect 498422 261258 505186 261494
rect 505422 261258 512186 261494
rect 512422 261258 519186 261494
rect 519422 261258 533186 261494
rect 533422 261258 540186 261494
rect 540422 261258 547186 261494
rect 547422 261258 554186 261494
rect 554422 261258 561186 261494
rect 561422 261258 568186 261494
rect 568422 261258 575186 261494
rect 575422 261258 582186 261494
rect 582422 261258 585818 261494
rect 586054 261258 586138 261494
rect 586374 261258 586458 261494
rect 586694 261258 586778 261494
rect 587014 261258 588874 261494
rect -4950 261216 588874 261258
rect -4950 255434 588874 255476
rect -4950 255198 -4842 255434
rect -4606 255198 -4522 255434
rect -4286 255198 -4202 255434
rect -3966 255198 -3882 255434
rect -3646 255198 2918 255434
rect 3154 255198 9918 255434
rect 10154 255198 16918 255434
rect 17154 255198 23918 255434
rect 24154 255198 30918 255434
rect 31154 255198 37918 255434
rect 38154 255198 44918 255434
rect 45154 255198 51918 255434
rect 52154 255198 58918 255434
rect 59154 255198 65918 255434
rect 66154 255198 72918 255434
rect 73154 255198 79918 255434
rect 80154 255198 86918 255434
rect 87154 255198 93918 255434
rect 94154 255198 100918 255434
rect 101154 255198 107918 255434
rect 108154 255198 114918 255434
rect 115154 255198 121918 255434
rect 122154 255198 128918 255434
rect 129154 255198 135918 255434
rect 136154 255198 142918 255434
rect 143154 255198 149918 255434
rect 150154 255198 156918 255434
rect 157154 255198 163918 255434
rect 164154 255198 170918 255434
rect 171154 255198 177918 255434
rect 178154 255198 184918 255434
rect 185154 255198 191918 255434
rect 192154 255198 198918 255434
rect 199154 255198 205918 255434
rect 206154 255198 212918 255434
rect 213154 255198 219918 255434
rect 220154 255198 226918 255434
rect 227154 255198 233918 255434
rect 234154 255198 240918 255434
rect 241154 255198 247918 255434
rect 248154 255198 254918 255434
rect 255154 255198 261918 255434
rect 262154 255198 268918 255434
rect 269154 255198 275918 255434
rect 276154 255198 282918 255434
rect 283154 255198 289918 255434
rect 290154 255198 296918 255434
rect 297154 255198 303918 255434
rect 304154 255198 310918 255434
rect 311154 255198 317918 255434
rect 318154 255198 324918 255434
rect 325154 255198 331918 255434
rect 332154 255198 338918 255434
rect 339154 255198 345918 255434
rect 346154 255198 352918 255434
rect 353154 255198 359918 255434
rect 360154 255198 366918 255434
rect 367154 255198 373918 255434
rect 374154 255198 380918 255434
rect 381154 255198 387918 255434
rect 388154 255198 394918 255434
rect 395154 255198 401918 255434
rect 402154 255198 408918 255434
rect 409154 255198 415918 255434
rect 416154 255198 422918 255434
rect 423154 255198 429918 255434
rect 430154 255198 436918 255434
rect 437154 255198 443918 255434
rect 444154 255198 450918 255434
rect 451154 255198 457918 255434
rect 458154 255198 464918 255434
rect 465154 255198 471918 255434
rect 472154 255198 478918 255434
rect 479154 255198 485918 255434
rect 486154 255198 492918 255434
rect 493154 255198 499918 255434
rect 500154 255198 506918 255434
rect 507154 255198 513918 255434
rect 514154 255198 520918 255434
rect 521154 255198 522850 255434
rect 523086 255198 524782 255434
rect 525018 255198 526714 255434
rect 526950 255198 527918 255434
rect 528154 255198 534918 255434
rect 535154 255198 541918 255434
rect 542154 255198 548918 255434
rect 549154 255198 555918 255434
rect 556154 255198 562918 255434
rect 563154 255198 569918 255434
rect 570154 255198 576918 255434
rect 577154 255198 587570 255434
rect 587806 255198 587890 255434
rect 588126 255198 588210 255434
rect 588446 255198 588530 255434
rect 588766 255198 588874 255434
rect -4950 255156 588874 255198
rect -4950 254494 588874 254536
rect -4950 254258 -3090 254494
rect -2854 254258 -2770 254494
rect -2534 254258 -2450 254494
rect -2214 254258 -2130 254494
rect -1894 254258 1186 254494
rect 1422 254258 8186 254494
rect 8422 254258 15186 254494
rect 15422 254258 22186 254494
rect 22422 254258 29186 254494
rect 29422 254258 36186 254494
rect 36422 254258 43186 254494
rect 43422 254258 50186 254494
rect 50422 254258 57186 254494
rect 57422 254258 64186 254494
rect 64422 254258 71186 254494
rect 71422 254258 78186 254494
rect 78422 254258 85186 254494
rect 85422 254258 92186 254494
rect 92422 254258 99186 254494
rect 99422 254258 106186 254494
rect 106422 254258 113186 254494
rect 113422 254258 120186 254494
rect 120422 254258 127186 254494
rect 127422 254258 134186 254494
rect 134422 254258 141186 254494
rect 141422 254258 148186 254494
rect 148422 254258 155186 254494
rect 155422 254258 162186 254494
rect 162422 254258 169186 254494
rect 169422 254258 176186 254494
rect 176422 254258 183186 254494
rect 183422 254258 190186 254494
rect 190422 254258 197186 254494
rect 197422 254258 204186 254494
rect 204422 254258 211186 254494
rect 211422 254258 218186 254494
rect 218422 254258 225186 254494
rect 225422 254258 232186 254494
rect 232422 254258 239186 254494
rect 239422 254258 246186 254494
rect 246422 254258 253186 254494
rect 253422 254258 260186 254494
rect 260422 254258 267186 254494
rect 267422 254258 274186 254494
rect 274422 254258 281186 254494
rect 281422 254258 288186 254494
rect 288422 254258 295186 254494
rect 295422 254258 302186 254494
rect 302422 254258 309186 254494
rect 309422 254258 316186 254494
rect 316422 254258 323186 254494
rect 323422 254258 330186 254494
rect 330422 254258 337186 254494
rect 337422 254258 344186 254494
rect 344422 254258 351186 254494
rect 351422 254258 358186 254494
rect 358422 254258 365186 254494
rect 365422 254258 372186 254494
rect 372422 254258 379186 254494
rect 379422 254258 386186 254494
rect 386422 254258 393186 254494
rect 393422 254258 400186 254494
rect 400422 254258 407186 254494
rect 407422 254258 414186 254494
rect 414422 254258 421186 254494
rect 421422 254258 428186 254494
rect 428422 254258 435186 254494
rect 435422 254258 442186 254494
rect 442422 254258 449186 254494
rect 449422 254258 456186 254494
rect 456422 254258 463186 254494
rect 463422 254258 470186 254494
rect 470422 254258 477186 254494
rect 477422 254258 484186 254494
rect 484422 254258 491186 254494
rect 491422 254258 498186 254494
rect 498422 254258 505186 254494
rect 505422 254258 512186 254494
rect 512422 254258 519186 254494
rect 519422 254258 519952 254494
rect 520188 254258 521884 254494
rect 522120 254258 523816 254494
rect 524052 254258 525748 254494
rect 525984 254258 533186 254494
rect 533422 254258 540186 254494
rect 540422 254258 547186 254494
rect 547422 254258 554186 254494
rect 554422 254258 561186 254494
rect 561422 254258 568186 254494
rect 568422 254258 575186 254494
rect 575422 254258 582186 254494
rect 582422 254258 585818 254494
rect 586054 254258 586138 254494
rect 586374 254258 586458 254494
rect 586694 254258 586778 254494
rect 587014 254258 588874 254494
rect -4950 254216 588874 254258
rect -4950 248434 588874 248476
rect -4950 248198 -4842 248434
rect -4606 248198 -4522 248434
rect -4286 248198 -4202 248434
rect -3966 248198 -3882 248434
rect -3646 248198 2918 248434
rect 3154 248198 9918 248434
rect 10154 248198 16918 248434
rect 17154 248198 23918 248434
rect 24154 248198 30918 248434
rect 31154 248198 37918 248434
rect 38154 248198 44918 248434
rect 45154 248198 51918 248434
rect 52154 248198 58918 248434
rect 59154 248198 65918 248434
rect 66154 248198 72918 248434
rect 73154 248198 79918 248434
rect 80154 248198 86918 248434
rect 87154 248198 93918 248434
rect 94154 248198 100918 248434
rect 101154 248198 107918 248434
rect 108154 248198 114918 248434
rect 115154 248198 121918 248434
rect 122154 248198 128918 248434
rect 129154 248198 135918 248434
rect 136154 248198 142918 248434
rect 143154 248198 149918 248434
rect 150154 248198 156918 248434
rect 157154 248198 163918 248434
rect 164154 248198 170918 248434
rect 171154 248198 177918 248434
rect 178154 248198 184918 248434
rect 185154 248198 191918 248434
rect 192154 248198 198918 248434
rect 199154 248198 205918 248434
rect 206154 248198 212918 248434
rect 213154 248198 219918 248434
rect 220154 248198 226918 248434
rect 227154 248198 233918 248434
rect 234154 248198 240918 248434
rect 241154 248198 247918 248434
rect 248154 248198 254918 248434
rect 255154 248198 261918 248434
rect 262154 248198 268918 248434
rect 269154 248198 275918 248434
rect 276154 248198 282918 248434
rect 283154 248198 289918 248434
rect 290154 248198 296918 248434
rect 297154 248198 303918 248434
rect 304154 248198 310918 248434
rect 311154 248198 317918 248434
rect 318154 248198 324918 248434
rect 325154 248198 331918 248434
rect 332154 248198 338918 248434
rect 339154 248198 345918 248434
rect 346154 248198 352918 248434
rect 353154 248198 359918 248434
rect 360154 248198 366918 248434
rect 367154 248198 373918 248434
rect 374154 248198 380918 248434
rect 381154 248198 387918 248434
rect 388154 248198 394918 248434
rect 395154 248198 401918 248434
rect 402154 248198 408918 248434
rect 409154 248198 415918 248434
rect 416154 248198 422918 248434
rect 423154 248198 429918 248434
rect 430154 248198 436918 248434
rect 437154 248198 443918 248434
rect 444154 248198 450918 248434
rect 451154 248198 457918 248434
rect 458154 248198 464918 248434
rect 465154 248198 471918 248434
rect 472154 248198 478918 248434
rect 479154 248198 485918 248434
rect 486154 248198 492918 248434
rect 493154 248198 499918 248434
rect 500154 248198 506918 248434
rect 507154 248198 513918 248434
rect 514154 248198 520918 248434
rect 521154 248198 522850 248434
rect 523086 248198 524782 248434
rect 525018 248198 526714 248434
rect 526950 248198 527918 248434
rect 528154 248198 534918 248434
rect 535154 248198 541918 248434
rect 542154 248198 548918 248434
rect 549154 248198 555918 248434
rect 556154 248198 562918 248434
rect 563154 248198 569918 248434
rect 570154 248198 576918 248434
rect 577154 248198 587570 248434
rect 587806 248198 587890 248434
rect 588126 248198 588210 248434
rect 588446 248198 588530 248434
rect 588766 248198 588874 248434
rect -4950 248156 588874 248198
rect -4950 247494 588874 247536
rect -4950 247258 -3090 247494
rect -2854 247258 -2770 247494
rect -2534 247258 -2450 247494
rect -2214 247258 -2130 247494
rect -1894 247258 1186 247494
rect 1422 247258 8186 247494
rect 8422 247258 15186 247494
rect 15422 247258 22186 247494
rect 22422 247258 29186 247494
rect 29422 247258 36186 247494
rect 36422 247258 43186 247494
rect 43422 247258 50186 247494
rect 50422 247258 57186 247494
rect 57422 247258 64186 247494
rect 64422 247258 71186 247494
rect 71422 247258 78186 247494
rect 78422 247258 85186 247494
rect 85422 247258 92186 247494
rect 92422 247258 99186 247494
rect 99422 247258 106186 247494
rect 106422 247258 113186 247494
rect 113422 247258 120186 247494
rect 120422 247258 127186 247494
rect 127422 247258 134186 247494
rect 134422 247258 141186 247494
rect 141422 247258 148186 247494
rect 148422 247258 155186 247494
rect 155422 247258 162186 247494
rect 162422 247258 169186 247494
rect 169422 247258 176186 247494
rect 176422 247258 183186 247494
rect 183422 247258 190186 247494
rect 190422 247258 197186 247494
rect 197422 247258 204186 247494
rect 204422 247258 211186 247494
rect 211422 247258 218186 247494
rect 218422 247258 225186 247494
rect 225422 247258 232186 247494
rect 232422 247258 239186 247494
rect 239422 247258 246186 247494
rect 246422 247258 253186 247494
rect 253422 247258 260186 247494
rect 260422 247258 267186 247494
rect 267422 247258 274186 247494
rect 274422 247258 281186 247494
rect 281422 247258 288186 247494
rect 288422 247258 295186 247494
rect 295422 247258 302186 247494
rect 302422 247258 309186 247494
rect 309422 247258 316186 247494
rect 316422 247258 323186 247494
rect 323422 247258 330186 247494
rect 330422 247258 337186 247494
rect 337422 247258 344186 247494
rect 344422 247258 351186 247494
rect 351422 247258 358186 247494
rect 358422 247258 365186 247494
rect 365422 247258 372186 247494
rect 372422 247258 379186 247494
rect 379422 247258 386186 247494
rect 386422 247258 393186 247494
rect 393422 247258 400186 247494
rect 400422 247258 407186 247494
rect 407422 247258 414186 247494
rect 414422 247258 421186 247494
rect 421422 247258 428186 247494
rect 428422 247258 435186 247494
rect 435422 247258 442186 247494
rect 442422 247258 449186 247494
rect 449422 247258 456186 247494
rect 456422 247258 463186 247494
rect 463422 247258 470186 247494
rect 470422 247258 477186 247494
rect 477422 247258 484186 247494
rect 484422 247258 491186 247494
rect 491422 247258 498186 247494
rect 498422 247258 505186 247494
rect 505422 247258 512186 247494
rect 512422 247258 519186 247494
rect 519422 247258 519952 247494
rect 520188 247258 521884 247494
rect 522120 247258 523816 247494
rect 524052 247258 525748 247494
rect 525984 247258 533186 247494
rect 533422 247258 540186 247494
rect 540422 247258 547186 247494
rect 547422 247258 554186 247494
rect 554422 247258 561186 247494
rect 561422 247258 568186 247494
rect 568422 247258 575186 247494
rect 575422 247258 582186 247494
rect 582422 247258 585818 247494
rect 586054 247258 586138 247494
rect 586374 247258 586458 247494
rect 586694 247258 586778 247494
rect 587014 247258 588874 247494
rect -4950 247216 588874 247258
rect -4950 241434 588874 241476
rect -4950 241198 -4842 241434
rect -4606 241198 -4522 241434
rect -4286 241198 -4202 241434
rect -3966 241198 -3882 241434
rect -3646 241198 2918 241434
rect 3154 241198 9918 241434
rect 10154 241198 16918 241434
rect 17154 241198 23918 241434
rect 24154 241198 30918 241434
rect 31154 241198 37918 241434
rect 38154 241198 44918 241434
rect 45154 241198 51918 241434
rect 52154 241198 58918 241434
rect 59154 241198 65918 241434
rect 66154 241198 72918 241434
rect 73154 241198 79918 241434
rect 80154 241198 86918 241434
rect 87154 241198 93918 241434
rect 94154 241198 100918 241434
rect 101154 241198 107918 241434
rect 108154 241198 114918 241434
rect 115154 241198 121918 241434
rect 122154 241198 128918 241434
rect 129154 241198 135918 241434
rect 136154 241198 142918 241434
rect 143154 241198 149918 241434
rect 150154 241198 156918 241434
rect 157154 241198 163918 241434
rect 164154 241198 170918 241434
rect 171154 241198 177918 241434
rect 178154 241198 184918 241434
rect 185154 241198 191918 241434
rect 192154 241198 198918 241434
rect 199154 241198 205918 241434
rect 206154 241198 212918 241434
rect 213154 241198 219918 241434
rect 220154 241198 226918 241434
rect 227154 241198 233918 241434
rect 234154 241198 240918 241434
rect 241154 241198 247918 241434
rect 248154 241198 254918 241434
rect 255154 241198 261918 241434
rect 262154 241198 268918 241434
rect 269154 241198 275918 241434
rect 276154 241198 282918 241434
rect 283154 241198 289918 241434
rect 290154 241198 296918 241434
rect 297154 241198 303918 241434
rect 304154 241198 310918 241434
rect 311154 241198 317918 241434
rect 318154 241198 324918 241434
rect 325154 241198 331918 241434
rect 332154 241198 338918 241434
rect 339154 241198 345918 241434
rect 346154 241198 352918 241434
rect 353154 241198 359918 241434
rect 360154 241198 366918 241434
rect 367154 241198 373918 241434
rect 374154 241198 380918 241434
rect 381154 241198 387918 241434
rect 388154 241198 394918 241434
rect 395154 241198 401918 241434
rect 402154 241198 408918 241434
rect 409154 241198 415918 241434
rect 416154 241198 422918 241434
rect 423154 241198 429918 241434
rect 430154 241198 436918 241434
rect 437154 241198 443918 241434
rect 444154 241198 450918 241434
rect 451154 241198 457918 241434
rect 458154 241198 464918 241434
rect 465154 241198 471918 241434
rect 472154 241198 478918 241434
rect 479154 241198 485918 241434
rect 486154 241198 492918 241434
rect 493154 241198 499918 241434
rect 500154 241198 506918 241434
rect 507154 241198 513918 241434
rect 514154 241198 527918 241434
rect 528154 241198 534918 241434
rect 535154 241198 541918 241434
rect 542154 241198 548918 241434
rect 549154 241198 555918 241434
rect 556154 241198 562918 241434
rect 563154 241198 569918 241434
rect 570154 241198 576918 241434
rect 577154 241198 587570 241434
rect 587806 241198 587890 241434
rect 588126 241198 588210 241434
rect 588446 241198 588530 241434
rect 588766 241198 588874 241434
rect -4950 241156 588874 241198
rect -4950 240494 588874 240536
rect -4950 240258 -3090 240494
rect -2854 240258 -2770 240494
rect -2534 240258 -2450 240494
rect -2214 240258 -2130 240494
rect -1894 240258 1186 240494
rect 1422 240258 8186 240494
rect 8422 240258 15186 240494
rect 15422 240258 22186 240494
rect 22422 240258 29186 240494
rect 29422 240258 36186 240494
rect 36422 240258 43186 240494
rect 43422 240258 50186 240494
rect 50422 240258 57186 240494
rect 57422 240258 64186 240494
rect 64422 240258 71186 240494
rect 71422 240258 78186 240494
rect 78422 240258 85186 240494
rect 85422 240258 92186 240494
rect 92422 240258 99186 240494
rect 99422 240258 106186 240494
rect 106422 240258 113186 240494
rect 113422 240258 120186 240494
rect 120422 240258 127186 240494
rect 127422 240258 134186 240494
rect 134422 240258 141186 240494
rect 141422 240258 148186 240494
rect 148422 240258 155186 240494
rect 155422 240258 162186 240494
rect 162422 240258 169186 240494
rect 169422 240258 176186 240494
rect 176422 240258 183186 240494
rect 183422 240258 190186 240494
rect 190422 240258 197186 240494
rect 197422 240258 204186 240494
rect 204422 240258 211186 240494
rect 211422 240258 218186 240494
rect 218422 240258 225186 240494
rect 225422 240258 232186 240494
rect 232422 240258 239186 240494
rect 239422 240258 246186 240494
rect 246422 240258 253186 240494
rect 253422 240258 260186 240494
rect 260422 240258 267186 240494
rect 267422 240258 274186 240494
rect 274422 240258 281186 240494
rect 281422 240258 288186 240494
rect 288422 240258 295186 240494
rect 295422 240258 302186 240494
rect 302422 240258 309186 240494
rect 309422 240258 316186 240494
rect 316422 240258 323186 240494
rect 323422 240258 330186 240494
rect 330422 240258 337186 240494
rect 337422 240258 344186 240494
rect 344422 240258 351186 240494
rect 351422 240258 358186 240494
rect 358422 240258 365186 240494
rect 365422 240258 372186 240494
rect 372422 240258 379186 240494
rect 379422 240258 386186 240494
rect 386422 240258 393186 240494
rect 393422 240258 400186 240494
rect 400422 240258 407186 240494
rect 407422 240258 414186 240494
rect 414422 240258 421186 240494
rect 421422 240258 428186 240494
rect 428422 240258 435186 240494
rect 435422 240258 442186 240494
rect 442422 240258 449186 240494
rect 449422 240258 456186 240494
rect 456422 240258 463186 240494
rect 463422 240258 470186 240494
rect 470422 240258 477186 240494
rect 477422 240258 484186 240494
rect 484422 240258 491186 240494
rect 491422 240258 498186 240494
rect 498422 240258 505186 240494
rect 505422 240258 512186 240494
rect 512422 240258 519186 240494
rect 519422 240258 533186 240494
rect 533422 240258 540186 240494
rect 540422 240258 547186 240494
rect 547422 240258 554186 240494
rect 554422 240258 561186 240494
rect 561422 240258 568186 240494
rect 568422 240258 575186 240494
rect 575422 240258 582186 240494
rect 582422 240258 585818 240494
rect 586054 240258 586138 240494
rect 586374 240258 586458 240494
rect 586694 240258 586778 240494
rect 587014 240258 588874 240494
rect -4950 240216 588874 240258
rect -4950 234434 588874 234476
rect -4950 234198 -4842 234434
rect -4606 234198 -4522 234434
rect -4286 234198 -4202 234434
rect -3966 234198 -3882 234434
rect -3646 234198 2918 234434
rect 3154 234198 9918 234434
rect 10154 234198 16918 234434
rect 17154 234198 23918 234434
rect 24154 234198 30918 234434
rect 31154 234198 37918 234434
rect 38154 234198 44918 234434
rect 45154 234198 51918 234434
rect 52154 234198 58918 234434
rect 59154 234198 65918 234434
rect 66154 234198 72918 234434
rect 73154 234198 79918 234434
rect 80154 234198 86918 234434
rect 87154 234198 93918 234434
rect 94154 234198 100918 234434
rect 101154 234198 107918 234434
rect 108154 234198 114918 234434
rect 115154 234198 121918 234434
rect 122154 234198 128918 234434
rect 129154 234198 135918 234434
rect 136154 234198 142918 234434
rect 143154 234198 149918 234434
rect 150154 234198 156918 234434
rect 157154 234198 163918 234434
rect 164154 234198 170918 234434
rect 171154 234198 177918 234434
rect 178154 234198 184918 234434
rect 185154 234198 191918 234434
rect 192154 234198 198918 234434
rect 199154 234198 205918 234434
rect 206154 234198 212918 234434
rect 213154 234198 219918 234434
rect 220154 234198 226918 234434
rect 227154 234198 233918 234434
rect 234154 234198 240918 234434
rect 241154 234198 247918 234434
rect 248154 234198 254918 234434
rect 255154 234198 261918 234434
rect 262154 234198 268918 234434
rect 269154 234198 275918 234434
rect 276154 234198 282918 234434
rect 283154 234198 289918 234434
rect 290154 234198 296918 234434
rect 297154 234198 303918 234434
rect 304154 234198 310918 234434
rect 311154 234198 317918 234434
rect 318154 234198 324918 234434
rect 325154 234198 331918 234434
rect 332154 234198 338918 234434
rect 339154 234198 345918 234434
rect 346154 234198 352918 234434
rect 353154 234198 359918 234434
rect 360154 234198 366918 234434
rect 367154 234198 373918 234434
rect 374154 234198 380918 234434
rect 381154 234198 387918 234434
rect 388154 234198 394918 234434
rect 395154 234198 401918 234434
rect 402154 234198 408918 234434
rect 409154 234198 415918 234434
rect 416154 234198 422918 234434
rect 423154 234198 429918 234434
rect 430154 234198 436918 234434
rect 437154 234198 443918 234434
rect 444154 234198 450918 234434
rect 451154 234198 457918 234434
rect 458154 234198 464918 234434
rect 465154 234198 471918 234434
rect 472154 234198 478918 234434
rect 479154 234198 485918 234434
rect 486154 234198 492918 234434
rect 493154 234198 499918 234434
rect 500154 234198 506918 234434
rect 507154 234198 513918 234434
rect 514154 234198 520918 234434
rect 521154 234198 527918 234434
rect 528154 234198 534918 234434
rect 535154 234198 541918 234434
rect 542154 234198 548918 234434
rect 549154 234198 555918 234434
rect 556154 234198 562918 234434
rect 563154 234198 569918 234434
rect 570154 234198 576918 234434
rect 577154 234198 587570 234434
rect 587806 234198 587890 234434
rect 588126 234198 588210 234434
rect 588446 234198 588530 234434
rect 588766 234198 588874 234434
rect -4950 234156 588874 234198
rect -4950 233494 588874 233536
rect -4950 233258 -3090 233494
rect -2854 233258 -2770 233494
rect -2534 233258 -2450 233494
rect -2214 233258 -2130 233494
rect -1894 233258 1186 233494
rect 1422 233258 8186 233494
rect 8422 233258 15186 233494
rect 15422 233258 22186 233494
rect 22422 233258 29186 233494
rect 29422 233258 36186 233494
rect 36422 233258 43186 233494
rect 43422 233258 50186 233494
rect 50422 233258 57186 233494
rect 57422 233258 64186 233494
rect 64422 233258 71186 233494
rect 71422 233258 78186 233494
rect 78422 233258 85186 233494
rect 85422 233258 92186 233494
rect 92422 233258 99186 233494
rect 99422 233258 106186 233494
rect 106422 233258 113186 233494
rect 113422 233258 120186 233494
rect 120422 233258 127186 233494
rect 127422 233258 134186 233494
rect 134422 233258 141186 233494
rect 141422 233258 148186 233494
rect 148422 233258 155186 233494
rect 155422 233258 162186 233494
rect 162422 233258 169186 233494
rect 169422 233258 176186 233494
rect 176422 233258 183186 233494
rect 183422 233258 190186 233494
rect 190422 233258 197186 233494
rect 197422 233258 204186 233494
rect 204422 233258 211186 233494
rect 211422 233258 218186 233494
rect 218422 233258 225186 233494
rect 225422 233258 232186 233494
rect 232422 233258 239186 233494
rect 239422 233258 246186 233494
rect 246422 233258 253186 233494
rect 253422 233258 260186 233494
rect 260422 233258 267186 233494
rect 267422 233258 274186 233494
rect 274422 233258 281186 233494
rect 281422 233258 288186 233494
rect 288422 233258 295186 233494
rect 295422 233258 302186 233494
rect 302422 233258 309186 233494
rect 309422 233258 316186 233494
rect 316422 233258 323186 233494
rect 323422 233258 330186 233494
rect 330422 233258 337186 233494
rect 337422 233258 344186 233494
rect 344422 233258 351186 233494
rect 351422 233258 358186 233494
rect 358422 233258 365186 233494
rect 365422 233258 372186 233494
rect 372422 233258 379186 233494
rect 379422 233258 386186 233494
rect 386422 233258 393186 233494
rect 393422 233258 400186 233494
rect 400422 233258 407186 233494
rect 407422 233258 414186 233494
rect 414422 233258 421186 233494
rect 421422 233258 428186 233494
rect 428422 233258 435186 233494
rect 435422 233258 442186 233494
rect 442422 233258 449186 233494
rect 449422 233258 456186 233494
rect 456422 233258 463186 233494
rect 463422 233258 470186 233494
rect 470422 233258 477186 233494
rect 477422 233258 484186 233494
rect 484422 233258 491186 233494
rect 491422 233258 498186 233494
rect 498422 233258 505186 233494
rect 505422 233258 512186 233494
rect 512422 233258 519186 233494
rect 519422 233258 526186 233494
rect 526422 233258 533186 233494
rect 533422 233258 540186 233494
rect 540422 233258 547186 233494
rect 547422 233258 554186 233494
rect 554422 233258 561186 233494
rect 561422 233258 568186 233494
rect 568422 233258 575186 233494
rect 575422 233258 582186 233494
rect 582422 233258 585818 233494
rect 586054 233258 586138 233494
rect 586374 233258 586458 233494
rect 586694 233258 586778 233494
rect 587014 233258 588874 233494
rect -4950 233216 588874 233258
rect -4950 227434 588874 227476
rect -4950 227198 -4842 227434
rect -4606 227198 -4522 227434
rect -4286 227198 -4202 227434
rect -3966 227198 -3882 227434
rect -3646 227198 2918 227434
rect 3154 227198 9918 227434
rect 10154 227198 16918 227434
rect 17154 227198 23918 227434
rect 24154 227198 30918 227434
rect 31154 227198 37918 227434
rect 38154 227198 44918 227434
rect 45154 227198 51918 227434
rect 52154 227198 58918 227434
rect 59154 227198 65918 227434
rect 66154 227198 72918 227434
rect 73154 227198 79918 227434
rect 80154 227198 86918 227434
rect 87154 227198 93918 227434
rect 94154 227198 100918 227434
rect 101154 227198 107918 227434
rect 108154 227198 114918 227434
rect 115154 227198 121918 227434
rect 122154 227198 128918 227434
rect 129154 227198 135918 227434
rect 136154 227198 142918 227434
rect 143154 227198 149918 227434
rect 150154 227198 156918 227434
rect 157154 227198 163918 227434
rect 164154 227198 170918 227434
rect 171154 227198 177918 227434
rect 178154 227198 184918 227434
rect 185154 227198 191918 227434
rect 192154 227198 198918 227434
rect 199154 227198 205918 227434
rect 206154 227198 212918 227434
rect 213154 227198 219918 227434
rect 220154 227198 226918 227434
rect 227154 227198 233918 227434
rect 234154 227198 240918 227434
rect 241154 227198 247918 227434
rect 248154 227198 254918 227434
rect 255154 227198 261918 227434
rect 262154 227198 268918 227434
rect 269154 227198 275918 227434
rect 276154 227198 282918 227434
rect 283154 227198 289918 227434
rect 290154 227198 296918 227434
rect 297154 227198 303918 227434
rect 304154 227198 310918 227434
rect 311154 227198 317918 227434
rect 318154 227198 324918 227434
rect 325154 227198 331918 227434
rect 332154 227198 338918 227434
rect 339154 227198 345918 227434
rect 346154 227198 352918 227434
rect 353154 227198 359918 227434
rect 360154 227198 366918 227434
rect 367154 227198 373918 227434
rect 374154 227198 380918 227434
rect 381154 227198 387918 227434
rect 388154 227198 394918 227434
rect 395154 227198 401918 227434
rect 402154 227198 408918 227434
rect 409154 227198 415918 227434
rect 416154 227198 422918 227434
rect 423154 227198 429918 227434
rect 430154 227198 436918 227434
rect 437154 227198 443918 227434
rect 444154 227198 450918 227434
rect 451154 227198 457918 227434
rect 458154 227198 464918 227434
rect 465154 227198 471918 227434
rect 472154 227198 478918 227434
rect 479154 227198 485918 227434
rect 486154 227198 492918 227434
rect 493154 227198 499918 227434
rect 500154 227198 506918 227434
rect 507154 227198 513918 227434
rect 514154 227198 520918 227434
rect 521154 227198 527918 227434
rect 528154 227198 534918 227434
rect 535154 227198 541918 227434
rect 542154 227198 548918 227434
rect 549154 227198 555918 227434
rect 556154 227198 562918 227434
rect 563154 227198 569918 227434
rect 570154 227198 576918 227434
rect 577154 227198 587570 227434
rect 587806 227198 587890 227434
rect 588126 227198 588210 227434
rect 588446 227198 588530 227434
rect 588766 227198 588874 227434
rect -4950 227156 588874 227198
rect -4950 226494 588874 226536
rect -4950 226258 -3090 226494
rect -2854 226258 -2770 226494
rect -2534 226258 -2450 226494
rect -2214 226258 -2130 226494
rect -1894 226258 1186 226494
rect 1422 226258 8186 226494
rect 8422 226258 15186 226494
rect 15422 226258 22186 226494
rect 22422 226258 29186 226494
rect 29422 226258 36186 226494
rect 36422 226258 43186 226494
rect 43422 226258 50186 226494
rect 50422 226258 57186 226494
rect 57422 226258 64186 226494
rect 64422 226258 71186 226494
rect 71422 226258 78186 226494
rect 78422 226258 85186 226494
rect 85422 226258 92186 226494
rect 92422 226258 99186 226494
rect 99422 226258 106186 226494
rect 106422 226258 113186 226494
rect 113422 226258 120186 226494
rect 120422 226258 127186 226494
rect 127422 226258 134186 226494
rect 134422 226258 141186 226494
rect 141422 226258 148186 226494
rect 148422 226258 155186 226494
rect 155422 226258 162186 226494
rect 162422 226258 169186 226494
rect 169422 226258 176186 226494
rect 176422 226258 183186 226494
rect 183422 226258 190186 226494
rect 190422 226258 197186 226494
rect 197422 226258 204186 226494
rect 204422 226258 211186 226494
rect 211422 226258 218186 226494
rect 218422 226258 225186 226494
rect 225422 226258 232186 226494
rect 232422 226258 239186 226494
rect 239422 226258 246186 226494
rect 246422 226258 253186 226494
rect 253422 226258 260186 226494
rect 260422 226258 267186 226494
rect 267422 226258 274186 226494
rect 274422 226258 281186 226494
rect 281422 226258 288186 226494
rect 288422 226258 295186 226494
rect 295422 226258 302186 226494
rect 302422 226258 309186 226494
rect 309422 226258 316186 226494
rect 316422 226258 323186 226494
rect 323422 226258 330186 226494
rect 330422 226258 337186 226494
rect 337422 226258 344186 226494
rect 344422 226258 351186 226494
rect 351422 226258 358186 226494
rect 358422 226258 365186 226494
rect 365422 226258 372186 226494
rect 372422 226258 379186 226494
rect 379422 226258 386186 226494
rect 386422 226258 393186 226494
rect 393422 226258 400186 226494
rect 400422 226258 407186 226494
rect 407422 226258 414186 226494
rect 414422 226258 421186 226494
rect 421422 226258 428186 226494
rect 428422 226258 435186 226494
rect 435422 226258 442186 226494
rect 442422 226258 449186 226494
rect 449422 226258 456186 226494
rect 456422 226258 463186 226494
rect 463422 226258 470186 226494
rect 470422 226258 477186 226494
rect 477422 226258 484186 226494
rect 484422 226258 491186 226494
rect 491422 226258 498186 226494
rect 498422 226258 505186 226494
rect 505422 226258 512186 226494
rect 512422 226258 519186 226494
rect 519422 226258 526186 226494
rect 526422 226258 533186 226494
rect 533422 226258 540186 226494
rect 540422 226258 547186 226494
rect 547422 226258 554186 226494
rect 554422 226258 561186 226494
rect 561422 226258 568186 226494
rect 568422 226258 575186 226494
rect 575422 226258 582186 226494
rect 582422 226258 585818 226494
rect 586054 226258 586138 226494
rect 586374 226258 586458 226494
rect 586694 226258 586778 226494
rect 587014 226258 588874 226494
rect -4950 226216 588874 226258
rect -4950 220434 588874 220476
rect -4950 220198 -4842 220434
rect -4606 220198 -4522 220434
rect -4286 220198 -4202 220434
rect -3966 220198 -3882 220434
rect -3646 220198 2918 220434
rect 3154 220198 9918 220434
rect 10154 220198 16918 220434
rect 17154 220198 23918 220434
rect 24154 220198 30918 220434
rect 31154 220198 37918 220434
rect 38154 220198 44918 220434
rect 45154 220198 51918 220434
rect 52154 220198 58918 220434
rect 59154 220198 65918 220434
rect 66154 220198 72918 220434
rect 73154 220198 79918 220434
rect 80154 220198 86918 220434
rect 87154 220198 93918 220434
rect 94154 220198 100918 220434
rect 101154 220198 107918 220434
rect 108154 220198 114918 220434
rect 115154 220198 121918 220434
rect 122154 220198 128918 220434
rect 129154 220198 135918 220434
rect 136154 220198 142918 220434
rect 143154 220198 149918 220434
rect 150154 220198 156918 220434
rect 157154 220198 163918 220434
rect 164154 220198 170918 220434
rect 171154 220198 177918 220434
rect 178154 220198 184918 220434
rect 185154 220198 191918 220434
rect 192154 220198 198918 220434
rect 199154 220198 205918 220434
rect 206154 220198 212918 220434
rect 213154 220198 219918 220434
rect 220154 220198 226918 220434
rect 227154 220198 233918 220434
rect 234154 220198 240918 220434
rect 241154 220198 247918 220434
rect 248154 220198 254918 220434
rect 255154 220198 261918 220434
rect 262154 220198 268918 220434
rect 269154 220198 275918 220434
rect 276154 220198 282918 220434
rect 283154 220198 289918 220434
rect 290154 220198 296918 220434
rect 297154 220198 303918 220434
rect 304154 220198 310918 220434
rect 311154 220198 317918 220434
rect 318154 220198 324918 220434
rect 325154 220198 331918 220434
rect 332154 220198 338918 220434
rect 339154 220198 345918 220434
rect 346154 220198 352918 220434
rect 353154 220198 359918 220434
rect 360154 220198 366918 220434
rect 367154 220198 373918 220434
rect 374154 220198 380918 220434
rect 381154 220198 387918 220434
rect 388154 220198 394918 220434
rect 395154 220198 401918 220434
rect 402154 220198 408918 220434
rect 409154 220198 415918 220434
rect 416154 220198 422918 220434
rect 423154 220198 429918 220434
rect 430154 220198 436918 220434
rect 437154 220198 443918 220434
rect 444154 220198 450918 220434
rect 451154 220198 457918 220434
rect 458154 220198 464918 220434
rect 465154 220198 471918 220434
rect 472154 220198 478918 220434
rect 479154 220198 485918 220434
rect 486154 220198 492918 220434
rect 493154 220198 499918 220434
rect 500154 220198 506918 220434
rect 507154 220198 513918 220434
rect 514154 220198 520918 220434
rect 521154 220198 527918 220434
rect 528154 220198 534918 220434
rect 535154 220198 541918 220434
rect 542154 220198 548918 220434
rect 549154 220198 555918 220434
rect 556154 220198 562918 220434
rect 563154 220198 569918 220434
rect 570154 220198 576918 220434
rect 577154 220198 587570 220434
rect 587806 220198 587890 220434
rect 588126 220198 588210 220434
rect 588446 220198 588530 220434
rect 588766 220198 588874 220434
rect -4950 220156 588874 220198
rect -4950 219494 588874 219536
rect -4950 219258 -3090 219494
rect -2854 219258 -2770 219494
rect -2534 219258 -2450 219494
rect -2214 219258 -2130 219494
rect -1894 219258 1186 219494
rect 1422 219258 8186 219494
rect 8422 219258 15186 219494
rect 15422 219258 22186 219494
rect 22422 219258 29186 219494
rect 29422 219258 36186 219494
rect 36422 219258 43186 219494
rect 43422 219258 50186 219494
rect 50422 219258 57186 219494
rect 57422 219258 64186 219494
rect 64422 219258 71186 219494
rect 71422 219258 78186 219494
rect 78422 219258 85186 219494
rect 85422 219258 92186 219494
rect 92422 219258 99186 219494
rect 99422 219258 106186 219494
rect 106422 219258 113186 219494
rect 113422 219258 120186 219494
rect 120422 219258 127186 219494
rect 127422 219258 134186 219494
rect 134422 219258 141186 219494
rect 141422 219258 148186 219494
rect 148422 219258 155186 219494
rect 155422 219258 162186 219494
rect 162422 219258 169186 219494
rect 169422 219258 176186 219494
rect 176422 219258 183186 219494
rect 183422 219258 190186 219494
rect 190422 219258 197186 219494
rect 197422 219258 204186 219494
rect 204422 219258 211186 219494
rect 211422 219258 218186 219494
rect 218422 219258 225186 219494
rect 225422 219258 232186 219494
rect 232422 219258 239186 219494
rect 239422 219258 246186 219494
rect 246422 219258 253186 219494
rect 253422 219258 260186 219494
rect 260422 219258 267186 219494
rect 267422 219258 274186 219494
rect 274422 219258 281186 219494
rect 281422 219258 288186 219494
rect 288422 219258 295186 219494
rect 295422 219258 302186 219494
rect 302422 219258 309186 219494
rect 309422 219258 316186 219494
rect 316422 219258 323186 219494
rect 323422 219258 330186 219494
rect 330422 219258 337186 219494
rect 337422 219258 344186 219494
rect 344422 219258 351186 219494
rect 351422 219258 358186 219494
rect 358422 219258 365186 219494
rect 365422 219258 372186 219494
rect 372422 219258 379186 219494
rect 379422 219258 386186 219494
rect 386422 219258 393186 219494
rect 393422 219258 400186 219494
rect 400422 219258 407186 219494
rect 407422 219258 414186 219494
rect 414422 219258 421186 219494
rect 421422 219258 428186 219494
rect 428422 219258 435186 219494
rect 435422 219258 442186 219494
rect 442422 219258 449186 219494
rect 449422 219258 456186 219494
rect 456422 219258 463186 219494
rect 463422 219258 470186 219494
rect 470422 219258 477186 219494
rect 477422 219258 484186 219494
rect 484422 219258 491186 219494
rect 491422 219258 498186 219494
rect 498422 219258 505186 219494
rect 505422 219258 512186 219494
rect 512422 219258 519186 219494
rect 519422 219258 526186 219494
rect 526422 219258 533186 219494
rect 533422 219258 540186 219494
rect 540422 219258 547186 219494
rect 547422 219258 554186 219494
rect 554422 219258 561186 219494
rect 561422 219258 568186 219494
rect 568422 219258 575186 219494
rect 575422 219258 582186 219494
rect 582422 219258 585818 219494
rect 586054 219258 586138 219494
rect 586374 219258 586458 219494
rect 586694 219258 586778 219494
rect 587014 219258 588874 219494
rect -4950 219216 588874 219258
rect -4950 213434 588874 213476
rect -4950 213198 -4842 213434
rect -4606 213198 -4522 213434
rect -4286 213198 -4202 213434
rect -3966 213198 -3882 213434
rect -3646 213198 2918 213434
rect 3154 213198 9918 213434
rect 10154 213198 16918 213434
rect 17154 213198 23918 213434
rect 24154 213198 30918 213434
rect 31154 213198 37918 213434
rect 38154 213198 44918 213434
rect 45154 213198 51918 213434
rect 52154 213198 58918 213434
rect 59154 213198 65918 213434
rect 66154 213198 72918 213434
rect 73154 213198 79918 213434
rect 80154 213198 86918 213434
rect 87154 213198 93918 213434
rect 94154 213198 100918 213434
rect 101154 213198 107918 213434
rect 108154 213198 114918 213434
rect 115154 213198 121918 213434
rect 122154 213198 128918 213434
rect 129154 213198 135918 213434
rect 136154 213198 142918 213434
rect 143154 213198 149918 213434
rect 150154 213198 156918 213434
rect 157154 213198 163918 213434
rect 164154 213198 170918 213434
rect 171154 213198 177918 213434
rect 178154 213198 184918 213434
rect 185154 213198 191918 213434
rect 192154 213198 198918 213434
rect 199154 213198 205918 213434
rect 206154 213198 212918 213434
rect 213154 213198 219918 213434
rect 220154 213198 226918 213434
rect 227154 213198 233918 213434
rect 234154 213198 240918 213434
rect 241154 213198 247918 213434
rect 248154 213198 254918 213434
rect 255154 213198 261918 213434
rect 262154 213198 268918 213434
rect 269154 213198 275918 213434
rect 276154 213198 282918 213434
rect 283154 213198 289918 213434
rect 290154 213198 296918 213434
rect 297154 213198 303918 213434
rect 304154 213198 310918 213434
rect 311154 213198 317918 213434
rect 318154 213198 324918 213434
rect 325154 213198 331918 213434
rect 332154 213198 338918 213434
rect 339154 213198 345918 213434
rect 346154 213198 352918 213434
rect 353154 213198 359918 213434
rect 360154 213198 366918 213434
rect 367154 213198 373918 213434
rect 374154 213198 380918 213434
rect 381154 213198 387918 213434
rect 388154 213198 394918 213434
rect 395154 213198 401918 213434
rect 402154 213198 408918 213434
rect 409154 213198 415918 213434
rect 416154 213198 422918 213434
rect 423154 213198 429918 213434
rect 430154 213198 436918 213434
rect 437154 213198 443918 213434
rect 444154 213198 450918 213434
rect 451154 213198 457918 213434
rect 458154 213198 464918 213434
rect 465154 213198 471918 213434
rect 472154 213198 478918 213434
rect 479154 213198 485918 213434
rect 486154 213198 492918 213434
rect 493154 213198 499918 213434
rect 500154 213198 506918 213434
rect 507154 213198 513918 213434
rect 514154 213198 520918 213434
rect 521154 213198 527918 213434
rect 528154 213198 534918 213434
rect 535154 213198 541918 213434
rect 542154 213198 548918 213434
rect 549154 213198 555918 213434
rect 556154 213198 562918 213434
rect 563154 213198 569918 213434
rect 570154 213198 576918 213434
rect 577154 213198 587570 213434
rect 587806 213198 587890 213434
rect 588126 213198 588210 213434
rect 588446 213198 588530 213434
rect 588766 213198 588874 213434
rect -4950 213156 588874 213198
rect -4950 212494 588874 212536
rect -4950 212258 -3090 212494
rect -2854 212258 -2770 212494
rect -2534 212258 -2450 212494
rect -2214 212258 -2130 212494
rect -1894 212258 1186 212494
rect 1422 212258 8186 212494
rect 8422 212258 15186 212494
rect 15422 212258 22186 212494
rect 22422 212258 29186 212494
rect 29422 212258 36186 212494
rect 36422 212258 43186 212494
rect 43422 212258 50186 212494
rect 50422 212258 57186 212494
rect 57422 212258 64186 212494
rect 64422 212258 71186 212494
rect 71422 212258 78186 212494
rect 78422 212258 85186 212494
rect 85422 212258 92186 212494
rect 92422 212258 99186 212494
rect 99422 212258 106186 212494
rect 106422 212258 113186 212494
rect 113422 212258 120186 212494
rect 120422 212258 127186 212494
rect 127422 212258 134186 212494
rect 134422 212258 141186 212494
rect 141422 212258 148186 212494
rect 148422 212258 155186 212494
rect 155422 212258 162186 212494
rect 162422 212258 169186 212494
rect 169422 212258 176186 212494
rect 176422 212258 183186 212494
rect 183422 212258 190186 212494
rect 190422 212258 197186 212494
rect 197422 212258 204186 212494
rect 204422 212258 211186 212494
rect 211422 212258 218186 212494
rect 218422 212258 225186 212494
rect 225422 212258 232186 212494
rect 232422 212258 239186 212494
rect 239422 212258 246186 212494
rect 246422 212258 253186 212494
rect 253422 212258 260186 212494
rect 260422 212258 267186 212494
rect 267422 212258 274186 212494
rect 274422 212258 281186 212494
rect 281422 212258 288186 212494
rect 288422 212258 295186 212494
rect 295422 212258 302186 212494
rect 302422 212258 309186 212494
rect 309422 212258 316186 212494
rect 316422 212258 323186 212494
rect 323422 212258 330186 212494
rect 330422 212258 337186 212494
rect 337422 212258 344186 212494
rect 344422 212258 351186 212494
rect 351422 212258 358186 212494
rect 358422 212258 365186 212494
rect 365422 212258 372186 212494
rect 372422 212258 379186 212494
rect 379422 212258 386186 212494
rect 386422 212258 393186 212494
rect 393422 212258 400186 212494
rect 400422 212258 407186 212494
rect 407422 212258 414186 212494
rect 414422 212258 421186 212494
rect 421422 212258 428186 212494
rect 428422 212258 435186 212494
rect 435422 212258 442186 212494
rect 442422 212258 449186 212494
rect 449422 212258 456186 212494
rect 456422 212258 463186 212494
rect 463422 212258 470186 212494
rect 470422 212258 477186 212494
rect 477422 212258 484186 212494
rect 484422 212258 491186 212494
rect 491422 212258 498186 212494
rect 498422 212258 505186 212494
rect 505422 212258 512186 212494
rect 512422 212258 519186 212494
rect 519422 212258 526186 212494
rect 526422 212258 533186 212494
rect 533422 212258 540186 212494
rect 540422 212258 547186 212494
rect 547422 212258 554186 212494
rect 554422 212258 561186 212494
rect 561422 212258 568186 212494
rect 568422 212258 575186 212494
rect 575422 212258 582186 212494
rect 582422 212258 585818 212494
rect 586054 212258 586138 212494
rect 586374 212258 586458 212494
rect 586694 212258 586778 212494
rect 587014 212258 588874 212494
rect -4950 212216 588874 212258
rect -4950 206434 588874 206476
rect -4950 206198 -4842 206434
rect -4606 206198 -4522 206434
rect -4286 206198 -4202 206434
rect -3966 206198 -3882 206434
rect -3646 206198 2918 206434
rect 3154 206198 9918 206434
rect 10154 206198 16918 206434
rect 17154 206198 23918 206434
rect 24154 206198 30918 206434
rect 31154 206198 37918 206434
rect 38154 206198 44918 206434
rect 45154 206198 51918 206434
rect 52154 206198 58918 206434
rect 59154 206198 65918 206434
rect 66154 206198 72918 206434
rect 73154 206198 79918 206434
rect 80154 206198 86918 206434
rect 87154 206198 93918 206434
rect 94154 206198 100918 206434
rect 101154 206198 107918 206434
rect 108154 206198 114918 206434
rect 115154 206198 121918 206434
rect 122154 206198 128918 206434
rect 129154 206198 135918 206434
rect 136154 206198 142918 206434
rect 143154 206198 149918 206434
rect 150154 206198 156918 206434
rect 157154 206198 163918 206434
rect 164154 206198 170918 206434
rect 171154 206198 177918 206434
rect 178154 206198 184918 206434
rect 185154 206198 191918 206434
rect 192154 206198 198918 206434
rect 199154 206198 205918 206434
rect 206154 206198 212918 206434
rect 213154 206198 219918 206434
rect 220154 206198 226918 206434
rect 227154 206198 233918 206434
rect 234154 206198 240918 206434
rect 241154 206198 247918 206434
rect 248154 206198 254918 206434
rect 255154 206198 261918 206434
rect 262154 206198 268918 206434
rect 269154 206198 275918 206434
rect 276154 206198 282918 206434
rect 283154 206198 289918 206434
rect 290154 206198 296918 206434
rect 297154 206198 303918 206434
rect 304154 206198 310918 206434
rect 311154 206198 317918 206434
rect 318154 206198 324918 206434
rect 325154 206198 331918 206434
rect 332154 206198 338918 206434
rect 339154 206198 345918 206434
rect 346154 206198 352918 206434
rect 353154 206198 359918 206434
rect 360154 206198 366918 206434
rect 367154 206198 373918 206434
rect 374154 206198 380918 206434
rect 381154 206198 387918 206434
rect 388154 206198 394918 206434
rect 395154 206198 401918 206434
rect 402154 206198 408918 206434
rect 409154 206198 415918 206434
rect 416154 206198 422918 206434
rect 423154 206198 429918 206434
rect 430154 206198 436918 206434
rect 437154 206198 443918 206434
rect 444154 206198 450918 206434
rect 451154 206198 457918 206434
rect 458154 206198 464918 206434
rect 465154 206198 471918 206434
rect 472154 206198 478918 206434
rect 479154 206198 485918 206434
rect 486154 206198 492918 206434
rect 493154 206198 499918 206434
rect 500154 206198 506918 206434
rect 507154 206198 513918 206434
rect 514154 206198 520918 206434
rect 521154 206198 527918 206434
rect 528154 206198 534918 206434
rect 535154 206198 541918 206434
rect 542154 206198 548918 206434
rect 549154 206198 555918 206434
rect 556154 206198 562918 206434
rect 563154 206198 569918 206434
rect 570154 206198 576918 206434
rect 577154 206198 587570 206434
rect 587806 206198 587890 206434
rect 588126 206198 588210 206434
rect 588446 206198 588530 206434
rect 588766 206198 588874 206434
rect -4950 206156 588874 206198
rect -4950 205494 588874 205536
rect -4950 205258 -3090 205494
rect -2854 205258 -2770 205494
rect -2534 205258 -2450 205494
rect -2214 205258 -2130 205494
rect -1894 205258 1186 205494
rect 1422 205258 8186 205494
rect 8422 205258 15186 205494
rect 15422 205258 22186 205494
rect 22422 205258 29186 205494
rect 29422 205258 36186 205494
rect 36422 205258 43186 205494
rect 43422 205258 50186 205494
rect 50422 205258 57186 205494
rect 57422 205258 64186 205494
rect 64422 205258 71186 205494
rect 71422 205258 78186 205494
rect 78422 205258 85186 205494
rect 85422 205258 92186 205494
rect 92422 205258 99186 205494
rect 99422 205258 106186 205494
rect 106422 205258 113186 205494
rect 113422 205258 120186 205494
rect 120422 205258 127186 205494
rect 127422 205258 134186 205494
rect 134422 205258 141186 205494
rect 141422 205258 148186 205494
rect 148422 205258 155186 205494
rect 155422 205258 162186 205494
rect 162422 205258 169186 205494
rect 169422 205258 176186 205494
rect 176422 205258 183186 205494
rect 183422 205258 190186 205494
rect 190422 205258 197186 205494
rect 197422 205258 204186 205494
rect 204422 205258 211186 205494
rect 211422 205258 218186 205494
rect 218422 205258 225186 205494
rect 225422 205258 232186 205494
rect 232422 205258 239186 205494
rect 239422 205258 246186 205494
rect 246422 205258 253186 205494
rect 253422 205258 260186 205494
rect 260422 205258 267186 205494
rect 267422 205258 274186 205494
rect 274422 205258 281186 205494
rect 281422 205258 288186 205494
rect 288422 205258 295186 205494
rect 295422 205258 302186 205494
rect 302422 205258 309186 205494
rect 309422 205258 316186 205494
rect 316422 205258 323186 205494
rect 323422 205258 330186 205494
rect 330422 205258 337186 205494
rect 337422 205258 344186 205494
rect 344422 205258 351186 205494
rect 351422 205258 358186 205494
rect 358422 205258 365186 205494
rect 365422 205258 372186 205494
rect 372422 205258 379186 205494
rect 379422 205258 386186 205494
rect 386422 205258 393186 205494
rect 393422 205258 400186 205494
rect 400422 205258 407186 205494
rect 407422 205258 414186 205494
rect 414422 205258 421186 205494
rect 421422 205258 428186 205494
rect 428422 205258 435186 205494
rect 435422 205258 442186 205494
rect 442422 205258 449186 205494
rect 449422 205258 456186 205494
rect 456422 205258 463186 205494
rect 463422 205258 470186 205494
rect 470422 205258 477186 205494
rect 477422 205258 484186 205494
rect 484422 205258 491186 205494
rect 491422 205258 498186 205494
rect 498422 205258 505186 205494
rect 505422 205258 512186 205494
rect 512422 205258 519186 205494
rect 519422 205258 526186 205494
rect 526422 205258 533186 205494
rect 533422 205258 540186 205494
rect 540422 205258 547186 205494
rect 547422 205258 554186 205494
rect 554422 205258 561186 205494
rect 561422 205258 568186 205494
rect 568422 205258 575186 205494
rect 575422 205258 582186 205494
rect 582422 205258 585818 205494
rect 586054 205258 586138 205494
rect 586374 205258 586458 205494
rect 586694 205258 586778 205494
rect 587014 205258 588874 205494
rect -4950 205216 588874 205258
rect -4950 199434 588874 199476
rect -4950 199198 -4842 199434
rect -4606 199198 -4522 199434
rect -4286 199198 -4202 199434
rect -3966 199198 -3882 199434
rect -3646 199198 2918 199434
rect 3154 199198 9918 199434
rect 10154 199198 16918 199434
rect 17154 199198 23918 199434
rect 24154 199198 30918 199434
rect 31154 199198 37918 199434
rect 38154 199198 44918 199434
rect 45154 199198 51918 199434
rect 52154 199198 58918 199434
rect 59154 199198 65918 199434
rect 66154 199198 72918 199434
rect 73154 199198 79918 199434
rect 80154 199198 86918 199434
rect 87154 199198 93918 199434
rect 94154 199198 100918 199434
rect 101154 199198 107918 199434
rect 108154 199198 114918 199434
rect 115154 199198 121918 199434
rect 122154 199198 128918 199434
rect 129154 199198 135918 199434
rect 136154 199198 142918 199434
rect 143154 199198 149918 199434
rect 150154 199198 156918 199434
rect 157154 199198 163918 199434
rect 164154 199198 170918 199434
rect 171154 199198 177918 199434
rect 178154 199198 184918 199434
rect 185154 199198 191918 199434
rect 192154 199198 198918 199434
rect 199154 199198 205918 199434
rect 206154 199198 212918 199434
rect 213154 199198 219918 199434
rect 220154 199198 226918 199434
rect 227154 199198 233918 199434
rect 234154 199198 240918 199434
rect 241154 199198 247918 199434
rect 248154 199198 254918 199434
rect 255154 199198 261918 199434
rect 262154 199198 268918 199434
rect 269154 199198 275918 199434
rect 276154 199198 282918 199434
rect 283154 199198 289918 199434
rect 290154 199198 310918 199434
rect 311154 199198 317918 199434
rect 318154 199198 324918 199434
rect 325154 199198 331918 199434
rect 332154 199198 338918 199434
rect 339154 199198 345918 199434
rect 346154 199198 352918 199434
rect 353154 199198 359918 199434
rect 360154 199198 366918 199434
rect 367154 199198 373918 199434
rect 374154 199198 380918 199434
rect 381154 199198 387918 199434
rect 388154 199198 394918 199434
rect 395154 199198 401918 199434
rect 402154 199198 408918 199434
rect 409154 199198 415918 199434
rect 416154 199198 422918 199434
rect 423154 199198 429918 199434
rect 430154 199198 436918 199434
rect 437154 199198 443918 199434
rect 444154 199198 450918 199434
rect 451154 199198 457918 199434
rect 458154 199198 464918 199434
rect 465154 199198 471918 199434
rect 472154 199198 478918 199434
rect 479154 199198 485918 199434
rect 486154 199198 492918 199434
rect 493154 199198 499918 199434
rect 500154 199198 506918 199434
rect 507154 199198 513918 199434
rect 514154 199198 520918 199434
rect 521154 199198 527918 199434
rect 528154 199198 534918 199434
rect 535154 199198 541918 199434
rect 542154 199198 548918 199434
rect 549154 199198 555918 199434
rect 556154 199198 562918 199434
rect 563154 199198 569918 199434
rect 570154 199198 576918 199434
rect 577154 199198 587570 199434
rect 587806 199198 587890 199434
rect 588126 199198 588210 199434
rect 588446 199198 588530 199434
rect 588766 199198 588874 199434
rect -4950 199156 588874 199198
rect -4950 198494 588874 198536
rect -4950 198258 -3090 198494
rect -2854 198258 -2770 198494
rect -2534 198258 -2450 198494
rect -2214 198258 -2130 198494
rect -1894 198258 1186 198494
rect 1422 198258 8186 198494
rect 8422 198258 15186 198494
rect 15422 198258 22186 198494
rect 22422 198258 29186 198494
rect 29422 198258 36186 198494
rect 36422 198258 43186 198494
rect 43422 198258 50186 198494
rect 50422 198258 57186 198494
rect 57422 198258 64186 198494
rect 64422 198258 71186 198494
rect 71422 198258 78186 198494
rect 78422 198258 85186 198494
rect 85422 198258 92186 198494
rect 92422 198258 99186 198494
rect 99422 198258 106186 198494
rect 106422 198258 113186 198494
rect 113422 198258 120186 198494
rect 120422 198258 127186 198494
rect 127422 198258 134186 198494
rect 134422 198258 141186 198494
rect 141422 198258 148186 198494
rect 148422 198258 155186 198494
rect 155422 198258 162186 198494
rect 162422 198258 169186 198494
rect 169422 198258 176186 198494
rect 176422 198258 183186 198494
rect 183422 198258 190186 198494
rect 190422 198258 197186 198494
rect 197422 198258 204186 198494
rect 204422 198258 211186 198494
rect 211422 198258 218186 198494
rect 218422 198258 225186 198494
rect 225422 198258 232186 198494
rect 232422 198258 239186 198494
rect 239422 198258 246186 198494
rect 246422 198258 253186 198494
rect 253422 198258 260186 198494
rect 260422 198258 267186 198494
rect 267422 198258 274186 198494
rect 274422 198258 281186 198494
rect 281422 198258 288186 198494
rect 288422 198258 309186 198494
rect 309422 198258 316186 198494
rect 316422 198258 323186 198494
rect 323422 198258 330186 198494
rect 330422 198258 337186 198494
rect 337422 198258 344186 198494
rect 344422 198258 351186 198494
rect 351422 198258 358186 198494
rect 358422 198258 365186 198494
rect 365422 198258 372186 198494
rect 372422 198258 379186 198494
rect 379422 198258 386186 198494
rect 386422 198258 393186 198494
rect 393422 198258 400186 198494
rect 400422 198258 407186 198494
rect 407422 198258 414186 198494
rect 414422 198258 421186 198494
rect 421422 198258 428186 198494
rect 428422 198258 435186 198494
rect 435422 198258 442186 198494
rect 442422 198258 449186 198494
rect 449422 198258 456186 198494
rect 456422 198258 463186 198494
rect 463422 198258 470186 198494
rect 470422 198258 477186 198494
rect 477422 198258 484186 198494
rect 484422 198258 491186 198494
rect 491422 198258 498186 198494
rect 498422 198258 505186 198494
rect 505422 198258 512186 198494
rect 512422 198258 519186 198494
rect 519422 198258 526186 198494
rect 526422 198258 533186 198494
rect 533422 198258 540186 198494
rect 540422 198258 547186 198494
rect 547422 198258 554186 198494
rect 554422 198258 561186 198494
rect 561422 198258 568186 198494
rect 568422 198258 575186 198494
rect 575422 198258 582186 198494
rect 582422 198258 585818 198494
rect 586054 198258 586138 198494
rect 586374 198258 586458 198494
rect 586694 198258 586778 198494
rect 587014 198258 588874 198494
rect -4950 198216 588874 198258
rect -4950 192434 588874 192476
rect -4950 192198 -4842 192434
rect -4606 192198 -4522 192434
rect -4286 192198 -4202 192434
rect -3966 192198 -3882 192434
rect -3646 192198 2918 192434
rect 3154 192198 9918 192434
rect 10154 192198 16918 192434
rect 17154 192198 23918 192434
rect 24154 192198 30918 192434
rect 31154 192198 37918 192434
rect 38154 192198 44918 192434
rect 45154 192198 51918 192434
rect 52154 192198 58918 192434
rect 59154 192198 65918 192434
rect 66154 192198 72918 192434
rect 73154 192198 79918 192434
rect 80154 192198 86918 192434
rect 87154 192198 93918 192434
rect 94154 192198 100918 192434
rect 101154 192198 107918 192434
rect 108154 192198 114918 192434
rect 115154 192198 121918 192434
rect 122154 192198 128918 192434
rect 129154 192198 135918 192434
rect 136154 192198 142918 192434
rect 143154 192198 149918 192434
rect 150154 192198 156918 192434
rect 157154 192198 163918 192434
rect 164154 192198 170918 192434
rect 171154 192198 177918 192434
rect 178154 192198 184918 192434
rect 185154 192198 191918 192434
rect 192154 192198 198918 192434
rect 199154 192198 205918 192434
rect 206154 192198 212918 192434
rect 213154 192198 219918 192434
rect 220154 192198 226918 192434
rect 227154 192198 233918 192434
rect 234154 192198 240918 192434
rect 241154 192198 247918 192434
rect 248154 192198 254918 192434
rect 255154 192198 261918 192434
rect 262154 192198 268918 192434
rect 269154 192198 275918 192434
rect 276154 192198 282918 192434
rect 283154 192198 289918 192434
rect 290154 192198 296918 192434
rect 297154 192198 303918 192434
rect 304154 192198 310918 192434
rect 311154 192198 317918 192434
rect 318154 192198 324918 192434
rect 325154 192198 331918 192434
rect 332154 192198 338918 192434
rect 339154 192198 345918 192434
rect 346154 192198 352918 192434
rect 353154 192198 359918 192434
rect 360154 192198 366918 192434
rect 367154 192198 373918 192434
rect 374154 192198 380918 192434
rect 381154 192198 387918 192434
rect 388154 192198 394918 192434
rect 395154 192198 401918 192434
rect 402154 192198 408918 192434
rect 409154 192198 415918 192434
rect 416154 192198 422918 192434
rect 423154 192198 429918 192434
rect 430154 192198 436918 192434
rect 437154 192198 443918 192434
rect 444154 192198 450918 192434
rect 451154 192198 457918 192434
rect 458154 192198 464918 192434
rect 465154 192198 471918 192434
rect 472154 192198 478918 192434
rect 479154 192198 485918 192434
rect 486154 192198 492918 192434
rect 493154 192198 499918 192434
rect 500154 192198 506918 192434
rect 507154 192198 513918 192434
rect 514154 192198 520918 192434
rect 521154 192198 527918 192434
rect 528154 192198 534918 192434
rect 535154 192198 541918 192434
rect 542154 192198 548918 192434
rect 549154 192198 555918 192434
rect 556154 192198 562918 192434
rect 563154 192198 569918 192434
rect 570154 192198 576918 192434
rect 577154 192198 587570 192434
rect 587806 192198 587890 192434
rect 588126 192198 588210 192434
rect 588446 192198 588530 192434
rect 588766 192198 588874 192434
rect -4950 192156 588874 192198
rect -4950 191494 588874 191536
rect -4950 191258 -3090 191494
rect -2854 191258 -2770 191494
rect -2534 191258 -2450 191494
rect -2214 191258 -2130 191494
rect -1894 191258 1186 191494
rect 1422 191258 8186 191494
rect 8422 191258 15186 191494
rect 15422 191258 22186 191494
rect 22422 191258 29186 191494
rect 29422 191258 36186 191494
rect 36422 191258 43186 191494
rect 43422 191258 50186 191494
rect 50422 191258 57186 191494
rect 57422 191258 64186 191494
rect 64422 191258 71186 191494
rect 71422 191258 78186 191494
rect 78422 191258 85186 191494
rect 85422 191258 92186 191494
rect 92422 191258 99186 191494
rect 99422 191258 106186 191494
rect 106422 191258 113186 191494
rect 113422 191258 120186 191494
rect 120422 191258 127186 191494
rect 127422 191258 134186 191494
rect 134422 191258 141186 191494
rect 141422 191258 148186 191494
rect 148422 191258 155186 191494
rect 155422 191258 162186 191494
rect 162422 191258 169186 191494
rect 169422 191258 176186 191494
rect 176422 191258 183186 191494
rect 183422 191258 190186 191494
rect 190422 191258 197186 191494
rect 197422 191258 204186 191494
rect 204422 191258 211186 191494
rect 211422 191258 218186 191494
rect 218422 191258 225186 191494
rect 225422 191258 232186 191494
rect 232422 191258 239186 191494
rect 239422 191258 246186 191494
rect 246422 191258 253186 191494
rect 253422 191258 260186 191494
rect 260422 191258 267186 191494
rect 267422 191258 274186 191494
rect 274422 191258 281186 191494
rect 281422 191258 288186 191494
rect 288422 191258 295186 191494
rect 295422 191258 302186 191494
rect 302422 191258 309186 191494
rect 309422 191258 316186 191494
rect 316422 191258 323186 191494
rect 323422 191258 330186 191494
rect 330422 191258 337186 191494
rect 337422 191258 344186 191494
rect 344422 191258 351186 191494
rect 351422 191258 358186 191494
rect 358422 191258 365186 191494
rect 365422 191258 372186 191494
rect 372422 191258 379186 191494
rect 379422 191258 386186 191494
rect 386422 191258 393186 191494
rect 393422 191258 400186 191494
rect 400422 191258 407186 191494
rect 407422 191258 414186 191494
rect 414422 191258 421186 191494
rect 421422 191258 428186 191494
rect 428422 191258 435186 191494
rect 435422 191258 442186 191494
rect 442422 191258 449186 191494
rect 449422 191258 456186 191494
rect 456422 191258 463186 191494
rect 463422 191258 470186 191494
rect 470422 191258 477186 191494
rect 477422 191258 484186 191494
rect 484422 191258 491186 191494
rect 491422 191258 498186 191494
rect 498422 191258 505186 191494
rect 505422 191258 512186 191494
rect 512422 191258 519186 191494
rect 519422 191258 526186 191494
rect 526422 191258 533186 191494
rect 533422 191258 540186 191494
rect 540422 191258 547186 191494
rect 547422 191258 554186 191494
rect 554422 191258 561186 191494
rect 561422 191258 568186 191494
rect 568422 191258 575186 191494
rect 575422 191258 582186 191494
rect 582422 191258 585818 191494
rect 586054 191258 586138 191494
rect 586374 191258 586458 191494
rect 586694 191258 586778 191494
rect 587014 191258 588874 191494
rect -4950 191216 588874 191258
rect -4950 185434 588874 185476
rect -4950 185198 -4842 185434
rect -4606 185198 -4522 185434
rect -4286 185198 -4202 185434
rect -3966 185198 -3882 185434
rect -3646 185198 2918 185434
rect 3154 185198 9918 185434
rect 10154 185198 16918 185434
rect 17154 185198 23918 185434
rect 24154 185198 30918 185434
rect 31154 185198 37918 185434
rect 38154 185198 44918 185434
rect 45154 185198 51918 185434
rect 52154 185198 58918 185434
rect 59154 185198 65918 185434
rect 66154 185198 72918 185434
rect 73154 185198 79918 185434
rect 80154 185198 86918 185434
rect 87154 185198 93918 185434
rect 94154 185198 100918 185434
rect 101154 185198 107918 185434
rect 108154 185198 114918 185434
rect 115154 185198 121918 185434
rect 122154 185198 128918 185434
rect 129154 185198 135918 185434
rect 136154 185198 142918 185434
rect 143154 185198 149918 185434
rect 150154 185198 156918 185434
rect 157154 185198 163918 185434
rect 164154 185198 170918 185434
rect 171154 185198 177918 185434
rect 178154 185198 184918 185434
rect 185154 185198 191918 185434
rect 192154 185198 198918 185434
rect 199154 185198 205918 185434
rect 206154 185198 212918 185434
rect 213154 185198 219918 185434
rect 220154 185198 226918 185434
rect 227154 185198 233918 185434
rect 234154 185198 240918 185434
rect 241154 185198 247918 185434
rect 248154 185198 254918 185434
rect 255154 185198 261918 185434
rect 262154 185198 268918 185434
rect 269154 185198 275918 185434
rect 276154 185198 282918 185434
rect 283154 185198 289918 185434
rect 290154 185198 296918 185434
rect 297154 185198 303918 185434
rect 304154 185198 310918 185434
rect 311154 185198 317918 185434
rect 318154 185198 324918 185434
rect 325154 185198 331918 185434
rect 332154 185198 338918 185434
rect 339154 185198 345918 185434
rect 346154 185198 352918 185434
rect 353154 185198 359918 185434
rect 360154 185198 366918 185434
rect 367154 185198 373918 185434
rect 374154 185198 380918 185434
rect 381154 185198 387918 185434
rect 388154 185198 394918 185434
rect 395154 185198 401918 185434
rect 402154 185198 408918 185434
rect 409154 185198 415918 185434
rect 416154 185198 422918 185434
rect 423154 185198 429918 185434
rect 430154 185198 436918 185434
rect 437154 185198 443918 185434
rect 444154 185198 450918 185434
rect 451154 185198 457918 185434
rect 458154 185198 464918 185434
rect 465154 185198 471918 185434
rect 472154 185198 478918 185434
rect 479154 185198 485918 185434
rect 486154 185198 492918 185434
rect 493154 185198 499918 185434
rect 500154 185198 506918 185434
rect 507154 185198 513918 185434
rect 514154 185198 520918 185434
rect 521154 185198 527918 185434
rect 528154 185198 534918 185434
rect 535154 185198 541918 185434
rect 542154 185198 548918 185434
rect 549154 185198 555918 185434
rect 556154 185198 562918 185434
rect 563154 185198 569918 185434
rect 570154 185198 576918 185434
rect 577154 185198 587570 185434
rect 587806 185198 587890 185434
rect 588126 185198 588210 185434
rect 588446 185198 588530 185434
rect 588766 185198 588874 185434
rect -4950 185156 588874 185198
rect -4950 184494 588874 184536
rect -4950 184258 -3090 184494
rect -2854 184258 -2770 184494
rect -2534 184258 -2450 184494
rect -2214 184258 -2130 184494
rect -1894 184258 1186 184494
rect 1422 184258 8186 184494
rect 8422 184258 15186 184494
rect 15422 184258 22186 184494
rect 22422 184258 29186 184494
rect 29422 184258 36186 184494
rect 36422 184258 43186 184494
rect 43422 184258 50186 184494
rect 50422 184258 57186 184494
rect 57422 184258 64186 184494
rect 64422 184258 71186 184494
rect 71422 184258 78186 184494
rect 78422 184258 85186 184494
rect 85422 184258 92186 184494
rect 92422 184258 99186 184494
rect 99422 184258 106186 184494
rect 106422 184258 113186 184494
rect 113422 184258 120186 184494
rect 120422 184258 127186 184494
rect 127422 184258 134186 184494
rect 134422 184258 141186 184494
rect 141422 184258 148186 184494
rect 148422 184258 155186 184494
rect 155422 184258 162186 184494
rect 162422 184258 169186 184494
rect 169422 184258 176186 184494
rect 176422 184258 183186 184494
rect 183422 184258 190186 184494
rect 190422 184258 197186 184494
rect 197422 184258 204186 184494
rect 204422 184258 211186 184494
rect 211422 184258 218186 184494
rect 218422 184258 225186 184494
rect 225422 184258 232186 184494
rect 232422 184258 239186 184494
rect 239422 184258 246186 184494
rect 246422 184258 253186 184494
rect 253422 184258 260186 184494
rect 260422 184258 267186 184494
rect 267422 184258 274186 184494
rect 274422 184258 281186 184494
rect 281422 184258 288186 184494
rect 288422 184258 295186 184494
rect 295422 184258 302186 184494
rect 302422 184258 309186 184494
rect 309422 184258 316186 184494
rect 316422 184258 323186 184494
rect 323422 184258 330186 184494
rect 330422 184258 337186 184494
rect 337422 184258 344186 184494
rect 344422 184258 351186 184494
rect 351422 184258 358186 184494
rect 358422 184258 365186 184494
rect 365422 184258 372186 184494
rect 372422 184258 379186 184494
rect 379422 184258 386186 184494
rect 386422 184258 393186 184494
rect 393422 184258 400186 184494
rect 400422 184258 407186 184494
rect 407422 184258 414186 184494
rect 414422 184258 421186 184494
rect 421422 184258 428186 184494
rect 428422 184258 435186 184494
rect 435422 184258 442186 184494
rect 442422 184258 449186 184494
rect 449422 184258 456186 184494
rect 456422 184258 463186 184494
rect 463422 184258 470186 184494
rect 470422 184258 477186 184494
rect 477422 184258 484186 184494
rect 484422 184258 491186 184494
rect 491422 184258 498186 184494
rect 498422 184258 505186 184494
rect 505422 184258 512186 184494
rect 512422 184258 519186 184494
rect 519422 184258 526186 184494
rect 526422 184258 533186 184494
rect 533422 184258 540186 184494
rect 540422 184258 547186 184494
rect 547422 184258 554186 184494
rect 554422 184258 561186 184494
rect 561422 184258 568186 184494
rect 568422 184258 575186 184494
rect 575422 184258 582186 184494
rect 582422 184258 585818 184494
rect 586054 184258 586138 184494
rect 586374 184258 586458 184494
rect 586694 184258 586778 184494
rect 587014 184258 588874 184494
rect -4950 184216 588874 184258
rect -4950 178434 588874 178476
rect -4950 178198 -4842 178434
rect -4606 178198 -4522 178434
rect -4286 178198 -4202 178434
rect -3966 178198 -3882 178434
rect -3646 178198 2918 178434
rect 3154 178198 9918 178434
rect 10154 178198 16918 178434
rect 17154 178198 23918 178434
rect 24154 178198 30918 178434
rect 31154 178198 37918 178434
rect 38154 178198 44918 178434
rect 45154 178198 51918 178434
rect 52154 178198 58918 178434
rect 59154 178198 65918 178434
rect 66154 178198 72918 178434
rect 73154 178198 79918 178434
rect 80154 178198 86918 178434
rect 87154 178198 93918 178434
rect 94154 178198 100918 178434
rect 101154 178198 107918 178434
rect 108154 178198 114918 178434
rect 115154 178198 121918 178434
rect 122154 178198 128918 178434
rect 129154 178198 135918 178434
rect 136154 178198 142918 178434
rect 143154 178198 149918 178434
rect 150154 178198 156918 178434
rect 157154 178198 163918 178434
rect 164154 178198 170918 178434
rect 171154 178198 177918 178434
rect 178154 178198 184918 178434
rect 185154 178198 191918 178434
rect 192154 178198 198918 178434
rect 199154 178198 205918 178434
rect 206154 178198 212918 178434
rect 213154 178198 219918 178434
rect 220154 178198 226918 178434
rect 227154 178198 233918 178434
rect 234154 178198 240918 178434
rect 241154 178198 247918 178434
rect 248154 178198 254918 178434
rect 255154 178198 261918 178434
rect 262154 178198 268918 178434
rect 269154 178198 275918 178434
rect 276154 178198 282918 178434
rect 283154 178198 289918 178434
rect 290154 178198 296918 178434
rect 297154 178198 303918 178434
rect 304154 178198 310918 178434
rect 311154 178198 317918 178434
rect 318154 178198 324918 178434
rect 325154 178198 331918 178434
rect 332154 178198 338918 178434
rect 339154 178198 345918 178434
rect 346154 178198 352918 178434
rect 353154 178198 359918 178434
rect 360154 178198 366918 178434
rect 367154 178198 373918 178434
rect 374154 178198 380918 178434
rect 381154 178198 387918 178434
rect 388154 178198 394918 178434
rect 395154 178198 401918 178434
rect 402154 178198 408918 178434
rect 409154 178198 415918 178434
rect 416154 178198 422918 178434
rect 423154 178198 429918 178434
rect 430154 178198 436918 178434
rect 437154 178198 443918 178434
rect 444154 178198 450918 178434
rect 451154 178198 457918 178434
rect 458154 178198 464918 178434
rect 465154 178198 471918 178434
rect 472154 178198 478918 178434
rect 479154 178198 485918 178434
rect 486154 178198 492918 178434
rect 493154 178198 499918 178434
rect 500154 178198 506918 178434
rect 507154 178198 513918 178434
rect 514154 178198 520918 178434
rect 521154 178198 527918 178434
rect 528154 178198 534918 178434
rect 535154 178198 541918 178434
rect 542154 178198 548918 178434
rect 549154 178198 555918 178434
rect 556154 178198 562918 178434
rect 563154 178198 569918 178434
rect 570154 178198 576918 178434
rect 577154 178198 587570 178434
rect 587806 178198 587890 178434
rect 588126 178198 588210 178434
rect 588446 178198 588530 178434
rect 588766 178198 588874 178434
rect -4950 178156 588874 178198
rect -4950 177494 588874 177536
rect -4950 177258 -3090 177494
rect -2854 177258 -2770 177494
rect -2534 177258 -2450 177494
rect -2214 177258 -2130 177494
rect -1894 177258 1186 177494
rect 1422 177258 8186 177494
rect 8422 177258 15186 177494
rect 15422 177258 22186 177494
rect 22422 177258 29186 177494
rect 29422 177258 36186 177494
rect 36422 177258 43186 177494
rect 43422 177258 50186 177494
rect 50422 177258 57186 177494
rect 57422 177258 64186 177494
rect 64422 177258 71186 177494
rect 71422 177258 78186 177494
rect 78422 177258 85186 177494
rect 85422 177258 92186 177494
rect 92422 177258 99186 177494
rect 99422 177258 106186 177494
rect 106422 177258 113186 177494
rect 113422 177258 120186 177494
rect 120422 177258 127186 177494
rect 127422 177258 134186 177494
rect 134422 177258 141186 177494
rect 141422 177258 148186 177494
rect 148422 177258 155186 177494
rect 155422 177258 162186 177494
rect 162422 177258 169186 177494
rect 169422 177258 176186 177494
rect 176422 177258 183186 177494
rect 183422 177258 190186 177494
rect 190422 177258 197186 177494
rect 197422 177258 204186 177494
rect 204422 177258 211186 177494
rect 211422 177258 218186 177494
rect 218422 177258 225186 177494
rect 225422 177258 232186 177494
rect 232422 177258 239186 177494
rect 239422 177258 246186 177494
rect 246422 177258 253186 177494
rect 253422 177258 260186 177494
rect 260422 177258 267186 177494
rect 267422 177258 274186 177494
rect 274422 177258 281186 177494
rect 281422 177258 288186 177494
rect 288422 177258 295186 177494
rect 295422 177258 302186 177494
rect 302422 177258 309186 177494
rect 309422 177258 316186 177494
rect 316422 177258 323186 177494
rect 323422 177258 330186 177494
rect 330422 177258 337186 177494
rect 337422 177258 344186 177494
rect 344422 177258 351186 177494
rect 351422 177258 358186 177494
rect 358422 177258 365186 177494
rect 365422 177258 372186 177494
rect 372422 177258 379186 177494
rect 379422 177258 386186 177494
rect 386422 177258 393186 177494
rect 393422 177258 400186 177494
rect 400422 177258 407186 177494
rect 407422 177258 414186 177494
rect 414422 177258 421186 177494
rect 421422 177258 428186 177494
rect 428422 177258 435186 177494
rect 435422 177258 442186 177494
rect 442422 177258 449186 177494
rect 449422 177258 456186 177494
rect 456422 177258 463186 177494
rect 463422 177258 470186 177494
rect 470422 177258 477186 177494
rect 477422 177258 484186 177494
rect 484422 177258 491186 177494
rect 491422 177258 498186 177494
rect 498422 177258 505186 177494
rect 505422 177258 512186 177494
rect 512422 177258 519186 177494
rect 519422 177258 526186 177494
rect 526422 177258 533186 177494
rect 533422 177258 540186 177494
rect 540422 177258 547186 177494
rect 547422 177258 554186 177494
rect 554422 177258 561186 177494
rect 561422 177258 568186 177494
rect 568422 177258 575186 177494
rect 575422 177258 582186 177494
rect 582422 177258 585818 177494
rect 586054 177258 586138 177494
rect 586374 177258 586458 177494
rect 586694 177258 586778 177494
rect 587014 177258 588874 177494
rect -4950 177216 588874 177258
rect -4950 171434 588874 171476
rect -4950 171198 -4842 171434
rect -4606 171198 -4522 171434
rect -4286 171198 -4202 171434
rect -3966 171198 -3882 171434
rect -3646 171198 2918 171434
rect 3154 171198 9918 171434
rect 10154 171198 16918 171434
rect 17154 171198 23918 171434
rect 24154 171198 30918 171434
rect 31154 171198 37918 171434
rect 38154 171198 44918 171434
rect 45154 171198 51918 171434
rect 52154 171198 58918 171434
rect 59154 171198 65918 171434
rect 66154 171198 72918 171434
rect 73154 171198 79918 171434
rect 80154 171198 86918 171434
rect 87154 171198 93918 171434
rect 94154 171198 100918 171434
rect 101154 171198 107918 171434
rect 108154 171198 114918 171434
rect 115154 171198 121918 171434
rect 122154 171198 128918 171434
rect 129154 171198 135918 171434
rect 136154 171198 142918 171434
rect 143154 171198 149918 171434
rect 150154 171198 156918 171434
rect 157154 171198 163918 171434
rect 164154 171198 170918 171434
rect 171154 171198 177918 171434
rect 178154 171198 184918 171434
rect 185154 171198 191918 171434
rect 192154 171198 198918 171434
rect 199154 171198 205918 171434
rect 206154 171198 212918 171434
rect 213154 171198 219918 171434
rect 220154 171198 226918 171434
rect 227154 171198 233918 171434
rect 234154 171198 240918 171434
rect 241154 171198 247918 171434
rect 248154 171198 254918 171434
rect 255154 171198 261918 171434
rect 262154 171198 268918 171434
rect 269154 171198 275918 171434
rect 276154 171198 282918 171434
rect 283154 171198 289918 171434
rect 290154 171198 296918 171434
rect 297154 171198 303918 171434
rect 304154 171198 310918 171434
rect 311154 171198 317918 171434
rect 318154 171198 324918 171434
rect 325154 171198 331918 171434
rect 332154 171198 338918 171434
rect 339154 171198 345918 171434
rect 346154 171198 352918 171434
rect 353154 171198 359918 171434
rect 360154 171198 366918 171434
rect 367154 171198 373918 171434
rect 374154 171198 380918 171434
rect 381154 171198 387918 171434
rect 388154 171198 394918 171434
rect 395154 171198 401918 171434
rect 402154 171198 408918 171434
rect 409154 171198 415918 171434
rect 416154 171198 422918 171434
rect 423154 171198 429918 171434
rect 430154 171198 436918 171434
rect 437154 171198 443918 171434
rect 444154 171198 450918 171434
rect 451154 171198 457918 171434
rect 458154 171198 464918 171434
rect 465154 171198 471918 171434
rect 472154 171198 478918 171434
rect 479154 171198 485918 171434
rect 486154 171198 492918 171434
rect 493154 171198 499918 171434
rect 500154 171198 506918 171434
rect 507154 171198 513918 171434
rect 514154 171198 520918 171434
rect 521154 171198 527918 171434
rect 528154 171198 534918 171434
rect 535154 171198 541918 171434
rect 542154 171198 548918 171434
rect 549154 171198 555918 171434
rect 556154 171198 562918 171434
rect 563154 171198 569918 171434
rect 570154 171198 576918 171434
rect 577154 171198 587570 171434
rect 587806 171198 587890 171434
rect 588126 171198 588210 171434
rect 588446 171198 588530 171434
rect 588766 171198 588874 171434
rect -4950 171156 588874 171198
rect -4950 170494 588874 170536
rect -4950 170258 -3090 170494
rect -2854 170258 -2770 170494
rect -2534 170258 -2450 170494
rect -2214 170258 -2130 170494
rect -1894 170258 1186 170494
rect 1422 170258 8186 170494
rect 8422 170258 15186 170494
rect 15422 170258 22186 170494
rect 22422 170258 29186 170494
rect 29422 170258 36186 170494
rect 36422 170258 43186 170494
rect 43422 170258 50186 170494
rect 50422 170258 57186 170494
rect 57422 170258 64186 170494
rect 64422 170258 71186 170494
rect 71422 170258 78186 170494
rect 78422 170258 85186 170494
rect 85422 170258 92186 170494
rect 92422 170258 99186 170494
rect 99422 170258 106186 170494
rect 106422 170258 113186 170494
rect 113422 170258 120186 170494
rect 120422 170258 127186 170494
rect 127422 170258 134186 170494
rect 134422 170258 141186 170494
rect 141422 170258 148186 170494
rect 148422 170258 155186 170494
rect 155422 170258 162186 170494
rect 162422 170258 169186 170494
rect 169422 170258 176186 170494
rect 176422 170258 183186 170494
rect 183422 170258 190186 170494
rect 190422 170258 197186 170494
rect 197422 170258 204186 170494
rect 204422 170258 211186 170494
rect 211422 170258 218186 170494
rect 218422 170258 225186 170494
rect 225422 170258 232186 170494
rect 232422 170258 239186 170494
rect 239422 170258 246186 170494
rect 246422 170258 253186 170494
rect 253422 170258 260186 170494
rect 260422 170258 267186 170494
rect 267422 170258 274186 170494
rect 274422 170258 281186 170494
rect 281422 170258 288186 170494
rect 288422 170258 295186 170494
rect 295422 170258 302186 170494
rect 302422 170258 309186 170494
rect 309422 170258 316186 170494
rect 316422 170258 323186 170494
rect 323422 170258 330186 170494
rect 330422 170258 337186 170494
rect 337422 170258 344186 170494
rect 344422 170258 351186 170494
rect 351422 170258 358186 170494
rect 358422 170258 365186 170494
rect 365422 170258 372186 170494
rect 372422 170258 379186 170494
rect 379422 170258 386186 170494
rect 386422 170258 393186 170494
rect 393422 170258 400186 170494
rect 400422 170258 407186 170494
rect 407422 170258 414186 170494
rect 414422 170258 421186 170494
rect 421422 170258 428186 170494
rect 428422 170258 435186 170494
rect 435422 170258 442186 170494
rect 442422 170258 449186 170494
rect 449422 170258 456186 170494
rect 456422 170258 463186 170494
rect 463422 170258 470186 170494
rect 470422 170258 477186 170494
rect 477422 170258 484186 170494
rect 484422 170258 491186 170494
rect 491422 170258 498186 170494
rect 498422 170258 505186 170494
rect 505422 170258 512186 170494
rect 512422 170258 519186 170494
rect 519422 170258 526186 170494
rect 526422 170258 533186 170494
rect 533422 170258 540186 170494
rect 540422 170258 547186 170494
rect 547422 170258 554186 170494
rect 554422 170258 561186 170494
rect 561422 170258 568186 170494
rect 568422 170258 575186 170494
rect 575422 170258 582186 170494
rect 582422 170258 585818 170494
rect 586054 170258 586138 170494
rect 586374 170258 586458 170494
rect 586694 170258 586778 170494
rect 587014 170258 588874 170494
rect -4950 170216 588874 170258
rect -4950 164434 588874 164476
rect -4950 164198 -4842 164434
rect -4606 164198 -4522 164434
rect -4286 164198 -4202 164434
rect -3966 164198 -3882 164434
rect -3646 164198 2918 164434
rect 3154 164198 9918 164434
rect 10154 164198 16918 164434
rect 17154 164198 23918 164434
rect 24154 164198 30918 164434
rect 31154 164198 37918 164434
rect 38154 164198 44918 164434
rect 45154 164198 51918 164434
rect 52154 164198 58918 164434
rect 59154 164198 65918 164434
rect 66154 164198 72918 164434
rect 73154 164198 79918 164434
rect 80154 164198 86918 164434
rect 87154 164198 93918 164434
rect 94154 164198 100918 164434
rect 101154 164198 107918 164434
rect 108154 164198 114918 164434
rect 115154 164198 121918 164434
rect 122154 164198 128918 164434
rect 129154 164198 135918 164434
rect 136154 164198 142918 164434
rect 143154 164198 149918 164434
rect 150154 164198 156918 164434
rect 157154 164198 163918 164434
rect 164154 164198 170918 164434
rect 171154 164198 177918 164434
rect 178154 164198 184918 164434
rect 185154 164198 191918 164434
rect 192154 164198 198918 164434
rect 199154 164198 205918 164434
rect 206154 164198 212918 164434
rect 213154 164198 219918 164434
rect 220154 164198 226918 164434
rect 227154 164198 233918 164434
rect 234154 164198 240918 164434
rect 241154 164198 247918 164434
rect 248154 164198 254918 164434
rect 255154 164198 261918 164434
rect 262154 164198 268918 164434
rect 269154 164198 275918 164434
rect 276154 164198 282918 164434
rect 283154 164198 289918 164434
rect 290154 164198 296918 164434
rect 297154 164198 303918 164434
rect 304154 164198 310918 164434
rect 311154 164198 317918 164434
rect 318154 164198 324918 164434
rect 325154 164198 331918 164434
rect 332154 164198 338918 164434
rect 339154 164198 345918 164434
rect 346154 164198 352918 164434
rect 353154 164198 359918 164434
rect 360154 164198 366918 164434
rect 367154 164198 373918 164434
rect 374154 164198 380918 164434
rect 381154 164198 387918 164434
rect 388154 164198 394918 164434
rect 395154 164198 401918 164434
rect 402154 164198 408918 164434
rect 409154 164198 415918 164434
rect 416154 164198 422918 164434
rect 423154 164198 429918 164434
rect 430154 164198 436918 164434
rect 437154 164198 443918 164434
rect 444154 164198 450918 164434
rect 451154 164198 457918 164434
rect 458154 164198 464918 164434
rect 465154 164198 471918 164434
rect 472154 164198 478918 164434
rect 479154 164198 485918 164434
rect 486154 164198 492918 164434
rect 493154 164198 499918 164434
rect 500154 164198 506918 164434
rect 507154 164198 513918 164434
rect 514154 164198 520918 164434
rect 521154 164198 527918 164434
rect 528154 164198 534918 164434
rect 535154 164198 541918 164434
rect 542154 164198 548918 164434
rect 549154 164198 555918 164434
rect 556154 164198 562918 164434
rect 563154 164198 569918 164434
rect 570154 164198 576918 164434
rect 577154 164198 587570 164434
rect 587806 164198 587890 164434
rect 588126 164198 588210 164434
rect 588446 164198 588530 164434
rect 588766 164198 588874 164434
rect -4950 164156 588874 164198
rect -4950 163494 588874 163536
rect -4950 163258 -3090 163494
rect -2854 163258 -2770 163494
rect -2534 163258 -2450 163494
rect -2214 163258 -2130 163494
rect -1894 163258 1186 163494
rect 1422 163258 8186 163494
rect 8422 163258 15186 163494
rect 15422 163258 22186 163494
rect 22422 163258 29186 163494
rect 29422 163258 36186 163494
rect 36422 163258 43186 163494
rect 43422 163258 50186 163494
rect 50422 163258 57186 163494
rect 57422 163258 64186 163494
rect 64422 163258 71186 163494
rect 71422 163258 78186 163494
rect 78422 163258 85186 163494
rect 85422 163258 92186 163494
rect 92422 163258 99186 163494
rect 99422 163258 106186 163494
rect 106422 163258 113186 163494
rect 113422 163258 120186 163494
rect 120422 163258 127186 163494
rect 127422 163258 134186 163494
rect 134422 163258 141186 163494
rect 141422 163258 148186 163494
rect 148422 163258 155186 163494
rect 155422 163258 162186 163494
rect 162422 163258 169186 163494
rect 169422 163258 176186 163494
rect 176422 163258 183186 163494
rect 183422 163258 190186 163494
rect 190422 163258 197186 163494
rect 197422 163258 204186 163494
rect 204422 163258 211186 163494
rect 211422 163258 218186 163494
rect 218422 163258 225186 163494
rect 225422 163258 232186 163494
rect 232422 163258 239186 163494
rect 239422 163258 246186 163494
rect 246422 163258 253186 163494
rect 253422 163258 260186 163494
rect 260422 163258 267186 163494
rect 267422 163258 274186 163494
rect 274422 163258 281186 163494
rect 281422 163258 288186 163494
rect 288422 163258 295186 163494
rect 295422 163258 302186 163494
rect 302422 163258 309186 163494
rect 309422 163258 316186 163494
rect 316422 163258 323186 163494
rect 323422 163258 330186 163494
rect 330422 163258 337186 163494
rect 337422 163258 344186 163494
rect 344422 163258 351186 163494
rect 351422 163258 358186 163494
rect 358422 163258 365186 163494
rect 365422 163258 372186 163494
rect 372422 163258 379186 163494
rect 379422 163258 386186 163494
rect 386422 163258 393186 163494
rect 393422 163258 400186 163494
rect 400422 163258 407186 163494
rect 407422 163258 414186 163494
rect 414422 163258 421186 163494
rect 421422 163258 428186 163494
rect 428422 163258 435186 163494
rect 435422 163258 442186 163494
rect 442422 163258 449186 163494
rect 449422 163258 456186 163494
rect 456422 163258 463186 163494
rect 463422 163258 470186 163494
rect 470422 163258 477186 163494
rect 477422 163258 484186 163494
rect 484422 163258 491186 163494
rect 491422 163258 498186 163494
rect 498422 163258 505186 163494
rect 505422 163258 512186 163494
rect 512422 163258 519186 163494
rect 519422 163258 526186 163494
rect 526422 163258 533186 163494
rect 533422 163258 540186 163494
rect 540422 163258 547186 163494
rect 547422 163258 554186 163494
rect 554422 163258 561186 163494
rect 561422 163258 568186 163494
rect 568422 163258 575186 163494
rect 575422 163258 582186 163494
rect 582422 163258 585818 163494
rect 586054 163258 586138 163494
rect 586374 163258 586458 163494
rect 586694 163258 586778 163494
rect 587014 163258 588874 163494
rect -4950 163216 588874 163258
rect -4950 157434 588874 157476
rect -4950 157198 -4842 157434
rect -4606 157198 -4522 157434
rect -4286 157198 -4202 157434
rect -3966 157198 -3882 157434
rect -3646 157198 2918 157434
rect 3154 157198 9918 157434
rect 10154 157198 16918 157434
rect 17154 157198 23918 157434
rect 24154 157198 30918 157434
rect 31154 157198 37918 157434
rect 38154 157198 44918 157434
rect 45154 157198 51918 157434
rect 52154 157198 58918 157434
rect 59154 157198 65918 157434
rect 66154 157198 72918 157434
rect 73154 157198 79918 157434
rect 80154 157198 86918 157434
rect 87154 157198 93918 157434
rect 94154 157198 100918 157434
rect 101154 157198 107918 157434
rect 108154 157198 114918 157434
rect 115154 157198 121918 157434
rect 122154 157198 128918 157434
rect 129154 157198 135918 157434
rect 136154 157198 142918 157434
rect 143154 157198 149918 157434
rect 150154 157198 156918 157434
rect 157154 157198 163918 157434
rect 164154 157198 170918 157434
rect 171154 157198 177918 157434
rect 178154 157198 184918 157434
rect 185154 157198 191918 157434
rect 192154 157198 198918 157434
rect 199154 157198 205918 157434
rect 206154 157198 212918 157434
rect 213154 157198 219918 157434
rect 220154 157198 226918 157434
rect 227154 157198 233918 157434
rect 234154 157198 240918 157434
rect 241154 157198 247918 157434
rect 248154 157198 254918 157434
rect 255154 157198 261918 157434
rect 262154 157198 268918 157434
rect 269154 157198 275918 157434
rect 276154 157198 282918 157434
rect 283154 157198 289918 157434
rect 290154 157198 296918 157434
rect 297154 157198 303918 157434
rect 304154 157198 310918 157434
rect 311154 157198 317918 157434
rect 318154 157198 324918 157434
rect 325154 157198 331918 157434
rect 332154 157198 338918 157434
rect 339154 157198 345918 157434
rect 346154 157198 352918 157434
rect 353154 157198 359918 157434
rect 360154 157198 366918 157434
rect 367154 157198 373918 157434
rect 374154 157198 380918 157434
rect 381154 157198 387918 157434
rect 388154 157198 394918 157434
rect 395154 157198 401918 157434
rect 402154 157198 408918 157434
rect 409154 157198 415918 157434
rect 416154 157198 422918 157434
rect 423154 157198 429918 157434
rect 430154 157198 436918 157434
rect 437154 157198 443918 157434
rect 444154 157198 450918 157434
rect 451154 157198 457918 157434
rect 458154 157198 464918 157434
rect 465154 157198 471918 157434
rect 472154 157198 478918 157434
rect 479154 157198 485918 157434
rect 486154 157198 492918 157434
rect 493154 157198 499918 157434
rect 500154 157198 506918 157434
rect 507154 157198 513918 157434
rect 514154 157198 520918 157434
rect 521154 157198 527918 157434
rect 528154 157198 534918 157434
rect 535154 157198 541918 157434
rect 542154 157198 548918 157434
rect 549154 157198 555918 157434
rect 556154 157198 562918 157434
rect 563154 157198 569918 157434
rect 570154 157198 576918 157434
rect 577154 157198 587570 157434
rect 587806 157198 587890 157434
rect 588126 157198 588210 157434
rect 588446 157198 588530 157434
rect 588766 157198 588874 157434
rect -4950 157156 588874 157198
rect -4950 156494 588874 156536
rect -4950 156258 -3090 156494
rect -2854 156258 -2770 156494
rect -2534 156258 -2450 156494
rect -2214 156258 -2130 156494
rect -1894 156258 1186 156494
rect 1422 156258 8186 156494
rect 8422 156258 15186 156494
rect 15422 156258 22186 156494
rect 22422 156258 29186 156494
rect 29422 156258 36186 156494
rect 36422 156258 43186 156494
rect 43422 156258 50186 156494
rect 50422 156258 57186 156494
rect 57422 156258 64186 156494
rect 64422 156258 71186 156494
rect 71422 156258 78186 156494
rect 78422 156258 85186 156494
rect 85422 156258 92186 156494
rect 92422 156258 99186 156494
rect 99422 156258 106186 156494
rect 106422 156258 113186 156494
rect 113422 156258 120186 156494
rect 120422 156258 127186 156494
rect 127422 156258 134186 156494
rect 134422 156258 141186 156494
rect 141422 156258 148186 156494
rect 148422 156258 155186 156494
rect 155422 156258 162186 156494
rect 162422 156258 169186 156494
rect 169422 156258 176186 156494
rect 176422 156258 183186 156494
rect 183422 156258 190186 156494
rect 190422 156258 197186 156494
rect 197422 156258 204186 156494
rect 204422 156258 211186 156494
rect 211422 156258 218186 156494
rect 218422 156258 225186 156494
rect 225422 156258 232186 156494
rect 232422 156258 239186 156494
rect 239422 156258 246186 156494
rect 246422 156258 253186 156494
rect 253422 156258 260186 156494
rect 260422 156258 267186 156494
rect 267422 156258 274186 156494
rect 274422 156258 281186 156494
rect 281422 156258 288186 156494
rect 288422 156258 295186 156494
rect 295422 156258 302186 156494
rect 302422 156258 309186 156494
rect 309422 156258 316186 156494
rect 316422 156258 323186 156494
rect 323422 156258 330186 156494
rect 330422 156258 337186 156494
rect 337422 156258 344186 156494
rect 344422 156258 351186 156494
rect 351422 156258 358186 156494
rect 358422 156258 365186 156494
rect 365422 156258 372186 156494
rect 372422 156258 379186 156494
rect 379422 156258 386186 156494
rect 386422 156258 393186 156494
rect 393422 156258 400186 156494
rect 400422 156258 407186 156494
rect 407422 156258 414186 156494
rect 414422 156258 421186 156494
rect 421422 156258 428186 156494
rect 428422 156258 435186 156494
rect 435422 156258 442186 156494
rect 442422 156258 449186 156494
rect 449422 156258 456186 156494
rect 456422 156258 463186 156494
rect 463422 156258 470186 156494
rect 470422 156258 477186 156494
rect 477422 156258 484186 156494
rect 484422 156258 491186 156494
rect 491422 156258 498186 156494
rect 498422 156258 505186 156494
rect 505422 156258 512186 156494
rect 512422 156258 519186 156494
rect 519422 156258 526186 156494
rect 526422 156258 533186 156494
rect 533422 156258 540186 156494
rect 540422 156258 547186 156494
rect 547422 156258 554186 156494
rect 554422 156258 561186 156494
rect 561422 156258 568186 156494
rect 568422 156258 575186 156494
rect 575422 156258 582186 156494
rect 582422 156258 585818 156494
rect 586054 156258 586138 156494
rect 586374 156258 586458 156494
rect 586694 156258 586778 156494
rect 587014 156258 588874 156494
rect -4950 156216 588874 156258
rect -4950 150434 588874 150476
rect -4950 150198 -4842 150434
rect -4606 150198 -4522 150434
rect -4286 150198 -4202 150434
rect -3966 150198 -3882 150434
rect -3646 150198 2918 150434
rect 3154 150198 9918 150434
rect 10154 150198 16918 150434
rect 17154 150198 23918 150434
rect 24154 150198 30918 150434
rect 31154 150198 37918 150434
rect 38154 150198 44918 150434
rect 45154 150198 51918 150434
rect 52154 150198 58918 150434
rect 59154 150198 65918 150434
rect 66154 150198 72918 150434
rect 73154 150198 79918 150434
rect 80154 150198 86918 150434
rect 87154 150198 93918 150434
rect 94154 150198 100918 150434
rect 101154 150198 107918 150434
rect 108154 150198 114918 150434
rect 115154 150198 121918 150434
rect 122154 150198 128918 150434
rect 129154 150198 135918 150434
rect 136154 150198 142918 150434
rect 143154 150198 149918 150434
rect 150154 150198 156918 150434
rect 157154 150198 163918 150434
rect 164154 150198 170918 150434
rect 171154 150198 177918 150434
rect 178154 150198 184918 150434
rect 185154 150198 191918 150434
rect 192154 150198 198918 150434
rect 199154 150198 205918 150434
rect 206154 150198 212918 150434
rect 213154 150198 219918 150434
rect 220154 150198 226918 150434
rect 227154 150198 233918 150434
rect 234154 150198 240918 150434
rect 241154 150198 247918 150434
rect 248154 150198 254918 150434
rect 255154 150198 261918 150434
rect 262154 150198 268918 150434
rect 269154 150198 275918 150434
rect 276154 150198 282918 150434
rect 283154 150198 289918 150434
rect 290154 150198 296918 150434
rect 297154 150198 303918 150434
rect 304154 150198 310918 150434
rect 311154 150198 317918 150434
rect 318154 150198 324918 150434
rect 325154 150198 331918 150434
rect 332154 150198 338918 150434
rect 339154 150198 345918 150434
rect 346154 150198 352918 150434
rect 353154 150198 359918 150434
rect 360154 150198 366918 150434
rect 367154 150198 373918 150434
rect 374154 150198 380918 150434
rect 381154 150198 387918 150434
rect 388154 150198 394918 150434
rect 395154 150198 401918 150434
rect 402154 150198 408918 150434
rect 409154 150198 415918 150434
rect 416154 150198 422918 150434
rect 423154 150198 429918 150434
rect 430154 150198 436918 150434
rect 437154 150198 443918 150434
rect 444154 150198 450918 150434
rect 451154 150198 457918 150434
rect 458154 150198 464918 150434
rect 465154 150198 471918 150434
rect 472154 150198 478918 150434
rect 479154 150198 485918 150434
rect 486154 150198 492918 150434
rect 493154 150198 499918 150434
rect 500154 150198 506918 150434
rect 507154 150198 513918 150434
rect 514154 150198 520918 150434
rect 521154 150198 527918 150434
rect 528154 150198 534918 150434
rect 535154 150198 541918 150434
rect 542154 150198 548918 150434
rect 549154 150198 555918 150434
rect 556154 150198 562918 150434
rect 563154 150198 569918 150434
rect 570154 150198 576918 150434
rect 577154 150198 587570 150434
rect 587806 150198 587890 150434
rect 588126 150198 588210 150434
rect 588446 150198 588530 150434
rect 588766 150198 588874 150434
rect -4950 150156 588874 150198
rect -4950 149494 588874 149536
rect -4950 149258 -3090 149494
rect -2854 149258 -2770 149494
rect -2534 149258 -2450 149494
rect -2214 149258 -2130 149494
rect -1894 149258 1186 149494
rect 1422 149258 8186 149494
rect 8422 149258 15186 149494
rect 15422 149258 22186 149494
rect 22422 149258 29186 149494
rect 29422 149258 36186 149494
rect 36422 149258 43186 149494
rect 43422 149258 50186 149494
rect 50422 149258 57186 149494
rect 57422 149258 64186 149494
rect 64422 149258 71186 149494
rect 71422 149258 78186 149494
rect 78422 149258 85186 149494
rect 85422 149258 92186 149494
rect 92422 149258 99186 149494
rect 99422 149258 106186 149494
rect 106422 149258 113186 149494
rect 113422 149258 120186 149494
rect 120422 149258 127186 149494
rect 127422 149258 134186 149494
rect 134422 149258 141186 149494
rect 141422 149258 148186 149494
rect 148422 149258 155186 149494
rect 155422 149258 162186 149494
rect 162422 149258 169186 149494
rect 169422 149258 176186 149494
rect 176422 149258 183186 149494
rect 183422 149258 190186 149494
rect 190422 149258 197186 149494
rect 197422 149258 204186 149494
rect 204422 149258 211186 149494
rect 211422 149258 218186 149494
rect 218422 149258 225186 149494
rect 225422 149258 232186 149494
rect 232422 149258 239186 149494
rect 239422 149258 246186 149494
rect 246422 149258 253186 149494
rect 253422 149258 260186 149494
rect 260422 149258 267186 149494
rect 267422 149258 274186 149494
rect 274422 149258 281186 149494
rect 281422 149258 288186 149494
rect 288422 149258 295186 149494
rect 295422 149258 302186 149494
rect 302422 149258 309186 149494
rect 309422 149258 316186 149494
rect 316422 149258 323186 149494
rect 323422 149258 330186 149494
rect 330422 149258 337186 149494
rect 337422 149258 344186 149494
rect 344422 149258 351186 149494
rect 351422 149258 358186 149494
rect 358422 149258 365186 149494
rect 365422 149258 372186 149494
rect 372422 149258 379186 149494
rect 379422 149258 386186 149494
rect 386422 149258 393186 149494
rect 393422 149258 400186 149494
rect 400422 149258 407186 149494
rect 407422 149258 414186 149494
rect 414422 149258 421186 149494
rect 421422 149258 428186 149494
rect 428422 149258 435186 149494
rect 435422 149258 442186 149494
rect 442422 149258 449186 149494
rect 449422 149258 456186 149494
rect 456422 149258 463186 149494
rect 463422 149258 470186 149494
rect 470422 149258 477186 149494
rect 477422 149258 484186 149494
rect 484422 149258 491186 149494
rect 491422 149258 498186 149494
rect 498422 149258 505186 149494
rect 505422 149258 512186 149494
rect 512422 149258 519186 149494
rect 519422 149258 526186 149494
rect 526422 149258 533186 149494
rect 533422 149258 540186 149494
rect 540422 149258 547186 149494
rect 547422 149258 554186 149494
rect 554422 149258 561186 149494
rect 561422 149258 568186 149494
rect 568422 149258 575186 149494
rect 575422 149258 582186 149494
rect 582422 149258 585818 149494
rect 586054 149258 586138 149494
rect 586374 149258 586458 149494
rect 586694 149258 586778 149494
rect 587014 149258 588874 149494
rect -4950 149216 588874 149258
rect -4950 143434 588874 143476
rect -4950 143198 -4842 143434
rect -4606 143198 -4522 143434
rect -4286 143198 -4202 143434
rect -3966 143198 -3882 143434
rect -3646 143198 2918 143434
rect 3154 143198 9918 143434
rect 10154 143198 16918 143434
rect 17154 143198 23918 143434
rect 24154 143198 30918 143434
rect 31154 143198 37918 143434
rect 38154 143198 44918 143434
rect 45154 143198 51918 143434
rect 52154 143198 58918 143434
rect 59154 143198 65918 143434
rect 66154 143198 72918 143434
rect 73154 143198 79918 143434
rect 80154 143198 86918 143434
rect 87154 143198 93918 143434
rect 94154 143198 100918 143434
rect 101154 143198 107918 143434
rect 108154 143198 114918 143434
rect 115154 143198 121918 143434
rect 122154 143198 128918 143434
rect 129154 143198 135918 143434
rect 136154 143198 142918 143434
rect 143154 143198 149918 143434
rect 150154 143198 156918 143434
rect 157154 143198 163918 143434
rect 164154 143198 170918 143434
rect 171154 143198 177918 143434
rect 178154 143198 184918 143434
rect 185154 143198 191918 143434
rect 192154 143198 198918 143434
rect 199154 143198 205918 143434
rect 206154 143198 212918 143434
rect 213154 143198 219918 143434
rect 220154 143198 226918 143434
rect 227154 143198 233918 143434
rect 234154 143198 240918 143434
rect 241154 143198 247918 143434
rect 248154 143198 254918 143434
rect 255154 143198 261918 143434
rect 262154 143198 268918 143434
rect 269154 143198 275918 143434
rect 276154 143198 282918 143434
rect 283154 143198 289918 143434
rect 290154 143198 296918 143434
rect 297154 143198 303918 143434
rect 304154 143198 310918 143434
rect 311154 143198 317918 143434
rect 318154 143198 324918 143434
rect 325154 143198 331918 143434
rect 332154 143198 338918 143434
rect 339154 143198 345918 143434
rect 346154 143198 352918 143434
rect 353154 143198 359918 143434
rect 360154 143198 366918 143434
rect 367154 143198 373918 143434
rect 374154 143198 380918 143434
rect 381154 143198 387918 143434
rect 388154 143198 394918 143434
rect 395154 143198 401918 143434
rect 402154 143198 408918 143434
rect 409154 143198 415918 143434
rect 416154 143198 422918 143434
rect 423154 143198 429918 143434
rect 430154 143198 436918 143434
rect 437154 143198 443918 143434
rect 444154 143198 450918 143434
rect 451154 143198 457918 143434
rect 458154 143198 464918 143434
rect 465154 143198 471918 143434
rect 472154 143198 478918 143434
rect 479154 143198 485918 143434
rect 486154 143198 492918 143434
rect 493154 143198 499918 143434
rect 500154 143198 506918 143434
rect 507154 143198 513918 143434
rect 514154 143198 520918 143434
rect 521154 143198 527918 143434
rect 528154 143198 534918 143434
rect 535154 143198 541918 143434
rect 542154 143198 548918 143434
rect 549154 143198 555918 143434
rect 556154 143198 562918 143434
rect 563154 143198 569918 143434
rect 570154 143198 576918 143434
rect 577154 143198 587570 143434
rect 587806 143198 587890 143434
rect 588126 143198 588210 143434
rect 588446 143198 588530 143434
rect 588766 143198 588874 143434
rect -4950 143156 588874 143198
rect -4950 142494 588874 142536
rect -4950 142258 -3090 142494
rect -2854 142258 -2770 142494
rect -2534 142258 -2450 142494
rect -2214 142258 -2130 142494
rect -1894 142258 1186 142494
rect 1422 142258 8186 142494
rect 8422 142258 15186 142494
rect 15422 142258 22186 142494
rect 22422 142258 29186 142494
rect 29422 142258 36186 142494
rect 36422 142258 43186 142494
rect 43422 142258 50186 142494
rect 50422 142258 57186 142494
rect 57422 142258 64186 142494
rect 64422 142258 71186 142494
rect 71422 142258 78186 142494
rect 78422 142258 85186 142494
rect 85422 142258 92186 142494
rect 92422 142258 99186 142494
rect 99422 142258 106186 142494
rect 106422 142258 113186 142494
rect 113422 142258 120186 142494
rect 120422 142258 127186 142494
rect 127422 142258 134186 142494
rect 134422 142258 141186 142494
rect 141422 142258 148186 142494
rect 148422 142258 155186 142494
rect 155422 142258 162186 142494
rect 162422 142258 169186 142494
rect 169422 142258 176186 142494
rect 176422 142258 183186 142494
rect 183422 142258 190186 142494
rect 190422 142258 197186 142494
rect 197422 142258 204186 142494
rect 204422 142258 211186 142494
rect 211422 142258 218186 142494
rect 218422 142258 225186 142494
rect 225422 142258 232186 142494
rect 232422 142258 239186 142494
rect 239422 142258 246186 142494
rect 246422 142258 253186 142494
rect 253422 142258 260186 142494
rect 260422 142258 267186 142494
rect 267422 142258 274186 142494
rect 274422 142258 281186 142494
rect 281422 142258 288186 142494
rect 288422 142258 295186 142494
rect 295422 142258 302186 142494
rect 302422 142258 309186 142494
rect 309422 142258 316186 142494
rect 316422 142258 323186 142494
rect 323422 142258 330186 142494
rect 330422 142258 337186 142494
rect 337422 142258 344186 142494
rect 344422 142258 351186 142494
rect 351422 142258 358186 142494
rect 358422 142258 365186 142494
rect 365422 142258 372186 142494
rect 372422 142258 379186 142494
rect 379422 142258 386186 142494
rect 386422 142258 393186 142494
rect 393422 142258 400186 142494
rect 400422 142258 407186 142494
rect 407422 142258 414186 142494
rect 414422 142258 421186 142494
rect 421422 142258 428186 142494
rect 428422 142258 435186 142494
rect 435422 142258 442186 142494
rect 442422 142258 449186 142494
rect 449422 142258 456186 142494
rect 456422 142258 463186 142494
rect 463422 142258 470186 142494
rect 470422 142258 477186 142494
rect 477422 142258 484186 142494
rect 484422 142258 491186 142494
rect 491422 142258 498186 142494
rect 498422 142258 505186 142494
rect 505422 142258 512186 142494
rect 512422 142258 519186 142494
rect 519422 142258 526186 142494
rect 526422 142258 533186 142494
rect 533422 142258 540186 142494
rect 540422 142258 547186 142494
rect 547422 142258 554186 142494
rect 554422 142258 561186 142494
rect 561422 142258 568186 142494
rect 568422 142258 575186 142494
rect 575422 142258 582186 142494
rect 582422 142258 585818 142494
rect 586054 142258 586138 142494
rect 586374 142258 586458 142494
rect 586694 142258 586778 142494
rect 587014 142258 588874 142494
rect -4950 142216 588874 142258
rect -4950 136434 588874 136476
rect -4950 136198 -4842 136434
rect -4606 136198 -4522 136434
rect -4286 136198 -4202 136434
rect -3966 136198 -3882 136434
rect -3646 136198 2918 136434
rect 3154 136198 9918 136434
rect 10154 136198 16918 136434
rect 17154 136198 23918 136434
rect 24154 136198 30918 136434
rect 31154 136198 37918 136434
rect 38154 136198 44918 136434
rect 45154 136198 51918 136434
rect 52154 136198 58918 136434
rect 59154 136198 65918 136434
rect 66154 136198 72918 136434
rect 73154 136198 79918 136434
rect 80154 136198 86918 136434
rect 87154 136198 93918 136434
rect 94154 136198 100918 136434
rect 101154 136198 107918 136434
rect 108154 136198 114918 136434
rect 115154 136198 121918 136434
rect 122154 136198 128918 136434
rect 129154 136198 135918 136434
rect 136154 136198 142918 136434
rect 143154 136198 149918 136434
rect 150154 136198 156918 136434
rect 157154 136198 163918 136434
rect 164154 136198 170918 136434
rect 171154 136198 177918 136434
rect 178154 136198 184918 136434
rect 185154 136198 191918 136434
rect 192154 136198 198918 136434
rect 199154 136198 205918 136434
rect 206154 136198 212918 136434
rect 213154 136198 219918 136434
rect 220154 136198 226918 136434
rect 227154 136198 233918 136434
rect 234154 136198 240918 136434
rect 241154 136198 247918 136434
rect 248154 136198 254918 136434
rect 255154 136198 261918 136434
rect 262154 136198 268918 136434
rect 269154 136198 275918 136434
rect 276154 136198 282918 136434
rect 283154 136198 289918 136434
rect 290154 136198 296918 136434
rect 297154 136198 303918 136434
rect 304154 136198 310918 136434
rect 311154 136198 317918 136434
rect 318154 136198 324918 136434
rect 325154 136198 331918 136434
rect 332154 136198 338918 136434
rect 339154 136198 345918 136434
rect 346154 136198 352918 136434
rect 353154 136198 359918 136434
rect 360154 136198 366918 136434
rect 367154 136198 373918 136434
rect 374154 136198 380918 136434
rect 381154 136198 387918 136434
rect 388154 136198 394918 136434
rect 395154 136198 401918 136434
rect 402154 136198 408918 136434
rect 409154 136198 415918 136434
rect 416154 136198 422918 136434
rect 423154 136198 429918 136434
rect 430154 136198 436918 136434
rect 437154 136198 443918 136434
rect 444154 136198 450918 136434
rect 451154 136198 457918 136434
rect 458154 136198 464918 136434
rect 465154 136198 471918 136434
rect 472154 136198 478918 136434
rect 479154 136198 485918 136434
rect 486154 136198 492918 136434
rect 493154 136198 499918 136434
rect 500154 136198 506918 136434
rect 507154 136198 513918 136434
rect 514154 136198 520918 136434
rect 521154 136198 527918 136434
rect 528154 136198 534918 136434
rect 535154 136198 541918 136434
rect 542154 136198 548918 136434
rect 549154 136198 555918 136434
rect 556154 136198 562918 136434
rect 563154 136198 569918 136434
rect 570154 136198 576918 136434
rect 577154 136198 587570 136434
rect 587806 136198 587890 136434
rect 588126 136198 588210 136434
rect 588446 136198 588530 136434
rect 588766 136198 588874 136434
rect -4950 136156 588874 136198
rect -4950 135494 588874 135536
rect -4950 135258 -3090 135494
rect -2854 135258 -2770 135494
rect -2534 135258 -2450 135494
rect -2214 135258 -2130 135494
rect -1894 135258 1186 135494
rect 1422 135258 8186 135494
rect 8422 135258 15186 135494
rect 15422 135258 22186 135494
rect 22422 135258 29186 135494
rect 29422 135258 36186 135494
rect 36422 135258 43186 135494
rect 43422 135258 50186 135494
rect 50422 135258 57186 135494
rect 57422 135258 64186 135494
rect 64422 135258 71186 135494
rect 71422 135258 78186 135494
rect 78422 135258 85186 135494
rect 85422 135258 92186 135494
rect 92422 135258 99186 135494
rect 99422 135258 106186 135494
rect 106422 135258 113186 135494
rect 113422 135258 120186 135494
rect 120422 135258 127186 135494
rect 127422 135258 134186 135494
rect 134422 135258 141186 135494
rect 141422 135258 148186 135494
rect 148422 135258 155186 135494
rect 155422 135258 162186 135494
rect 162422 135258 169186 135494
rect 169422 135258 176186 135494
rect 176422 135258 183186 135494
rect 183422 135258 190186 135494
rect 190422 135258 197186 135494
rect 197422 135258 204186 135494
rect 204422 135258 211186 135494
rect 211422 135258 218186 135494
rect 218422 135258 225186 135494
rect 225422 135258 232186 135494
rect 232422 135258 239186 135494
rect 239422 135258 246186 135494
rect 246422 135258 253186 135494
rect 253422 135258 260186 135494
rect 260422 135258 267186 135494
rect 267422 135258 274186 135494
rect 274422 135258 281186 135494
rect 281422 135258 288186 135494
rect 288422 135258 295186 135494
rect 295422 135258 302186 135494
rect 302422 135258 309186 135494
rect 309422 135258 316186 135494
rect 316422 135258 323186 135494
rect 323422 135258 330186 135494
rect 330422 135258 337186 135494
rect 337422 135258 344186 135494
rect 344422 135258 351186 135494
rect 351422 135258 358186 135494
rect 358422 135258 365186 135494
rect 365422 135258 372186 135494
rect 372422 135258 379186 135494
rect 379422 135258 386186 135494
rect 386422 135258 393186 135494
rect 393422 135258 400186 135494
rect 400422 135258 407186 135494
rect 407422 135258 414186 135494
rect 414422 135258 421186 135494
rect 421422 135258 428186 135494
rect 428422 135258 435186 135494
rect 435422 135258 442186 135494
rect 442422 135258 449186 135494
rect 449422 135258 456186 135494
rect 456422 135258 463186 135494
rect 463422 135258 470186 135494
rect 470422 135258 477186 135494
rect 477422 135258 484186 135494
rect 484422 135258 491186 135494
rect 491422 135258 498186 135494
rect 498422 135258 505186 135494
rect 505422 135258 512186 135494
rect 512422 135258 519186 135494
rect 519422 135258 526186 135494
rect 526422 135258 533186 135494
rect 533422 135258 540186 135494
rect 540422 135258 547186 135494
rect 547422 135258 554186 135494
rect 554422 135258 561186 135494
rect 561422 135258 568186 135494
rect 568422 135258 575186 135494
rect 575422 135258 582186 135494
rect 582422 135258 585818 135494
rect 586054 135258 586138 135494
rect 586374 135258 586458 135494
rect 586694 135258 586778 135494
rect 587014 135258 588874 135494
rect -4950 135216 588874 135258
rect -4950 129434 588874 129476
rect -4950 129198 -4842 129434
rect -4606 129198 -4522 129434
rect -4286 129198 -4202 129434
rect -3966 129198 -3882 129434
rect -3646 129198 2918 129434
rect 3154 129198 9918 129434
rect 10154 129198 16918 129434
rect 17154 129198 23918 129434
rect 24154 129198 30918 129434
rect 31154 129198 37918 129434
rect 38154 129198 44918 129434
rect 45154 129198 51918 129434
rect 52154 129198 58918 129434
rect 59154 129198 65918 129434
rect 66154 129198 72918 129434
rect 73154 129198 79918 129434
rect 80154 129198 86918 129434
rect 87154 129198 93918 129434
rect 94154 129198 100918 129434
rect 101154 129198 107918 129434
rect 108154 129198 114918 129434
rect 115154 129198 121918 129434
rect 122154 129198 128918 129434
rect 129154 129198 135918 129434
rect 136154 129198 142918 129434
rect 143154 129198 149918 129434
rect 150154 129198 156918 129434
rect 157154 129198 163918 129434
rect 164154 129198 170918 129434
rect 171154 129198 177918 129434
rect 178154 129198 184918 129434
rect 185154 129198 191918 129434
rect 192154 129198 198918 129434
rect 199154 129198 205918 129434
rect 206154 129198 212918 129434
rect 213154 129198 219918 129434
rect 220154 129198 226918 129434
rect 227154 129198 233918 129434
rect 234154 129198 240918 129434
rect 241154 129198 247918 129434
rect 248154 129198 254918 129434
rect 255154 129198 261918 129434
rect 262154 129198 268918 129434
rect 269154 129198 275918 129434
rect 276154 129198 282918 129434
rect 283154 129198 289918 129434
rect 290154 129198 296918 129434
rect 297154 129198 303918 129434
rect 304154 129198 310918 129434
rect 311154 129198 317918 129434
rect 318154 129198 324918 129434
rect 325154 129198 331918 129434
rect 332154 129198 338918 129434
rect 339154 129198 345918 129434
rect 346154 129198 352918 129434
rect 353154 129198 359918 129434
rect 360154 129198 366918 129434
rect 367154 129198 373918 129434
rect 374154 129198 380918 129434
rect 381154 129198 387918 129434
rect 388154 129198 394918 129434
rect 395154 129198 401918 129434
rect 402154 129198 408918 129434
rect 409154 129198 415918 129434
rect 416154 129198 422918 129434
rect 423154 129198 429918 129434
rect 430154 129198 436918 129434
rect 437154 129198 443918 129434
rect 444154 129198 450918 129434
rect 451154 129198 457918 129434
rect 458154 129198 464918 129434
rect 465154 129198 471918 129434
rect 472154 129198 478918 129434
rect 479154 129198 485918 129434
rect 486154 129198 492918 129434
rect 493154 129198 499918 129434
rect 500154 129198 506918 129434
rect 507154 129198 513918 129434
rect 514154 129198 520918 129434
rect 521154 129198 527918 129434
rect 528154 129198 534918 129434
rect 535154 129198 541918 129434
rect 542154 129198 548918 129434
rect 549154 129198 555918 129434
rect 556154 129198 562918 129434
rect 563154 129198 569918 129434
rect 570154 129198 576918 129434
rect 577154 129198 587570 129434
rect 587806 129198 587890 129434
rect 588126 129198 588210 129434
rect 588446 129198 588530 129434
rect 588766 129198 588874 129434
rect -4950 129156 588874 129198
rect -4950 128494 588874 128536
rect -4950 128258 -3090 128494
rect -2854 128258 -2770 128494
rect -2534 128258 -2450 128494
rect -2214 128258 -2130 128494
rect -1894 128258 1186 128494
rect 1422 128258 8186 128494
rect 8422 128258 15186 128494
rect 15422 128258 22186 128494
rect 22422 128258 29186 128494
rect 29422 128258 36186 128494
rect 36422 128258 43186 128494
rect 43422 128258 50186 128494
rect 50422 128258 57186 128494
rect 57422 128258 64186 128494
rect 64422 128258 71186 128494
rect 71422 128258 78186 128494
rect 78422 128258 85186 128494
rect 85422 128258 92186 128494
rect 92422 128258 99186 128494
rect 99422 128258 106186 128494
rect 106422 128258 113186 128494
rect 113422 128258 120186 128494
rect 120422 128258 127186 128494
rect 127422 128258 134186 128494
rect 134422 128258 141186 128494
rect 141422 128258 148186 128494
rect 148422 128258 155186 128494
rect 155422 128258 162186 128494
rect 162422 128258 169186 128494
rect 169422 128258 176186 128494
rect 176422 128258 183186 128494
rect 183422 128258 190186 128494
rect 190422 128258 197186 128494
rect 197422 128258 204186 128494
rect 204422 128258 211186 128494
rect 211422 128258 218186 128494
rect 218422 128258 225186 128494
rect 225422 128258 232186 128494
rect 232422 128258 239186 128494
rect 239422 128258 246186 128494
rect 246422 128258 253186 128494
rect 253422 128258 260186 128494
rect 260422 128258 267186 128494
rect 267422 128258 274186 128494
rect 274422 128258 281186 128494
rect 281422 128258 288186 128494
rect 288422 128258 295186 128494
rect 295422 128258 302186 128494
rect 302422 128258 309186 128494
rect 309422 128258 316186 128494
rect 316422 128258 323186 128494
rect 323422 128258 330186 128494
rect 330422 128258 337186 128494
rect 337422 128258 344186 128494
rect 344422 128258 351186 128494
rect 351422 128258 358186 128494
rect 358422 128258 365186 128494
rect 365422 128258 372186 128494
rect 372422 128258 379186 128494
rect 379422 128258 386186 128494
rect 386422 128258 393186 128494
rect 393422 128258 400186 128494
rect 400422 128258 407186 128494
rect 407422 128258 414186 128494
rect 414422 128258 421186 128494
rect 421422 128258 428186 128494
rect 428422 128258 435186 128494
rect 435422 128258 442186 128494
rect 442422 128258 449186 128494
rect 449422 128258 456186 128494
rect 456422 128258 463186 128494
rect 463422 128258 470186 128494
rect 470422 128258 477186 128494
rect 477422 128258 484186 128494
rect 484422 128258 491186 128494
rect 491422 128258 498186 128494
rect 498422 128258 505186 128494
rect 505422 128258 512186 128494
rect 512422 128258 519186 128494
rect 519422 128258 526186 128494
rect 526422 128258 533186 128494
rect 533422 128258 540186 128494
rect 540422 128258 547186 128494
rect 547422 128258 554186 128494
rect 554422 128258 561186 128494
rect 561422 128258 568186 128494
rect 568422 128258 575186 128494
rect 575422 128258 582186 128494
rect 582422 128258 585818 128494
rect 586054 128258 586138 128494
rect 586374 128258 586458 128494
rect 586694 128258 586778 128494
rect 587014 128258 588874 128494
rect -4950 128216 588874 128258
rect -4950 122434 588874 122476
rect -4950 122198 -4842 122434
rect -4606 122198 -4522 122434
rect -4286 122198 -4202 122434
rect -3966 122198 -3882 122434
rect -3646 122198 2918 122434
rect 3154 122198 9918 122434
rect 10154 122198 16918 122434
rect 17154 122198 23918 122434
rect 24154 122198 30918 122434
rect 31154 122198 37918 122434
rect 38154 122198 44918 122434
rect 45154 122198 51918 122434
rect 52154 122198 58918 122434
rect 59154 122198 65918 122434
rect 66154 122198 72918 122434
rect 73154 122198 79918 122434
rect 80154 122198 86918 122434
rect 87154 122198 93918 122434
rect 94154 122198 100918 122434
rect 101154 122198 107918 122434
rect 108154 122198 114918 122434
rect 115154 122198 121918 122434
rect 122154 122198 128918 122434
rect 129154 122198 135918 122434
rect 136154 122198 142918 122434
rect 143154 122198 149918 122434
rect 150154 122198 156918 122434
rect 157154 122198 163918 122434
rect 164154 122198 170918 122434
rect 171154 122198 177918 122434
rect 178154 122198 184918 122434
rect 185154 122198 191918 122434
rect 192154 122198 198918 122434
rect 199154 122198 205918 122434
rect 206154 122198 212918 122434
rect 213154 122198 219918 122434
rect 220154 122198 226918 122434
rect 227154 122198 233918 122434
rect 234154 122198 240918 122434
rect 241154 122198 247918 122434
rect 248154 122198 254918 122434
rect 255154 122198 261918 122434
rect 262154 122198 268918 122434
rect 269154 122198 275918 122434
rect 276154 122198 282918 122434
rect 283154 122198 289918 122434
rect 290154 122198 296918 122434
rect 297154 122198 303918 122434
rect 304154 122198 310918 122434
rect 311154 122198 317918 122434
rect 318154 122198 324918 122434
rect 325154 122198 331918 122434
rect 332154 122198 338918 122434
rect 339154 122198 345918 122434
rect 346154 122198 352918 122434
rect 353154 122198 359918 122434
rect 360154 122198 366918 122434
rect 367154 122198 373918 122434
rect 374154 122198 380918 122434
rect 381154 122198 387918 122434
rect 388154 122198 394918 122434
rect 395154 122198 401918 122434
rect 402154 122198 408918 122434
rect 409154 122198 415918 122434
rect 416154 122198 422918 122434
rect 423154 122198 429918 122434
rect 430154 122198 436918 122434
rect 437154 122198 443918 122434
rect 444154 122198 450918 122434
rect 451154 122198 457918 122434
rect 458154 122198 464918 122434
rect 465154 122198 471918 122434
rect 472154 122198 478918 122434
rect 479154 122198 485918 122434
rect 486154 122198 492918 122434
rect 493154 122198 499918 122434
rect 500154 122198 506918 122434
rect 507154 122198 513918 122434
rect 514154 122198 520918 122434
rect 521154 122198 527918 122434
rect 528154 122198 534918 122434
rect 535154 122198 541918 122434
rect 542154 122198 548918 122434
rect 549154 122198 555918 122434
rect 556154 122198 562918 122434
rect 563154 122198 569918 122434
rect 570154 122198 576918 122434
rect 577154 122198 587570 122434
rect 587806 122198 587890 122434
rect 588126 122198 588210 122434
rect 588446 122198 588530 122434
rect 588766 122198 588874 122434
rect -4950 122156 588874 122198
rect -4950 121494 588874 121536
rect -4950 121258 -3090 121494
rect -2854 121258 -2770 121494
rect -2534 121258 -2450 121494
rect -2214 121258 -2130 121494
rect -1894 121258 1186 121494
rect 1422 121258 8186 121494
rect 8422 121258 15186 121494
rect 15422 121258 22186 121494
rect 22422 121258 29186 121494
rect 29422 121258 36186 121494
rect 36422 121258 43186 121494
rect 43422 121258 50186 121494
rect 50422 121258 57186 121494
rect 57422 121258 64186 121494
rect 64422 121258 71186 121494
rect 71422 121258 78186 121494
rect 78422 121258 85186 121494
rect 85422 121258 92186 121494
rect 92422 121258 99186 121494
rect 99422 121258 106186 121494
rect 106422 121258 113186 121494
rect 113422 121258 120186 121494
rect 120422 121258 127186 121494
rect 127422 121258 134186 121494
rect 134422 121258 141186 121494
rect 141422 121258 148186 121494
rect 148422 121258 155186 121494
rect 155422 121258 162186 121494
rect 162422 121258 169186 121494
rect 169422 121258 176186 121494
rect 176422 121258 183186 121494
rect 183422 121258 190186 121494
rect 190422 121258 197186 121494
rect 197422 121258 204186 121494
rect 204422 121258 211186 121494
rect 211422 121258 218186 121494
rect 218422 121258 225186 121494
rect 225422 121258 232186 121494
rect 232422 121258 239186 121494
rect 239422 121258 246186 121494
rect 246422 121258 253186 121494
rect 253422 121258 260186 121494
rect 260422 121258 267186 121494
rect 267422 121258 274186 121494
rect 274422 121258 281186 121494
rect 281422 121258 288186 121494
rect 288422 121258 295186 121494
rect 295422 121258 302186 121494
rect 302422 121258 309186 121494
rect 309422 121258 316186 121494
rect 316422 121258 323186 121494
rect 323422 121258 330186 121494
rect 330422 121258 337186 121494
rect 337422 121258 344186 121494
rect 344422 121258 351186 121494
rect 351422 121258 358186 121494
rect 358422 121258 365186 121494
rect 365422 121258 372186 121494
rect 372422 121258 379186 121494
rect 379422 121258 386186 121494
rect 386422 121258 393186 121494
rect 393422 121258 400186 121494
rect 400422 121258 407186 121494
rect 407422 121258 414186 121494
rect 414422 121258 421186 121494
rect 421422 121258 428186 121494
rect 428422 121258 435186 121494
rect 435422 121258 442186 121494
rect 442422 121258 449186 121494
rect 449422 121258 456186 121494
rect 456422 121258 463186 121494
rect 463422 121258 470186 121494
rect 470422 121258 477186 121494
rect 477422 121258 484186 121494
rect 484422 121258 491186 121494
rect 491422 121258 498186 121494
rect 498422 121258 505186 121494
rect 505422 121258 512186 121494
rect 512422 121258 519186 121494
rect 519422 121258 526186 121494
rect 526422 121258 533186 121494
rect 533422 121258 540186 121494
rect 540422 121258 547186 121494
rect 547422 121258 554186 121494
rect 554422 121258 561186 121494
rect 561422 121258 568186 121494
rect 568422 121258 575186 121494
rect 575422 121258 582186 121494
rect 582422 121258 585818 121494
rect 586054 121258 586138 121494
rect 586374 121258 586458 121494
rect 586694 121258 586778 121494
rect 587014 121258 588874 121494
rect -4950 121216 588874 121258
rect -4950 115434 588874 115476
rect -4950 115198 -4842 115434
rect -4606 115198 -4522 115434
rect -4286 115198 -4202 115434
rect -3966 115198 -3882 115434
rect -3646 115198 2918 115434
rect 3154 115198 9918 115434
rect 10154 115198 16918 115434
rect 17154 115198 23918 115434
rect 24154 115198 30918 115434
rect 31154 115198 37918 115434
rect 38154 115198 44918 115434
rect 45154 115198 51918 115434
rect 52154 115198 58918 115434
rect 59154 115198 65918 115434
rect 66154 115198 72918 115434
rect 73154 115198 79918 115434
rect 80154 115198 86918 115434
rect 87154 115198 93918 115434
rect 94154 115198 100918 115434
rect 101154 115198 107918 115434
rect 108154 115198 114918 115434
rect 115154 115198 121918 115434
rect 122154 115198 128918 115434
rect 129154 115198 135918 115434
rect 136154 115198 142918 115434
rect 143154 115198 149918 115434
rect 150154 115198 156918 115434
rect 157154 115198 163918 115434
rect 164154 115198 170918 115434
rect 171154 115198 177918 115434
rect 178154 115198 184918 115434
rect 185154 115198 191918 115434
rect 192154 115198 198918 115434
rect 199154 115198 205918 115434
rect 206154 115198 212918 115434
rect 213154 115198 219918 115434
rect 220154 115198 226918 115434
rect 227154 115198 233918 115434
rect 234154 115198 240918 115434
rect 241154 115198 247918 115434
rect 248154 115198 254918 115434
rect 255154 115198 261918 115434
rect 262154 115198 268918 115434
rect 269154 115198 275918 115434
rect 276154 115198 282918 115434
rect 283154 115198 289918 115434
rect 290154 115198 296918 115434
rect 297154 115198 303918 115434
rect 304154 115198 310918 115434
rect 311154 115198 317918 115434
rect 318154 115198 324918 115434
rect 325154 115198 331918 115434
rect 332154 115198 338918 115434
rect 339154 115198 345918 115434
rect 346154 115198 352918 115434
rect 353154 115198 359918 115434
rect 360154 115198 366918 115434
rect 367154 115198 373918 115434
rect 374154 115198 380918 115434
rect 381154 115198 387918 115434
rect 388154 115198 394918 115434
rect 395154 115198 401918 115434
rect 402154 115198 408918 115434
rect 409154 115198 415918 115434
rect 416154 115198 422918 115434
rect 423154 115198 429918 115434
rect 430154 115198 436918 115434
rect 437154 115198 443918 115434
rect 444154 115198 450918 115434
rect 451154 115198 457918 115434
rect 458154 115198 464918 115434
rect 465154 115198 471918 115434
rect 472154 115198 478918 115434
rect 479154 115198 485918 115434
rect 486154 115198 492918 115434
rect 493154 115198 499918 115434
rect 500154 115198 506918 115434
rect 507154 115198 513918 115434
rect 514154 115198 520918 115434
rect 521154 115198 527918 115434
rect 528154 115198 534918 115434
rect 535154 115198 541918 115434
rect 542154 115198 548918 115434
rect 549154 115198 555918 115434
rect 556154 115198 562918 115434
rect 563154 115198 569918 115434
rect 570154 115198 576918 115434
rect 577154 115198 587570 115434
rect 587806 115198 587890 115434
rect 588126 115198 588210 115434
rect 588446 115198 588530 115434
rect 588766 115198 588874 115434
rect -4950 115156 588874 115198
rect -4950 114494 588874 114536
rect -4950 114258 -3090 114494
rect -2854 114258 -2770 114494
rect -2534 114258 -2450 114494
rect -2214 114258 -2130 114494
rect -1894 114258 1186 114494
rect 1422 114258 8186 114494
rect 8422 114258 15186 114494
rect 15422 114258 22186 114494
rect 22422 114258 29186 114494
rect 29422 114258 36186 114494
rect 36422 114258 43186 114494
rect 43422 114258 50186 114494
rect 50422 114258 57186 114494
rect 57422 114258 64186 114494
rect 64422 114258 71186 114494
rect 71422 114258 78186 114494
rect 78422 114258 85186 114494
rect 85422 114258 92186 114494
rect 92422 114258 99186 114494
rect 99422 114258 106186 114494
rect 106422 114258 113186 114494
rect 113422 114258 120186 114494
rect 120422 114258 127186 114494
rect 127422 114258 134186 114494
rect 134422 114258 141186 114494
rect 141422 114258 148186 114494
rect 148422 114258 155186 114494
rect 155422 114258 162186 114494
rect 162422 114258 169186 114494
rect 169422 114258 176186 114494
rect 176422 114258 183186 114494
rect 183422 114258 190186 114494
rect 190422 114258 197186 114494
rect 197422 114258 204186 114494
rect 204422 114258 211186 114494
rect 211422 114258 218186 114494
rect 218422 114258 225186 114494
rect 225422 114258 232186 114494
rect 232422 114258 239186 114494
rect 239422 114258 246186 114494
rect 246422 114258 253186 114494
rect 253422 114258 260186 114494
rect 260422 114258 267186 114494
rect 267422 114258 274186 114494
rect 274422 114258 281186 114494
rect 281422 114258 288186 114494
rect 288422 114258 295186 114494
rect 295422 114258 302186 114494
rect 302422 114258 309186 114494
rect 309422 114258 316186 114494
rect 316422 114258 323186 114494
rect 323422 114258 330186 114494
rect 330422 114258 337186 114494
rect 337422 114258 344186 114494
rect 344422 114258 351186 114494
rect 351422 114258 358186 114494
rect 358422 114258 365186 114494
rect 365422 114258 372186 114494
rect 372422 114258 379186 114494
rect 379422 114258 386186 114494
rect 386422 114258 393186 114494
rect 393422 114258 400186 114494
rect 400422 114258 407186 114494
rect 407422 114258 414186 114494
rect 414422 114258 421186 114494
rect 421422 114258 428186 114494
rect 428422 114258 435186 114494
rect 435422 114258 442186 114494
rect 442422 114258 449186 114494
rect 449422 114258 456186 114494
rect 456422 114258 463186 114494
rect 463422 114258 470186 114494
rect 470422 114258 477186 114494
rect 477422 114258 484186 114494
rect 484422 114258 491186 114494
rect 491422 114258 498186 114494
rect 498422 114258 505186 114494
rect 505422 114258 512186 114494
rect 512422 114258 519186 114494
rect 519422 114258 526186 114494
rect 526422 114258 533186 114494
rect 533422 114258 540186 114494
rect 540422 114258 547186 114494
rect 547422 114258 554186 114494
rect 554422 114258 561186 114494
rect 561422 114258 568186 114494
rect 568422 114258 575186 114494
rect 575422 114258 582186 114494
rect 582422 114258 585818 114494
rect 586054 114258 586138 114494
rect 586374 114258 586458 114494
rect 586694 114258 586778 114494
rect 587014 114258 588874 114494
rect -4950 114216 588874 114258
rect -4950 108434 588874 108476
rect -4950 108198 -4842 108434
rect -4606 108198 -4522 108434
rect -4286 108198 -4202 108434
rect -3966 108198 -3882 108434
rect -3646 108198 2918 108434
rect 3154 108198 9918 108434
rect 10154 108198 16918 108434
rect 17154 108198 23918 108434
rect 24154 108198 30918 108434
rect 31154 108198 37918 108434
rect 38154 108198 44918 108434
rect 45154 108198 51918 108434
rect 52154 108198 58918 108434
rect 59154 108198 65918 108434
rect 66154 108198 72918 108434
rect 73154 108198 79918 108434
rect 80154 108198 86918 108434
rect 87154 108198 93918 108434
rect 94154 108198 100918 108434
rect 101154 108198 107918 108434
rect 108154 108198 114918 108434
rect 115154 108198 121918 108434
rect 122154 108198 128918 108434
rect 129154 108198 135918 108434
rect 136154 108198 142918 108434
rect 143154 108198 149918 108434
rect 150154 108198 156918 108434
rect 157154 108198 163918 108434
rect 164154 108198 170918 108434
rect 171154 108198 177918 108434
rect 178154 108198 184918 108434
rect 185154 108198 191918 108434
rect 192154 108198 198918 108434
rect 199154 108198 205918 108434
rect 206154 108198 212918 108434
rect 213154 108198 219918 108434
rect 220154 108198 226918 108434
rect 227154 108198 233918 108434
rect 234154 108198 240918 108434
rect 241154 108198 247918 108434
rect 248154 108198 254918 108434
rect 255154 108198 261918 108434
rect 262154 108198 268918 108434
rect 269154 108198 275918 108434
rect 276154 108198 282918 108434
rect 283154 108198 289918 108434
rect 290154 108198 296918 108434
rect 297154 108198 303918 108434
rect 304154 108198 310918 108434
rect 311154 108198 317918 108434
rect 318154 108198 324918 108434
rect 325154 108198 331918 108434
rect 332154 108198 338918 108434
rect 339154 108198 345918 108434
rect 346154 108198 352918 108434
rect 353154 108198 359918 108434
rect 360154 108198 366918 108434
rect 367154 108198 373918 108434
rect 374154 108198 380918 108434
rect 381154 108198 387918 108434
rect 388154 108198 394918 108434
rect 395154 108198 401918 108434
rect 402154 108198 408918 108434
rect 409154 108198 415918 108434
rect 416154 108198 422918 108434
rect 423154 108198 429918 108434
rect 430154 108198 436918 108434
rect 437154 108198 443918 108434
rect 444154 108198 450918 108434
rect 451154 108198 457918 108434
rect 458154 108198 464918 108434
rect 465154 108198 471918 108434
rect 472154 108198 478918 108434
rect 479154 108198 485918 108434
rect 486154 108198 492918 108434
rect 493154 108198 499918 108434
rect 500154 108198 506918 108434
rect 507154 108198 513918 108434
rect 514154 108198 520918 108434
rect 521154 108198 527918 108434
rect 528154 108198 534918 108434
rect 535154 108198 541918 108434
rect 542154 108198 548918 108434
rect 549154 108198 555918 108434
rect 556154 108198 562918 108434
rect 563154 108198 569918 108434
rect 570154 108198 576918 108434
rect 577154 108198 587570 108434
rect 587806 108198 587890 108434
rect 588126 108198 588210 108434
rect 588446 108198 588530 108434
rect 588766 108198 588874 108434
rect -4950 108156 588874 108198
rect -4950 107494 588874 107536
rect -4950 107258 -3090 107494
rect -2854 107258 -2770 107494
rect -2534 107258 -2450 107494
rect -2214 107258 -2130 107494
rect -1894 107258 1186 107494
rect 1422 107258 8186 107494
rect 8422 107258 15186 107494
rect 15422 107258 22186 107494
rect 22422 107258 29186 107494
rect 29422 107258 36186 107494
rect 36422 107258 43186 107494
rect 43422 107258 50186 107494
rect 50422 107258 57186 107494
rect 57422 107258 64186 107494
rect 64422 107258 71186 107494
rect 71422 107258 78186 107494
rect 78422 107258 85186 107494
rect 85422 107258 92186 107494
rect 92422 107258 99186 107494
rect 99422 107258 106186 107494
rect 106422 107258 113186 107494
rect 113422 107258 120186 107494
rect 120422 107258 127186 107494
rect 127422 107258 134186 107494
rect 134422 107258 141186 107494
rect 141422 107258 148186 107494
rect 148422 107258 155186 107494
rect 155422 107258 162186 107494
rect 162422 107258 169186 107494
rect 169422 107258 176186 107494
rect 176422 107258 183186 107494
rect 183422 107258 190186 107494
rect 190422 107258 197186 107494
rect 197422 107258 204186 107494
rect 204422 107258 211186 107494
rect 211422 107258 218186 107494
rect 218422 107258 225186 107494
rect 225422 107258 232186 107494
rect 232422 107258 239186 107494
rect 239422 107258 246186 107494
rect 246422 107258 253186 107494
rect 253422 107258 260186 107494
rect 260422 107258 267186 107494
rect 267422 107258 274186 107494
rect 274422 107258 281186 107494
rect 281422 107258 288186 107494
rect 288422 107258 295186 107494
rect 295422 107258 302186 107494
rect 302422 107258 309186 107494
rect 309422 107258 316186 107494
rect 316422 107258 323186 107494
rect 323422 107258 330186 107494
rect 330422 107258 337186 107494
rect 337422 107258 344186 107494
rect 344422 107258 351186 107494
rect 351422 107258 358186 107494
rect 358422 107258 365186 107494
rect 365422 107258 372186 107494
rect 372422 107258 379186 107494
rect 379422 107258 386186 107494
rect 386422 107258 393186 107494
rect 393422 107258 400186 107494
rect 400422 107258 407186 107494
rect 407422 107258 414186 107494
rect 414422 107258 421186 107494
rect 421422 107258 428186 107494
rect 428422 107258 435186 107494
rect 435422 107258 442186 107494
rect 442422 107258 449186 107494
rect 449422 107258 456186 107494
rect 456422 107258 463186 107494
rect 463422 107258 470186 107494
rect 470422 107258 477186 107494
rect 477422 107258 484186 107494
rect 484422 107258 491186 107494
rect 491422 107258 498186 107494
rect 498422 107258 505186 107494
rect 505422 107258 512186 107494
rect 512422 107258 519186 107494
rect 519422 107258 526186 107494
rect 526422 107258 533186 107494
rect 533422 107258 540186 107494
rect 540422 107258 547186 107494
rect 547422 107258 554186 107494
rect 554422 107258 561186 107494
rect 561422 107258 568186 107494
rect 568422 107258 575186 107494
rect 575422 107258 582186 107494
rect 582422 107258 585818 107494
rect 586054 107258 586138 107494
rect 586374 107258 586458 107494
rect 586694 107258 586778 107494
rect 587014 107258 588874 107494
rect -4950 107216 588874 107258
rect -4950 101434 588874 101476
rect -4950 101198 -4842 101434
rect -4606 101198 -4522 101434
rect -4286 101198 -4202 101434
rect -3966 101198 -3882 101434
rect -3646 101198 2918 101434
rect 3154 101198 9918 101434
rect 10154 101198 16918 101434
rect 17154 101198 23918 101434
rect 24154 101198 30918 101434
rect 31154 101198 37918 101434
rect 38154 101198 44918 101434
rect 45154 101198 51918 101434
rect 52154 101198 58918 101434
rect 59154 101198 65918 101434
rect 66154 101198 72918 101434
rect 73154 101198 79918 101434
rect 80154 101198 86918 101434
rect 87154 101198 93918 101434
rect 94154 101198 100918 101434
rect 101154 101198 107918 101434
rect 108154 101198 114918 101434
rect 115154 101198 121918 101434
rect 122154 101198 128918 101434
rect 129154 101198 135918 101434
rect 136154 101198 142918 101434
rect 143154 101198 149918 101434
rect 150154 101198 156918 101434
rect 157154 101198 163918 101434
rect 164154 101198 170918 101434
rect 171154 101198 177918 101434
rect 178154 101198 184918 101434
rect 185154 101198 191918 101434
rect 192154 101198 198918 101434
rect 199154 101198 205918 101434
rect 206154 101198 212918 101434
rect 213154 101198 219918 101434
rect 220154 101198 226918 101434
rect 227154 101198 233918 101434
rect 234154 101198 240918 101434
rect 241154 101198 247918 101434
rect 248154 101198 254918 101434
rect 255154 101198 261918 101434
rect 262154 101198 268918 101434
rect 269154 101198 275918 101434
rect 276154 101198 282918 101434
rect 283154 101198 289918 101434
rect 290154 101198 296918 101434
rect 297154 101198 303918 101434
rect 304154 101198 310918 101434
rect 311154 101198 317918 101434
rect 318154 101198 324918 101434
rect 325154 101198 331918 101434
rect 332154 101198 338918 101434
rect 339154 101198 345918 101434
rect 346154 101198 352918 101434
rect 353154 101198 359918 101434
rect 360154 101198 366918 101434
rect 367154 101198 373918 101434
rect 374154 101198 380918 101434
rect 381154 101198 387918 101434
rect 388154 101198 394918 101434
rect 395154 101198 401918 101434
rect 402154 101198 408918 101434
rect 409154 101198 415918 101434
rect 416154 101198 422918 101434
rect 423154 101198 429918 101434
rect 430154 101198 436918 101434
rect 437154 101198 443918 101434
rect 444154 101198 450918 101434
rect 451154 101198 457918 101434
rect 458154 101198 464918 101434
rect 465154 101198 471918 101434
rect 472154 101198 478918 101434
rect 479154 101198 485918 101434
rect 486154 101198 492918 101434
rect 493154 101198 499918 101434
rect 500154 101198 506918 101434
rect 507154 101198 513918 101434
rect 514154 101198 520918 101434
rect 521154 101198 527918 101434
rect 528154 101198 534918 101434
rect 535154 101198 541918 101434
rect 542154 101198 548918 101434
rect 549154 101198 555918 101434
rect 556154 101198 562918 101434
rect 563154 101198 569918 101434
rect 570154 101198 576918 101434
rect 577154 101198 587570 101434
rect 587806 101198 587890 101434
rect 588126 101198 588210 101434
rect 588446 101198 588530 101434
rect 588766 101198 588874 101434
rect -4950 101156 588874 101198
rect -4950 100494 588874 100536
rect -4950 100258 -3090 100494
rect -2854 100258 -2770 100494
rect -2534 100258 -2450 100494
rect -2214 100258 -2130 100494
rect -1894 100258 1186 100494
rect 1422 100258 8186 100494
rect 8422 100258 15186 100494
rect 15422 100258 22186 100494
rect 22422 100258 29186 100494
rect 29422 100258 36186 100494
rect 36422 100258 43186 100494
rect 43422 100258 50186 100494
rect 50422 100258 57186 100494
rect 57422 100258 64186 100494
rect 64422 100258 71186 100494
rect 71422 100258 78186 100494
rect 78422 100258 85186 100494
rect 85422 100258 92186 100494
rect 92422 100258 99186 100494
rect 99422 100258 106186 100494
rect 106422 100258 113186 100494
rect 113422 100258 120186 100494
rect 120422 100258 127186 100494
rect 127422 100258 134186 100494
rect 134422 100258 141186 100494
rect 141422 100258 148186 100494
rect 148422 100258 155186 100494
rect 155422 100258 162186 100494
rect 162422 100258 169186 100494
rect 169422 100258 176186 100494
rect 176422 100258 183186 100494
rect 183422 100258 190186 100494
rect 190422 100258 197186 100494
rect 197422 100258 204186 100494
rect 204422 100258 211186 100494
rect 211422 100258 218186 100494
rect 218422 100258 225186 100494
rect 225422 100258 232186 100494
rect 232422 100258 239186 100494
rect 239422 100258 246186 100494
rect 246422 100258 253186 100494
rect 253422 100258 260186 100494
rect 260422 100258 267186 100494
rect 267422 100258 274186 100494
rect 274422 100258 281186 100494
rect 281422 100258 288186 100494
rect 288422 100258 295186 100494
rect 295422 100258 302186 100494
rect 302422 100258 309186 100494
rect 309422 100258 316186 100494
rect 316422 100258 323186 100494
rect 323422 100258 330186 100494
rect 330422 100258 337186 100494
rect 337422 100258 344186 100494
rect 344422 100258 351186 100494
rect 351422 100258 358186 100494
rect 358422 100258 365186 100494
rect 365422 100258 372186 100494
rect 372422 100258 379186 100494
rect 379422 100258 386186 100494
rect 386422 100258 393186 100494
rect 393422 100258 400186 100494
rect 400422 100258 407186 100494
rect 407422 100258 414186 100494
rect 414422 100258 421186 100494
rect 421422 100258 428186 100494
rect 428422 100258 435186 100494
rect 435422 100258 442186 100494
rect 442422 100258 449186 100494
rect 449422 100258 456186 100494
rect 456422 100258 463186 100494
rect 463422 100258 470186 100494
rect 470422 100258 477186 100494
rect 477422 100258 484186 100494
rect 484422 100258 491186 100494
rect 491422 100258 498186 100494
rect 498422 100258 505186 100494
rect 505422 100258 512186 100494
rect 512422 100258 519186 100494
rect 519422 100258 526186 100494
rect 526422 100258 533186 100494
rect 533422 100258 540186 100494
rect 540422 100258 547186 100494
rect 547422 100258 554186 100494
rect 554422 100258 561186 100494
rect 561422 100258 568186 100494
rect 568422 100258 575186 100494
rect 575422 100258 582186 100494
rect 582422 100258 585818 100494
rect 586054 100258 586138 100494
rect 586374 100258 586458 100494
rect 586694 100258 586778 100494
rect 587014 100258 588874 100494
rect -4950 100216 588874 100258
rect -4950 94434 588874 94476
rect -4950 94198 -4842 94434
rect -4606 94198 -4522 94434
rect -4286 94198 -4202 94434
rect -3966 94198 -3882 94434
rect -3646 94198 2918 94434
rect 3154 94198 9918 94434
rect 10154 94198 16918 94434
rect 17154 94198 23918 94434
rect 24154 94198 30918 94434
rect 31154 94198 37918 94434
rect 38154 94198 44918 94434
rect 45154 94198 51918 94434
rect 52154 94198 58918 94434
rect 59154 94198 65918 94434
rect 66154 94198 72918 94434
rect 73154 94198 79918 94434
rect 80154 94198 86918 94434
rect 87154 94198 93918 94434
rect 94154 94198 100918 94434
rect 101154 94198 107918 94434
rect 108154 94198 114918 94434
rect 115154 94198 121918 94434
rect 122154 94198 128918 94434
rect 129154 94198 135918 94434
rect 136154 94198 142918 94434
rect 143154 94198 149918 94434
rect 150154 94198 156918 94434
rect 157154 94198 163918 94434
rect 164154 94198 170918 94434
rect 171154 94198 177918 94434
rect 178154 94198 184918 94434
rect 185154 94198 191918 94434
rect 192154 94198 198918 94434
rect 199154 94198 205918 94434
rect 206154 94198 212918 94434
rect 213154 94198 219918 94434
rect 220154 94198 226918 94434
rect 227154 94198 233918 94434
rect 234154 94198 240918 94434
rect 241154 94198 247918 94434
rect 248154 94198 254918 94434
rect 255154 94198 261918 94434
rect 262154 94198 268918 94434
rect 269154 94198 275918 94434
rect 276154 94198 282918 94434
rect 283154 94198 289918 94434
rect 290154 94198 296918 94434
rect 297154 94198 303918 94434
rect 304154 94198 310918 94434
rect 311154 94198 317918 94434
rect 318154 94198 324918 94434
rect 325154 94198 331918 94434
rect 332154 94198 338918 94434
rect 339154 94198 345918 94434
rect 346154 94198 352918 94434
rect 353154 94198 359918 94434
rect 360154 94198 366918 94434
rect 367154 94198 373918 94434
rect 374154 94198 380918 94434
rect 381154 94198 387918 94434
rect 388154 94198 394918 94434
rect 395154 94198 401918 94434
rect 402154 94198 408918 94434
rect 409154 94198 415918 94434
rect 416154 94198 422918 94434
rect 423154 94198 429918 94434
rect 430154 94198 436918 94434
rect 437154 94198 443918 94434
rect 444154 94198 450918 94434
rect 451154 94198 457918 94434
rect 458154 94198 464918 94434
rect 465154 94198 471918 94434
rect 472154 94198 478918 94434
rect 479154 94198 485918 94434
rect 486154 94198 492918 94434
rect 493154 94198 499918 94434
rect 500154 94198 506918 94434
rect 507154 94198 513918 94434
rect 514154 94198 520918 94434
rect 521154 94198 527918 94434
rect 528154 94198 534918 94434
rect 535154 94198 541918 94434
rect 542154 94198 548918 94434
rect 549154 94198 555918 94434
rect 556154 94198 562918 94434
rect 563154 94198 569918 94434
rect 570154 94198 576918 94434
rect 577154 94198 587570 94434
rect 587806 94198 587890 94434
rect 588126 94198 588210 94434
rect 588446 94198 588530 94434
rect 588766 94198 588874 94434
rect -4950 94156 588874 94198
rect -4950 93494 588874 93536
rect -4950 93258 -3090 93494
rect -2854 93258 -2770 93494
rect -2534 93258 -2450 93494
rect -2214 93258 -2130 93494
rect -1894 93258 1186 93494
rect 1422 93258 8186 93494
rect 8422 93258 15186 93494
rect 15422 93258 22186 93494
rect 22422 93258 29186 93494
rect 29422 93258 36186 93494
rect 36422 93258 43186 93494
rect 43422 93258 50186 93494
rect 50422 93258 57186 93494
rect 57422 93258 64186 93494
rect 64422 93258 71186 93494
rect 71422 93258 78186 93494
rect 78422 93258 85186 93494
rect 85422 93258 92186 93494
rect 92422 93258 99186 93494
rect 99422 93258 106186 93494
rect 106422 93258 113186 93494
rect 113422 93258 120186 93494
rect 120422 93258 127186 93494
rect 127422 93258 134186 93494
rect 134422 93258 141186 93494
rect 141422 93258 148186 93494
rect 148422 93258 155186 93494
rect 155422 93258 162186 93494
rect 162422 93258 169186 93494
rect 169422 93258 176186 93494
rect 176422 93258 183186 93494
rect 183422 93258 190186 93494
rect 190422 93258 197186 93494
rect 197422 93258 204186 93494
rect 204422 93258 211186 93494
rect 211422 93258 218186 93494
rect 218422 93258 225186 93494
rect 225422 93258 232186 93494
rect 232422 93258 239186 93494
rect 239422 93258 246186 93494
rect 246422 93258 253186 93494
rect 253422 93258 260186 93494
rect 260422 93258 267186 93494
rect 267422 93258 274186 93494
rect 274422 93258 281186 93494
rect 281422 93258 288186 93494
rect 288422 93258 295186 93494
rect 295422 93258 302186 93494
rect 302422 93258 309186 93494
rect 309422 93258 316186 93494
rect 316422 93258 323186 93494
rect 323422 93258 330186 93494
rect 330422 93258 337186 93494
rect 337422 93258 344186 93494
rect 344422 93258 351186 93494
rect 351422 93258 358186 93494
rect 358422 93258 365186 93494
rect 365422 93258 372186 93494
rect 372422 93258 379186 93494
rect 379422 93258 386186 93494
rect 386422 93258 393186 93494
rect 393422 93258 400186 93494
rect 400422 93258 407186 93494
rect 407422 93258 414186 93494
rect 414422 93258 421186 93494
rect 421422 93258 428186 93494
rect 428422 93258 435186 93494
rect 435422 93258 442186 93494
rect 442422 93258 449186 93494
rect 449422 93258 456186 93494
rect 456422 93258 463186 93494
rect 463422 93258 470186 93494
rect 470422 93258 477186 93494
rect 477422 93258 484186 93494
rect 484422 93258 491186 93494
rect 491422 93258 498186 93494
rect 498422 93258 505186 93494
rect 505422 93258 512186 93494
rect 512422 93258 519186 93494
rect 519422 93258 526186 93494
rect 526422 93258 533186 93494
rect 533422 93258 540186 93494
rect 540422 93258 547186 93494
rect 547422 93258 554186 93494
rect 554422 93258 561186 93494
rect 561422 93258 568186 93494
rect 568422 93258 575186 93494
rect 575422 93258 582186 93494
rect 582422 93258 585818 93494
rect 586054 93258 586138 93494
rect 586374 93258 586458 93494
rect 586694 93258 586778 93494
rect 587014 93258 588874 93494
rect -4950 93216 588874 93258
rect -4950 87434 588874 87476
rect -4950 87198 -4842 87434
rect -4606 87198 -4522 87434
rect -4286 87198 -4202 87434
rect -3966 87198 -3882 87434
rect -3646 87198 2918 87434
rect 3154 87198 9918 87434
rect 10154 87198 16918 87434
rect 17154 87198 23918 87434
rect 24154 87198 30918 87434
rect 31154 87198 37918 87434
rect 38154 87198 44918 87434
rect 45154 87198 51918 87434
rect 52154 87198 58918 87434
rect 59154 87198 65918 87434
rect 66154 87198 72918 87434
rect 73154 87198 79918 87434
rect 80154 87198 86918 87434
rect 87154 87198 93918 87434
rect 94154 87198 100918 87434
rect 101154 87198 107918 87434
rect 108154 87198 114918 87434
rect 115154 87198 121918 87434
rect 122154 87198 128918 87434
rect 129154 87198 135918 87434
rect 136154 87198 142918 87434
rect 143154 87198 149918 87434
rect 150154 87198 156918 87434
rect 157154 87198 163918 87434
rect 164154 87198 170918 87434
rect 171154 87198 177918 87434
rect 178154 87198 184918 87434
rect 185154 87198 191918 87434
rect 192154 87198 198918 87434
rect 199154 87198 205918 87434
rect 206154 87198 212918 87434
rect 213154 87198 219918 87434
rect 220154 87198 226918 87434
rect 227154 87198 233918 87434
rect 234154 87198 240918 87434
rect 241154 87198 247918 87434
rect 248154 87198 254918 87434
rect 255154 87198 261918 87434
rect 262154 87198 268918 87434
rect 269154 87198 275918 87434
rect 276154 87198 282918 87434
rect 283154 87198 289918 87434
rect 290154 87198 296918 87434
rect 297154 87198 303918 87434
rect 304154 87198 310918 87434
rect 311154 87198 317918 87434
rect 318154 87198 324918 87434
rect 325154 87198 331918 87434
rect 332154 87198 338918 87434
rect 339154 87198 345918 87434
rect 346154 87198 352918 87434
rect 353154 87198 359918 87434
rect 360154 87198 366918 87434
rect 367154 87198 373918 87434
rect 374154 87198 380918 87434
rect 381154 87198 387918 87434
rect 388154 87198 394918 87434
rect 395154 87198 401918 87434
rect 402154 87198 408918 87434
rect 409154 87198 415918 87434
rect 416154 87198 422918 87434
rect 423154 87198 429918 87434
rect 430154 87198 436918 87434
rect 437154 87198 443918 87434
rect 444154 87198 450918 87434
rect 451154 87198 457918 87434
rect 458154 87198 464918 87434
rect 465154 87198 471918 87434
rect 472154 87198 478918 87434
rect 479154 87198 485918 87434
rect 486154 87198 492918 87434
rect 493154 87198 499918 87434
rect 500154 87198 506918 87434
rect 507154 87198 513918 87434
rect 514154 87198 520918 87434
rect 521154 87198 527918 87434
rect 528154 87198 534918 87434
rect 535154 87198 541918 87434
rect 542154 87198 548918 87434
rect 549154 87198 555918 87434
rect 556154 87198 562918 87434
rect 563154 87198 569918 87434
rect 570154 87198 576918 87434
rect 577154 87198 587570 87434
rect 587806 87198 587890 87434
rect 588126 87198 588210 87434
rect 588446 87198 588530 87434
rect 588766 87198 588874 87434
rect -4950 87156 588874 87198
rect -4950 86494 588874 86536
rect -4950 86258 -3090 86494
rect -2854 86258 -2770 86494
rect -2534 86258 -2450 86494
rect -2214 86258 -2130 86494
rect -1894 86258 1186 86494
rect 1422 86258 8186 86494
rect 8422 86258 15186 86494
rect 15422 86258 22186 86494
rect 22422 86258 29186 86494
rect 29422 86258 36186 86494
rect 36422 86258 43186 86494
rect 43422 86258 50186 86494
rect 50422 86258 57186 86494
rect 57422 86258 64186 86494
rect 64422 86258 71186 86494
rect 71422 86258 78186 86494
rect 78422 86258 85186 86494
rect 85422 86258 92186 86494
rect 92422 86258 99186 86494
rect 99422 86258 106186 86494
rect 106422 86258 113186 86494
rect 113422 86258 120186 86494
rect 120422 86258 127186 86494
rect 127422 86258 134186 86494
rect 134422 86258 141186 86494
rect 141422 86258 148186 86494
rect 148422 86258 155186 86494
rect 155422 86258 162186 86494
rect 162422 86258 169186 86494
rect 169422 86258 176186 86494
rect 176422 86258 183186 86494
rect 183422 86258 190186 86494
rect 190422 86258 197186 86494
rect 197422 86258 204186 86494
rect 204422 86258 211186 86494
rect 211422 86258 218186 86494
rect 218422 86258 225186 86494
rect 225422 86258 232186 86494
rect 232422 86258 239186 86494
rect 239422 86258 246186 86494
rect 246422 86258 253186 86494
rect 253422 86258 260186 86494
rect 260422 86258 267186 86494
rect 267422 86258 274186 86494
rect 274422 86258 281186 86494
rect 281422 86258 288186 86494
rect 288422 86258 295186 86494
rect 295422 86258 302186 86494
rect 302422 86258 309186 86494
rect 309422 86258 316186 86494
rect 316422 86258 323186 86494
rect 323422 86258 330186 86494
rect 330422 86258 337186 86494
rect 337422 86258 344186 86494
rect 344422 86258 351186 86494
rect 351422 86258 358186 86494
rect 358422 86258 365186 86494
rect 365422 86258 372186 86494
rect 372422 86258 379186 86494
rect 379422 86258 386186 86494
rect 386422 86258 393186 86494
rect 393422 86258 400186 86494
rect 400422 86258 407186 86494
rect 407422 86258 414186 86494
rect 414422 86258 421186 86494
rect 421422 86258 428186 86494
rect 428422 86258 435186 86494
rect 435422 86258 442186 86494
rect 442422 86258 449186 86494
rect 449422 86258 456186 86494
rect 456422 86258 463186 86494
rect 463422 86258 470186 86494
rect 470422 86258 477186 86494
rect 477422 86258 484186 86494
rect 484422 86258 491186 86494
rect 491422 86258 498186 86494
rect 498422 86258 505186 86494
rect 505422 86258 512186 86494
rect 512422 86258 519186 86494
rect 519422 86258 526186 86494
rect 526422 86258 533186 86494
rect 533422 86258 540186 86494
rect 540422 86258 547186 86494
rect 547422 86258 554186 86494
rect 554422 86258 561186 86494
rect 561422 86258 568186 86494
rect 568422 86258 575186 86494
rect 575422 86258 582186 86494
rect 582422 86258 585818 86494
rect 586054 86258 586138 86494
rect 586374 86258 586458 86494
rect 586694 86258 586778 86494
rect 587014 86258 588874 86494
rect -4950 86216 588874 86258
rect -4950 80434 588874 80476
rect -4950 80198 -4842 80434
rect -4606 80198 -4522 80434
rect -4286 80198 -4202 80434
rect -3966 80198 -3882 80434
rect -3646 80198 2918 80434
rect 3154 80198 9918 80434
rect 10154 80198 16918 80434
rect 17154 80198 23918 80434
rect 24154 80198 30918 80434
rect 31154 80198 37918 80434
rect 38154 80198 44918 80434
rect 45154 80198 51918 80434
rect 52154 80198 58918 80434
rect 59154 80198 65918 80434
rect 66154 80198 72918 80434
rect 73154 80198 79918 80434
rect 80154 80198 86918 80434
rect 87154 80198 93918 80434
rect 94154 80198 100918 80434
rect 101154 80198 107918 80434
rect 108154 80198 114918 80434
rect 115154 80198 121918 80434
rect 122154 80198 128918 80434
rect 129154 80198 135918 80434
rect 136154 80198 142918 80434
rect 143154 80198 149918 80434
rect 150154 80198 156918 80434
rect 157154 80198 163918 80434
rect 164154 80198 170918 80434
rect 171154 80198 177918 80434
rect 178154 80198 184918 80434
rect 185154 80198 191918 80434
rect 192154 80198 198918 80434
rect 199154 80198 205918 80434
rect 206154 80198 212918 80434
rect 213154 80198 219918 80434
rect 220154 80198 226918 80434
rect 227154 80198 233918 80434
rect 234154 80198 240918 80434
rect 241154 80198 247918 80434
rect 248154 80198 254918 80434
rect 255154 80198 261918 80434
rect 262154 80198 268918 80434
rect 269154 80198 275918 80434
rect 276154 80198 282918 80434
rect 283154 80198 289918 80434
rect 290154 80198 296918 80434
rect 297154 80198 303918 80434
rect 304154 80198 310918 80434
rect 311154 80198 317918 80434
rect 318154 80198 324918 80434
rect 325154 80198 331918 80434
rect 332154 80198 338918 80434
rect 339154 80198 345918 80434
rect 346154 80198 352918 80434
rect 353154 80198 359918 80434
rect 360154 80198 366918 80434
rect 367154 80198 373918 80434
rect 374154 80198 380918 80434
rect 381154 80198 387918 80434
rect 388154 80198 394918 80434
rect 395154 80198 401918 80434
rect 402154 80198 408918 80434
rect 409154 80198 415918 80434
rect 416154 80198 422918 80434
rect 423154 80198 429918 80434
rect 430154 80198 436918 80434
rect 437154 80198 443918 80434
rect 444154 80198 450918 80434
rect 451154 80198 457918 80434
rect 458154 80198 464918 80434
rect 465154 80198 471918 80434
rect 472154 80198 478918 80434
rect 479154 80198 485918 80434
rect 486154 80198 492918 80434
rect 493154 80198 499918 80434
rect 500154 80198 506918 80434
rect 507154 80198 513918 80434
rect 514154 80198 520918 80434
rect 521154 80198 527918 80434
rect 528154 80198 534918 80434
rect 535154 80198 541918 80434
rect 542154 80198 548918 80434
rect 549154 80198 555918 80434
rect 556154 80198 562918 80434
rect 563154 80198 569918 80434
rect 570154 80198 576918 80434
rect 577154 80198 587570 80434
rect 587806 80198 587890 80434
rect 588126 80198 588210 80434
rect 588446 80198 588530 80434
rect 588766 80198 588874 80434
rect -4950 80156 588874 80198
rect -4950 79494 588874 79536
rect -4950 79258 -3090 79494
rect -2854 79258 -2770 79494
rect -2534 79258 -2450 79494
rect -2214 79258 -2130 79494
rect -1894 79258 1186 79494
rect 1422 79258 8186 79494
rect 8422 79258 15186 79494
rect 15422 79258 22186 79494
rect 22422 79258 29186 79494
rect 29422 79258 36186 79494
rect 36422 79258 43186 79494
rect 43422 79258 50186 79494
rect 50422 79258 57186 79494
rect 57422 79258 64186 79494
rect 64422 79258 71186 79494
rect 71422 79258 78186 79494
rect 78422 79258 85186 79494
rect 85422 79258 92186 79494
rect 92422 79258 99186 79494
rect 99422 79258 106186 79494
rect 106422 79258 113186 79494
rect 113422 79258 120186 79494
rect 120422 79258 127186 79494
rect 127422 79258 134186 79494
rect 134422 79258 141186 79494
rect 141422 79258 148186 79494
rect 148422 79258 155186 79494
rect 155422 79258 162186 79494
rect 162422 79258 169186 79494
rect 169422 79258 176186 79494
rect 176422 79258 183186 79494
rect 183422 79258 190186 79494
rect 190422 79258 197186 79494
rect 197422 79258 204186 79494
rect 204422 79258 211186 79494
rect 211422 79258 218186 79494
rect 218422 79258 225186 79494
rect 225422 79258 232186 79494
rect 232422 79258 239186 79494
rect 239422 79258 246186 79494
rect 246422 79258 253186 79494
rect 253422 79258 260186 79494
rect 260422 79258 267186 79494
rect 267422 79258 274186 79494
rect 274422 79258 281186 79494
rect 281422 79258 288186 79494
rect 288422 79258 295186 79494
rect 295422 79258 302186 79494
rect 302422 79258 309186 79494
rect 309422 79258 316186 79494
rect 316422 79258 323186 79494
rect 323422 79258 330186 79494
rect 330422 79258 337186 79494
rect 337422 79258 344186 79494
rect 344422 79258 351186 79494
rect 351422 79258 358186 79494
rect 358422 79258 365186 79494
rect 365422 79258 372186 79494
rect 372422 79258 379186 79494
rect 379422 79258 386186 79494
rect 386422 79258 393186 79494
rect 393422 79258 400186 79494
rect 400422 79258 407186 79494
rect 407422 79258 414186 79494
rect 414422 79258 421186 79494
rect 421422 79258 428186 79494
rect 428422 79258 435186 79494
rect 435422 79258 442186 79494
rect 442422 79258 449186 79494
rect 449422 79258 456186 79494
rect 456422 79258 463186 79494
rect 463422 79258 470186 79494
rect 470422 79258 477186 79494
rect 477422 79258 484186 79494
rect 484422 79258 491186 79494
rect 491422 79258 498186 79494
rect 498422 79258 505186 79494
rect 505422 79258 512186 79494
rect 512422 79258 519186 79494
rect 519422 79258 526186 79494
rect 526422 79258 533186 79494
rect 533422 79258 540186 79494
rect 540422 79258 547186 79494
rect 547422 79258 554186 79494
rect 554422 79258 561186 79494
rect 561422 79258 568186 79494
rect 568422 79258 575186 79494
rect 575422 79258 582186 79494
rect 582422 79258 585818 79494
rect 586054 79258 586138 79494
rect 586374 79258 586458 79494
rect 586694 79258 586778 79494
rect 587014 79258 588874 79494
rect -4950 79216 588874 79258
rect -4950 73434 588874 73476
rect -4950 73198 -4842 73434
rect -4606 73198 -4522 73434
rect -4286 73198 -4202 73434
rect -3966 73198 -3882 73434
rect -3646 73198 2918 73434
rect 3154 73198 9918 73434
rect 10154 73198 16918 73434
rect 17154 73198 23918 73434
rect 24154 73198 30918 73434
rect 31154 73198 37918 73434
rect 38154 73198 44918 73434
rect 45154 73198 51918 73434
rect 52154 73198 58918 73434
rect 59154 73198 65918 73434
rect 66154 73198 72918 73434
rect 73154 73198 79918 73434
rect 80154 73198 86918 73434
rect 87154 73198 93918 73434
rect 94154 73198 100918 73434
rect 101154 73198 107918 73434
rect 108154 73198 114918 73434
rect 115154 73198 121918 73434
rect 122154 73198 128918 73434
rect 129154 73198 135918 73434
rect 136154 73198 142918 73434
rect 143154 73198 149918 73434
rect 150154 73198 156918 73434
rect 157154 73198 163918 73434
rect 164154 73198 170918 73434
rect 171154 73198 177918 73434
rect 178154 73198 184918 73434
rect 185154 73198 191918 73434
rect 192154 73198 198918 73434
rect 199154 73198 205918 73434
rect 206154 73198 212918 73434
rect 213154 73198 219918 73434
rect 220154 73198 226918 73434
rect 227154 73198 233918 73434
rect 234154 73198 240918 73434
rect 241154 73198 247918 73434
rect 248154 73198 254918 73434
rect 255154 73198 261918 73434
rect 262154 73198 268918 73434
rect 269154 73198 275918 73434
rect 276154 73198 282918 73434
rect 283154 73198 289918 73434
rect 290154 73198 296918 73434
rect 297154 73198 303918 73434
rect 304154 73198 310918 73434
rect 311154 73198 317918 73434
rect 318154 73198 324918 73434
rect 325154 73198 331918 73434
rect 332154 73198 338918 73434
rect 339154 73198 345918 73434
rect 346154 73198 352918 73434
rect 353154 73198 359918 73434
rect 360154 73198 366918 73434
rect 367154 73198 373918 73434
rect 374154 73198 380918 73434
rect 381154 73198 387918 73434
rect 388154 73198 394918 73434
rect 395154 73198 401918 73434
rect 402154 73198 408918 73434
rect 409154 73198 415918 73434
rect 416154 73198 422918 73434
rect 423154 73198 429918 73434
rect 430154 73198 436918 73434
rect 437154 73198 443918 73434
rect 444154 73198 450918 73434
rect 451154 73198 457918 73434
rect 458154 73198 464918 73434
rect 465154 73198 471918 73434
rect 472154 73198 478918 73434
rect 479154 73198 485918 73434
rect 486154 73198 492918 73434
rect 493154 73198 499918 73434
rect 500154 73198 506918 73434
rect 507154 73198 513918 73434
rect 514154 73198 520918 73434
rect 521154 73198 527918 73434
rect 528154 73198 534918 73434
rect 535154 73198 541918 73434
rect 542154 73198 548918 73434
rect 549154 73198 555918 73434
rect 556154 73198 562918 73434
rect 563154 73198 569918 73434
rect 570154 73198 576918 73434
rect 577154 73198 587570 73434
rect 587806 73198 587890 73434
rect 588126 73198 588210 73434
rect 588446 73198 588530 73434
rect 588766 73198 588874 73434
rect -4950 73156 588874 73198
rect -4950 72494 588874 72536
rect -4950 72258 -3090 72494
rect -2854 72258 -2770 72494
rect -2534 72258 -2450 72494
rect -2214 72258 -2130 72494
rect -1894 72258 1186 72494
rect 1422 72258 8186 72494
rect 8422 72258 15186 72494
rect 15422 72258 22186 72494
rect 22422 72258 29186 72494
rect 29422 72258 36186 72494
rect 36422 72258 43186 72494
rect 43422 72258 50186 72494
rect 50422 72258 57186 72494
rect 57422 72258 64186 72494
rect 64422 72258 71186 72494
rect 71422 72258 78186 72494
rect 78422 72258 85186 72494
rect 85422 72258 92186 72494
rect 92422 72258 99186 72494
rect 99422 72258 106186 72494
rect 106422 72258 113186 72494
rect 113422 72258 120186 72494
rect 120422 72258 127186 72494
rect 127422 72258 134186 72494
rect 134422 72258 141186 72494
rect 141422 72258 148186 72494
rect 148422 72258 155186 72494
rect 155422 72258 162186 72494
rect 162422 72258 169186 72494
rect 169422 72258 176186 72494
rect 176422 72258 183186 72494
rect 183422 72258 190186 72494
rect 190422 72258 197186 72494
rect 197422 72258 204186 72494
rect 204422 72258 211186 72494
rect 211422 72258 218186 72494
rect 218422 72258 225186 72494
rect 225422 72258 232186 72494
rect 232422 72258 239186 72494
rect 239422 72258 246186 72494
rect 246422 72258 253186 72494
rect 253422 72258 260186 72494
rect 260422 72258 267186 72494
rect 267422 72258 274186 72494
rect 274422 72258 281186 72494
rect 281422 72258 288186 72494
rect 288422 72258 295186 72494
rect 295422 72258 302186 72494
rect 302422 72258 309186 72494
rect 309422 72258 316186 72494
rect 316422 72258 323186 72494
rect 323422 72258 330186 72494
rect 330422 72258 337186 72494
rect 337422 72258 344186 72494
rect 344422 72258 351186 72494
rect 351422 72258 358186 72494
rect 358422 72258 365186 72494
rect 365422 72258 372186 72494
rect 372422 72258 379186 72494
rect 379422 72258 386186 72494
rect 386422 72258 393186 72494
rect 393422 72258 400186 72494
rect 400422 72258 407186 72494
rect 407422 72258 414186 72494
rect 414422 72258 421186 72494
rect 421422 72258 428186 72494
rect 428422 72258 435186 72494
rect 435422 72258 442186 72494
rect 442422 72258 449186 72494
rect 449422 72258 456186 72494
rect 456422 72258 463186 72494
rect 463422 72258 470186 72494
rect 470422 72258 477186 72494
rect 477422 72258 484186 72494
rect 484422 72258 491186 72494
rect 491422 72258 498186 72494
rect 498422 72258 505186 72494
rect 505422 72258 512186 72494
rect 512422 72258 519186 72494
rect 519422 72258 526186 72494
rect 526422 72258 533186 72494
rect 533422 72258 540186 72494
rect 540422 72258 547186 72494
rect 547422 72258 554186 72494
rect 554422 72258 561186 72494
rect 561422 72258 568186 72494
rect 568422 72258 575186 72494
rect 575422 72258 582186 72494
rect 582422 72258 585818 72494
rect 586054 72258 586138 72494
rect 586374 72258 586458 72494
rect 586694 72258 586778 72494
rect 587014 72258 588874 72494
rect -4950 72216 588874 72258
rect -4950 66434 588874 66476
rect -4950 66198 -4842 66434
rect -4606 66198 -4522 66434
rect -4286 66198 -4202 66434
rect -3966 66198 -3882 66434
rect -3646 66198 2918 66434
rect 3154 66198 9918 66434
rect 10154 66198 16918 66434
rect 17154 66198 23918 66434
rect 24154 66198 30918 66434
rect 31154 66198 37918 66434
rect 38154 66198 44918 66434
rect 45154 66198 51918 66434
rect 52154 66198 58918 66434
rect 59154 66198 65918 66434
rect 66154 66198 72918 66434
rect 73154 66198 79918 66434
rect 80154 66198 86918 66434
rect 87154 66198 93918 66434
rect 94154 66198 100918 66434
rect 101154 66198 107918 66434
rect 108154 66198 114918 66434
rect 115154 66198 121918 66434
rect 122154 66198 128918 66434
rect 129154 66198 135918 66434
rect 136154 66198 142918 66434
rect 143154 66198 149918 66434
rect 150154 66198 156918 66434
rect 157154 66198 163918 66434
rect 164154 66198 170918 66434
rect 171154 66198 177918 66434
rect 178154 66198 184918 66434
rect 185154 66198 191918 66434
rect 192154 66198 198918 66434
rect 199154 66198 205918 66434
rect 206154 66198 212918 66434
rect 213154 66198 219918 66434
rect 220154 66198 226918 66434
rect 227154 66198 233918 66434
rect 234154 66198 240918 66434
rect 241154 66198 247918 66434
rect 248154 66198 254918 66434
rect 255154 66198 261918 66434
rect 262154 66198 268918 66434
rect 269154 66198 275918 66434
rect 276154 66198 282918 66434
rect 283154 66198 289918 66434
rect 290154 66198 296918 66434
rect 297154 66198 303918 66434
rect 304154 66198 310918 66434
rect 311154 66198 317918 66434
rect 318154 66198 324918 66434
rect 325154 66198 331918 66434
rect 332154 66198 338918 66434
rect 339154 66198 345918 66434
rect 346154 66198 352918 66434
rect 353154 66198 359918 66434
rect 360154 66198 366918 66434
rect 367154 66198 373918 66434
rect 374154 66198 380918 66434
rect 381154 66198 387918 66434
rect 388154 66198 394918 66434
rect 395154 66198 401918 66434
rect 402154 66198 408918 66434
rect 409154 66198 415918 66434
rect 416154 66198 422918 66434
rect 423154 66198 429918 66434
rect 430154 66198 436918 66434
rect 437154 66198 443918 66434
rect 444154 66198 450918 66434
rect 451154 66198 457918 66434
rect 458154 66198 464918 66434
rect 465154 66198 471918 66434
rect 472154 66198 478918 66434
rect 479154 66198 485918 66434
rect 486154 66198 492918 66434
rect 493154 66198 499918 66434
rect 500154 66198 506918 66434
rect 507154 66198 513918 66434
rect 514154 66198 520918 66434
rect 521154 66198 527918 66434
rect 528154 66198 534918 66434
rect 535154 66198 541918 66434
rect 542154 66198 548918 66434
rect 549154 66198 555918 66434
rect 556154 66198 562918 66434
rect 563154 66198 569918 66434
rect 570154 66198 576918 66434
rect 577154 66198 587570 66434
rect 587806 66198 587890 66434
rect 588126 66198 588210 66434
rect 588446 66198 588530 66434
rect 588766 66198 588874 66434
rect -4950 66156 588874 66198
rect -4950 65494 588874 65536
rect -4950 65258 -3090 65494
rect -2854 65258 -2770 65494
rect -2534 65258 -2450 65494
rect -2214 65258 -2130 65494
rect -1894 65258 1186 65494
rect 1422 65258 8186 65494
rect 8422 65258 15186 65494
rect 15422 65258 22186 65494
rect 22422 65258 29186 65494
rect 29422 65258 36186 65494
rect 36422 65258 43186 65494
rect 43422 65258 50186 65494
rect 50422 65258 57186 65494
rect 57422 65258 64186 65494
rect 64422 65258 71186 65494
rect 71422 65258 78186 65494
rect 78422 65258 85186 65494
rect 85422 65258 92186 65494
rect 92422 65258 99186 65494
rect 99422 65258 106186 65494
rect 106422 65258 113186 65494
rect 113422 65258 120186 65494
rect 120422 65258 127186 65494
rect 127422 65258 134186 65494
rect 134422 65258 141186 65494
rect 141422 65258 148186 65494
rect 148422 65258 155186 65494
rect 155422 65258 162186 65494
rect 162422 65258 169186 65494
rect 169422 65258 176186 65494
rect 176422 65258 183186 65494
rect 183422 65258 190186 65494
rect 190422 65258 197186 65494
rect 197422 65258 204186 65494
rect 204422 65258 211186 65494
rect 211422 65258 218186 65494
rect 218422 65258 225186 65494
rect 225422 65258 232186 65494
rect 232422 65258 239186 65494
rect 239422 65258 246186 65494
rect 246422 65258 253186 65494
rect 253422 65258 260186 65494
rect 260422 65258 267186 65494
rect 267422 65258 274186 65494
rect 274422 65258 281186 65494
rect 281422 65258 288186 65494
rect 288422 65258 295186 65494
rect 295422 65258 302186 65494
rect 302422 65258 309186 65494
rect 309422 65258 316186 65494
rect 316422 65258 323186 65494
rect 323422 65258 330186 65494
rect 330422 65258 337186 65494
rect 337422 65258 344186 65494
rect 344422 65258 351186 65494
rect 351422 65258 358186 65494
rect 358422 65258 365186 65494
rect 365422 65258 372186 65494
rect 372422 65258 379186 65494
rect 379422 65258 386186 65494
rect 386422 65258 393186 65494
rect 393422 65258 400186 65494
rect 400422 65258 407186 65494
rect 407422 65258 414186 65494
rect 414422 65258 421186 65494
rect 421422 65258 428186 65494
rect 428422 65258 435186 65494
rect 435422 65258 442186 65494
rect 442422 65258 449186 65494
rect 449422 65258 456186 65494
rect 456422 65258 463186 65494
rect 463422 65258 470186 65494
rect 470422 65258 477186 65494
rect 477422 65258 484186 65494
rect 484422 65258 491186 65494
rect 491422 65258 498186 65494
rect 498422 65258 505186 65494
rect 505422 65258 512186 65494
rect 512422 65258 519186 65494
rect 519422 65258 526186 65494
rect 526422 65258 533186 65494
rect 533422 65258 540186 65494
rect 540422 65258 547186 65494
rect 547422 65258 554186 65494
rect 554422 65258 561186 65494
rect 561422 65258 568186 65494
rect 568422 65258 575186 65494
rect 575422 65258 582186 65494
rect 582422 65258 585818 65494
rect 586054 65258 586138 65494
rect 586374 65258 586458 65494
rect 586694 65258 586778 65494
rect 587014 65258 588874 65494
rect -4950 65216 588874 65258
rect -4950 59434 588874 59476
rect -4950 59198 -4842 59434
rect -4606 59198 -4522 59434
rect -4286 59198 -4202 59434
rect -3966 59198 -3882 59434
rect -3646 59198 2918 59434
rect 3154 59198 9918 59434
rect 10154 59198 16918 59434
rect 17154 59198 23918 59434
rect 24154 59198 30918 59434
rect 31154 59198 37918 59434
rect 38154 59198 44918 59434
rect 45154 59198 51918 59434
rect 52154 59198 58918 59434
rect 59154 59198 65918 59434
rect 66154 59198 72918 59434
rect 73154 59198 79918 59434
rect 80154 59198 86918 59434
rect 87154 59198 93918 59434
rect 94154 59198 100918 59434
rect 101154 59198 107918 59434
rect 108154 59198 114918 59434
rect 115154 59198 121918 59434
rect 122154 59198 128918 59434
rect 129154 59198 135918 59434
rect 136154 59198 142918 59434
rect 143154 59198 149918 59434
rect 150154 59198 156918 59434
rect 157154 59198 163918 59434
rect 164154 59198 170918 59434
rect 171154 59198 177918 59434
rect 178154 59198 184918 59434
rect 185154 59198 191918 59434
rect 192154 59198 198918 59434
rect 199154 59198 205918 59434
rect 206154 59198 212918 59434
rect 213154 59198 219918 59434
rect 220154 59198 226918 59434
rect 227154 59198 233918 59434
rect 234154 59198 240918 59434
rect 241154 59198 247918 59434
rect 248154 59198 254918 59434
rect 255154 59198 261918 59434
rect 262154 59198 268918 59434
rect 269154 59198 275918 59434
rect 276154 59198 282918 59434
rect 283154 59198 289918 59434
rect 290154 59198 296918 59434
rect 297154 59198 303918 59434
rect 304154 59198 310918 59434
rect 311154 59198 317918 59434
rect 318154 59198 324918 59434
rect 325154 59198 331918 59434
rect 332154 59198 338918 59434
rect 339154 59198 345918 59434
rect 346154 59198 352918 59434
rect 353154 59198 359918 59434
rect 360154 59198 366918 59434
rect 367154 59198 373918 59434
rect 374154 59198 380918 59434
rect 381154 59198 387918 59434
rect 388154 59198 394918 59434
rect 395154 59198 401918 59434
rect 402154 59198 408918 59434
rect 409154 59198 415918 59434
rect 416154 59198 422918 59434
rect 423154 59198 429918 59434
rect 430154 59198 436918 59434
rect 437154 59198 443918 59434
rect 444154 59198 450918 59434
rect 451154 59198 457918 59434
rect 458154 59198 464918 59434
rect 465154 59198 471918 59434
rect 472154 59198 478918 59434
rect 479154 59198 485918 59434
rect 486154 59198 492918 59434
rect 493154 59198 499918 59434
rect 500154 59198 506918 59434
rect 507154 59198 513918 59434
rect 514154 59198 520918 59434
rect 521154 59198 527918 59434
rect 528154 59198 534918 59434
rect 535154 59198 541918 59434
rect 542154 59198 548918 59434
rect 549154 59198 555918 59434
rect 556154 59198 562918 59434
rect 563154 59198 569918 59434
rect 570154 59198 576918 59434
rect 577154 59198 587570 59434
rect 587806 59198 587890 59434
rect 588126 59198 588210 59434
rect 588446 59198 588530 59434
rect 588766 59198 588874 59434
rect -4950 59156 588874 59198
rect -4950 58494 588874 58536
rect -4950 58258 -3090 58494
rect -2854 58258 -2770 58494
rect -2534 58258 -2450 58494
rect -2214 58258 -2130 58494
rect -1894 58258 1186 58494
rect 1422 58258 8186 58494
rect 8422 58258 15186 58494
rect 15422 58258 22186 58494
rect 22422 58258 29186 58494
rect 29422 58258 36186 58494
rect 36422 58258 43186 58494
rect 43422 58258 50186 58494
rect 50422 58258 57186 58494
rect 57422 58258 64186 58494
rect 64422 58258 71186 58494
rect 71422 58258 78186 58494
rect 78422 58258 85186 58494
rect 85422 58258 92186 58494
rect 92422 58258 99186 58494
rect 99422 58258 106186 58494
rect 106422 58258 113186 58494
rect 113422 58258 120186 58494
rect 120422 58258 127186 58494
rect 127422 58258 134186 58494
rect 134422 58258 141186 58494
rect 141422 58258 148186 58494
rect 148422 58258 155186 58494
rect 155422 58258 162186 58494
rect 162422 58258 169186 58494
rect 169422 58258 176186 58494
rect 176422 58258 183186 58494
rect 183422 58258 190186 58494
rect 190422 58258 197186 58494
rect 197422 58258 204186 58494
rect 204422 58258 211186 58494
rect 211422 58258 218186 58494
rect 218422 58258 225186 58494
rect 225422 58258 232186 58494
rect 232422 58258 239186 58494
rect 239422 58258 246186 58494
rect 246422 58258 253186 58494
rect 253422 58258 260186 58494
rect 260422 58258 267186 58494
rect 267422 58258 274186 58494
rect 274422 58258 281186 58494
rect 281422 58258 288186 58494
rect 288422 58258 295186 58494
rect 295422 58258 302186 58494
rect 302422 58258 309186 58494
rect 309422 58258 316186 58494
rect 316422 58258 323186 58494
rect 323422 58258 330186 58494
rect 330422 58258 337186 58494
rect 337422 58258 344186 58494
rect 344422 58258 351186 58494
rect 351422 58258 358186 58494
rect 358422 58258 365186 58494
rect 365422 58258 372186 58494
rect 372422 58258 379186 58494
rect 379422 58258 386186 58494
rect 386422 58258 393186 58494
rect 393422 58258 400186 58494
rect 400422 58258 407186 58494
rect 407422 58258 414186 58494
rect 414422 58258 421186 58494
rect 421422 58258 428186 58494
rect 428422 58258 435186 58494
rect 435422 58258 442186 58494
rect 442422 58258 449186 58494
rect 449422 58258 456186 58494
rect 456422 58258 463186 58494
rect 463422 58258 470186 58494
rect 470422 58258 477186 58494
rect 477422 58258 484186 58494
rect 484422 58258 491186 58494
rect 491422 58258 498186 58494
rect 498422 58258 505186 58494
rect 505422 58258 512186 58494
rect 512422 58258 519186 58494
rect 519422 58258 526186 58494
rect 526422 58258 533186 58494
rect 533422 58258 540186 58494
rect 540422 58258 547186 58494
rect 547422 58258 554186 58494
rect 554422 58258 561186 58494
rect 561422 58258 568186 58494
rect 568422 58258 575186 58494
rect 575422 58258 582186 58494
rect 582422 58258 585818 58494
rect 586054 58258 586138 58494
rect 586374 58258 586458 58494
rect 586694 58258 586778 58494
rect 587014 58258 588874 58494
rect -4950 58216 588874 58258
rect -4950 52434 588874 52476
rect -4950 52198 -4842 52434
rect -4606 52198 -4522 52434
rect -4286 52198 -4202 52434
rect -3966 52198 -3882 52434
rect -3646 52198 2918 52434
rect 3154 52198 9918 52434
rect 10154 52198 16918 52434
rect 17154 52198 23918 52434
rect 24154 52198 30918 52434
rect 31154 52198 37918 52434
rect 38154 52198 44918 52434
rect 45154 52198 51918 52434
rect 52154 52198 58918 52434
rect 59154 52198 65918 52434
rect 66154 52198 72918 52434
rect 73154 52198 79918 52434
rect 80154 52198 86918 52434
rect 87154 52198 93918 52434
rect 94154 52198 100918 52434
rect 101154 52198 107918 52434
rect 108154 52198 114918 52434
rect 115154 52198 121918 52434
rect 122154 52198 128918 52434
rect 129154 52198 135918 52434
rect 136154 52198 142918 52434
rect 143154 52198 149918 52434
rect 150154 52198 156918 52434
rect 157154 52198 163918 52434
rect 164154 52198 170918 52434
rect 171154 52198 177918 52434
rect 178154 52198 184918 52434
rect 185154 52198 191918 52434
rect 192154 52198 198918 52434
rect 199154 52198 205918 52434
rect 206154 52198 212918 52434
rect 213154 52198 219918 52434
rect 220154 52198 226918 52434
rect 227154 52198 233918 52434
rect 234154 52198 240918 52434
rect 241154 52198 247918 52434
rect 248154 52198 254918 52434
rect 255154 52198 261918 52434
rect 262154 52198 268918 52434
rect 269154 52198 275918 52434
rect 276154 52198 282918 52434
rect 283154 52198 289918 52434
rect 290154 52198 296918 52434
rect 297154 52198 303918 52434
rect 304154 52198 310918 52434
rect 311154 52198 317918 52434
rect 318154 52198 324918 52434
rect 325154 52198 331918 52434
rect 332154 52198 338918 52434
rect 339154 52198 345918 52434
rect 346154 52198 352918 52434
rect 353154 52198 359918 52434
rect 360154 52198 366918 52434
rect 367154 52198 373918 52434
rect 374154 52198 380918 52434
rect 381154 52198 387918 52434
rect 388154 52198 394918 52434
rect 395154 52198 401918 52434
rect 402154 52198 408918 52434
rect 409154 52198 415918 52434
rect 416154 52198 422918 52434
rect 423154 52198 429918 52434
rect 430154 52198 436918 52434
rect 437154 52198 443918 52434
rect 444154 52198 450918 52434
rect 451154 52198 457918 52434
rect 458154 52198 464918 52434
rect 465154 52198 471918 52434
rect 472154 52198 478918 52434
rect 479154 52198 485918 52434
rect 486154 52198 492918 52434
rect 493154 52198 499918 52434
rect 500154 52198 506918 52434
rect 507154 52198 513918 52434
rect 514154 52198 520918 52434
rect 521154 52198 527918 52434
rect 528154 52198 534918 52434
rect 535154 52198 541918 52434
rect 542154 52198 548918 52434
rect 549154 52198 555918 52434
rect 556154 52198 562918 52434
rect 563154 52198 569918 52434
rect 570154 52198 576918 52434
rect 577154 52198 587570 52434
rect 587806 52198 587890 52434
rect 588126 52198 588210 52434
rect 588446 52198 588530 52434
rect 588766 52198 588874 52434
rect -4950 52156 588874 52198
rect -4950 51494 588874 51536
rect -4950 51258 -3090 51494
rect -2854 51258 -2770 51494
rect -2534 51258 -2450 51494
rect -2214 51258 -2130 51494
rect -1894 51258 1186 51494
rect 1422 51258 8186 51494
rect 8422 51258 15186 51494
rect 15422 51258 22186 51494
rect 22422 51258 29186 51494
rect 29422 51258 36186 51494
rect 36422 51258 43186 51494
rect 43422 51258 50186 51494
rect 50422 51258 57186 51494
rect 57422 51258 64186 51494
rect 64422 51258 71186 51494
rect 71422 51258 78186 51494
rect 78422 51258 85186 51494
rect 85422 51258 92186 51494
rect 92422 51258 99186 51494
rect 99422 51258 106186 51494
rect 106422 51258 113186 51494
rect 113422 51258 120186 51494
rect 120422 51258 127186 51494
rect 127422 51258 134186 51494
rect 134422 51258 141186 51494
rect 141422 51258 148186 51494
rect 148422 51258 155186 51494
rect 155422 51258 162186 51494
rect 162422 51258 169186 51494
rect 169422 51258 176186 51494
rect 176422 51258 183186 51494
rect 183422 51258 190186 51494
rect 190422 51258 197186 51494
rect 197422 51258 204186 51494
rect 204422 51258 211186 51494
rect 211422 51258 218186 51494
rect 218422 51258 225186 51494
rect 225422 51258 232186 51494
rect 232422 51258 239186 51494
rect 239422 51258 246186 51494
rect 246422 51258 253186 51494
rect 253422 51258 260186 51494
rect 260422 51258 267186 51494
rect 267422 51258 274186 51494
rect 274422 51258 281186 51494
rect 281422 51258 288186 51494
rect 288422 51258 295186 51494
rect 295422 51258 302186 51494
rect 302422 51258 309186 51494
rect 309422 51258 316186 51494
rect 316422 51258 323186 51494
rect 323422 51258 330186 51494
rect 330422 51258 337186 51494
rect 337422 51258 344186 51494
rect 344422 51258 351186 51494
rect 351422 51258 358186 51494
rect 358422 51258 365186 51494
rect 365422 51258 372186 51494
rect 372422 51258 379186 51494
rect 379422 51258 386186 51494
rect 386422 51258 393186 51494
rect 393422 51258 400186 51494
rect 400422 51258 407186 51494
rect 407422 51258 414186 51494
rect 414422 51258 421186 51494
rect 421422 51258 428186 51494
rect 428422 51258 435186 51494
rect 435422 51258 442186 51494
rect 442422 51258 449186 51494
rect 449422 51258 456186 51494
rect 456422 51258 463186 51494
rect 463422 51258 470186 51494
rect 470422 51258 477186 51494
rect 477422 51258 484186 51494
rect 484422 51258 491186 51494
rect 491422 51258 498186 51494
rect 498422 51258 505186 51494
rect 505422 51258 512186 51494
rect 512422 51258 519186 51494
rect 519422 51258 526186 51494
rect 526422 51258 533186 51494
rect 533422 51258 540186 51494
rect 540422 51258 547186 51494
rect 547422 51258 554186 51494
rect 554422 51258 561186 51494
rect 561422 51258 568186 51494
rect 568422 51258 575186 51494
rect 575422 51258 582186 51494
rect 582422 51258 585818 51494
rect 586054 51258 586138 51494
rect 586374 51258 586458 51494
rect 586694 51258 586778 51494
rect 587014 51258 588874 51494
rect -4950 51216 588874 51258
rect -4950 45434 588874 45476
rect -4950 45198 -4842 45434
rect -4606 45198 -4522 45434
rect -4286 45198 -4202 45434
rect -3966 45198 -3882 45434
rect -3646 45198 2918 45434
rect 3154 45198 9918 45434
rect 10154 45198 16918 45434
rect 17154 45198 23918 45434
rect 24154 45198 30918 45434
rect 31154 45198 37918 45434
rect 38154 45198 44918 45434
rect 45154 45198 51918 45434
rect 52154 45198 58918 45434
rect 59154 45198 65918 45434
rect 66154 45198 72918 45434
rect 73154 45198 79918 45434
rect 80154 45198 86918 45434
rect 87154 45198 93918 45434
rect 94154 45198 100918 45434
rect 101154 45198 107918 45434
rect 108154 45198 114918 45434
rect 115154 45198 121918 45434
rect 122154 45198 128918 45434
rect 129154 45198 135918 45434
rect 136154 45198 142918 45434
rect 143154 45198 149918 45434
rect 150154 45198 156918 45434
rect 157154 45198 163918 45434
rect 164154 45198 170918 45434
rect 171154 45198 177918 45434
rect 178154 45198 184918 45434
rect 185154 45198 191918 45434
rect 192154 45198 198918 45434
rect 199154 45198 205918 45434
rect 206154 45198 212918 45434
rect 213154 45198 219918 45434
rect 220154 45198 226918 45434
rect 227154 45198 233918 45434
rect 234154 45198 240918 45434
rect 241154 45198 247918 45434
rect 248154 45198 254918 45434
rect 255154 45198 261918 45434
rect 262154 45198 268918 45434
rect 269154 45198 275918 45434
rect 276154 45198 282918 45434
rect 283154 45198 289918 45434
rect 290154 45198 296918 45434
rect 297154 45198 303918 45434
rect 304154 45198 310918 45434
rect 311154 45198 317918 45434
rect 318154 45198 324918 45434
rect 325154 45198 331918 45434
rect 332154 45198 338918 45434
rect 339154 45198 345918 45434
rect 346154 45198 352918 45434
rect 353154 45198 359918 45434
rect 360154 45198 366918 45434
rect 367154 45198 373918 45434
rect 374154 45198 380918 45434
rect 381154 45198 387918 45434
rect 388154 45198 394918 45434
rect 395154 45198 401918 45434
rect 402154 45198 408918 45434
rect 409154 45198 415918 45434
rect 416154 45198 422918 45434
rect 423154 45198 429918 45434
rect 430154 45198 436918 45434
rect 437154 45198 443918 45434
rect 444154 45198 450918 45434
rect 451154 45198 457918 45434
rect 458154 45198 464918 45434
rect 465154 45198 471918 45434
rect 472154 45198 478918 45434
rect 479154 45198 485918 45434
rect 486154 45198 492918 45434
rect 493154 45198 499918 45434
rect 500154 45198 506918 45434
rect 507154 45198 513918 45434
rect 514154 45198 520918 45434
rect 521154 45198 527918 45434
rect 528154 45198 534918 45434
rect 535154 45198 541918 45434
rect 542154 45198 548918 45434
rect 549154 45198 555918 45434
rect 556154 45198 562918 45434
rect 563154 45198 569918 45434
rect 570154 45198 576918 45434
rect 577154 45198 587570 45434
rect 587806 45198 587890 45434
rect 588126 45198 588210 45434
rect 588446 45198 588530 45434
rect 588766 45198 588874 45434
rect -4950 45156 588874 45198
rect -4950 44494 588874 44536
rect -4950 44258 -3090 44494
rect -2854 44258 -2770 44494
rect -2534 44258 -2450 44494
rect -2214 44258 -2130 44494
rect -1894 44258 1186 44494
rect 1422 44258 8186 44494
rect 8422 44258 15186 44494
rect 15422 44258 22186 44494
rect 22422 44258 29186 44494
rect 29422 44258 36186 44494
rect 36422 44258 43186 44494
rect 43422 44258 50186 44494
rect 50422 44258 57186 44494
rect 57422 44258 64186 44494
rect 64422 44258 71186 44494
rect 71422 44258 78186 44494
rect 78422 44258 85186 44494
rect 85422 44258 92186 44494
rect 92422 44258 99186 44494
rect 99422 44258 106186 44494
rect 106422 44258 113186 44494
rect 113422 44258 120186 44494
rect 120422 44258 127186 44494
rect 127422 44258 134186 44494
rect 134422 44258 141186 44494
rect 141422 44258 148186 44494
rect 148422 44258 155186 44494
rect 155422 44258 162186 44494
rect 162422 44258 169186 44494
rect 169422 44258 176186 44494
rect 176422 44258 183186 44494
rect 183422 44258 190186 44494
rect 190422 44258 197186 44494
rect 197422 44258 204186 44494
rect 204422 44258 211186 44494
rect 211422 44258 218186 44494
rect 218422 44258 225186 44494
rect 225422 44258 232186 44494
rect 232422 44258 239186 44494
rect 239422 44258 246186 44494
rect 246422 44258 253186 44494
rect 253422 44258 260186 44494
rect 260422 44258 267186 44494
rect 267422 44258 274186 44494
rect 274422 44258 281186 44494
rect 281422 44258 288186 44494
rect 288422 44258 295186 44494
rect 295422 44258 302186 44494
rect 302422 44258 309186 44494
rect 309422 44258 316186 44494
rect 316422 44258 323186 44494
rect 323422 44258 330186 44494
rect 330422 44258 337186 44494
rect 337422 44258 344186 44494
rect 344422 44258 351186 44494
rect 351422 44258 358186 44494
rect 358422 44258 365186 44494
rect 365422 44258 372186 44494
rect 372422 44258 379186 44494
rect 379422 44258 386186 44494
rect 386422 44258 393186 44494
rect 393422 44258 400186 44494
rect 400422 44258 407186 44494
rect 407422 44258 414186 44494
rect 414422 44258 421186 44494
rect 421422 44258 428186 44494
rect 428422 44258 435186 44494
rect 435422 44258 442186 44494
rect 442422 44258 449186 44494
rect 449422 44258 456186 44494
rect 456422 44258 463186 44494
rect 463422 44258 470186 44494
rect 470422 44258 477186 44494
rect 477422 44258 484186 44494
rect 484422 44258 491186 44494
rect 491422 44258 498186 44494
rect 498422 44258 505186 44494
rect 505422 44258 512186 44494
rect 512422 44258 519186 44494
rect 519422 44258 526186 44494
rect 526422 44258 533186 44494
rect 533422 44258 540186 44494
rect 540422 44258 547186 44494
rect 547422 44258 554186 44494
rect 554422 44258 561186 44494
rect 561422 44258 568186 44494
rect 568422 44258 575186 44494
rect 575422 44258 582186 44494
rect 582422 44258 585818 44494
rect 586054 44258 586138 44494
rect 586374 44258 586458 44494
rect 586694 44258 586778 44494
rect 587014 44258 588874 44494
rect -4950 44216 588874 44258
rect -4950 38434 588874 38476
rect -4950 38198 -4842 38434
rect -4606 38198 -4522 38434
rect -4286 38198 -4202 38434
rect -3966 38198 -3882 38434
rect -3646 38198 2918 38434
rect 3154 38198 9918 38434
rect 10154 38198 16918 38434
rect 17154 38198 23918 38434
rect 24154 38198 30918 38434
rect 31154 38198 37918 38434
rect 38154 38198 44918 38434
rect 45154 38198 51918 38434
rect 52154 38198 58918 38434
rect 59154 38198 65918 38434
rect 66154 38198 72918 38434
rect 73154 38198 79918 38434
rect 80154 38198 86918 38434
rect 87154 38198 93918 38434
rect 94154 38198 100918 38434
rect 101154 38198 107918 38434
rect 108154 38198 114918 38434
rect 115154 38198 121918 38434
rect 122154 38198 128918 38434
rect 129154 38198 135918 38434
rect 136154 38198 142918 38434
rect 143154 38198 149918 38434
rect 150154 38198 156918 38434
rect 157154 38198 163918 38434
rect 164154 38198 170918 38434
rect 171154 38198 177918 38434
rect 178154 38198 184918 38434
rect 185154 38198 191918 38434
rect 192154 38198 198918 38434
rect 199154 38198 205918 38434
rect 206154 38198 212918 38434
rect 213154 38198 219918 38434
rect 220154 38198 226918 38434
rect 227154 38198 233918 38434
rect 234154 38198 240918 38434
rect 241154 38198 247918 38434
rect 248154 38198 254918 38434
rect 255154 38198 261918 38434
rect 262154 38198 268918 38434
rect 269154 38198 275918 38434
rect 276154 38198 282918 38434
rect 283154 38198 289918 38434
rect 290154 38198 296918 38434
rect 297154 38198 303918 38434
rect 304154 38198 310918 38434
rect 311154 38198 317918 38434
rect 318154 38198 324918 38434
rect 325154 38198 331918 38434
rect 332154 38198 338918 38434
rect 339154 38198 345918 38434
rect 346154 38198 352918 38434
rect 353154 38198 359918 38434
rect 360154 38198 366918 38434
rect 367154 38198 373918 38434
rect 374154 38198 380918 38434
rect 381154 38198 387918 38434
rect 388154 38198 394918 38434
rect 395154 38198 401918 38434
rect 402154 38198 408918 38434
rect 409154 38198 415918 38434
rect 416154 38198 422918 38434
rect 423154 38198 429918 38434
rect 430154 38198 436918 38434
rect 437154 38198 443918 38434
rect 444154 38198 450918 38434
rect 451154 38198 457918 38434
rect 458154 38198 464918 38434
rect 465154 38198 471918 38434
rect 472154 38198 478918 38434
rect 479154 38198 485918 38434
rect 486154 38198 492918 38434
rect 493154 38198 499918 38434
rect 500154 38198 506918 38434
rect 507154 38198 513918 38434
rect 514154 38198 520918 38434
rect 521154 38198 527918 38434
rect 528154 38198 534918 38434
rect 535154 38198 541918 38434
rect 542154 38198 548918 38434
rect 549154 38198 555918 38434
rect 556154 38198 562918 38434
rect 563154 38198 569918 38434
rect 570154 38198 576918 38434
rect 577154 38198 587570 38434
rect 587806 38198 587890 38434
rect 588126 38198 588210 38434
rect 588446 38198 588530 38434
rect 588766 38198 588874 38434
rect -4950 38156 588874 38198
rect -4950 37494 588874 37536
rect -4950 37258 -3090 37494
rect -2854 37258 -2770 37494
rect -2534 37258 -2450 37494
rect -2214 37258 -2130 37494
rect -1894 37258 1186 37494
rect 1422 37258 8186 37494
rect 8422 37258 15186 37494
rect 15422 37258 22186 37494
rect 22422 37258 29186 37494
rect 29422 37258 36186 37494
rect 36422 37258 43186 37494
rect 43422 37258 50186 37494
rect 50422 37258 57186 37494
rect 57422 37258 64186 37494
rect 64422 37258 71186 37494
rect 71422 37258 78186 37494
rect 78422 37258 85186 37494
rect 85422 37258 92186 37494
rect 92422 37258 99186 37494
rect 99422 37258 106186 37494
rect 106422 37258 113186 37494
rect 113422 37258 120186 37494
rect 120422 37258 127186 37494
rect 127422 37258 134186 37494
rect 134422 37258 141186 37494
rect 141422 37258 148186 37494
rect 148422 37258 155186 37494
rect 155422 37258 162186 37494
rect 162422 37258 169186 37494
rect 169422 37258 176186 37494
rect 176422 37258 183186 37494
rect 183422 37258 190186 37494
rect 190422 37258 197186 37494
rect 197422 37258 204186 37494
rect 204422 37258 211186 37494
rect 211422 37258 218186 37494
rect 218422 37258 225186 37494
rect 225422 37258 232186 37494
rect 232422 37258 239186 37494
rect 239422 37258 246186 37494
rect 246422 37258 253186 37494
rect 253422 37258 260186 37494
rect 260422 37258 267186 37494
rect 267422 37258 274186 37494
rect 274422 37258 281186 37494
rect 281422 37258 288186 37494
rect 288422 37258 295186 37494
rect 295422 37258 302186 37494
rect 302422 37258 309186 37494
rect 309422 37258 316186 37494
rect 316422 37258 323186 37494
rect 323422 37258 330186 37494
rect 330422 37258 337186 37494
rect 337422 37258 344186 37494
rect 344422 37258 351186 37494
rect 351422 37258 358186 37494
rect 358422 37258 365186 37494
rect 365422 37258 372186 37494
rect 372422 37258 379186 37494
rect 379422 37258 386186 37494
rect 386422 37258 393186 37494
rect 393422 37258 400186 37494
rect 400422 37258 407186 37494
rect 407422 37258 414186 37494
rect 414422 37258 421186 37494
rect 421422 37258 428186 37494
rect 428422 37258 435186 37494
rect 435422 37258 442186 37494
rect 442422 37258 449186 37494
rect 449422 37258 456186 37494
rect 456422 37258 463186 37494
rect 463422 37258 470186 37494
rect 470422 37258 477186 37494
rect 477422 37258 484186 37494
rect 484422 37258 491186 37494
rect 491422 37258 498186 37494
rect 498422 37258 505186 37494
rect 505422 37258 512186 37494
rect 512422 37258 519186 37494
rect 519422 37258 526186 37494
rect 526422 37258 533186 37494
rect 533422 37258 540186 37494
rect 540422 37258 547186 37494
rect 547422 37258 554186 37494
rect 554422 37258 561186 37494
rect 561422 37258 568186 37494
rect 568422 37258 575186 37494
rect 575422 37258 582186 37494
rect 582422 37258 585818 37494
rect 586054 37258 586138 37494
rect 586374 37258 586458 37494
rect 586694 37258 586778 37494
rect 587014 37258 588874 37494
rect -4950 37216 588874 37258
rect -4950 31434 588874 31476
rect -4950 31198 -4842 31434
rect -4606 31198 -4522 31434
rect -4286 31198 -4202 31434
rect -3966 31198 -3882 31434
rect -3646 31198 2918 31434
rect 3154 31198 9918 31434
rect 10154 31198 16918 31434
rect 17154 31198 23918 31434
rect 24154 31198 30918 31434
rect 31154 31198 37918 31434
rect 38154 31198 44918 31434
rect 45154 31198 51918 31434
rect 52154 31198 58918 31434
rect 59154 31198 65918 31434
rect 66154 31198 72918 31434
rect 73154 31198 79918 31434
rect 80154 31198 86918 31434
rect 87154 31198 93918 31434
rect 94154 31198 100918 31434
rect 101154 31198 107918 31434
rect 108154 31198 114918 31434
rect 115154 31198 121918 31434
rect 122154 31198 128918 31434
rect 129154 31198 135918 31434
rect 136154 31198 142918 31434
rect 143154 31198 149918 31434
rect 150154 31198 156918 31434
rect 157154 31198 163918 31434
rect 164154 31198 170918 31434
rect 171154 31198 177918 31434
rect 178154 31198 184918 31434
rect 185154 31198 191918 31434
rect 192154 31198 198918 31434
rect 199154 31198 205918 31434
rect 206154 31198 212918 31434
rect 213154 31198 219918 31434
rect 220154 31198 226918 31434
rect 227154 31198 233918 31434
rect 234154 31198 240918 31434
rect 241154 31198 247918 31434
rect 248154 31198 254918 31434
rect 255154 31198 261918 31434
rect 262154 31198 268918 31434
rect 269154 31198 275918 31434
rect 276154 31198 282918 31434
rect 283154 31198 289918 31434
rect 290154 31198 296918 31434
rect 297154 31198 303918 31434
rect 304154 31198 310918 31434
rect 311154 31198 317918 31434
rect 318154 31198 324918 31434
rect 325154 31198 331918 31434
rect 332154 31198 338918 31434
rect 339154 31198 345918 31434
rect 346154 31198 352918 31434
rect 353154 31198 359918 31434
rect 360154 31198 366918 31434
rect 367154 31198 373918 31434
rect 374154 31198 380918 31434
rect 381154 31198 387918 31434
rect 388154 31198 394918 31434
rect 395154 31198 401918 31434
rect 402154 31198 408918 31434
rect 409154 31198 415918 31434
rect 416154 31198 422918 31434
rect 423154 31198 429918 31434
rect 430154 31198 436918 31434
rect 437154 31198 443918 31434
rect 444154 31198 450918 31434
rect 451154 31198 457918 31434
rect 458154 31198 464918 31434
rect 465154 31198 471918 31434
rect 472154 31198 478918 31434
rect 479154 31198 485918 31434
rect 486154 31198 492918 31434
rect 493154 31198 499918 31434
rect 500154 31198 506918 31434
rect 507154 31198 513918 31434
rect 514154 31198 520918 31434
rect 521154 31198 527918 31434
rect 528154 31198 534918 31434
rect 535154 31198 541918 31434
rect 542154 31198 548918 31434
rect 549154 31198 555918 31434
rect 556154 31198 562918 31434
rect 563154 31198 569918 31434
rect 570154 31198 576918 31434
rect 577154 31198 587570 31434
rect 587806 31198 587890 31434
rect 588126 31198 588210 31434
rect 588446 31198 588530 31434
rect 588766 31198 588874 31434
rect -4950 31156 588874 31198
rect -4950 30494 588874 30536
rect -4950 30258 -3090 30494
rect -2854 30258 -2770 30494
rect -2534 30258 -2450 30494
rect -2214 30258 -2130 30494
rect -1894 30258 1186 30494
rect 1422 30258 8186 30494
rect 8422 30258 15186 30494
rect 15422 30258 22186 30494
rect 22422 30258 29186 30494
rect 29422 30258 36186 30494
rect 36422 30258 43186 30494
rect 43422 30258 50186 30494
rect 50422 30258 57186 30494
rect 57422 30258 64186 30494
rect 64422 30258 71186 30494
rect 71422 30258 78186 30494
rect 78422 30258 85186 30494
rect 85422 30258 92186 30494
rect 92422 30258 99186 30494
rect 99422 30258 106186 30494
rect 106422 30258 113186 30494
rect 113422 30258 120186 30494
rect 120422 30258 127186 30494
rect 127422 30258 134186 30494
rect 134422 30258 141186 30494
rect 141422 30258 148186 30494
rect 148422 30258 155186 30494
rect 155422 30258 162186 30494
rect 162422 30258 169186 30494
rect 169422 30258 176186 30494
rect 176422 30258 183186 30494
rect 183422 30258 190186 30494
rect 190422 30258 197186 30494
rect 197422 30258 204186 30494
rect 204422 30258 211186 30494
rect 211422 30258 218186 30494
rect 218422 30258 225186 30494
rect 225422 30258 232186 30494
rect 232422 30258 239186 30494
rect 239422 30258 246186 30494
rect 246422 30258 253186 30494
rect 253422 30258 260186 30494
rect 260422 30258 267186 30494
rect 267422 30258 274186 30494
rect 274422 30258 281186 30494
rect 281422 30258 288186 30494
rect 288422 30258 295186 30494
rect 295422 30258 302186 30494
rect 302422 30258 309186 30494
rect 309422 30258 316186 30494
rect 316422 30258 323186 30494
rect 323422 30258 330186 30494
rect 330422 30258 337186 30494
rect 337422 30258 344186 30494
rect 344422 30258 351186 30494
rect 351422 30258 358186 30494
rect 358422 30258 365186 30494
rect 365422 30258 372186 30494
rect 372422 30258 379186 30494
rect 379422 30258 386186 30494
rect 386422 30258 393186 30494
rect 393422 30258 400186 30494
rect 400422 30258 407186 30494
rect 407422 30258 414186 30494
rect 414422 30258 421186 30494
rect 421422 30258 428186 30494
rect 428422 30258 435186 30494
rect 435422 30258 442186 30494
rect 442422 30258 449186 30494
rect 449422 30258 456186 30494
rect 456422 30258 463186 30494
rect 463422 30258 470186 30494
rect 470422 30258 477186 30494
rect 477422 30258 484186 30494
rect 484422 30258 491186 30494
rect 491422 30258 498186 30494
rect 498422 30258 505186 30494
rect 505422 30258 512186 30494
rect 512422 30258 519186 30494
rect 519422 30258 526186 30494
rect 526422 30258 533186 30494
rect 533422 30258 540186 30494
rect 540422 30258 547186 30494
rect 547422 30258 554186 30494
rect 554422 30258 561186 30494
rect 561422 30258 568186 30494
rect 568422 30258 575186 30494
rect 575422 30258 582186 30494
rect 582422 30258 585818 30494
rect 586054 30258 586138 30494
rect 586374 30258 586458 30494
rect 586694 30258 586778 30494
rect 587014 30258 588874 30494
rect -4950 30216 588874 30258
rect -4950 24434 588874 24476
rect -4950 24198 -4842 24434
rect -4606 24198 -4522 24434
rect -4286 24198 -4202 24434
rect -3966 24198 -3882 24434
rect -3646 24198 2918 24434
rect 3154 24198 9918 24434
rect 10154 24198 16918 24434
rect 17154 24198 23918 24434
rect 24154 24198 30918 24434
rect 31154 24198 37918 24434
rect 38154 24198 44918 24434
rect 45154 24198 51918 24434
rect 52154 24198 58918 24434
rect 59154 24198 65918 24434
rect 66154 24198 72918 24434
rect 73154 24198 79918 24434
rect 80154 24198 86918 24434
rect 87154 24198 93918 24434
rect 94154 24198 100918 24434
rect 101154 24198 107918 24434
rect 108154 24198 114918 24434
rect 115154 24198 121918 24434
rect 122154 24198 128918 24434
rect 129154 24198 135918 24434
rect 136154 24198 142918 24434
rect 143154 24198 149918 24434
rect 150154 24198 156918 24434
rect 157154 24198 163918 24434
rect 164154 24198 170918 24434
rect 171154 24198 177918 24434
rect 178154 24198 184918 24434
rect 185154 24198 191918 24434
rect 192154 24198 198918 24434
rect 199154 24198 205918 24434
rect 206154 24198 212918 24434
rect 213154 24198 219918 24434
rect 220154 24198 226918 24434
rect 227154 24198 233918 24434
rect 234154 24198 240918 24434
rect 241154 24198 247918 24434
rect 248154 24198 254918 24434
rect 255154 24198 261918 24434
rect 262154 24198 268918 24434
rect 269154 24198 275918 24434
rect 276154 24198 282918 24434
rect 283154 24198 289918 24434
rect 290154 24198 296918 24434
rect 297154 24198 303918 24434
rect 304154 24198 310918 24434
rect 311154 24198 317918 24434
rect 318154 24198 324918 24434
rect 325154 24198 331918 24434
rect 332154 24198 338918 24434
rect 339154 24198 345918 24434
rect 346154 24198 352918 24434
rect 353154 24198 359918 24434
rect 360154 24198 366918 24434
rect 367154 24198 373918 24434
rect 374154 24198 380918 24434
rect 381154 24198 387918 24434
rect 388154 24198 394918 24434
rect 395154 24198 401918 24434
rect 402154 24198 408918 24434
rect 409154 24198 415918 24434
rect 416154 24198 422918 24434
rect 423154 24198 429918 24434
rect 430154 24198 436918 24434
rect 437154 24198 443918 24434
rect 444154 24198 450918 24434
rect 451154 24198 457918 24434
rect 458154 24198 464918 24434
rect 465154 24198 471918 24434
rect 472154 24198 478918 24434
rect 479154 24198 485918 24434
rect 486154 24198 492918 24434
rect 493154 24198 499918 24434
rect 500154 24198 506918 24434
rect 507154 24198 513918 24434
rect 514154 24198 520918 24434
rect 521154 24198 527918 24434
rect 528154 24198 534918 24434
rect 535154 24198 541918 24434
rect 542154 24198 548918 24434
rect 549154 24198 555918 24434
rect 556154 24198 562918 24434
rect 563154 24198 569918 24434
rect 570154 24198 576918 24434
rect 577154 24198 587570 24434
rect 587806 24198 587890 24434
rect 588126 24198 588210 24434
rect 588446 24198 588530 24434
rect 588766 24198 588874 24434
rect -4950 24156 588874 24198
rect -4950 23494 588874 23536
rect -4950 23258 -3090 23494
rect -2854 23258 -2770 23494
rect -2534 23258 -2450 23494
rect -2214 23258 -2130 23494
rect -1894 23258 1186 23494
rect 1422 23258 8186 23494
rect 8422 23258 15186 23494
rect 15422 23258 22186 23494
rect 22422 23258 29186 23494
rect 29422 23258 36186 23494
rect 36422 23258 43186 23494
rect 43422 23258 50186 23494
rect 50422 23258 57186 23494
rect 57422 23258 64186 23494
rect 64422 23258 71186 23494
rect 71422 23258 78186 23494
rect 78422 23258 85186 23494
rect 85422 23258 92186 23494
rect 92422 23258 99186 23494
rect 99422 23258 106186 23494
rect 106422 23258 113186 23494
rect 113422 23258 120186 23494
rect 120422 23258 127186 23494
rect 127422 23258 134186 23494
rect 134422 23258 141186 23494
rect 141422 23258 148186 23494
rect 148422 23258 155186 23494
rect 155422 23258 162186 23494
rect 162422 23258 169186 23494
rect 169422 23258 176186 23494
rect 176422 23258 183186 23494
rect 183422 23258 190186 23494
rect 190422 23258 197186 23494
rect 197422 23258 204186 23494
rect 204422 23258 211186 23494
rect 211422 23258 218186 23494
rect 218422 23258 225186 23494
rect 225422 23258 232186 23494
rect 232422 23258 239186 23494
rect 239422 23258 246186 23494
rect 246422 23258 253186 23494
rect 253422 23258 260186 23494
rect 260422 23258 267186 23494
rect 267422 23258 274186 23494
rect 274422 23258 281186 23494
rect 281422 23258 288186 23494
rect 288422 23258 295186 23494
rect 295422 23258 302186 23494
rect 302422 23258 309186 23494
rect 309422 23258 316186 23494
rect 316422 23258 323186 23494
rect 323422 23258 330186 23494
rect 330422 23258 337186 23494
rect 337422 23258 344186 23494
rect 344422 23258 351186 23494
rect 351422 23258 358186 23494
rect 358422 23258 365186 23494
rect 365422 23258 372186 23494
rect 372422 23258 379186 23494
rect 379422 23258 386186 23494
rect 386422 23258 393186 23494
rect 393422 23258 400186 23494
rect 400422 23258 407186 23494
rect 407422 23258 414186 23494
rect 414422 23258 421186 23494
rect 421422 23258 428186 23494
rect 428422 23258 435186 23494
rect 435422 23258 442186 23494
rect 442422 23258 449186 23494
rect 449422 23258 456186 23494
rect 456422 23258 463186 23494
rect 463422 23258 470186 23494
rect 470422 23258 477186 23494
rect 477422 23258 484186 23494
rect 484422 23258 491186 23494
rect 491422 23258 498186 23494
rect 498422 23258 505186 23494
rect 505422 23258 512186 23494
rect 512422 23258 519186 23494
rect 519422 23258 526186 23494
rect 526422 23258 533186 23494
rect 533422 23258 540186 23494
rect 540422 23258 547186 23494
rect 547422 23258 554186 23494
rect 554422 23258 561186 23494
rect 561422 23258 568186 23494
rect 568422 23258 575186 23494
rect 575422 23258 582186 23494
rect 582422 23258 585818 23494
rect 586054 23258 586138 23494
rect 586374 23258 586458 23494
rect 586694 23258 586778 23494
rect 587014 23258 588874 23494
rect -4950 23216 588874 23258
rect -4950 17434 588874 17476
rect -4950 17198 -4842 17434
rect -4606 17198 -4522 17434
rect -4286 17198 -4202 17434
rect -3966 17198 -3882 17434
rect -3646 17198 2918 17434
rect 3154 17198 9918 17434
rect 10154 17198 16918 17434
rect 17154 17198 23918 17434
rect 24154 17198 30918 17434
rect 31154 17198 37918 17434
rect 38154 17198 44918 17434
rect 45154 17198 51918 17434
rect 52154 17198 58918 17434
rect 59154 17198 65918 17434
rect 66154 17198 72918 17434
rect 73154 17198 79918 17434
rect 80154 17198 86918 17434
rect 87154 17198 93918 17434
rect 94154 17198 100918 17434
rect 101154 17198 107918 17434
rect 108154 17198 114918 17434
rect 115154 17198 121918 17434
rect 122154 17198 128918 17434
rect 129154 17198 135918 17434
rect 136154 17198 142918 17434
rect 143154 17198 149918 17434
rect 150154 17198 156918 17434
rect 157154 17198 163918 17434
rect 164154 17198 170918 17434
rect 171154 17198 177918 17434
rect 178154 17198 184918 17434
rect 185154 17198 191918 17434
rect 192154 17198 198918 17434
rect 199154 17198 205918 17434
rect 206154 17198 212918 17434
rect 213154 17198 219918 17434
rect 220154 17198 226918 17434
rect 227154 17198 233918 17434
rect 234154 17198 240918 17434
rect 241154 17198 247918 17434
rect 248154 17198 254918 17434
rect 255154 17198 261918 17434
rect 262154 17198 268918 17434
rect 269154 17198 275918 17434
rect 276154 17198 282918 17434
rect 283154 17198 289918 17434
rect 290154 17198 296918 17434
rect 297154 17198 303918 17434
rect 304154 17198 310918 17434
rect 311154 17198 317918 17434
rect 318154 17198 324918 17434
rect 325154 17198 331918 17434
rect 332154 17198 338918 17434
rect 339154 17198 345918 17434
rect 346154 17198 352918 17434
rect 353154 17198 359918 17434
rect 360154 17198 366918 17434
rect 367154 17198 373918 17434
rect 374154 17198 380918 17434
rect 381154 17198 387918 17434
rect 388154 17198 394918 17434
rect 395154 17198 401918 17434
rect 402154 17198 408918 17434
rect 409154 17198 415918 17434
rect 416154 17198 422918 17434
rect 423154 17198 429918 17434
rect 430154 17198 436918 17434
rect 437154 17198 443918 17434
rect 444154 17198 450918 17434
rect 451154 17198 457918 17434
rect 458154 17198 464918 17434
rect 465154 17198 471918 17434
rect 472154 17198 478918 17434
rect 479154 17198 485918 17434
rect 486154 17198 492918 17434
rect 493154 17198 499918 17434
rect 500154 17198 506918 17434
rect 507154 17198 513918 17434
rect 514154 17198 520918 17434
rect 521154 17198 527918 17434
rect 528154 17198 534918 17434
rect 535154 17198 541918 17434
rect 542154 17198 548918 17434
rect 549154 17198 555918 17434
rect 556154 17198 562918 17434
rect 563154 17198 569918 17434
rect 570154 17198 576918 17434
rect 577154 17198 587570 17434
rect 587806 17198 587890 17434
rect 588126 17198 588210 17434
rect 588446 17198 588530 17434
rect 588766 17198 588874 17434
rect -4950 17156 588874 17198
rect -4950 16494 588874 16536
rect -4950 16258 -3090 16494
rect -2854 16258 -2770 16494
rect -2534 16258 -2450 16494
rect -2214 16258 -2130 16494
rect -1894 16258 1186 16494
rect 1422 16258 8186 16494
rect 8422 16258 15186 16494
rect 15422 16258 22186 16494
rect 22422 16258 29186 16494
rect 29422 16258 36186 16494
rect 36422 16258 43186 16494
rect 43422 16258 50186 16494
rect 50422 16258 57186 16494
rect 57422 16258 64186 16494
rect 64422 16258 71186 16494
rect 71422 16258 78186 16494
rect 78422 16258 85186 16494
rect 85422 16258 92186 16494
rect 92422 16258 99186 16494
rect 99422 16258 106186 16494
rect 106422 16258 113186 16494
rect 113422 16258 120186 16494
rect 120422 16258 127186 16494
rect 127422 16258 134186 16494
rect 134422 16258 141186 16494
rect 141422 16258 148186 16494
rect 148422 16258 155186 16494
rect 155422 16258 162186 16494
rect 162422 16258 169186 16494
rect 169422 16258 176186 16494
rect 176422 16258 183186 16494
rect 183422 16258 190186 16494
rect 190422 16258 197186 16494
rect 197422 16258 204186 16494
rect 204422 16258 211186 16494
rect 211422 16258 218186 16494
rect 218422 16258 225186 16494
rect 225422 16258 232186 16494
rect 232422 16258 239186 16494
rect 239422 16258 246186 16494
rect 246422 16258 253186 16494
rect 253422 16258 260186 16494
rect 260422 16258 267186 16494
rect 267422 16258 274186 16494
rect 274422 16258 281186 16494
rect 281422 16258 288186 16494
rect 288422 16258 295186 16494
rect 295422 16258 302186 16494
rect 302422 16258 309186 16494
rect 309422 16258 316186 16494
rect 316422 16258 323186 16494
rect 323422 16258 330186 16494
rect 330422 16258 337186 16494
rect 337422 16258 344186 16494
rect 344422 16258 351186 16494
rect 351422 16258 358186 16494
rect 358422 16258 365186 16494
rect 365422 16258 372186 16494
rect 372422 16258 379186 16494
rect 379422 16258 386186 16494
rect 386422 16258 393186 16494
rect 393422 16258 400186 16494
rect 400422 16258 407186 16494
rect 407422 16258 414186 16494
rect 414422 16258 421186 16494
rect 421422 16258 428186 16494
rect 428422 16258 435186 16494
rect 435422 16258 442186 16494
rect 442422 16258 449186 16494
rect 449422 16258 456186 16494
rect 456422 16258 463186 16494
rect 463422 16258 470186 16494
rect 470422 16258 477186 16494
rect 477422 16258 484186 16494
rect 484422 16258 491186 16494
rect 491422 16258 498186 16494
rect 498422 16258 505186 16494
rect 505422 16258 512186 16494
rect 512422 16258 519186 16494
rect 519422 16258 526186 16494
rect 526422 16258 533186 16494
rect 533422 16258 540186 16494
rect 540422 16258 547186 16494
rect 547422 16258 554186 16494
rect 554422 16258 561186 16494
rect 561422 16258 568186 16494
rect 568422 16258 575186 16494
rect 575422 16258 582186 16494
rect 582422 16258 585818 16494
rect 586054 16258 586138 16494
rect 586374 16258 586458 16494
rect 586694 16258 586778 16494
rect 587014 16258 588874 16494
rect -4950 16216 588874 16258
rect -4950 10434 588874 10476
rect -4950 10198 -4842 10434
rect -4606 10198 -4522 10434
rect -4286 10198 -4202 10434
rect -3966 10198 -3882 10434
rect -3646 10198 2918 10434
rect 3154 10198 9918 10434
rect 10154 10198 16918 10434
rect 17154 10198 23918 10434
rect 24154 10198 30918 10434
rect 31154 10198 37918 10434
rect 38154 10198 44918 10434
rect 45154 10198 51918 10434
rect 52154 10198 58918 10434
rect 59154 10198 65918 10434
rect 66154 10198 72918 10434
rect 73154 10198 79918 10434
rect 80154 10198 86918 10434
rect 87154 10198 93918 10434
rect 94154 10198 100918 10434
rect 101154 10198 107918 10434
rect 108154 10198 114918 10434
rect 115154 10198 121918 10434
rect 122154 10198 128918 10434
rect 129154 10198 135918 10434
rect 136154 10198 142918 10434
rect 143154 10198 149918 10434
rect 150154 10198 156918 10434
rect 157154 10198 163918 10434
rect 164154 10198 170918 10434
rect 171154 10198 177918 10434
rect 178154 10198 184918 10434
rect 185154 10198 191918 10434
rect 192154 10198 198918 10434
rect 199154 10198 205918 10434
rect 206154 10198 212918 10434
rect 213154 10198 219918 10434
rect 220154 10198 226918 10434
rect 227154 10198 233918 10434
rect 234154 10198 240918 10434
rect 241154 10198 247918 10434
rect 248154 10198 254918 10434
rect 255154 10198 261918 10434
rect 262154 10198 268918 10434
rect 269154 10198 275918 10434
rect 276154 10198 282918 10434
rect 283154 10198 289918 10434
rect 290154 10198 296918 10434
rect 297154 10198 303918 10434
rect 304154 10198 310918 10434
rect 311154 10198 317918 10434
rect 318154 10198 324918 10434
rect 325154 10198 331918 10434
rect 332154 10198 338918 10434
rect 339154 10198 345918 10434
rect 346154 10198 352918 10434
rect 353154 10198 359918 10434
rect 360154 10198 366918 10434
rect 367154 10198 373918 10434
rect 374154 10198 380918 10434
rect 381154 10198 387918 10434
rect 388154 10198 394918 10434
rect 395154 10198 401918 10434
rect 402154 10198 408918 10434
rect 409154 10198 415918 10434
rect 416154 10198 422918 10434
rect 423154 10198 429918 10434
rect 430154 10198 436918 10434
rect 437154 10198 443918 10434
rect 444154 10198 450918 10434
rect 451154 10198 457918 10434
rect 458154 10198 464918 10434
rect 465154 10198 471918 10434
rect 472154 10198 478918 10434
rect 479154 10198 485918 10434
rect 486154 10198 492918 10434
rect 493154 10198 499918 10434
rect 500154 10198 506918 10434
rect 507154 10198 513918 10434
rect 514154 10198 520918 10434
rect 521154 10198 527918 10434
rect 528154 10198 534918 10434
rect 535154 10198 541918 10434
rect 542154 10198 548918 10434
rect 549154 10198 555918 10434
rect 556154 10198 562918 10434
rect 563154 10198 569918 10434
rect 570154 10198 576918 10434
rect 577154 10198 587570 10434
rect 587806 10198 587890 10434
rect 588126 10198 588210 10434
rect 588446 10198 588530 10434
rect 588766 10198 588874 10434
rect -4950 10156 588874 10198
rect -4950 9494 588874 9536
rect -4950 9258 -3090 9494
rect -2854 9258 -2770 9494
rect -2534 9258 -2450 9494
rect -2214 9258 -2130 9494
rect -1894 9258 1186 9494
rect 1422 9258 8186 9494
rect 8422 9258 15186 9494
rect 15422 9258 22186 9494
rect 22422 9258 29186 9494
rect 29422 9258 36186 9494
rect 36422 9258 43186 9494
rect 43422 9258 50186 9494
rect 50422 9258 57186 9494
rect 57422 9258 64186 9494
rect 64422 9258 71186 9494
rect 71422 9258 78186 9494
rect 78422 9258 85186 9494
rect 85422 9258 92186 9494
rect 92422 9258 99186 9494
rect 99422 9258 106186 9494
rect 106422 9258 113186 9494
rect 113422 9258 120186 9494
rect 120422 9258 127186 9494
rect 127422 9258 134186 9494
rect 134422 9258 141186 9494
rect 141422 9258 148186 9494
rect 148422 9258 155186 9494
rect 155422 9258 162186 9494
rect 162422 9258 169186 9494
rect 169422 9258 176186 9494
rect 176422 9258 183186 9494
rect 183422 9258 190186 9494
rect 190422 9258 197186 9494
rect 197422 9258 204186 9494
rect 204422 9258 211186 9494
rect 211422 9258 218186 9494
rect 218422 9258 225186 9494
rect 225422 9258 232186 9494
rect 232422 9258 239186 9494
rect 239422 9258 246186 9494
rect 246422 9258 253186 9494
rect 253422 9258 260186 9494
rect 260422 9258 267186 9494
rect 267422 9258 274186 9494
rect 274422 9258 281186 9494
rect 281422 9258 288186 9494
rect 288422 9258 295186 9494
rect 295422 9258 302186 9494
rect 302422 9258 309186 9494
rect 309422 9258 316186 9494
rect 316422 9258 323186 9494
rect 323422 9258 330186 9494
rect 330422 9258 337186 9494
rect 337422 9258 344186 9494
rect 344422 9258 351186 9494
rect 351422 9258 358186 9494
rect 358422 9258 365186 9494
rect 365422 9258 372186 9494
rect 372422 9258 379186 9494
rect 379422 9258 386186 9494
rect 386422 9258 393186 9494
rect 393422 9258 400186 9494
rect 400422 9258 407186 9494
rect 407422 9258 414186 9494
rect 414422 9258 421186 9494
rect 421422 9258 428186 9494
rect 428422 9258 435186 9494
rect 435422 9258 442186 9494
rect 442422 9258 449186 9494
rect 449422 9258 456186 9494
rect 456422 9258 463186 9494
rect 463422 9258 470186 9494
rect 470422 9258 477186 9494
rect 477422 9258 484186 9494
rect 484422 9258 491186 9494
rect 491422 9258 498186 9494
rect 498422 9258 505186 9494
rect 505422 9258 512186 9494
rect 512422 9258 519186 9494
rect 519422 9258 526186 9494
rect 526422 9258 533186 9494
rect 533422 9258 540186 9494
rect 540422 9258 547186 9494
rect 547422 9258 554186 9494
rect 554422 9258 561186 9494
rect 561422 9258 568186 9494
rect 568422 9258 575186 9494
rect 575422 9258 582186 9494
rect 582422 9258 585818 9494
rect 586054 9258 586138 9494
rect 586374 9258 586458 9494
rect 586694 9258 586778 9494
rect 587014 9258 588874 9494
rect -4950 9216 588874 9258
rect -4950 3434 588874 3476
rect -4950 3198 -4842 3434
rect -4606 3198 -4522 3434
rect -4286 3198 -4202 3434
rect -3966 3198 -3882 3434
rect -3646 3198 2918 3434
rect 3154 3198 9918 3434
rect 10154 3198 16918 3434
rect 17154 3198 23918 3434
rect 24154 3198 30918 3434
rect 31154 3198 37918 3434
rect 38154 3198 44918 3434
rect 45154 3198 51918 3434
rect 52154 3198 58918 3434
rect 59154 3198 65918 3434
rect 66154 3198 72918 3434
rect 73154 3198 79918 3434
rect 80154 3198 86918 3434
rect 87154 3198 93918 3434
rect 94154 3198 100918 3434
rect 101154 3198 107918 3434
rect 108154 3198 114918 3434
rect 115154 3198 121918 3434
rect 122154 3198 128918 3434
rect 129154 3198 135918 3434
rect 136154 3198 142918 3434
rect 143154 3198 149918 3434
rect 150154 3198 156918 3434
rect 157154 3198 163918 3434
rect 164154 3198 170918 3434
rect 171154 3198 177918 3434
rect 178154 3198 184918 3434
rect 185154 3198 191918 3434
rect 192154 3198 198918 3434
rect 199154 3198 205918 3434
rect 206154 3198 212918 3434
rect 213154 3198 219918 3434
rect 220154 3198 226918 3434
rect 227154 3198 233918 3434
rect 234154 3198 240918 3434
rect 241154 3198 247918 3434
rect 248154 3198 254918 3434
rect 255154 3198 261918 3434
rect 262154 3198 268918 3434
rect 269154 3198 275918 3434
rect 276154 3198 282918 3434
rect 283154 3198 289918 3434
rect 290154 3198 296918 3434
rect 297154 3198 303918 3434
rect 304154 3198 310918 3434
rect 311154 3198 317918 3434
rect 318154 3198 324918 3434
rect 325154 3198 331918 3434
rect 332154 3198 338918 3434
rect 339154 3198 345918 3434
rect 346154 3198 352918 3434
rect 353154 3198 359918 3434
rect 360154 3198 366918 3434
rect 367154 3198 373918 3434
rect 374154 3198 380918 3434
rect 381154 3198 387918 3434
rect 388154 3198 394918 3434
rect 395154 3198 401918 3434
rect 402154 3198 408918 3434
rect 409154 3198 415918 3434
rect 416154 3198 422918 3434
rect 423154 3198 429918 3434
rect 430154 3198 436918 3434
rect 437154 3198 443918 3434
rect 444154 3198 450918 3434
rect 451154 3198 457918 3434
rect 458154 3198 464918 3434
rect 465154 3198 471918 3434
rect 472154 3198 478918 3434
rect 479154 3198 485918 3434
rect 486154 3198 492918 3434
rect 493154 3198 499918 3434
rect 500154 3198 506918 3434
rect 507154 3198 513918 3434
rect 514154 3198 520918 3434
rect 521154 3198 527918 3434
rect 528154 3198 534918 3434
rect 535154 3198 541918 3434
rect 542154 3198 548918 3434
rect 549154 3198 555918 3434
rect 556154 3198 562918 3434
rect 563154 3198 569918 3434
rect 570154 3198 576918 3434
rect 577154 3198 587570 3434
rect 587806 3198 587890 3434
rect 588126 3198 588210 3434
rect 588446 3198 588530 3434
rect 588766 3198 588874 3434
rect -4950 3156 588874 3198
rect -4950 2494 588874 2536
rect -4950 2258 -3090 2494
rect -2854 2258 -2770 2494
rect -2534 2258 -2450 2494
rect -2214 2258 -2130 2494
rect -1894 2258 1186 2494
rect 1422 2258 8186 2494
rect 8422 2258 15186 2494
rect 15422 2258 22186 2494
rect 22422 2258 29186 2494
rect 29422 2258 36186 2494
rect 36422 2258 43186 2494
rect 43422 2258 50186 2494
rect 50422 2258 57186 2494
rect 57422 2258 64186 2494
rect 64422 2258 71186 2494
rect 71422 2258 78186 2494
rect 78422 2258 85186 2494
rect 85422 2258 92186 2494
rect 92422 2258 99186 2494
rect 99422 2258 106186 2494
rect 106422 2258 113186 2494
rect 113422 2258 120186 2494
rect 120422 2258 127186 2494
rect 127422 2258 134186 2494
rect 134422 2258 141186 2494
rect 141422 2258 148186 2494
rect 148422 2258 155186 2494
rect 155422 2258 162186 2494
rect 162422 2258 169186 2494
rect 169422 2258 176186 2494
rect 176422 2258 183186 2494
rect 183422 2258 190186 2494
rect 190422 2258 197186 2494
rect 197422 2258 204186 2494
rect 204422 2258 211186 2494
rect 211422 2258 218186 2494
rect 218422 2258 225186 2494
rect 225422 2258 232186 2494
rect 232422 2258 239186 2494
rect 239422 2258 246186 2494
rect 246422 2258 253186 2494
rect 253422 2258 260186 2494
rect 260422 2258 267186 2494
rect 267422 2258 274186 2494
rect 274422 2258 281186 2494
rect 281422 2258 288186 2494
rect 288422 2258 295186 2494
rect 295422 2258 302186 2494
rect 302422 2258 309186 2494
rect 309422 2258 316186 2494
rect 316422 2258 323186 2494
rect 323422 2258 330186 2494
rect 330422 2258 337186 2494
rect 337422 2258 344186 2494
rect 344422 2258 351186 2494
rect 351422 2258 358186 2494
rect 358422 2258 365186 2494
rect 365422 2258 372186 2494
rect 372422 2258 379186 2494
rect 379422 2258 386186 2494
rect 386422 2258 393186 2494
rect 393422 2258 400186 2494
rect 400422 2258 407186 2494
rect 407422 2258 414186 2494
rect 414422 2258 421186 2494
rect 421422 2258 428186 2494
rect 428422 2258 435186 2494
rect 435422 2258 442186 2494
rect 442422 2258 449186 2494
rect 449422 2258 456186 2494
rect 456422 2258 463186 2494
rect 463422 2258 470186 2494
rect 470422 2258 477186 2494
rect 477422 2258 484186 2494
rect 484422 2258 491186 2494
rect 491422 2258 498186 2494
rect 498422 2258 505186 2494
rect 505422 2258 512186 2494
rect 512422 2258 519186 2494
rect 519422 2258 526186 2494
rect 526422 2258 533186 2494
rect 533422 2258 540186 2494
rect 540422 2258 547186 2494
rect 547422 2258 554186 2494
rect 554422 2258 561186 2494
rect 561422 2258 568186 2494
rect 568422 2258 575186 2494
rect 575422 2258 582186 2494
rect 582422 2258 585818 2494
rect 586054 2258 586138 2494
rect 586374 2258 586458 2494
rect 586694 2258 586778 2494
rect 587014 2258 588874 2494
rect -4950 2216 588874 2258
rect -2406 -746 587122 -714
rect -2406 -982 -2374 -746
rect -2138 -982 -2054 -746
rect -1818 -982 1186 -746
rect 1422 -982 8186 -746
rect 8422 -982 15186 -746
rect 15422 -982 22186 -746
rect 22422 -982 29186 -746
rect 29422 -982 36186 -746
rect 36422 -982 43186 -746
rect 43422 -982 50186 -746
rect 50422 -982 57186 -746
rect 57422 -982 64186 -746
rect 64422 -982 71186 -746
rect 71422 -982 78186 -746
rect 78422 -982 85186 -746
rect 85422 -982 92186 -746
rect 92422 -982 99186 -746
rect 99422 -982 106186 -746
rect 106422 -982 113186 -746
rect 113422 -982 120186 -746
rect 120422 -982 127186 -746
rect 127422 -982 134186 -746
rect 134422 -982 141186 -746
rect 141422 -982 148186 -746
rect 148422 -982 155186 -746
rect 155422 -982 162186 -746
rect 162422 -982 169186 -746
rect 169422 -982 176186 -746
rect 176422 -982 183186 -746
rect 183422 -982 190186 -746
rect 190422 -982 197186 -746
rect 197422 -982 204186 -746
rect 204422 -982 211186 -746
rect 211422 -982 218186 -746
rect 218422 -982 225186 -746
rect 225422 -982 232186 -746
rect 232422 -982 239186 -746
rect 239422 -982 246186 -746
rect 246422 -982 253186 -746
rect 253422 -982 260186 -746
rect 260422 -982 267186 -746
rect 267422 -982 274186 -746
rect 274422 -982 281186 -746
rect 281422 -982 288186 -746
rect 288422 -982 295186 -746
rect 295422 -982 302186 -746
rect 302422 -982 309186 -746
rect 309422 -982 316186 -746
rect 316422 -982 323186 -746
rect 323422 -982 330186 -746
rect 330422 -982 337186 -746
rect 337422 -982 344186 -746
rect 344422 -982 351186 -746
rect 351422 -982 358186 -746
rect 358422 -982 365186 -746
rect 365422 -982 372186 -746
rect 372422 -982 379186 -746
rect 379422 -982 386186 -746
rect 386422 -982 393186 -746
rect 393422 -982 400186 -746
rect 400422 -982 407186 -746
rect 407422 -982 414186 -746
rect 414422 -982 421186 -746
rect 421422 -982 428186 -746
rect 428422 -982 435186 -746
rect 435422 -982 442186 -746
rect 442422 -982 449186 -746
rect 449422 -982 456186 -746
rect 456422 -982 463186 -746
rect 463422 -982 470186 -746
rect 470422 -982 477186 -746
rect 477422 -982 484186 -746
rect 484422 -982 491186 -746
rect 491422 -982 498186 -746
rect 498422 -982 505186 -746
rect 505422 -982 512186 -746
rect 512422 -982 519186 -746
rect 519422 -982 526186 -746
rect 526422 -982 533186 -746
rect 533422 -982 540186 -746
rect 540422 -982 547186 -746
rect 547422 -982 554186 -746
rect 554422 -982 561186 -746
rect 561422 -982 568186 -746
rect 568422 -982 575186 -746
rect 575422 -982 582186 -746
rect 582422 -982 585818 -746
rect 586054 -982 586138 -746
rect 586374 -982 586458 -746
rect 586694 -982 586778 -746
rect 587014 -982 587122 -746
rect -2406 -1066 587122 -982
rect -2406 -1302 -2374 -1066
rect -2138 -1302 -2054 -1066
rect -1818 -1302 1186 -1066
rect 1422 -1302 8186 -1066
rect 8422 -1302 15186 -1066
rect 15422 -1302 22186 -1066
rect 22422 -1302 29186 -1066
rect 29422 -1302 36186 -1066
rect 36422 -1302 43186 -1066
rect 43422 -1302 50186 -1066
rect 50422 -1302 57186 -1066
rect 57422 -1302 64186 -1066
rect 64422 -1302 71186 -1066
rect 71422 -1302 78186 -1066
rect 78422 -1302 85186 -1066
rect 85422 -1302 92186 -1066
rect 92422 -1302 99186 -1066
rect 99422 -1302 106186 -1066
rect 106422 -1302 113186 -1066
rect 113422 -1302 120186 -1066
rect 120422 -1302 127186 -1066
rect 127422 -1302 134186 -1066
rect 134422 -1302 141186 -1066
rect 141422 -1302 148186 -1066
rect 148422 -1302 155186 -1066
rect 155422 -1302 162186 -1066
rect 162422 -1302 169186 -1066
rect 169422 -1302 176186 -1066
rect 176422 -1302 183186 -1066
rect 183422 -1302 190186 -1066
rect 190422 -1302 197186 -1066
rect 197422 -1302 204186 -1066
rect 204422 -1302 211186 -1066
rect 211422 -1302 218186 -1066
rect 218422 -1302 225186 -1066
rect 225422 -1302 232186 -1066
rect 232422 -1302 239186 -1066
rect 239422 -1302 246186 -1066
rect 246422 -1302 253186 -1066
rect 253422 -1302 260186 -1066
rect 260422 -1302 267186 -1066
rect 267422 -1302 274186 -1066
rect 274422 -1302 281186 -1066
rect 281422 -1302 288186 -1066
rect 288422 -1302 295186 -1066
rect 295422 -1302 302186 -1066
rect 302422 -1302 309186 -1066
rect 309422 -1302 316186 -1066
rect 316422 -1302 323186 -1066
rect 323422 -1302 330186 -1066
rect 330422 -1302 337186 -1066
rect 337422 -1302 344186 -1066
rect 344422 -1302 351186 -1066
rect 351422 -1302 358186 -1066
rect 358422 -1302 365186 -1066
rect 365422 -1302 372186 -1066
rect 372422 -1302 379186 -1066
rect 379422 -1302 386186 -1066
rect 386422 -1302 393186 -1066
rect 393422 -1302 400186 -1066
rect 400422 -1302 407186 -1066
rect 407422 -1302 414186 -1066
rect 414422 -1302 421186 -1066
rect 421422 -1302 428186 -1066
rect 428422 -1302 435186 -1066
rect 435422 -1302 442186 -1066
rect 442422 -1302 449186 -1066
rect 449422 -1302 456186 -1066
rect 456422 -1302 463186 -1066
rect 463422 -1302 470186 -1066
rect 470422 -1302 477186 -1066
rect 477422 -1302 484186 -1066
rect 484422 -1302 491186 -1066
rect 491422 -1302 498186 -1066
rect 498422 -1302 505186 -1066
rect 505422 -1302 512186 -1066
rect 512422 -1302 519186 -1066
rect 519422 -1302 526186 -1066
rect 526422 -1302 533186 -1066
rect 533422 -1302 540186 -1066
rect 540422 -1302 547186 -1066
rect 547422 -1302 554186 -1066
rect 554422 -1302 561186 -1066
rect 561422 -1302 568186 -1066
rect 568422 -1302 575186 -1066
rect 575422 -1302 582186 -1066
rect 582422 -1302 585818 -1066
rect 586054 -1302 586138 -1066
rect 586374 -1302 586458 -1066
rect 586694 -1302 586778 -1066
rect 587014 -1302 587122 -1066
rect -2406 -1334 587122 -1302
rect -3366 -1706 587290 -1674
rect -3366 -1942 2918 -1706
rect 3154 -1942 9918 -1706
rect 10154 -1942 16918 -1706
rect 17154 -1942 23918 -1706
rect 24154 -1942 30918 -1706
rect 31154 -1942 37918 -1706
rect 38154 -1942 44918 -1706
rect 45154 -1942 51918 -1706
rect 52154 -1942 58918 -1706
rect 59154 -1942 65918 -1706
rect 66154 -1942 72918 -1706
rect 73154 -1942 79918 -1706
rect 80154 -1942 86918 -1706
rect 87154 -1942 93918 -1706
rect 94154 -1942 100918 -1706
rect 101154 -1942 107918 -1706
rect 108154 -1942 114918 -1706
rect 115154 -1942 121918 -1706
rect 122154 -1942 128918 -1706
rect 129154 -1942 135918 -1706
rect 136154 -1942 142918 -1706
rect 143154 -1942 149918 -1706
rect 150154 -1942 156918 -1706
rect 157154 -1942 163918 -1706
rect 164154 -1942 170918 -1706
rect 171154 -1942 177918 -1706
rect 178154 -1942 184918 -1706
rect 185154 -1942 191918 -1706
rect 192154 -1942 198918 -1706
rect 199154 -1942 205918 -1706
rect 206154 -1942 212918 -1706
rect 213154 -1942 219918 -1706
rect 220154 -1942 226918 -1706
rect 227154 -1942 233918 -1706
rect 234154 -1942 240918 -1706
rect 241154 -1942 247918 -1706
rect 248154 -1942 254918 -1706
rect 255154 -1942 261918 -1706
rect 262154 -1942 268918 -1706
rect 269154 -1942 275918 -1706
rect 276154 -1942 282918 -1706
rect 283154 -1942 289918 -1706
rect 290154 -1942 296918 -1706
rect 297154 -1942 303918 -1706
rect 304154 -1942 310918 -1706
rect 311154 -1942 317918 -1706
rect 318154 -1942 324918 -1706
rect 325154 -1942 331918 -1706
rect 332154 -1942 338918 -1706
rect 339154 -1942 345918 -1706
rect 346154 -1942 352918 -1706
rect 353154 -1942 359918 -1706
rect 360154 -1942 366918 -1706
rect 367154 -1942 373918 -1706
rect 374154 -1942 380918 -1706
rect 381154 -1942 387918 -1706
rect 388154 -1942 394918 -1706
rect 395154 -1942 401918 -1706
rect 402154 -1942 408918 -1706
rect 409154 -1942 415918 -1706
rect 416154 -1942 422918 -1706
rect 423154 -1942 429918 -1706
rect 430154 -1942 436918 -1706
rect 437154 -1942 443918 -1706
rect 444154 -1942 450918 -1706
rect 451154 -1942 457918 -1706
rect 458154 -1942 464918 -1706
rect 465154 -1942 471918 -1706
rect 472154 -1942 478918 -1706
rect 479154 -1942 485918 -1706
rect 486154 -1942 492918 -1706
rect 493154 -1942 499918 -1706
rect 500154 -1942 506918 -1706
rect 507154 -1942 513918 -1706
rect 514154 -1942 520918 -1706
rect 521154 -1942 527918 -1706
rect 528154 -1942 534918 -1706
rect 535154 -1942 541918 -1706
rect 542154 -1942 548918 -1706
rect 549154 -1942 555918 -1706
rect 556154 -1942 562918 -1706
rect 563154 -1942 569918 -1706
rect 570154 -1942 576918 -1706
rect 577154 -1942 587290 -1706
rect -3366 -2026 587290 -1942
rect -3366 -2262 2918 -2026
rect 3154 -2262 9918 -2026
rect 10154 -2262 16918 -2026
rect 17154 -2262 23918 -2026
rect 24154 -2262 30918 -2026
rect 31154 -2262 37918 -2026
rect 38154 -2262 44918 -2026
rect 45154 -2262 51918 -2026
rect 52154 -2262 58918 -2026
rect 59154 -2262 65918 -2026
rect 66154 -2262 72918 -2026
rect 73154 -2262 79918 -2026
rect 80154 -2262 86918 -2026
rect 87154 -2262 93918 -2026
rect 94154 -2262 100918 -2026
rect 101154 -2262 107918 -2026
rect 108154 -2262 114918 -2026
rect 115154 -2262 121918 -2026
rect 122154 -2262 128918 -2026
rect 129154 -2262 135918 -2026
rect 136154 -2262 142918 -2026
rect 143154 -2262 149918 -2026
rect 150154 -2262 156918 -2026
rect 157154 -2262 163918 -2026
rect 164154 -2262 170918 -2026
rect 171154 -2262 177918 -2026
rect 178154 -2262 184918 -2026
rect 185154 -2262 191918 -2026
rect 192154 -2262 198918 -2026
rect 199154 -2262 205918 -2026
rect 206154 -2262 212918 -2026
rect 213154 -2262 219918 -2026
rect 220154 -2262 226918 -2026
rect 227154 -2262 233918 -2026
rect 234154 -2262 240918 -2026
rect 241154 -2262 247918 -2026
rect 248154 -2262 254918 -2026
rect 255154 -2262 261918 -2026
rect 262154 -2262 268918 -2026
rect 269154 -2262 275918 -2026
rect 276154 -2262 282918 -2026
rect 283154 -2262 289918 -2026
rect 290154 -2262 296918 -2026
rect 297154 -2262 303918 -2026
rect 304154 -2262 310918 -2026
rect 311154 -2262 317918 -2026
rect 318154 -2262 324918 -2026
rect 325154 -2262 331918 -2026
rect 332154 -2262 338918 -2026
rect 339154 -2262 345918 -2026
rect 346154 -2262 352918 -2026
rect 353154 -2262 359918 -2026
rect 360154 -2262 366918 -2026
rect 367154 -2262 373918 -2026
rect 374154 -2262 380918 -2026
rect 381154 -2262 387918 -2026
rect 388154 -2262 394918 -2026
rect 395154 -2262 401918 -2026
rect 402154 -2262 408918 -2026
rect 409154 -2262 415918 -2026
rect 416154 -2262 422918 -2026
rect 423154 -2262 429918 -2026
rect 430154 -2262 436918 -2026
rect 437154 -2262 443918 -2026
rect 444154 -2262 450918 -2026
rect 451154 -2262 457918 -2026
rect 458154 -2262 464918 -2026
rect 465154 -2262 471918 -2026
rect 472154 -2262 478918 -2026
rect 479154 -2262 485918 -2026
rect 486154 -2262 492918 -2026
rect 493154 -2262 499918 -2026
rect 500154 -2262 506918 -2026
rect 507154 -2262 513918 -2026
rect 514154 -2262 520918 -2026
rect 521154 -2262 527918 -2026
rect 528154 -2262 534918 -2026
rect 535154 -2262 541918 -2026
rect 542154 -2262 548918 -2026
rect 549154 -2262 555918 -2026
rect 556154 -2262 562918 -2026
rect 563154 -2262 569918 -2026
rect 570154 -2262 576918 -2026
rect 577154 -2262 587290 -2026
rect -3366 -2294 587290 -2262
use mux16x1_project  mprj1
timestamp 0
transform 1 0 518000 0 1 400000
box 0 552 10000 22000
use mux16x1_project  mprj2
timestamp 0
transform 1 0 518000 0 1 360000
box 0 552 10000 22000
use mux16x1_project  mprj3
timestamp 0
transform 1 0 518000 0 1 320000
box 0 552 10000 22000
use mux16x1_project  mprj4
timestamp 0
transform 1 0 518000 0 1 280000
box 0 552 10000 22000
use mux16x1_project  mprj5
timestamp 0
transform 1 0 518000 0 1 240000
box 0 552 10000 22000
use sky130_osu_ring_oscillator_mpr2aa_8_b0r1  ro1
timestamp 0
transform 1 0 292001 0 1 491600
box -1 0 16356 1776
use sky130_osu_ring_oscillator_mpr2at_8_b0r1  ro2
timestamp 0
transform 1 0 291708 0 1 470600
box 292 0 18779 1776
use sky130_osu_ring_oscillator_mpr2ca_8_b0r1  ro3
timestamp 0
transform 1 0 292000 0 1 449600
box 0 0 17151 1776
use sky130_osu_ring_oscillator_mpr2ct_8_b0r1  ro4
timestamp 0
transform 1 0 292000 0 1 428600
box 0 0 17782 1776
use sky130_osu_ring_oscillator_mpr2ea_8_b0r1  ro5
timestamp 0
transform 1 0 292000 0 1 407600
box 0 0 16885 1776
use sky130_osu_ring_oscillator_mpr2et_8_b0r1  ro6
timestamp 0
transform 1 0 292000 0 1 386600
box 0 0 19119 1776
use sky130_osu_ring_oscillator_mpr2xa_8_b0r1  ro7
timestamp 0
transform 1 0 292000 0 1 365600
box 2 0 15820 1776
use sky130_osu_ring_oscillator_mpr2ya_8_b0r1  ro8
timestamp 0
transform 1 0 292000 0 1 344600
box 0 0 15819 1778
use sky130_osu_ring_oscillator_mpr2aa_8_b0r2  ro9
timestamp 0
transform 1 0 292000 0 1 323600
box 0 0 16353 1776
use sky130_osu_ring_oscillator_mpr2at_8_b0r2  ro10
timestamp 0
transform 1 0 292000 0 1 302600
box 0 0 18515 1776
use sky130_osu_ring_oscillator_mpr2ca_8_b0r2  ro11
timestamp 0
transform 1 0 292000 0 1 281600
box 0 0 17176 1776
use sky130_osu_ring_oscillator_mpr2ct_8_b0r2  ro12
timestamp 0
transform 1 0 292000 0 1 260600
box 0 0 17780 1776
use sky130_osu_ring_oscillator_mpr2ea_8_b0r2  ro13
timestamp 0
transform 1 0 292000 0 1 239600
box 0 0 16884 1776
use sky130_osu_ring_oscillator_mpr2et_8_b0r2  ro14
timestamp 0
transform 1 0 292000 0 1 218600
box 0 0 19119 1776
use sky130_osu_ring_oscillator_mpr2xa_8_b0r2  ro15
timestamp 0
transform 1 0 292000 0 1 197600
box 0 0 15819 1776
use sky130_osu_ring_oscillator_mpr2ya_8_b0r2  ro16
timestamp 0
transform 1 0 292000 0 1 176800
box 0 0 15819 1776
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal4 s -3198 -2126 -1786 706062 0 FreeSans 7680 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -2406 -1334 587122 -714 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -2406 704650 587122 705270 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 585710 -2126 587122 706062 0 FreeSans 7680 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 1144 -2294 1464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 8144 -2294 8464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 15144 -2294 15464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 22144 -2294 22464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 29144 -2294 29464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 36144 -2294 36464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 43144 -2294 43464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 50144 -2294 50464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 57144 -2294 57464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 64144 -2294 64464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 71144 -2294 71464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 78144 -2294 78464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 85144 -2294 85464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 92144 -2294 92464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 99144 -2294 99464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 106144 -2294 106464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 113144 -2294 113464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 120144 -2294 120464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 127144 -2294 127464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 134144 -2294 134464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 141144 -2294 141464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 148144 -2294 148464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 155144 -2294 155464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 162144 -2294 162464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 169144 -2294 169464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 176144 -2294 176464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 183144 -2294 183464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 190144 -2294 190464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 197144 -2294 197464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 204144 -2294 204464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 211144 -2294 211464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 218144 -2294 218464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 225144 -2294 225464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 232144 -2294 232464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 239144 -2294 239464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 246144 -2294 246464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 253144 -2294 253464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 260144 -2294 260464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 267144 -2294 267464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 274144 -2294 274464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 281144 -2294 281464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 288144 -2294 288464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 295144 -2294 295464 195976 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 295144 200380 295464 363976 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 295144 368380 295464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 302144 -2294 302464 195976 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 302144 200380 302464 363976 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 302144 368380 302464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 309144 -2294 309464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 316144 -2294 316464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 323144 -2294 323464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 330144 -2294 330464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 337144 -2294 337464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 344144 -2294 344464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 351144 -2294 351464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 358144 -2294 358464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 365144 -2294 365464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 372144 -2294 372464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 379144 -2294 379464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 386144 -2294 386464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 393144 -2294 393464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 400144 -2294 400464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 407144 -2294 407464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 414144 -2294 414464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 421144 -2294 421464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 428144 -2294 428464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 435144 -2294 435464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 442144 -2294 442464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 449144 -2294 449464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 456144 -2294 456464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 463144 -2294 463464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 470144 -2294 470464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 477144 -2294 477464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 484144 -2294 484464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 491144 -2294 491464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 498144 -2294 498464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 505144 -2294 505464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 512144 -2294 512464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 519144 -2294 519464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 -2294 526464 240008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 261752 526464 280008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 301752 526464 320008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 341752 526464 360008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 381752 526464 400008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 421752 526464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 533144 -2294 533464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 540144 -2294 540464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 547144 -2294 547464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 554144 -2294 554464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 561144 -2294 561464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 568144 -2294 568464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 575144 -2294 575464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 582144 -2294 582464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 2216 588874 2536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 9216 588874 9536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 16216 588874 16536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 23216 588874 23536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 30216 588874 30536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 37216 588874 37536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 44216 588874 44536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 51216 588874 51536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 58216 588874 58536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 65216 588874 65536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 72216 588874 72536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 79216 588874 79536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 86216 588874 86536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 93216 588874 93536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 100216 588874 100536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 107216 588874 107536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 114216 588874 114536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 121216 588874 121536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 128216 588874 128536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 135216 588874 135536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 142216 588874 142536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 149216 588874 149536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 156216 588874 156536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 163216 588874 163536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 170216 588874 170536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 177216 588874 177536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 184216 588874 184536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 191216 588874 191536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 198216 588874 198536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 205216 588874 205536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 212216 588874 212536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 219216 588874 219536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 226216 588874 226536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 233216 588874 233536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 240216 588874 240536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 247216 588874 247536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 254216 588874 254536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 261216 588874 261536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 268216 588874 268536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 275216 588874 275536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 282216 588874 282536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 289216 588874 289536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 296216 588874 296536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 303216 588874 303536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 310216 588874 310536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 317216 588874 317536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 324216 588874 324536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 331216 588874 331536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 338216 588874 338536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 345216 588874 345536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 352216 588874 352536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 359216 588874 359536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 366216 588874 366536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 373216 588874 373536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 380216 588874 380536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 387216 588874 387536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 394216 588874 394536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 401216 588874 401536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 408216 588874 408536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 415216 588874 415536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 422216 588874 422536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 429216 588874 429536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 436216 588874 436536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 443216 588874 443536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 450216 588874 450536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 457216 588874 457536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 464216 588874 464536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 471216 588874 471536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 478216 588874 478536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 485216 588874 485536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 492216 588874 492536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 499216 588874 499536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 506216 588874 506536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 513216 588874 513536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 520216 588874 520536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 527216 588874 527536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 534216 588874 534536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 541216 588874 541536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 548216 588874 548536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 555216 588874 555536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 562216 588874 562536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 569216 588874 569536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 576216 588874 576536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 583216 588874 583536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 590216 588874 590536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 597216 588874 597536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 604216 588874 604536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 611216 588874 611536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 618216 588874 618536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 625216 588874 625536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 632216 588874 632536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 639216 588874 639536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 646216 588874 646536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 653216 588874 653536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 660216 588874 660536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 667216 588874 667536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 674216 588874 674536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 681216 588874 681536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 688216 588874 688536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 695216 588874 695536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s -4950 -3878 -3538 707814 0 FreeSans 7680 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3366 -2294 587290 -1674 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3366 705610 587290 706230 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 587462 -3878 588874 707814 0 FreeSans 7680 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 2876 -2294 3196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 9876 -2294 10196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 16876 -2294 17196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 23876 -2294 24196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 30876 -2294 31196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 37876 -2294 38196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 44876 -2294 45196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 51876 -2294 52196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 58876 -2294 59196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 65876 -2294 66196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 72876 -2294 73196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 79876 -2294 80196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 86876 -2294 87196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 93876 -2294 94196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 100876 -2294 101196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 107876 -2294 108196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 114876 -2294 115196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 121876 -2294 122196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 128876 -2294 129196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 135876 -2294 136196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 142876 -2294 143196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 149876 -2294 150196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 156876 -2294 157196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 163876 -2294 164196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 170876 -2294 171196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 177876 -2294 178196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 184876 -2294 185196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 191876 -2294 192196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 198876 -2294 199196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 205876 -2294 206196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 212876 -2294 213196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 219876 -2294 220196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 226876 -2294 227196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 233876 -2294 234196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 240876 -2294 241196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 247876 -2294 248196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 254876 -2294 255196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 261876 -2294 262196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 268876 -2294 269196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 275876 -2294 276196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 282876 -2294 283196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 289876 -2294 290196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 296876 -2294 297196 195976 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 296876 200380 297196 363976 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 296876 368380 297196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 303876 -2294 304196 195976 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 303876 200380 304196 363976 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 303876 368380 304196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 310876 -2294 311196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 317876 -2294 318196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 324876 -2294 325196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 331876 -2294 332196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 338876 -2294 339196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 345876 -2294 346196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 352876 -2294 353196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 359876 -2294 360196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 366876 -2294 367196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 373876 -2294 374196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 380876 -2294 381196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 387876 -2294 388196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 394876 -2294 395196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 401876 -2294 402196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 408876 -2294 409196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 415876 -2294 416196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 422876 -2294 423196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 429876 -2294 430196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 436876 -2294 437196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 443876 -2294 444196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 450876 -2294 451196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 457876 -2294 458196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 464876 -2294 465196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 471876 -2294 472196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 478876 -2294 479196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 485876 -2294 486196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 492876 -2294 493196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 499876 -2294 500196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 506876 -2294 507196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 513876 -2294 514196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 -2294 521196 240008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 261752 521196 280008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 301752 521196 320008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 341752 521196 360008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 381752 521196 400008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 421752 521196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 527876 -2294 528196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 534876 -2294 535196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 541876 -2294 542196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 548876 -2294 549196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 555876 -2294 556196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 562876 -2294 563196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 569876 -2294 570196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 576876 -2294 577196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 3156 588874 3476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 10156 588874 10476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 17156 588874 17476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 24156 588874 24476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 31156 588874 31476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 38156 588874 38476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 45156 588874 45476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 52156 588874 52476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 59156 588874 59476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 66156 588874 66476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 73156 588874 73476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 80156 588874 80476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 87156 588874 87476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 94156 588874 94476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 101156 588874 101476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 108156 588874 108476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 115156 588874 115476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 122156 588874 122476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 129156 588874 129476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 136156 588874 136476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 143156 588874 143476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 150156 588874 150476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 157156 588874 157476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 164156 588874 164476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 171156 588874 171476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 178156 588874 178476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 185156 588874 185476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 192156 588874 192476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 199156 588874 199476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 206156 588874 206476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 213156 588874 213476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 220156 588874 220476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 227156 588874 227476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 234156 588874 234476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 241156 588874 241476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 248156 588874 248476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 255156 588874 255476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 262156 588874 262476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 269156 588874 269476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 276156 588874 276476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 283156 588874 283476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 290156 588874 290476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 297156 588874 297476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 304156 588874 304476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 311156 588874 311476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 318156 588874 318476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 325156 588874 325476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 332156 588874 332476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 339156 588874 339476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 346156 588874 346476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 353156 588874 353476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 360156 588874 360476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 367156 588874 367476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 374156 588874 374476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 381156 588874 381476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 388156 588874 388476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 395156 588874 395476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 402156 588874 402476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 409156 588874 409476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 416156 588874 416476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 423156 588874 423476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 430156 588874 430476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 437156 588874 437476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 444156 588874 444476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 451156 588874 451476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 458156 588874 458476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 465156 588874 465476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 472156 588874 472476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 479156 588874 479476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 486156 588874 486476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 493156 588874 493476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 500156 588874 500476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 507156 588874 507476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 514156 588874 514476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 521156 588874 521476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 528156 588874 528476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 535156 588874 535476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 542156 588874 542476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 549156 588874 549476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 556156 588874 556476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 563156 588874 563476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 570156 588874 570476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 577156 588874 577476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 584156 588874 584476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 591156 588874 591476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 598156 588874 598476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 605156 588874 605476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 612156 588874 612476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 619156 588874 619476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 626156 588874 626476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 633156 588874 633476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 640156 588874 640476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 647156 588874 647476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 654156 588874 654476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 661156 588874 661476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 668156 588874 668476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 675156 588874 675476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 682156 588874 682476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 689156 588874 689476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 696156 588874 696476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 145 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 146 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 147 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 148 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 149 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 150 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 151 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 152 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 153 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 154 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 155 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 156 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 157 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 158 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 159 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 160 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 161 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 162 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 163 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 164 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 165 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 166 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 167 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 168 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 169 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 170 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 171 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 172 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 173 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 174 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 175 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 176 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 177 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 178 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 179 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 180 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 181 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 182 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 183 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 184 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 185 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 186 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 187 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 188 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 189 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 190 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 191 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 192 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 193 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 194 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 195 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 196 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 197 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 198 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 199 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 200 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 201 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 202 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 203 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 204 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 205 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 206 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 207 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 208 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 209 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 210 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 211 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 212 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 213 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 214 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 215 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 216 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 217 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 218 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 219 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 220 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 221 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 222 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 223 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 224 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 225 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 226 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 227 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 228 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 229 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 230 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 231 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 232 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 233 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 234 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 235 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 236 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 237 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 238 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 239 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 240 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 241 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 242 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 243 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 244 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 245 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 246 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 247 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 248 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 249 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 250 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
