magic
tech sky130A
magscale 1 2
timestamp 1604095907
<< checkpaint >>
rect -1269 2461 1615 2601
rect -1760 -1129 6260 2461
rect -1269 -1260 1615 -1129
<< nwell >>
rect -9 485 355 897
<< locali >>
rect 0 827 352 888
rect 0 0 352 61
<< metal1 >>
rect 0 827 352 888
rect 0 0 352 61
<< labels >>
rlabel metal1 199 856 199 856 1 vccd1
rlabel metal1 196 30 196 30 1 vssd1
<< end >>
