magic
tech sky130A
magscale 1 2
timestamp 1707510517
<< error_s >>
rect 1380 1037 1523 1039
rect 321 1023 422 1034
rect 608 1033 872 1034
rect 872 1023 927 1033
rect 1030 1027 1039 1036
rect 1077 1027 1086 1036
rect 1380 1034 1502 1037
rect 1352 1033 1369 1034
rect 1182 1027 1352 1033
rect 306 1021 321 1023
rect 300 1019 306 1021
rect 929 1019 934 1021
rect 296 1014 300 1019
rect 934 1014 941 1019
rect 1021 1018 1030 1027
rect 1086 1024 1182 1027
rect 1523 1023 1631 1037
rect 1381 1015 1397 1022
rect 1399 1015 1415 1022
rect 941 1007 953 1014
rect 1371 1013 1383 1015
rect 1393 1013 1405 1015
rect 1411 1013 1415 1015
rect 1599 1013 1615 1022
rect 1631 1021 1649 1023
rect 1650 1017 1657 1020
rect 1657 1013 1663 1017
rect 1371 1008 1415 1013
rect 1558 1008 1595 1009
rect 1663 1008 1666 1013
rect 1367 1006 1369 1008
rect 1371 1006 1503 1008
rect 422 1005 776 1006
rect 402 1003 420 1005
rect 862 1003 875 1005
rect 954 1003 957 1005
rect 1365 1003 1503 1006
rect 346 1000 402 1003
rect 220 992 232 1000
rect 242 992 254 1000
rect 318 994 402 1000
rect 875 994 885 1003
rect 318 993 346 994
rect 216 989 218 992
rect 318 991 337 993
rect 886 991 889 993
rect 258 988 262 989
rect 208 977 216 988
rect 219 986 254 988
rect 217 977 219 983
rect 208 976 217 977
rect 216 972 217 976
rect 215 971 216 972
rect 213 966 215 969
rect 88 964 153 965
rect 80 956 88 964
rect 153 956 157 964
rect 79 950 80 956
rect 208 954 216 966
rect 220 956 222 986
rect 251 985 254 986
rect 253 979 254 985
rect 258 981 266 988
rect 262 980 270 981
rect 294 980 295 990
rect 318 980 333 991
rect 592 981 629 983
rect 270 979 276 980
rect 293 979 294 980
rect 318 979 325 980
rect 276 969 338 979
rect 346 972 352 978
rect 392 972 398 978
rect 592 977 618 981
rect 629 977 634 981
rect 889 980 902 991
rect 865 979 879 980
rect 586 972 592 977
rect 634 972 643 977
rect 847 972 865 979
rect 879 977 886 979
rect 957 977 978 1003
rect 1359 996 1503 1003
rect 1519 1006 1620 1008
rect 1519 996 1631 1006
rect 1320 990 1381 996
rect 1285 987 1320 990
rect 1098 981 1285 987
rect 1371 986 1381 990
rect 886 972 901 977
rect 340 969 346 972
rect 347 970 404 972
rect 643 971 644 972
rect 481 970 484 971
rect 502 970 505 971
rect 584 970 585 971
rect 644 970 647 971
rect 347 969 355 970
rect 318 968 355 969
rect 220 954 254 956
rect 209 951 211 954
rect 205 938 209 950
rect 220 942 232 950
rect 245 945 254 954
rect 292 952 293 955
rect 318 951 323 968
rect 340 966 355 968
rect 398 966 404 970
rect 477 967 481 970
rect 505 967 510 970
rect 647 968 648 970
rect 839 969 847 972
rect 876 971 901 972
rect 910 971 914 972
rect 872 970 876 971
rect 886 970 923 971
rect 648 967 651 968
rect 346 964 355 966
rect 346 951 351 964
rect 399 955 418 958
rect 453 955 477 967
rect 510 959 528 967
rect 583 959 584 967
rect 255 949 260 950
rect 260 948 265 949
rect 265 947 268 948
rect 270 945 279 947
rect 243 942 245 945
rect 279 944 284 945
rect 284 943 290 944
rect 291 943 292 951
rect 318 943 324 951
rect 242 939 243 942
rect 290 938 324 943
rect 203 931 205 937
rect 240 930 242 938
rect 291 932 292 938
rect 318 935 346 938
rect 318 933 348 935
rect 318 931 349 933
rect 350 931 351 951
rect 418 946 480 955
rect 528 952 536 959
rect 582 951 583 958
rect 651 954 655 967
rect 831 966 839 969
rect 869 968 872 970
rect 865 967 869 968
rect 860 965 865 967
rect 886 965 901 970
rect 910 969 914 970
rect 923 969 924 970
rect 980 969 985 975
rect 1021 971 1030 980
rect 1086 978 1098 981
rect 1086 971 1095 978
rect 1365 972 1381 986
rect 1404 972 1405 996
rect 1410 991 1431 996
rect 1415 990 1431 991
rect 1548 989 1554 996
rect 1600 989 1606 996
rect 1620 990 1631 996
rect 1666 990 1675 1008
rect 1415 972 1431 988
rect 1548 985 1556 989
rect 1554 983 1556 985
rect 1464 974 1492 978
rect 1494 974 1505 978
rect 914 965 919 969
rect 924 965 926 968
rect 985 965 988 969
rect 826 964 830 965
rect 901 964 904 965
rect 926 964 927 965
rect 822 962 826 964
rect 436 945 446 946
rect 468 945 469 946
rect 432 943 436 945
rect 480 943 500 946
rect 581 943 582 950
rect 654 943 655 950
rect 789 949 822 962
rect 906 959 910 962
rect 921 960 925 963
rect 1030 962 1039 971
rect 1063 961 1066 963
rect 1077 962 1086 971
rect 1371 970 1405 972
rect 1414 971 1415 972
rect 1461 971 1464 974
rect 1410 970 1415 971
rect 1460 970 1461 971
rect 1371 968 1415 970
rect 1458 969 1460 970
rect 1367 965 1368 967
rect 1141 961 1150 963
rect 1058 959 1063 961
rect 703 943 709 949
rect 749 948 755 949
rect 786 948 789 949
rect 749 947 786 948
rect 749 943 755 947
rect 841 946 847 952
rect 887 946 893 952
rect 909 949 910 959
rect 1056 958 1058 959
rect 1152 958 1158 961
rect 927 955 931 958
rect 995 955 997 958
rect 931 946 941 955
rect 420 931 428 943
rect 432 941 466 943
rect 156 924 157 929
rect 106 915 115 924
rect 153 920 162 924
rect 153 915 167 920
rect 97 912 106 915
rect 97 911 100 912
rect 90 908 99 911
rect 78 907 99 908
rect 78 905 96 907
rect 136 905 142 911
rect 156 906 171 915
rect 196 908 203 929
rect 78 900 90 905
rect 74 898 77 900
rect 78 899 79 900
rect 84 899 90 900
rect 142 899 148 905
rect 155 904 167 906
rect 194 904 196 908
rect 234 907 240 929
rect 291 926 292 929
rect 318 928 379 931
rect 318 917 324 928
rect 346 926 379 928
rect 340 925 379 926
rect 398 925 404 926
rect 340 921 404 925
rect 340 920 426 921
rect 318 913 327 917
rect 346 914 352 920
rect 392 914 398 920
rect 401 917 426 920
rect 410 913 426 917
rect 432 913 434 941
rect 463 939 466 941
rect 318 909 333 913
rect 420 909 434 913
rect 464 909 466 939
rect 470 931 478 943
rect 500 934 563 943
rect 697 938 703 943
rect 715 941 751 943
rect 715 938 720 941
rect 656 937 703 938
rect 717 937 720 938
rect 755 937 761 943
rect 835 940 841 946
rect 893 940 899 946
rect 656 936 699 937
rect 580 934 581 936
rect 602 934 656 936
rect 536 922 551 934
rect 563 933 602 934
rect 580 929 581 933
rect 712 929 715 936
rect 839 933 841 934
rect 837 929 839 933
rect 233 904 234 906
rect 293 905 294 909
rect 153 899 155 904
rect 299 903 305 909
rect 318 903 337 909
rect 345 903 351 909
rect 193 899 194 903
rect 152 897 153 899
rect 192 897 193 899
rect 66 884 74 896
rect 78 894 96 896
rect 151 895 152 896
rect 231 895 233 903
rect 293 897 299 903
rect 318 897 357 903
rect 359 897 371 905
rect 432 904 449 909
rect 440 899 447 904
rect 449 903 453 904
rect 469 903 470 905
rect 536 904 551 920
rect 578 906 580 928
rect 453 900 472 903
rect 577 900 589 905
rect 599 900 611 905
rect 652 904 654 928
rect 703 904 712 928
rect 748 904 751 909
rect 789 908 824 910
rect 835 908 837 929
rect 859 909 860 929
rect 907 928 909 944
rect 941 942 946 946
rect 997 942 1009 955
rect 1158 951 1171 958
rect 1381 956 1397 968
rect 1399 956 1415 968
rect 1454 965 1458 968
rect 1452 963 1454 965
rect 1450 961 1452 963
rect 1505 961 1518 974
rect 1554 967 1557 983
rect 1556 961 1557 967
rect 1560 967 1561 989
rect 1599 985 1606 989
rect 1627 987 1629 990
rect 1599 983 1600 985
rect 1620 984 1621 986
rect 1560 963 1562 967
rect 1593 963 1594 966
rect 1598 965 1600 983
rect 1629 981 1632 987
rect 1632 979 1633 981
rect 1634 975 1635 977
rect 1635 972 1636 975
rect 1675 973 1683 990
rect 1637 965 1640 969
rect 1560 961 1564 963
rect 1598 962 1599 965
rect 1640 963 1641 965
rect 1446 958 1449 961
rect 1518 959 1521 961
rect 1444 953 1446 958
rect 1521 957 1523 959
rect 1279 952 1316 953
rect 1443 952 1444 953
rect 1523 952 1525 957
rect 1551 955 1557 961
rect 1564 959 1570 961
rect 1571 957 1577 959
rect 1597 957 1603 961
rect 1641 960 1642 963
rect 1642 958 1643 960
rect 1577 956 1603 957
rect 1279 951 1304 952
rect 1316 951 1317 952
rect 1173 948 1177 951
rect 1244 948 1271 951
rect 1319 948 1326 951
rect 1371 949 1372 952
rect 1442 951 1443 952
rect 1326 943 1337 948
rect 1372 945 1374 949
rect 1407 947 1408 949
rect 1440 948 1442 951
rect 1337 942 1341 943
rect 1009 939 1010 942
rect 1341 938 1348 942
rect 951 929 961 938
rect 1011 931 1017 938
rect 1348 937 1350 938
rect 1350 933 1366 937
rect 1366 932 1371 933
rect 1374 932 1382 944
rect 1371 929 1382 932
rect 1408 929 1412 944
rect 1438 943 1440 948
rect 1525 944 1528 951
rect 1545 949 1551 955
rect 1577 951 1621 956
rect 1643 955 1645 958
rect 1603 949 1609 951
rect 1645 948 1648 955
rect 1437 942 1438 943
rect 1648 942 1651 948
rect 1683 943 1684 973
rect 1791 951 1807 954
rect 1719 943 1742 951
rect 1797 943 1814 951
rect 1436 940 1437 942
rect 1435 939 1436 940
rect 1651 939 1652 942
rect 1434 937 1435 938
rect 1431 933 1434 937
rect 1429 932 1431 933
rect 1427 929 1429 932
rect 1652 931 1653 938
rect 1682 929 1683 942
rect 1711 938 1719 943
rect 1797 938 1821 943
rect 1701 932 1711 938
rect 1694 929 1701 932
rect 904 917 906 920
rect 900 914 903 916
rect 898 913 900 914
rect 895 911 898 913
rect 893 910 895 911
rect 779 906 789 908
rect 824 906 841 908
rect 768 904 779 906
rect 702 900 703 903
rect 746 900 748 904
rect 760 902 768 904
rect 756 901 760 902
rect 835 900 837 906
rect 859 904 860 906
rect 927 904 943 920
rect 961 910 983 929
rect 1021 920 1029 927
rect 1029 918 1036 920
rect 1036 914 1052 918
rect 1055 914 1056 929
rect 1374 928 1387 929
rect 1380 927 1387 928
rect 1412 927 1413 928
rect 1426 927 1427 929
rect 1550 927 1551 929
rect 1382 923 1383 926
rect 1387 924 1424 927
rect 1114 921 1145 922
rect 1105 920 1114 921
rect 1145 920 1152 921
rect 1412 920 1413 924
rect 1076 917 1105 920
rect 1152 917 1167 920
rect 1074 916 1076 917
rect 1067 914 1074 916
rect 1167 914 1179 917
rect 1384 915 1385 917
rect 1413 915 1414 920
rect 1418 915 1427 924
rect 1465 915 1474 924
rect 1549 922 1550 927
rect 1548 920 1549 922
rect 1547 918 1548 920
rect 1546 916 1547 918
rect 1409 914 1418 915
rect 1052 911 1418 914
rect 1055 910 1056 911
rect 1058 910 1060 911
rect 1194 910 1202 911
rect 983 909 985 910
rect 860 900 864 904
rect 914 900 927 904
rect 985 903 993 909
rect 1054 908 1058 910
rect 1202 906 1220 910
rect 1385 906 1386 909
rect 1415 906 1416 909
rect 1047 904 1052 906
rect 318 895 373 897
rect 447 895 453 899
rect 467 898 468 900
rect 466 895 467 897
rect 472 896 641 900
rect 700 897 702 900
rect 697 896 703 897
rect 743 896 746 900
rect 577 895 578 896
rect 641 895 703 896
rect 66 862 74 874
rect 78 865 80 894
rect 150 893 151 894
rect 191 893 192 894
rect 318 893 375 895
rect 453 893 454 895
rect 145 889 151 893
rect 190 889 191 893
rect 230 889 231 893
rect 286 889 293 893
rect 318 892 383 893
rect 131 888 151 889
rect 131 878 145 888
rect 187 879 190 889
rect 228 878 230 889
rect 283 879 286 889
rect 115 866 131 878
rect 78 862 81 865
rect 112 862 115 866
rect 162 859 171 868
rect 183 866 187 878
rect 227 875 228 878
rect 282 875 283 878
rect 182 862 183 866
rect 77 857 79 858
rect 84 857 90 859
rect 78 853 90 857
rect 142 853 148 859
rect 154 857 162 859
rect 181 858 182 862
rect 223 859 227 875
rect 277 859 282 875
rect 295 864 298 892
rect 345 891 371 892
rect 369 861 371 891
rect 375 881 383 892
rect 454 879 474 893
rect 522 879 536 894
rect 565 881 573 893
rect 577 891 611 893
rect 430 876 431 879
rect 460 876 461 879
rect 474 877 486 879
rect 520 877 522 879
rect 474 875 520 877
rect 345 859 371 861
rect 375 859 383 871
rect 428 869 430 875
rect 458 870 460 875
rect 426 862 428 869
rect 455 862 458 869
rect 425 859 426 862
rect 454 859 455 862
rect 577 859 579 891
rect 609 875 611 891
rect 615 881 623 893
rect 697 891 703 895
rect 741 891 743 895
rect 755 891 761 897
rect 835 894 841 900
rect 864 896 879 900
rect 879 895 880 896
rect 893 895 927 900
rect 993 899 999 903
rect 1044 902 1047 904
rect 1220 902 1240 906
rect 1311 902 1324 903
rect 651 881 652 889
rect 695 881 698 891
rect 703 885 709 891
rect 735 881 741 891
rect 749 885 755 891
rect 838 883 839 891
rect 841 888 847 894
rect 880 893 899 895
rect 610 865 611 874
rect 615 872 616 875
rect 645 870 651 880
rect 690 870 695 881
rect 633 866 645 870
rect 689 867 690 870
rect 728 867 735 881
rect 878 872 881 892
rect 887 888 893 893
rect 911 888 927 895
rect 999 894 1010 899
rect 1038 898 1042 900
rect 1035 897 1038 898
rect 1032 895 1035 897
rect 1055 895 1058 900
rect 1240 897 1265 902
rect 1290 900 1308 902
rect 1329 900 1352 902
rect 1288 899 1300 900
rect 1352 899 1361 900
rect 1361 898 1362 899
rect 1386 898 1387 902
rect 1265 895 1270 897
rect 1281 895 1288 898
rect 1010 885 1041 894
rect 1058 893 1060 895
rect 1060 891 1062 893
rect 1270 891 1288 895
rect 1362 894 1369 898
rect 1416 897 1417 902
rect 1474 901 1483 915
rect 1544 911 1545 914
rect 1571 909 1603 913
rect 1538 903 1542 906
rect 1545 903 1551 909
rect 1571 904 1609 909
rect 1640 904 1694 929
rect 1797 922 1823 938
rect 1568 903 1609 904
rect 1525 901 1537 902
rect 1483 899 1487 901
rect 1505 900 1525 901
rect 1499 899 1505 900
rect 1525 895 1527 900
rect 1551 897 1557 903
rect 1585 899 1586 901
rect 1369 891 1375 894
rect 1387 891 1388 895
rect 1000 880 1041 885
rect 1062 888 1135 891
rect 1270 889 1287 891
rect 1062 885 1142 888
rect 1062 881 1135 885
rect 1142 881 1212 885
rect 1273 882 1281 889
rect 1287 887 1292 889
rect 1292 885 1296 887
rect 1375 885 1388 891
rect 1417 887 1419 895
rect 1523 892 1525 895
rect 1522 891 1523 892
rect 1000 876 1016 880
rect 1041 876 1059 880
rect 1062 876 1080 881
rect 1135 876 1240 881
rect 1059 875 1240 876
rect 1266 875 1273 882
rect 1296 876 1318 885
rect 1375 882 1389 885
rect 1388 881 1391 882
rect 1388 878 1389 881
rect 1391 880 1392 881
rect 1392 879 1401 880
rect 1419 879 1421 885
rect 1510 882 1522 891
rect 1504 881 1510 882
rect 1476 880 1492 881
rect 1500 880 1504 881
rect 1569 880 1584 899
rect 1597 897 1603 903
rect 1634 901 1640 904
rect 1648 903 1649 904
rect 1623 895 1634 901
rect 1647 899 1648 901
rect 1620 892 1623 895
rect 1619 891 1620 892
rect 1611 885 1619 891
rect 1448 879 1471 880
rect 1318 875 1321 876
rect 727 866 728 867
rect 632 865 633 866
rect 610 862 632 865
rect 686 862 689 866
rect 611 859 632 862
rect 683 859 689 862
rect 153 855 162 857
rect 78 852 87 853
rect 78 850 88 852
rect 90 850 96 853
rect 88 847 96 850
rect 88 842 92 847
rect 141 840 142 853
rect 151 852 162 855
rect 149 851 151 852
rect 146 850 149 851
rect 153 850 162 852
rect 177 845 181 858
rect 220 846 223 858
rect 273 846 277 858
rect 293 851 299 857
rect 322 856 326 859
rect 616 858 617 859
rect 299 845 305 851
rect 317 845 322 856
rect 351 851 357 857
rect 424 855 425 858
rect 453 855 454 858
rect 683 857 686 859
rect 685 856 686 857
rect 681 855 685 856
rect 345 845 351 851
rect 359 847 371 855
rect 575 853 576 855
rect 173 841 177 845
rect 219 841 220 845
rect 271 842 273 845
rect 171 840 173 841
rect 315 840 317 845
rect 419 841 422 850
rect 449 841 452 850
rect 576 841 578 849
rect 617 842 618 849
rect 678 847 685 855
rect 672 845 679 847
rect 681 845 685 847
rect 715 845 727 865
rect 839 859 841 872
rect 672 840 681 845
rect 712 844 719 845
rect 874 844 878 870
rect 989 869 999 875
rect 1052 872 1252 875
rect 1263 872 1266 875
rect 1321 872 1331 875
rect 1337 872 1349 878
rect 1392 875 1471 879
rect 1599 876 1631 885
rect 1644 880 1647 898
rect 1643 876 1644 880
rect 1679 878 1681 904
rect 1797 895 1820 922
rect 1852 895 1853 929
rect 1797 881 1819 895
rect 1831 889 1853 895
rect 1052 871 1060 872
rect 1047 869 1051 871
rect 987 868 989 869
rect 984 866 987 868
rect 1042 866 1046 868
rect 1135 867 1359 872
rect 1389 871 1390 875
rect 1401 871 1448 875
rect 1562 872 1565 876
rect 1596 875 1631 876
rect 1407 869 1448 871
rect 1413 868 1438 869
rect 1151 866 1359 867
rect 977 862 984 866
rect 1032 862 1042 866
rect 1151 863 1361 866
rect 1264 862 1273 863
rect 1347 862 1369 863
rect 1390 862 1391 868
rect 1414 867 1438 868
rect 1554 863 1562 872
rect 1609 869 1610 874
rect 971 858 977 862
rect 1273 858 1280 862
rect 969 857 971 858
rect 960 852 969 857
rect 1280 852 1291 858
rect 1347 854 1361 862
rect 1369 856 1402 862
rect 1421 859 1422 862
rect 1550 857 1554 862
rect 1477 856 1489 857
rect 1402 855 1408 856
rect 1426 855 1448 856
rect 1408 854 1448 855
rect 1469 854 1489 856
rect 955 850 960 852
rect 1291 850 1295 852
rect 920 849 926 850
rect 953 849 955 850
rect 902 844 953 849
rect 966 844 972 850
rect 1016 845 1019 849
rect 1296 845 1304 849
rect 1347 846 1359 854
rect 1477 852 1509 854
rect 1392 850 1393 852
rect 1422 850 1423 852
rect 1478 847 1509 852
rect 1547 849 1549 856
rect 1547 847 1548 849
rect 712 840 716 844
rect 93 836 94 840
rect 94 833 95 836
rect 141 832 143 840
rect 159 832 171 840
rect 218 838 219 840
rect 270 838 271 840
rect 217 832 218 838
rect 269 833 270 838
rect 312 832 315 840
rect 418 837 419 840
rect 417 833 418 836
rect 446 834 448 840
rect 618 837 619 840
rect 579 832 583 837
rect 670 832 679 840
rect 708 834 716 840
rect 708 832 712 834
rect 95 817 103 832
rect 141 825 145 832
rect 157 828 159 832
rect 216 828 217 832
rect 267 828 268 832
rect 143 817 145 825
rect 154 819 157 828
rect 214 819 216 828
rect 265 824 267 827
rect 261 820 267 824
rect 103 809 107 817
rect 145 811 146 817
rect 153 815 154 819
rect 213 815 214 819
rect 261 815 265 820
rect 307 819 312 832
rect 152 809 153 814
rect 211 809 213 814
rect 261 809 263 815
rect 304 814 307 818
rect 357 814 373 824
rect 375 814 391 824
rect 411 817 417 832
rect 300 809 304 814
rect 344 809 351 814
rect 396 808 404 814
rect 409 811 411 817
rect 439 811 446 832
rect 580 827 584 832
rect 619 827 625 832
rect 438 809 439 811
rect 453 808 469 824
rect 569 822 635 827
rect 655 824 670 832
rect 569 821 625 822
rect 560 814 569 821
rect 580 818 584 821
rect 476 808 495 809
rect 501 808 503 809
rect 108 804 109 807
rect 109 799 111 803
rect 146 799 147 803
rect 149 800 152 808
rect 209 800 211 808
rect 111 794 113 798
rect 149 794 151 800
rect 207 794 209 798
rect 114 785 117 793
rect 148 790 150 793
rect 151 790 165 794
rect 148 786 165 790
rect 117 775 122 785
rect 122 771 123 775
rect 149 774 165 786
rect 199 790 207 794
rect 245 792 261 808
rect 295 801 300 808
rect 340 801 344 808
rect 396 807 407 808
rect 437 807 453 808
rect 503 807 504 808
rect 552 807 560 814
rect 583 811 584 817
rect 619 811 625 821
rect 635 814 639 821
rect 653 819 670 824
rect 701 819 708 832
rect 710 828 712 832
rect 841 832 843 844
rect 853 840 865 844
rect 881 842 902 844
rect 872 841 881 842
rect 867 840 874 841
rect 853 836 867 840
rect 653 818 655 819
rect 653 815 654 818
rect 699 817 701 819
rect 698 816 699 817
rect 639 812 643 814
rect 652 812 653 813
rect 698 812 701 816
rect 731 812 743 815
rect 625 809 626 811
rect 580 808 582 809
rect 639 808 650 812
rect 697 808 698 812
rect 731 808 747 812
rect 749 808 765 824
rect 767 808 783 824
rect 841 820 849 832
rect 853 831 869 832
rect 853 830 863 831
rect 785 808 794 812
rect 844 810 845 814
rect 569 807 579 808
rect 396 806 408 807
rect 403 804 408 806
rect 436 804 453 807
rect 504 806 507 807
rect 295 792 299 801
rect 199 774 215 790
rect 245 774 261 790
rect 295 787 311 790
rect 290 781 311 787
rect 331 787 340 801
rect 403 792 407 804
rect 435 799 436 803
rect 433 794 435 798
rect 437 792 453 804
rect 476 798 488 806
rect 507 804 510 806
rect 540 804 569 807
rect 491 799 540 804
rect 541 799 547 804
rect 552 799 560 804
rect 626 799 628 804
rect 637 803 652 808
rect 697 806 702 808
rect 731 807 748 808
rect 753 807 765 808
rect 331 785 342 787
rect 351 785 363 791
rect 403 785 404 792
rect 431 788 433 792
rect 320 783 342 785
rect 352 783 363 785
rect 402 783 407 785
rect 314 781 319 783
rect 284 775 290 781
rect 295 774 311 781
rect 329 779 331 783
rect 336 781 342 783
rect 363 781 367 783
rect 342 775 348 781
rect 351 778 363 779
rect 151 771 155 774
rect 123 754 131 771
rect 155 754 162 771
rect 165 758 181 774
rect 183 758 199 774
rect 261 772 269 774
rect 287 772 295 774
rect 361 772 363 778
rect 367 772 375 779
rect 400 778 402 783
rect 403 778 407 783
rect 400 774 407 778
rect 400 772 402 774
rect 261 758 277 772
rect 279 758 295 772
rect 342 757 405 772
rect 429 760 431 786
rect 437 774 453 790
rect 464 782 472 794
rect 476 793 497 794
rect 535 793 541 799
rect 476 792 494 793
rect 453 763 457 767
rect 464 763 472 772
rect 476 763 478 792
rect 629 788 631 796
rect 637 794 659 803
rect 637 792 652 794
rect 689 792 702 806
rect 727 804 729 807
rect 733 806 747 807
rect 731 803 747 806
rect 783 805 799 808
rect 781 803 799 805
rect 689 790 697 792
rect 719 791 727 803
rect 729 801 765 803
rect 729 793 749 801
rect 762 800 765 801
rect 763 793 765 800
rect 769 799 777 803
rect 781 799 803 803
rect 783 794 803 799
rect 841 798 849 810
rect 853 800 855 830
rect 872 826 874 840
rect 914 838 920 844
rect 972 838 978 844
rect 1011 841 1016 845
rect 1304 841 1309 845
rect 1303 832 1311 841
rect 1315 834 1317 839
rect 1347 834 1349 846
rect 1607 845 1609 865
rect 1641 863 1643 872
rect 1678 863 1679 872
rect 1797 868 1814 881
rect 1842 868 1847 872
rect 1797 866 1806 868
rect 1797 865 1805 866
rect 1831 865 1839 866
rect 1640 857 1641 862
rect 1638 849 1639 855
rect 1359 844 1367 845
rect 1315 832 1349 834
rect 1353 832 1367 844
rect 887 826 888 832
rect 1359 830 1367 832
rect 998 829 1001 830
rect 974 827 1009 829
rect 872 818 873 826
rect 970 825 974 827
rect 873 800 876 814
rect 888 812 890 825
rect 941 808 970 825
rect 972 814 974 817
rect 982 812 998 827
rect 977 811 998 812
rect 1009 824 1169 827
rect 853 798 887 800
rect 873 795 876 798
rect 631 778 634 788
rect 634 769 636 778
rect 637 774 652 790
rect 689 774 703 790
rect 726 781 727 788
rect 636 765 637 769
rect 453 762 478 763
rect 507 762 510 763
rect 453 760 510 762
rect 453 758 469 760
rect 637 759 638 763
rect 131 746 134 754
rect 162 748 167 754
rect 167 745 171 748
rect 361 745 363 757
rect 366 745 400 757
rect 405 756 407 757
rect 514 756 541 759
rect 638 757 639 759
rect 653 758 669 772
rect 671 758 687 772
rect 719 769 727 781
rect 731 774 749 793
rect 783 792 799 794
rect 783 774 799 790
rect 829 774 844 790
rect 846 775 848 789
rect 853 786 865 794
rect 875 786 887 794
rect 889 790 890 808
rect 976 805 986 811
rect 1009 808 1175 824
rect 1237 808 1253 824
rect 1255 808 1271 824
rect 1315 820 1327 828
rect 1337 820 1349 828
rect 1315 810 1317 820
rect 1367 816 1371 830
rect 1393 828 1395 845
rect 1395 819 1396 828
rect 1423 819 1426 845
rect 1428 843 1477 845
rect 1512 843 1514 844
rect 1428 833 1470 843
rect 1548 838 1549 843
rect 1515 827 1516 836
rect 1549 827 1550 836
rect 1606 834 1607 844
rect 1637 843 1638 847
rect 1636 837 1637 843
rect 1465 811 1470 823
rect 1517 817 1518 820
rect 1550 816 1551 820
rect 1605 819 1606 832
rect 1634 827 1636 836
rect 1676 829 1678 862
rect 1789 855 1805 865
rect 1842 864 1846 868
rect 1726 845 1789 855
rect 1834 851 1842 864
rect 1717 844 1726 845
rect 1711 842 1717 844
rect 1701 834 1711 842
rect 1633 821 1634 826
rect 1674 820 1676 827
rect 1518 811 1519 814
rect 1551 811 1552 814
rect 1604 811 1605 818
rect 1618 811 1624 817
rect 1632 816 1633 820
rect 1673 818 1674 820
rect 1681 818 1701 834
rect 1631 814 1632 816
rect 1630 812 1631 814
rect 1664 811 1670 817
rect 1672 813 1681 818
rect 1671 811 1681 813
rect 1427 808 1428 810
rect 1519 808 1520 810
rect 981 803 986 805
rect 1106 803 1115 808
rect 1153 803 1162 808
rect 893 802 902 803
rect 891 798 899 802
rect 902 799 917 802
rect 917 798 920 799
rect 914 792 920 798
rect 972 792 978 798
rect 986 794 995 803
rect 1097 794 1106 803
rect 1162 794 1171 803
rect 1088 792 1095 793
rect 920 790 926 792
rect 731 772 765 774
rect 778 772 783 774
rect 876 772 879 786
rect 889 774 895 790
rect 920 786 941 790
rect 966 786 972 792
rect 1082 791 1088 792
rect 1139 791 1143 793
rect 1175 792 1191 808
rect 1221 792 1237 808
rect 1248 803 1254 808
rect 1248 802 1263 803
rect 1242 796 1248 802
rect 1271 798 1287 808
rect 1294 802 1300 808
rect 1247 791 1248 793
rect 1280 791 1285 798
rect 1300 796 1306 802
rect 1318 800 1319 808
rect 1080 790 1082 791
rect 1079 787 1080 790
rect 1144 789 1146 790
rect 925 774 941 786
rect 992 778 1019 781
rect 975 774 992 778
rect 1019 774 1027 778
rect 731 769 783 772
rect 844 769 850 772
rect 879 771 883 772
rect 731 757 735 765
rect 767 758 783 769
rect 845 762 862 769
rect 879 762 889 771
rect 845 758 861 762
rect 862 760 867 762
rect 871 760 883 762
rect 867 759 883 760
rect 863 758 883 759
rect 941 758 957 774
rect 1027 772 1030 774
rect 1095 772 1101 778
rect 1104 772 1106 779
rect 1146 772 1147 778
rect 1175 774 1191 790
rect 1221 774 1237 790
rect 1239 779 1248 791
rect 1030 763 1050 772
rect 1079 767 1080 769
rect 1089 766 1095 772
rect 1147 766 1153 772
rect 1168 763 1175 774
rect 1050 762 1052 763
rect 1052 759 1058 762
rect 407 751 428 756
rect 428 747 444 751
rect 476 748 488 756
rect 639 754 640 756
rect 535 747 541 753
rect 566 747 621 753
rect 640 750 641 754
rect 641 747 643 748
rect 650 747 659 756
rect 729 747 735 756
rect 787 747 793 753
rect 794 747 803 756
rect 848 751 851 758
rect 134 741 136 745
rect 171 740 179 745
rect 397 742 398 745
rect 444 742 464 747
rect 464 741 469 742
rect 541 741 547 747
rect 587 741 593 747
rect 363 740 365 741
rect 136 737 138 740
rect 179 737 184 740
rect 353 739 363 740
rect 342 738 363 739
rect 469 738 473 741
rect 594 738 603 747
rect 641 745 650 747
rect 641 742 656 745
rect 641 738 650 742
rect 656 740 660 742
rect 735 741 747 747
rect 781 741 794 747
rect 850 744 851 751
rect 660 739 663 740
rect 184 736 186 737
rect 351 736 370 738
rect 139 733 140 736
rect 186 733 190 736
rect 140 727 143 733
rect 190 731 194 733
rect 194 729 197 731
rect 284 729 290 735
rect 342 729 348 735
rect 351 733 388 736
rect 395 733 396 736
rect 362 729 388 733
rect 391 729 395 731
rect 427 729 428 730
rect 197 726 201 729
rect 143 720 147 726
rect 201 720 211 726
rect 214 720 226 724
rect 290 723 296 729
rect 336 723 342 729
rect 388 726 428 729
rect 388 723 427 726
rect 473 725 490 738
rect 594 737 595 738
rect 663 736 670 739
rect 738 738 747 741
rect 785 738 794 741
rect 844 739 851 744
rect 879 742 883 758
rect 921 747 930 756
rect 986 747 995 756
rect 1058 754 1069 759
rect 1162 758 1175 763
rect 1237 769 1246 774
rect 1247 769 1248 779
rect 1237 763 1248 769
rect 1251 763 1253 791
rect 1319 790 1321 791
rect 1317 785 1321 790
rect 1370 790 1371 808
rect 1477 799 1489 804
rect 1521 796 1522 799
rect 1552 796 1553 805
rect 1603 799 1604 808
rect 1612 805 1618 811
rect 1670 808 1676 811
rect 1725 808 1741 824
rect 1668 805 1676 808
rect 1668 804 1670 805
rect 1671 800 1672 802
rect 1672 797 1674 800
rect 1237 758 1253 763
rect 1302 773 1363 785
rect 1370 779 1383 790
rect 1369 774 1383 779
rect 1413 774 1428 790
rect 1429 777 1431 793
rect 1522 789 1523 793
rect 1553 789 1554 795
rect 1302 759 1367 773
rect 1333 758 1349 759
rect 1351 758 1367 759
rect 1394 758 1395 760
rect 1429 758 1445 774
rect 1523 767 1527 785
rect 1554 779 1555 788
rect 1603 787 1605 794
rect 1668 790 1669 794
rect 1674 791 1677 797
rect 1709 792 1725 808
rect 1759 802 1787 808
rect 1753 794 1787 802
rect 1749 791 1751 794
rect 1759 790 1787 794
rect 1605 781 1606 787
rect 1668 782 1685 790
rect 1555 766 1560 779
rect 1607 774 1615 780
rect 1669 776 1685 782
rect 1741 779 1749 790
rect 1738 778 1749 779
rect 1753 788 1787 790
rect 1669 774 1679 776
rect 1615 773 1617 774
rect 1527 760 1528 766
rect 1560 759 1562 766
rect 1617 765 1631 773
rect 1669 766 1670 774
rect 1685 768 1690 776
rect 1738 770 1747 778
rect 1666 765 1670 766
rect 1612 764 1645 765
rect 1666 764 1676 765
rect 1612 759 1618 764
rect 1162 756 1168 758
rect 1239 757 1253 758
rect 1365 757 1368 758
rect 1247 756 1300 757
rect 1080 754 1081 756
rect 1162 754 1171 756
rect 844 738 850 739
rect 890 738 896 744
rect 930 738 939 747
rect 977 738 986 747
rect 1069 746 1083 754
rect 1157 747 1171 754
rect 1242 750 1306 756
rect 1369 750 1384 756
rect 1391 754 1392 756
rect 1433 752 1434 753
rect 1157 746 1162 747
rect 1083 745 1086 746
rect 596 734 597 736
rect 598 727 601 733
rect 670 731 685 736
rect 838 732 844 738
rect 896 733 902 738
rect 950 734 962 738
rect 1003 734 1019 744
rect 1081 742 1082 745
rect 1086 742 1125 745
rect 1155 743 1162 746
rect 1248 745 1263 750
rect 1294 747 1303 750
rect 1248 744 1254 745
rect 1294 744 1300 747
rect 1082 740 1125 742
rect 1086 737 1125 740
rect 1148 739 1155 743
rect 1157 739 1162 743
rect 1303 742 1317 747
rect 1384 745 1397 750
rect 1433 747 1441 752
rect 1529 751 1530 756
rect 1563 750 1566 756
rect 1618 753 1624 759
rect 1629 758 1645 764
rect 1647 758 1663 764
rect 1670 759 1676 764
rect 1690 762 1693 768
rect 1729 761 1738 770
rect 1664 753 1670 759
rect 1695 756 1697 760
rect 1725 757 1726 758
rect 1383 742 1385 745
rect 1397 742 1403 745
rect 1434 744 1441 747
rect 1530 746 1531 750
rect 1566 744 1568 750
rect 1652 745 1655 747
rect 1443 742 1444 744
rect 1697 743 1705 756
rect 1726 754 1729 757
rect 1741 756 1749 768
rect 1753 758 1755 788
rect 1784 787 1787 788
rect 1791 779 1834 791
rect 1785 776 1834 779
rect 1785 770 1794 776
rect 1805 774 1821 776
rect 1834 774 1855 776
rect 1794 764 1803 770
rect 1797 763 1803 764
rect 1821 768 1855 774
rect 1798 759 1801 763
rect 1821 758 1837 768
rect 1855 762 1872 768
rect 1858 758 1864 762
rect 1872 760 1878 762
rect 1878 758 1882 760
rect 1904 758 1910 764
rect 1753 757 1768 758
rect 1753 756 1772 757
rect 1729 750 1734 754
rect 1769 752 1787 756
rect 1804 753 1810 756
rect 1852 753 1858 758
rect 1753 750 1787 752
rect 1810 751 1858 753
rect 1910 752 1916 758
rect 1734 749 1770 750
rect 1753 744 1765 749
rect 1820 744 1831 749
rect 1831 743 1833 744
rect 1317 739 1326 742
rect 1403 741 1405 742
rect 1705 741 1706 743
rect 1148 738 1162 739
rect 1135 737 1148 738
rect 1155 735 1157 738
rect 1326 735 1337 739
rect 1380 737 1381 739
rect 1337 734 1340 735
rect 946 733 1028 734
rect 896 732 962 733
rect 939 731 962 732
rect 685 726 697 731
rect 939 729 946 731
rect 950 730 962 731
rect 1028 729 1031 732
rect 1147 731 1154 734
rect 1340 731 1349 734
rect 1377 733 1379 736
rect 1349 729 1356 731
rect 1372 729 1376 731
rect 935 728 939 729
rect 928 726 935 728
rect 965 727 966 729
rect 1031 728 1033 729
rect 387 721 458 723
rect 211 719 226 720
rect 388 719 458 721
rect 490 719 494 725
rect 601 723 603 726
rect 214 716 226 719
rect 150 712 155 716
rect 227 714 230 716
rect 379 712 387 719
rect 389 717 399 719
rect 389 712 393 717
rect 155 696 176 712
rect 220 710 244 712
rect 224 705 244 710
rect 379 707 389 712
rect 386 705 389 707
rect 176 695 178 696
rect 182 689 183 692
rect 180 678 187 687
rect 224 680 226 705
rect 230 700 238 705
rect 244 699 250 705
rect 384 701 386 705
rect 378 699 386 701
rect 250 694 256 699
rect 378 695 384 699
rect 256 692 259 694
rect 192 678 226 680
rect 230 678 238 690
rect 259 688 260 692
rect 372 689 378 695
rect 382 692 383 694
rect 381 688 382 691
rect 391 689 393 712
rect 423 715 478 719
rect 423 701 446 715
rect 454 713 478 715
rect 498 713 499 715
rect 459 708 478 713
rect 499 708 503 713
rect 603 710 610 723
rect 697 722 727 726
rect 946 724 962 726
rect 697 714 739 722
rect 466 701 478 708
rect 503 706 504 708
rect 610 705 613 710
rect 691 709 740 710
rect 423 695 430 701
rect 423 693 436 695
rect 423 689 425 693
rect 430 689 436 693
rect 441 691 450 700
rect 469 696 478 701
rect 509 696 512 701
rect 472 691 478 696
rect 380 685 381 687
rect 424 685 425 689
rect 442 687 459 691
rect 475 689 478 691
rect 512 689 518 696
rect 613 695 650 705
rect 691 702 705 709
rect 721 708 740 709
rect 737 703 740 708
rect 690 699 691 701
rect 650 693 656 695
rect 688 694 690 699
rect 656 692 661 693
rect 687 692 688 694
rect 477 687 478 689
rect 443 686 459 687
rect 518 686 520 689
rect 661 688 677 692
rect 677 687 679 688
rect 260 680 262 685
rect 379 680 380 685
rect 445 682 448 686
rect 450 682 459 686
rect 451 680 452 682
rect 187 676 188 678
rect 191 676 192 678
rect 378 676 379 678
rect 452 677 453 680
rect 187 660 191 676
rect 227 674 230 676
rect 192 666 204 674
rect 214 666 226 674
rect 262 660 266 676
rect 186 654 187 658
rect 266 657 267 660
rect 186 630 188 654
rect 266 630 267 654
rect 378 649 430 663
rect 451 662 453 675
rect 480 672 492 685
rect 520 672 532 686
rect 682 685 688 687
rect 688 683 696 685
rect 693 681 697 683
rect 693 676 700 681
rect 737 678 739 703
rect 740 697 741 702
rect 743 698 751 710
rect 896 694 924 695
rect 960 694 962 724
rect 966 714 974 726
rect 1033 712 1035 728
rect 1356 727 1362 729
rect 1369 727 1372 729
rect 1089 720 1095 726
rect 1147 720 1153 726
rect 1353 723 1373 727
rect 1405 723 1426 741
rect 1431 738 1442 740
rect 1353 721 1369 723
rect 1348 720 1353 721
rect 1373 720 1381 723
rect 1095 714 1101 720
rect 1141 714 1147 720
rect 1341 717 1348 720
rect 1381 719 1384 720
rect 1426 719 1431 723
rect 1336 716 1341 717
rect 1384 716 1390 719
rect 1431 716 1435 719
rect 1439 716 1441 738
rect 1442 737 1443 738
rect 1445 737 1453 740
rect 1443 734 1453 737
rect 1445 729 1453 734
rect 1532 733 1533 741
rect 1569 737 1572 741
rect 1533 729 1534 733
rect 1562 729 1574 737
rect 1584 729 1596 737
rect 1659 729 1672 741
rect 1445 728 1454 729
rect 1450 726 1454 728
rect 1445 716 1453 718
rect 1327 713 1336 716
rect 1322 711 1327 713
rect 741 693 742 694
rect 916 692 924 694
rect 928 692 962 694
rect 966 692 974 704
rect 1033 694 1035 710
rect 1306 706 1322 711
rect 1390 706 1401 716
rect 1435 707 1453 716
rect 1417 706 1453 707
rect 1454 706 1477 726
rect 1534 724 1541 729
rect 1558 727 1561 729
rect 1574 725 1575 729
rect 1581 725 1587 729
rect 1535 723 1541 724
rect 1550 723 1558 725
rect 1562 723 1608 725
rect 1529 717 1535 723
rect 1562 717 1564 723
rect 1587 717 1593 723
rect 1594 717 1608 723
rect 1533 713 1535 714
rect 1531 709 1533 713
rect 1290 701 1306 706
rect 1401 705 1408 706
rect 1446 705 1479 706
rect 1401 702 1409 705
rect 1383 701 1417 702
rect 1443 701 1504 705
rect 1594 702 1596 717
rect 1600 713 1615 717
rect 1603 705 1615 713
rect 1672 712 1691 729
rect 1706 715 1740 741
rect 1835 723 1858 741
rect 1694 706 1704 709
rect 1705 706 1717 715
rect 1740 714 1742 715
rect 1742 709 1782 714
rect 1804 709 1816 714
rect 1782 707 1816 709
rect 1782 706 1830 707
rect 1852 706 1858 712
rect 1910 706 1916 712
rect 1279 698 1290 701
rect 1373 698 1381 701
rect 1401 700 1409 701
rect 742 688 743 692
rect 705 676 739 678
rect 743 676 751 688
rect 838 686 844 692
rect 896 686 902 692
rect 928 688 935 692
rect 1044 691 1050 697
rect 1090 691 1096 697
rect 1136 691 1279 698
rect 1351 691 1373 698
rect 1407 692 1409 700
rect 1410 693 1416 698
rect 1429 694 1441 701
rect 1031 688 1033 691
rect 928 687 940 688
rect 844 680 850 686
rect 890 680 896 686
rect 928 685 943 687
rect 950 685 962 688
rect 1030 687 1031 688
rect 1029 685 1030 687
rect 1038 685 1044 691
rect 1096 685 1102 691
rect 1103 689 1124 691
rect 1346 689 1351 691
rect 1340 687 1346 689
rect 1409 688 1410 692
rect 1418 689 1421 691
rect 1107 685 1142 687
rect 928 680 940 685
rect 943 680 965 685
rect 1027 683 1029 685
rect 965 676 978 680
rect 978 675 983 676
rect 992 675 1042 683
rect 1095 682 1107 685
rect 1086 680 1095 682
rect 1147 680 1149 685
rect 1330 684 1338 687
rect 1410 686 1411 687
rect 1323 682 1330 684
rect 1085 676 1086 680
rect 1316 679 1323 682
rect 1411 680 1413 682
rect 1311 678 1316 679
rect 1305 676 1311 678
rect 1413 676 1415 680
rect 1427 678 1434 684
rect 1446 682 1504 701
rect 1531 692 1532 698
rect 1595 692 1596 701
rect 1600 693 1608 703
rect 1615 702 1619 705
rect 1680 702 1705 706
rect 1802 704 1815 706
rect 1603 691 1608 693
rect 1619 692 1630 702
rect 1446 678 1479 682
rect 741 672 743 675
rect 983 674 1042 675
rect 992 672 1042 674
rect 448 656 451 662
rect 372 643 436 649
rect 446 648 448 656
rect 492 652 509 672
rect 532 666 539 672
rect 705 666 717 672
rect 727 666 739 672
rect 969 666 992 672
rect 539 664 745 666
rect 958 664 969 666
rect 378 637 405 643
rect 424 637 430 643
rect 440 642 446 647
rect 450 642 459 644
rect 509 643 517 652
rect 686 642 687 660
rect 188 626 191 630
rect 381 626 405 637
rect 440 635 459 642
rect 518 639 522 642
rect 522 636 527 639
rect 527 635 535 636
rect 440 630 455 635
rect 535 631 571 635
rect 439 626 455 630
rect 571 628 591 631
rect 685 630 687 642
rect 745 654 904 664
rect 916 654 958 664
rect 1082 663 1085 674
rect 1149 663 1152 676
rect 1300 674 1305 676
rect 1297 673 1300 674
rect 1292 672 1297 673
rect 1286 670 1292 672
rect 1415 670 1418 676
rect 1434 671 1442 678
rect 1479 671 1487 678
rect 1504 676 1510 682
rect 1533 679 1534 682
rect 1535 677 1536 687
rect 1587 681 1600 682
rect 1587 679 1596 681
rect 1630 679 1635 692
rect 1680 688 1729 702
rect 1754 698 1800 704
rect 1818 703 1820 706
rect 1830 704 1850 706
rect 1858 704 1877 706
rect 1801 700 1816 702
rect 1746 694 1754 698
rect 1680 687 1705 688
rect 1729 687 1735 688
rect 1737 687 1746 694
rect 1662 678 1680 687
rect 1729 686 1737 687
rect 1735 685 1739 686
rect 1725 677 1732 683
rect 1739 682 1747 685
rect 1747 681 1752 682
rect 1752 680 1757 681
rect 1758 678 1761 679
rect 1529 676 1550 677
rect 1587 676 1593 677
rect 1510 673 1514 676
rect 1267 668 1286 670
rect 1230 664 1267 668
rect 1153 663 1230 664
rect 1044 655 1230 663
rect 1418 660 1431 670
rect 1442 660 1464 671
rect 1487 663 1497 671
rect 1514 663 1518 673
rect 1529 671 1535 676
rect 1536 672 1550 676
rect 1576 671 1593 676
rect 1634 671 1635 676
rect 1645 671 1660 677
rect 1535 665 1541 671
rect 1581 665 1587 671
rect 1625 663 1645 671
rect 1716 669 1725 677
rect 1764 676 1769 678
rect 1770 674 1776 676
rect 745 652 916 654
rect 1044 653 1159 655
rect 745 642 747 652
rect 1044 651 1156 653
rect 1044 649 1149 651
rect 1044 648 1112 649
rect 1044 645 1096 648
rect 1038 644 1102 645
rect 1016 642 1102 644
rect 745 634 751 642
rect 1010 639 1027 642
rect 1038 639 1102 642
rect 1135 641 1147 649
rect 1152 643 1156 651
rect 992 636 1010 639
rect 746 630 751 634
rect 973 633 992 636
rect 1044 633 1050 639
rect 1076 636 1082 639
rect 1090 633 1096 639
rect 1154 636 1156 643
rect 1431 642 1477 660
rect 1497 652 1527 663
rect 1507 647 1541 652
rect 1561 647 1562 660
rect 1598 652 1625 663
rect 1634 660 1635 663
rect 1507 646 1578 647
rect 1586 646 1615 652
rect 1507 643 1615 646
rect 1513 642 1518 643
rect 1431 641 1479 642
rect 958 631 973 633
rect 762 630 802 631
rect 956 630 958 631
rect 601 628 762 630
rect 802 628 831 630
rect 685 626 688 628
rect 744 626 751 628
rect 191 618 199 626
rect 259 618 266 625
rect 199 617 259 618
rect 423 610 439 626
rect 688 615 694 626
rect 741 618 744 625
rect 831 622 892 628
rect 902 622 952 630
rect 1152 627 1154 636
rect 733 615 741 618
rect 694 613 735 615
rect 1076 613 1089 624
rect 1130 616 1152 627
rect 1431 626 1477 641
rect 1481 637 1484 639
rect 1484 636 1486 637
rect 1486 633 1493 636
rect 1513 634 1527 642
rect 1561 634 1562 643
rect 1633 637 1634 653
rect 1675 652 1716 669
rect 1770 668 1778 674
rect 1782 670 1784 672
rect 1814 670 1816 700
rect 1820 690 1828 702
rect 1858 700 1864 704
rect 1904 700 1910 706
rect 1928 693 1939 702
rect 1782 668 1816 670
rect 1820 668 1828 680
rect 1939 678 1942 692
rect 1942 676 1943 678
rect 1778 664 1781 666
rect 1782 656 1794 664
rect 1804 656 1816 664
rect 1943 661 1946 676
rect 1660 646 1675 652
rect 1782 648 1791 656
rect 1945 648 1946 661
rect 1646 641 1658 646
rect 1637 637 1646 641
rect 1493 631 1499 633
rect 1511 630 1527 634
rect 1502 626 1527 630
rect 1561 626 1563 630
rect 1495 622 1520 626
rect 1090 613 1130 616
rect 701 610 717 613
rect 719 610 735 613
rect 1495 610 1511 622
rect 1520 619 1528 622
rect 1528 618 1537 619
rect 1563 615 1568 626
rect 1595 620 1637 637
rect 1592 619 1595 620
rect 1586 618 1592 619
rect 1624 618 1631 620
rect 1620 615 1624 618
rect 1568 611 1589 615
rect 1611 611 1620 615
rect 1761 606 1785 629
rect 1791 626 1830 648
rect 1830 621 1839 626
rect 1936 622 1945 643
rect 1935 621 1936 622
rect 1839 615 1856 621
rect 1931 616 1935 621
rect 1928 615 1931 616
rect 1856 611 1928 615
rect 117 557 167 606
rect 197 557 263 606
rect 293 557 359 606
rect 389 557 455 606
rect 485 557 535 606
rect 605 557 655 606
rect 685 557 751 606
rect 781 557 847 606
rect 877 557 943 606
rect 973 557 1023 606
rect 1093 557 1143 606
rect 1173 557 1239 606
rect 1269 557 1335 606
rect 1365 557 1431 606
rect 1461 557 1511 606
rect 1581 557 1631 606
rect 1661 557 1727 606
rect 1757 557 1823 606
rect 1853 557 1903 606
<< nwell >>
rect 1 820 3170 1748
rect 1980 744 2194 820
rect 2976 772 3006 807
rect 3125 744 3170 820
<< ndiff >>
rect 3061 441 3095 475
<< locali >>
rect 0 2172 3171 2492
rect 1 1086 3170 1406
rect 1428 774 1511 845
rect 1831 834 1903 929
rect 1821 774 1903 834
rect 2027 829 2101 903
rect 51 320 2017 577
rect 0 0 3171 320
<< viali >>
rect 3061 1721 3095 1755
rect 3062 1461 3096 1495
rect 3061 441 3095 475
<< metal1 >>
rect 0 2172 3171 2492
rect 1388 1754 1422 2172
rect 1532 1931 1600 1937
rect 1532 1874 1538 1931
rect 1594 1874 1600 1931
rect 2539 1908 2823 1915
rect 2551 1902 2823 1908
rect 1532 1868 1600 1874
rect 2505 1881 2823 1902
rect 2505 1868 2551 1881
rect 2584 1846 2649 1853
rect 2584 1828 2591 1846
rect 1625 1794 2591 1828
rect 2643 1794 2649 1846
rect 2584 1788 2649 1794
rect 1388 1720 1462 1754
rect 2424 1708 2430 1766
rect 2482 1708 2488 1766
rect 2214 1692 2284 1698
rect 2214 1680 2220 1692
rect 1321 1646 2220 1680
rect 2214 1634 2220 1646
rect 2278 1634 2284 1692
rect 2789 1645 2823 1881
rect 3062 1848 3095 1906
rect 2898 1722 3021 1754
rect 2898 1721 2930 1722
rect 2988 1686 3021 1722
rect 2990 1646 3021 1686
rect 2214 1628 2284 1634
rect 3044 1508 3118 1517
rect 3044 1452 3053 1508
rect 3109 1452 3118 1508
rect 3044 1443 3118 1452
rect 1 1086 3170 1406
rect 1831 944 1903 949
rect 1821 914 1903 944
rect 1659 913 1903 914
rect 1651 902 1903 913
rect 1638 895 1903 902
rect 1631 885 1903 895
rect 1599 876 1903 885
rect 1596 875 1903 876
rect 1574 869 1903 875
rect 1551 866 1903 869
rect 2027 894 2101 903
rect 1551 862 1976 866
rect 1538 858 1976 862
rect 1510 852 1976 858
rect 1470 847 1673 852
rect 1470 843 1643 847
rect 1470 841 1519 843
rect 1528 841 1620 843
rect 1470 839 1620 841
rect 1470 833 1595 839
rect 1802 833 1976 852
rect 1470 826 1577 833
rect 1821 829 1976 833
rect 2027 838 2036 894
rect 2092 838 2101 894
rect 2027 829 2101 838
rect 2213 864 2283 870
rect 1470 815 1556 826
rect 1821 815 1903 829
rect 1470 810 1551 815
rect 1834 814 1903 815
rect 1470 807 1519 810
rect 1470 804 1516 807
rect 1939 577 1976 829
rect 2213 806 2219 864
rect 2277 806 2283 864
rect 2790 819 2824 846
rect 2968 845 3032 852
rect 2790 812 2825 819
rect 2791 809 2825 812
rect 2213 800 2283 806
rect 2790 806 2825 809
rect 2968 807 2989 845
rect 2424 790 2488 796
rect 2424 772 2430 790
rect 2404 738 2430 772
rect 2482 738 2488 790
rect 2424 732 2488 738
rect 2579 716 2649 722
rect 2579 698 2585 716
rect 2112 664 2585 698
rect 2112 597 2146 664
rect 2579 658 2585 664
rect 2643 658 2649 716
rect 2579 652 2649 658
rect 2790 624 2823 806
rect 2968 772 3006 807
rect 2897 738 3006 772
rect 2505 623 2539 624
rect 2551 623 2823 624
rect 2092 591 2162 597
rect 51 320 2017 577
rect 2092 533 2098 591
rect 2156 533 2162 591
rect 2505 590 2823 623
rect 3118 545 3124 603
rect 2092 527 2162 533
rect 0 0 3171 320
<< via1 >>
rect 1538 1874 1594 1931
rect 2591 1794 2643 1846
rect 2430 1708 2482 1766
rect 2220 1634 2278 1692
rect 3053 1495 3109 1508
rect 3053 1461 3062 1495
rect 3062 1461 3096 1495
rect 3096 1461 3109 1495
rect 3053 1452 3109 1461
rect 2036 838 2092 894
rect 2219 806 2277 864
rect 2430 738 2482 790
rect 2585 658 2643 716
rect 2098 533 2156 591
rect 3060 545 3118 603
<< metal2 >>
rect 1529 1931 1603 1939
rect 1529 1874 1538 1931
rect 1594 1874 1603 1931
rect 1529 1865 1603 1874
rect 2584 1846 2649 1853
rect 2584 1840 2591 1846
rect 2361 1806 2591 1840
rect 2214 1692 2284 1698
rect 2214 1634 2220 1692
rect 2278 1634 2284 1692
rect 2214 1628 2284 1634
rect 98 559 132 854
rect 1828 814 1903 929
rect 2027 894 2101 903
rect 2027 838 2036 894
rect 2092 838 2101 894
rect 2228 870 2263 1628
rect 2027 829 2101 838
rect 2213 864 2283 870
rect 1834 789 1903 814
rect 2044 742 2078 829
rect 2213 806 2219 864
rect 2277 806 2283 864
rect 2213 800 2283 806
rect 1869 706 2078 742
rect 2361 772 2393 1806
rect 2584 1794 2591 1806
rect 2643 1794 2649 1846
rect 2584 1788 2649 1794
rect 2424 1708 2430 1766
rect 2482 1708 2488 1766
rect 2424 1701 2488 1708
rect 2430 1666 2464 1701
rect 2430 1631 2465 1666
rect 2430 1596 2625 1631
rect 2424 790 2488 796
rect 2424 772 2430 790
rect 2361 738 2430 772
rect 2482 738 2488 790
rect 2424 732 2488 738
rect 2590 722 2625 1596
rect 3044 1508 3118 1517
rect 3044 1452 3053 1508
rect 3109 1452 3118 1508
rect 3044 1443 3118 1452
rect 2579 716 2649 722
rect 2579 658 2585 716
rect 2643 658 2649 716
rect 2579 652 2649 658
rect 3051 603 3127 612
rect 2092 591 2162 597
rect 2092 578 2098 591
rect 2091 559 2098 578
rect 98 533 2098 559
rect 2156 533 2162 591
rect 3051 545 3060 603
rect 3118 545 3127 603
rect 3051 536 3127 545
rect 98 527 2162 533
rect 98 525 2140 527
<< via2 >>
rect 1538 1874 1594 1930
rect 2036 838 2092 894
rect 3053 1452 3109 1508
rect 3060 545 3118 603
<< metal3 >>
rect 1529 1930 1603 1939
rect 1529 1874 1538 1930
rect 1594 1874 1603 1930
rect 1529 1865 1603 1874
rect 1537 1862 1603 1865
rect 1537 1801 2095 1862
rect 2034 903 2095 1801
rect 3044 1508 3114 2492
rect 3044 1452 3053 1508
rect 3109 1452 3114 1508
rect 3044 1443 3114 1452
rect 2027 894 2101 903
rect 2027 838 2036 894
rect 2092 838 2101 894
rect 2027 829 2101 838
rect 927 703 988 771
rect 1100 703 1174 789
rect 1736 703 1797 723
rect 927 629 1799 703
rect 3051 603 3127 612
rect 3051 545 3060 603
rect 3118 545 3127 603
rect 3051 0 3127 545
use scs130hd_mpr2aa_8  scs130hd_mpr2aa_8_0
timestamp 1697204803
transform 1 0 51 0 1 559
box -38 -48 1970 592
use sky130_osu_sc_12T_hs__fill_2  sky130_osu_sc_12T_hs__fill_2_0
timestamp 1604095901
transform 1 0 1631 0 -1 2233
box -7 0 161 1341
use sky130_osu_sc_12T_hs__fill_8  sky130_osu_sc_12T_hs__fill_8_0
timestamp 1604095905
transform 1 0 1802 0 -1 2233
box -9 0 179 897
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1706264206
transform 1 0 2743 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1706264206
transform 1 0 2940 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1706264206
transform 1 0 2941 0 -1 2233
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1706264206
transform 1 0 2743 0 -1 2233
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1698882961
transform 1 0 2194 0 1 259
box -9 0 553 903
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1698882961
transform 1 0 1238 0 -1 2233
box -9 0 553 903
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1698882961
transform 1 0 2194 0 -1 2233
box -9 0 553 903
<< labels >>
rlabel metal2 2242 840 2242 840 1 sel
port 7 n
rlabel metal1 51 292 51 292 1 vssd1
port 5 n
rlabel metal1 43 1158 43 1158 1 vccd1
port 6 n
rlabel viali 3061 441 3095 475 1 Y1
port 10 n
rlabel metal1 1625 1794 1645 1828 1 in
port 8 n
rlabel viali 3061 1721 3095 1755 1 Y0
port 9 n
<< end >>
