magic
tech sky130A
magscale 1 2
timestamp 1712684262
<< nwell >>
rect 3000 1407 6401 1748
rect 8015 1635 8073 1693
rect 11280 1635 11338 1693
rect 14545 1635 14603 1693
rect 17810 1635 17868 1693
rect 3000 1087 19884 1407
rect 3000 1018 6401 1087
rect 3000 800 4617 1018
rect 6703 974 6761 1032
rect 9968 974 10026 1032
rect 13233 974 13291 1032
rect 16498 974 16556 1032
rect 19763 974 19821 1032
rect 6815 799 6939 826
rect 10082 800 10206 827
rect 13348 800 13472 827
rect 16615 800 16739 829
<< ndiff >>
rect 6715 442 6750 476
rect 9980 442 10015 476
rect 13245 442 13280 476
rect 16510 442 16545 476
rect 19775 442 19810 476
rect 6718 441 6749 442
rect 9983 441 10014 442
rect 13248 441 13279 442
rect 16513 441 16544 442
rect 19778 441 19809 442
<< pdiff >>
rect 3045 1647 3079 1681
rect 4750 1635 4808 1693
rect 8015 1635 8073 1693
rect 11280 1635 11338 1693
rect 14545 1635 14603 1693
rect 17810 1635 17868 1693
rect 6703 974 6761 1032
<< locali >>
rect 0 2172 19884 2492
rect 3406 1407 3440 1472
rect 0 1087 19884 1407
rect 6703 974 6761 1032
rect 0 0 19884 320
<< viali >>
rect 3045 1647 3079 1681
rect 6715 442 6750 476
rect 9980 442 10015 476
rect 13245 442 13280 476
rect 16510 442 16545 476
rect 19775 442 19810 476
<< metal1 >>
rect 0 2172 19884 2492
rect 19808 1982 19811 2012
rect 19770 1976 19840 1982
rect 3302 1862 3308 1920
rect 3366 1862 3372 1920
rect 19770 1918 19776 1976
rect 19834 1918 19840 1976
rect 19770 1912 19840 1918
rect 6714 1852 6784 1858
rect 5317 1842 5387 1848
rect 5317 1784 5323 1842
rect 5381 1784 5387 1842
rect 6714 1794 6720 1852
rect 6778 1794 6784 1852
rect 9978 1853 10049 1860
rect 6714 1788 6784 1794
rect 8415 1843 8485 1849
rect 5317 1778 5387 1784
rect 8415 1785 8421 1843
rect 8479 1785 8485 1843
rect 9978 1795 9985 1853
rect 10043 1795 10049 1853
rect 13235 1852 13305 1858
rect 9978 1789 10049 1795
rect 11680 1844 11750 1850
rect 8415 1779 8485 1785
rect 11680 1786 11686 1844
rect 11744 1786 11750 1844
rect 13235 1794 13241 1852
rect 13299 1794 13305 1852
rect 16500 1852 16570 1858
rect 13235 1788 13305 1794
rect 14945 1843 15015 1849
rect 11680 1780 11750 1786
rect 14945 1785 14951 1843
rect 15009 1785 15015 1843
rect 16500 1794 16506 1852
rect 16564 1794 16570 1852
rect 16500 1788 16570 1794
rect 18211 1843 18281 1849
rect 14945 1779 15015 1785
rect 18211 1785 18217 1843
rect 18275 1785 18281 1843
rect 18211 1779 18281 1785
rect 3227 1714 3233 1772
rect 3291 1714 3297 1772
rect 3034 1681 3092 1686
rect 3034 1647 3045 1681
rect 3079 1647 3092 1681
rect 3034 1640 3092 1647
rect 0 1087 19884 1407
rect 6715 441 6749 442
rect 9980 441 10014 442
rect 13245 441 13279 442
rect 16510 441 16544 442
rect 19775 441 19809 442
rect 0 0 19884 320
<< via1 >>
rect 3308 1862 3366 1920
rect 19776 1918 19834 1976
rect 5323 1784 5381 1842
rect 6720 1794 6778 1852
rect 8421 1785 8479 1843
rect 9985 1795 10043 1853
rect 11686 1786 11744 1844
rect 13241 1794 13299 1852
rect 14951 1785 15009 1843
rect 16506 1794 16564 1852
rect 18217 1785 18275 1843
rect 3233 1714 3291 1772
rect 4750 1635 4808 1693
rect 8015 1635 8073 1693
rect 11280 1635 11338 1693
rect 14545 1635 14603 1693
rect 17810 1635 17868 1693
rect 6703 974 6761 1032
rect 9968 974 10026 1032
rect 13233 974 13291 1032
rect 16498 974 16556 1032
rect 19763 974 19821 1032
<< metal2 >>
rect 3245 2137 19810 2171
rect 3245 1778 3279 2137
rect 19776 1982 19810 2137
rect 19770 1976 19840 1982
rect 3308 1920 3366 1926
rect 19770 1918 19776 1976
rect 19834 1918 19840 1976
rect 19770 1912 19840 1918
rect 3366 1867 3576 1901
rect 3308 1856 3366 1862
rect 3542 1828 3576 1867
rect 6714 1852 6784 1858
rect 5317 1842 5387 1848
rect 5317 1828 5323 1842
rect 3542 1794 5323 1828
rect 5317 1784 5323 1794
rect 5381 1784 5387 1842
rect 6714 1794 6720 1852
rect 6778 1834 6784 1852
rect 9979 1853 10049 1859
rect 8415 1843 8485 1849
rect 8415 1834 8421 1843
rect 6778 1794 8421 1834
rect 6714 1788 6784 1794
rect 5317 1778 5387 1784
rect 8415 1785 8421 1794
rect 8479 1785 8485 1843
rect 9979 1795 9985 1853
rect 10043 1835 10049 1853
rect 13235 1852 13305 1858
rect 11680 1844 11750 1850
rect 11680 1835 11686 1844
rect 10043 1795 11686 1835
rect 9979 1789 10049 1795
rect 8415 1779 8485 1785
rect 11680 1786 11686 1795
rect 11744 1786 11750 1844
rect 13235 1794 13241 1852
rect 13299 1834 13305 1852
rect 16500 1852 16570 1858
rect 14945 1843 15015 1849
rect 14945 1834 14951 1843
rect 13299 1794 14951 1834
rect 13235 1788 13305 1794
rect 11680 1780 11750 1786
rect 14945 1785 14951 1794
rect 15009 1785 15015 1843
rect 16500 1794 16506 1852
rect 16564 1834 16570 1852
rect 18211 1843 18281 1849
rect 18211 1834 18217 1843
rect 16564 1794 18217 1834
rect 16500 1788 16570 1794
rect 14945 1779 15015 1785
rect 18211 1785 18217 1794
rect 18275 1785 18281 1843
rect 18211 1779 18281 1785
rect 3233 1772 3291 1778
rect 3233 1708 3291 1714
<< via2 >>
rect 4750 1635 4808 1693
rect 8015 1635 8073 1693
rect 11280 1635 11338 1693
rect 14545 1635 14603 1693
rect 17810 1635 17868 1693
rect 6703 974 6761 1032
rect 9968 974 10026 1032
rect 13233 974 13291 1032
rect 16498 974 16556 1032
rect 19763 974 19821 1032
<< metal3 >>
rect 8008 1693 8078 2492
rect 11273 1693 11343 2492
rect 14538 1693 14608 2492
rect 17803 1693 17873 2492
rect 6697 0 6767 974
rect 9962 0 10032 974
rect 13227 0 13297 974
rect 16492 0 16562 974
rect 19757 0 19827 974
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1710278372
transform 1 0 3009 0 -1 2233
box -10 0 552 902
use sky130_osu_single_mpr2ea_8_b0r2  sky130_osu_single_mpr2ea_8_b0r2_0
timestamp 1712684262
transform 1 0 16617 0 1 0
box 0 0 3268 2492
use sky130_osu_single_mpr2ea_8_b0r2  sky130_osu_single_mpr2ea_8_b0r2_1
timestamp 1712684262
transform 1 0 3557 0 1 0
box 0 0 3268 2492
use sky130_osu_single_mpr2ea_8_b0r2  sky130_osu_single_mpr2ea_8_b0r2_2
timestamp 1712684262
transform 1 0 6822 0 1 0
box 0 0 3268 2492
use sky130_osu_single_mpr2ea_8_b0r2  sky130_osu_single_mpr2ea_8_b0r2_3
timestamp 1712684262
transform 1 0 10087 0 1 0
box 0 0 3268 2492
use sky130_osu_single_mpr2ea_8_b0r2  sky130_osu_single_mpr2ea_8_b0r2_4
timestamp 1712684262
transform 1 0 13352 0 1 0
box 0 0 3268 2492
<< labels >>
flabel metal1 s 3034 1640 3092 1686 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 0 1087 19884 1407 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 0 0 19884 320 0 FreeSans 100 0 0 0 vssd1
port 16 nsew ground bidirectional
flabel metal1 s 0 2172 19884 2492 0 FreeSans 100 0 0 0 vssd1
port 16 nsew ground bidirectional
flabel metal1 s 4761 1647 4795 1681 0 FreeSans 100 0 0 0 s1
port 1 n signal input
flabel metal1 s 8026 1647 8060 1681 0 FreeSans 100 0 0 0 s2
port 2 n signal input
flabel metal1 s 11291 1647 11325 1681 0 FreeSans 100 0 0 0 s3
port 3 n signal input
flabel metal1 s 14556 1647 14590 1681 0 FreeSans 100 0 0 0 s4
port 4 n signal input
flabel metal1 s 17821 1647 17855 1681 0 FreeSans 100 0 0 0 s5
port 5 n signal input
flabel metal1 s 19775 442 19810 476 0 FreeSans 100 0 0 0 X5_Y1
port 10 s signal output
flabel metal1 s 16510 442 16545 476 0 FreeSans 100 0 0 0 X4_Y1
port 9 s signal output
flabel metal1 s 13245 442 13280 476 0 FreeSans 100 0 0 0 X3_Y1
port 8 s signal output
flabel metal1 s 9980 442 10015 476 0 FreeSans 100 0 0 0 X2_Y1
port 7 s signal output
flabel metal1 s 6715 442 6750 476 0 FreeSans 100 0 0 0 X1_Y1
port 6 s signal output
<< end >>
