magic
tech sky130A
magscale 1 2
timestamp 1713897945
<< nwell >>
rect 2937 1749 2979 1750
rect 0 1087 3052 1749
rect 0 829 109 1087
rect 1860 1086 2086 1087
rect 0 819 110 829
rect 1862 744 2076 1086
rect 2097 800 2165 870
rect 2858 772 2888 807
rect 3007 744 3052 1087
<< ndiff >>
rect 2942 441 2977 475
<< pdiff >>
rect 1032 1647 1038 1650
<< locali >>
rect 0 2173 3052 2493
rect 2627 1870 2678 1886
rect 2581 1852 2678 1870
rect 2765 1722 2881 1756
rect 2779 1690 2780 1722
rect 2944 1462 2978 1496
rect 0 1087 3052 1407
rect 1860 1086 2086 1087
rect 3016 1086 3052 1087
rect 2943 997 2977 1031
rect 2745 725 2902 759
rect 2581 623 2707 641
rect 420 559 459 578
rect 787 559 826 572
rect 1155 559 1194 578
rect 2627 607 2707 623
rect 1525 559 1565 576
rect 1859 559 1898 576
rect 175 544 1898 559
rect 150 320 1898 544
rect 0 0 3052 320
<< viali >>
rect 2581 1870 2627 1916
rect 2943 1744 2977 1778
rect 2581 577 2627 623
rect 2943 441 2977 475
<< metal1 >>
rect 0 2173 3052 2493
rect 1144 1721 1178 2173
rect 1244 1934 1318 1943
rect 1244 1878 1253 1934
rect 1309 1878 1318 1934
rect 2569 1916 2639 1922
rect 2421 1909 2581 1916
rect 2433 1903 2581 1909
rect 1244 1869 1318 1878
rect 2387 1882 2581 1903
rect 2387 1869 2433 1882
rect 2569 1870 2581 1882
rect 2627 1870 2639 1916
rect 2569 1864 2639 1870
rect 2466 1847 2531 1854
rect 2466 1829 2473 1847
rect 1316 1795 2473 1829
rect 2525 1795 2531 1847
rect 2466 1789 2531 1795
rect 2306 1709 2312 1767
rect 2364 1709 2370 1767
rect 2097 1694 2165 1700
rect 971 1681 1041 1694
rect 2097 1681 2103 1694
rect 971 1674 1042 1681
rect 2093 1674 2103 1681
rect 971 1647 2103 1674
rect 971 1641 2094 1647
rect 971 1636 1041 1641
rect 2097 1636 2103 1647
rect 2161 1636 2165 1694
rect 2097 1630 2165 1636
rect 0 1087 3052 1407
rect 1860 1086 2086 1087
rect 3016 1086 3052 1087
rect 1985 863 2053 869
rect 1985 805 1991 863
rect 2049 805 2053 863
rect 1985 799 2053 805
rect 2097 864 2165 870
rect 2097 806 2103 864
rect 2161 806 2165 864
rect 2097 800 2165 806
rect 2003 698 2037 799
rect 2306 790 2370 796
rect 2306 772 2312 790
rect 2299 738 2312 772
rect 2364 738 2370 790
rect 2306 732 2370 738
rect 2461 716 2531 722
rect 2461 698 2467 716
rect 347 564 405 670
rect 2003 664 2467 698
rect 2461 658 2467 664
rect 2525 658 2531 716
rect 2461 652 2531 658
rect 2569 624 2639 629
rect 2387 623 2421 624
rect 2433 623 2639 624
rect 2387 590 2581 623
rect 1859 583 1898 584
rect 420 559 459 578
rect 787 559 826 572
rect 1155 559 1194 578
rect 1859 576 1884 583
rect 2569 577 2581 590
rect 2627 577 2639 623
rect 1525 568 1565 576
rect 1859 559 1898 576
rect 2569 571 2639 577
rect 175 544 1898 559
rect 150 320 1898 544
rect 0 0 3052 320
<< via1 >>
rect 1253 1878 1309 1934
rect 2473 1795 2525 1847
rect 2312 1709 2364 1767
rect 2103 1636 2161 1694
rect 1991 805 2049 863
rect 2103 806 2161 864
rect 2312 738 2364 790
rect 2467 658 2525 716
<< metal2 >>
rect 1244 1934 1318 1943
rect 1244 1878 1253 1934
rect 1309 1878 1318 1934
rect 1244 1869 1318 1878
rect 2466 1847 2531 1854
rect 2466 1841 2473 1847
rect 2243 1807 2473 1841
rect 2097 1694 2165 1700
rect 2097 1636 2103 1694
rect 2161 1636 2165 1694
rect 2097 1630 2165 1636
rect 2113 870 2147 1630
rect 1985 863 2053 869
rect 1985 853 1991 863
rect 1860 813 1991 853
rect 1860 687 1900 813
rect 1985 805 1991 813
rect 2049 805 2053 863
rect 1985 799 2053 805
rect 2097 864 2165 870
rect 2097 806 2103 864
rect 2161 806 2165 864
rect 2097 800 2165 806
rect 2003 798 2037 799
rect 2243 772 2275 1807
rect 2466 1795 2473 1807
rect 2525 1795 2531 1847
rect 2466 1789 2531 1795
rect 2306 1709 2312 1767
rect 2364 1709 2370 1767
rect 2306 1702 2370 1709
rect 2312 1667 2346 1702
rect 2312 1632 2347 1667
rect 2312 1597 2507 1632
rect 2306 790 2370 796
rect 2306 772 2312 790
rect 2243 738 2312 772
rect 2364 738 2370 790
rect 2306 732 2370 738
rect 2472 722 2507 1597
rect 1776 647 1900 687
rect 2461 716 2531 722
rect 2461 658 2467 716
rect 2525 658 2531 716
rect 2461 652 2531 658
<< via2 >>
rect 1253 1878 1309 1934
<< metal3 >>
rect 1244 1934 1318 1943
rect 1244 1878 1253 1934
rect 1309 1878 1318 1934
rect 1244 1869 1318 1878
rect 1251 1306 1311 1869
rect 1250 1235 1311 1306
rect 1250 1154 1310 1235
rect 404 1094 1310 1154
rect 404 862 464 1094
rect 963 762 1023 1094
use scs130hd_mpr2xa_8  scs130hd_mpr2xa_8_0
timestamp 1713289166
transform 1 0 150 0 1 559
box -48 -48 1796 592
use sky130_osu_sc_12T_hs__fill_8  sky130_osu_sc_12T_hs__fill_8_0
timestamp 1713287902
transform 1 0 1684 0 -1 2234
box -9 0 179 897
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1713887963
transform 1 0 2625 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1713887963
transform 1 0 2822 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1713887963
transform 1 0 2823 0 -1 2234
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1713887963
transform 1 0 2625 0 -1 2234
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1713481735
transform 1 0 2076 0 1 259
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1713481735
transform 1 0 953 0 -1 2234
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1713481735
transform 1 0 2076 0 -1 2234
box -10 0 552 902
<< labels >>
rlabel metal1 50 1145 50 1145 1 vccd1
port 6 n
rlabel metal1 40 284 40 284 1 vssd1
port 5 n
rlabel metal2 2130 835 2130 835 1 sel
port 7 n
rlabel metal1 40 2206 40 2206 1 vssd1
port 5 n
rlabel metal1 1316 1795 1344 1829 1 in
port 11 n
rlabel viali 2943 441 2977 475 1 Y1
port 10 n
rlabel viali 2943 1744 2977 1778 1 Y0
port 9 n
<< end >>
