magic
tech sky130A
magscale 1 2
timestamp 1712692843
<< nwell >>
rect 2938 1749 2981 1750
rect 0 1087 3052 1749
rect 0 820 109 1087
rect 1860 1086 2086 1087
rect 0 819 106 820
rect 1862 744 2076 1086
rect 2097 800 2165 870
rect 2858 772 2888 807
rect 3007 744 3052 1087
<< ndiff >>
rect 2942 441 2976 475
<< locali >>
rect 0 2173 3052 2493
rect 0 1087 3052 1407
rect 1860 1086 2086 1087
rect 3016 1086 3052 1087
rect 420 559 459 578
rect 787 559 826 572
rect 1155 559 1194 578
rect 1525 559 1565 576
rect 1859 559 1898 576
rect 175 544 1898 559
rect 150 320 1898 544
rect 0 0 3052 320
<< viali >>
rect 2943 1722 2977 1756
rect 2944 1462 2978 1496
rect 2943 997 2977 1031
rect 2942 441 2977 475
<< metal1 >>
rect 0 2173 3052 2493
rect 1144 1721 1178 2173
rect 1244 1934 1318 1943
rect 1244 1878 1253 1934
rect 1309 1878 1318 1934
rect 2421 1909 2705 1916
rect 2433 1903 2705 1909
rect 1244 1869 1318 1878
rect 2387 1882 2705 1903
rect 2387 1869 2433 1882
rect 2466 1847 2531 1854
rect 2466 1829 2473 1847
rect 1316 1795 2473 1829
rect 2525 1795 2531 1847
rect 2466 1789 2531 1795
rect 2306 1709 2312 1767
rect 2364 1709 2370 1767
rect 2097 1694 2165 1700
rect 971 1636 977 1694
rect 1035 1681 1041 1694
rect 2097 1681 2103 1694
rect 1035 1647 2103 1681
rect 1035 1636 1041 1647
rect 2097 1636 2103 1647
rect 2161 1636 2165 1694
rect 2671 1646 2705 1882
rect 2780 1723 2903 1755
rect 2780 1722 2812 1723
rect 2870 1688 2903 1723
rect 2870 1687 2904 1688
rect 2872 1647 2904 1687
rect 2097 1630 2165 1636
rect 2926 1450 2932 1508
rect 2990 1450 2996 1508
rect 0 1087 3052 1407
rect 1860 1086 2086 1087
rect 3016 1086 3052 1087
rect 2925 985 2931 1043
rect 2989 985 2995 1043
rect 1985 863 2053 869
rect 1985 805 1991 863
rect 2049 805 2053 863
rect 1985 799 2053 805
rect 2097 864 2165 870
rect 2097 806 2103 864
rect 2161 806 2165 864
rect 2850 846 2914 852
rect 2672 819 2706 846
rect 2672 812 2707 819
rect 2673 809 2707 812
rect 2097 800 2165 806
rect 2672 806 2707 809
rect 2850 807 2871 846
rect 2003 698 2037 799
rect 2306 790 2370 796
rect 2306 772 2312 790
rect 2299 738 2312 772
rect 2364 738 2370 790
rect 2306 732 2370 738
rect 2461 716 2531 722
rect 2461 698 2467 716
rect 347 582 405 670
rect 2003 664 2467 698
rect 2461 658 2467 664
rect 2525 658 2531 716
rect 2461 652 2531 658
rect 2672 624 2705 806
rect 2850 772 2888 807
rect 2779 738 2888 772
rect 2387 623 2421 624
rect 2433 623 2705 624
rect 2387 590 2705 623
rect 420 559 459 578
rect 787 559 826 572
rect 1155 559 1194 578
rect 1859 576 1884 583
rect 1525 568 1565 576
rect 1859 559 1898 576
rect 175 544 1898 559
rect 150 320 1898 544
rect 0 0 3052 320
<< via1 >>
rect 1253 1878 1309 1934
rect 2473 1795 2525 1847
rect 2312 1709 2364 1767
rect 977 1636 1035 1694
rect 2103 1636 2161 1694
rect 2932 1496 2990 1508
rect 2932 1462 2944 1496
rect 2944 1462 2978 1496
rect 2978 1462 2990 1496
rect 2932 1450 2990 1462
rect 2931 1031 2989 1043
rect 2931 997 2943 1031
rect 2943 997 2977 1031
rect 2977 997 2989 1031
rect 2931 985 2989 997
rect 1991 805 2049 863
rect 2103 806 2161 864
rect 2312 738 2364 790
rect 2467 658 2525 716
<< metal2 >>
rect 1244 1934 1318 1943
rect 1244 1878 1253 1934
rect 1309 1878 1318 1934
rect 1244 1869 1318 1878
rect 2466 1847 2531 1854
rect 2466 1841 2473 1847
rect 2243 1807 2473 1841
rect 977 1694 1035 1703
rect 977 1627 1035 1636
rect 2097 1694 2165 1700
rect 2097 1636 2103 1694
rect 2161 1636 2165 1694
rect 2097 1630 2165 1636
rect 1991 869 2049 872
rect 2113 870 2147 1630
rect 1985 863 2053 869
rect 1985 805 1991 863
rect 2049 805 2053 863
rect 1985 799 2053 805
rect 2097 864 2165 870
rect 2097 806 2103 864
rect 2161 806 2165 864
rect 2097 800 2165 806
rect 1991 796 2049 799
rect 2243 772 2275 1807
rect 2466 1795 2473 1807
rect 2525 1795 2531 1847
rect 2466 1789 2531 1795
rect 2306 1709 2312 1767
rect 2364 1709 2370 1767
rect 2306 1702 2370 1709
rect 2312 1667 2346 1702
rect 2312 1632 2347 1667
rect 2312 1597 2507 1632
rect 2306 790 2370 796
rect 2306 772 2312 790
rect 2243 738 2312 772
rect 2364 738 2370 790
rect 2306 732 2370 738
rect 2472 722 2507 1597
rect 2923 1508 2999 1517
rect 2923 1450 2932 1508
rect 2990 1450 2999 1508
rect 2923 1441 2999 1450
rect 2922 1043 2998 1052
rect 2922 985 2931 1043
rect 2989 985 2998 1043
rect 2922 976 2998 985
rect 2461 716 2531 722
rect 1776 647 1787 687
rect 2461 658 2467 716
rect 2525 658 2531 716
rect 2461 652 2531 658
<< via2 >>
rect 1253 1878 1309 1934
rect 977 1636 1035 1694
rect 1991 805 2049 863
rect 2932 1450 2990 1508
rect 2931 985 2989 1043
<< metal3 >>
rect 971 1694 1041 2493
rect 1244 1934 1318 1943
rect 1244 1878 1253 1934
rect 1309 1878 1318 1934
rect 1244 1869 1318 1878
rect 971 1636 977 1694
rect 1035 1636 1041 1694
rect 971 1627 1041 1636
rect 1251 1214 1311 1869
rect 2923 1508 2999 2493
rect 2923 1450 2932 1508
rect 2990 1450 2999 1508
rect 2923 1441 2999 1450
rect 404 1154 1311 1214
rect 404 1110 1023 1154
rect 404 862 464 1110
rect 963 762 1023 1110
rect 2922 1043 2998 1052
rect 2922 985 2931 1043
rect 2989 985 2998 1043
rect 1985 863 2057 873
rect 1985 805 1991 863
rect 2049 805 2057 863
rect 1985 788 2057 805
rect 867 664 923 683
rect 867 540 927 664
rect 1985 540 2053 788
rect 867 480 2053 540
rect 2922 0 2998 985
use scs130hd_mpr2xa_8  scs130hd_mpr2xa_8_0
timestamp 1712675931
transform 1 0 150 0 1 559
box -48 -48 1796 592
use sky130_osu_sc_12T_hs__fill_8  sky130_osu_sc_12T_hs__fill_8_0
timestamp 1604095905
transform 1 0 1684 0 -1 2234
box -9 0 179 897
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1712691322
transform 1 0 2625 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1712691322
transform 1 0 2822 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1712691322
transform 1 0 2823 0 -1 2234
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1712691322
transform 1 0 2625 0 -1 2234
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1710278372
transform 1 0 2076 0 1 259
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1710278372
transform 1 0 953 0 -1 2234
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1710278372
transform 1 0 2076 0 -1 2234
box -10 0 552 902
<< labels >>
rlabel metal1 50 1145 50 1145 1 vccd1
port 6 n
rlabel metal1 40 284 40 284 1 vssd1
port 5 n
rlabel metal2 2130 835 2130 835 1 sel
port 7 n
rlabel metal1 40 2206 40 2206 1 vssd1
port 5 n
rlabel metal1 1316 1795 1344 1829 1 in
port 11 n
rlabel viali 2943 1722 2977 1756 1 Y0
port 9 n
rlabel viali 2942 441 2976 475 1 Y1
port 10 n
<< end >>
