magic
tech sky130A
magscale 1 2
timestamp 1714057206
<< nwell >>
rect -10 484 552 902
<< pmos >>
rect 80 520 110 772
rect 271 520 301 772
rect 357 520 387 772
<< nmoslvt >>
rect 80 114 110 224
rect 271 114 301 224
rect 357 114 387 224
<< ndiff >>
rect 26 170 80 224
rect 26 130 34 170
rect 68 130 80 170
rect 26 114 80 130
rect 110 170 163 224
rect 110 130 121 170
rect 155 130 163 170
rect 110 114 163 130
rect 217 170 271 224
rect 217 130 225 170
rect 259 130 271 170
rect 217 114 271 130
rect 301 170 357 224
rect 301 130 312 170
rect 346 130 357 170
rect 301 114 357 130
rect 387 170 440 224
rect 387 130 398 170
rect 432 130 440 170
rect 387 114 440 130
<< pdiff >>
rect 26 756 80 772
rect 26 696 34 756
rect 68 696 80 756
rect 26 520 80 696
rect 110 756 163 772
rect 110 560 121 756
rect 155 560 163 756
rect 110 520 163 560
rect 217 756 271 772
rect 217 560 225 756
rect 259 560 271 756
rect 217 520 271 560
rect 301 756 357 772
rect 301 560 312 756
rect 346 560 357 756
rect 301 520 357 560
rect 387 756 440 772
rect 387 560 398 756
rect 432 560 440 756
rect 387 520 440 560
<< ndiffc >>
rect 34 130 68 170
rect 121 130 155 170
rect 225 130 259 170
rect 312 130 346 170
rect 398 130 432 170
<< pdiffc >>
rect 34 696 68 756
rect 121 560 155 756
rect 225 560 259 756
rect 312 560 346 756
rect 398 560 432 756
<< psubdiff >>
rect 26 26 50 60
rect 84 26 108 60
rect 26 20 108 26
rect 162 26 186 60
rect 220 26 244 60
rect 162 20 244 26
rect 298 26 322 60
rect 356 26 380 60
rect 298 20 380 26
rect 434 26 458 60
rect 492 26 516 60
rect 434 20 516 26
<< nsubdiff >>
rect 434 860 516 866
rect 434 826 458 860
rect 492 826 516 860
<< psubdiffcont >>
rect 50 26 84 60
rect 186 26 220 60
rect 322 26 356 60
rect 458 26 492 60
<< nsubdiffcont >>
rect 458 826 492 860
<< poly >>
rect 80 788 301 818
rect 80 772 110 788
rect 271 772 301 788
rect 357 772 387 798
rect 80 398 110 520
rect 271 494 301 520
rect 152 464 219 474
rect 152 430 168 464
rect 202 450 219 464
rect 357 450 387 520
rect 202 430 387 450
rect 152 420 387 430
rect 26 382 110 398
rect 26 348 36 382
rect 70 378 110 382
rect 70 348 387 378
rect 26 332 110 348
rect 80 224 110 332
rect 152 296 219 306
rect 152 262 168 296
rect 202 282 219 296
rect 202 262 301 282
rect 152 252 301 262
rect 271 224 301 252
rect 357 224 387 348
rect 80 88 110 114
rect 271 88 301 114
rect 357 88 387 114
<< polycont >>
rect 168 430 202 464
rect 36 348 70 382
rect 168 262 202 296
<< locali >>
rect 0 866 550 888
rect 0 826 458 866
rect 492 826 550 866
rect 34 756 68 826
rect 34 680 68 696
rect 120 756 155 772
rect 36 382 70 552
rect 36 332 70 348
rect 120 560 121 756
rect 120 520 155 560
rect 225 756 259 772
rect 311 756 346 772
rect 311 560 312 756
rect 225 526 271 560
rect 120 480 154 520
rect 237 510 271 526
rect 120 464 202 480
rect 120 430 168 464
rect 120 414 202 430
rect 120 312 154 414
rect 120 296 202 312
rect 120 262 168 296
rect 120 246 202 262
rect 120 212 154 246
rect 34 170 68 186
rect 34 60 68 130
rect 120 170 155 212
rect 237 204 271 476
rect 311 520 346 560
rect 397 756 432 772
rect 397 560 398 756
rect 397 544 432 560
rect 311 364 345 520
rect 397 438 431 544
rect 397 224 431 404
rect 120 130 121 170
rect 120 114 155 130
rect 225 170 271 204
rect 345 182 346 216
rect 311 170 346 182
rect 225 114 259 130
rect 311 130 312 170
rect 311 114 346 130
rect 397 170 432 224
rect 397 130 398 170
rect 397 114 432 130
rect 0 20 50 60
rect 84 20 186 60
rect 220 20 322 60
rect 356 20 458 60
rect 492 20 550 60
rect 0 0 550 20
<< viali >>
rect 458 860 492 866
rect 458 832 492 860
rect 36 552 70 586
rect 237 476 271 510
rect 311 330 345 364
rect 397 404 431 438
rect 311 182 345 216
rect 50 26 84 54
rect 50 20 84 26
rect 186 26 220 54
rect 186 20 220 26
rect 322 26 356 54
rect 322 20 356 26
rect 458 26 492 54
rect 458 20 492 26
<< metal1 >>
rect 0 866 550 888
rect 0 832 458 866
rect 492 832 550 866
rect 0 826 550 832
rect 24 586 82 592
rect 24 552 36 586
rect 70 552 116 586
rect 24 546 82 552
rect 225 510 283 516
rect 190 476 237 510
rect 271 476 283 510
rect 225 470 283 476
rect 385 438 443 444
rect 351 404 397 438
rect 431 404 443 438
rect 385 398 443 404
rect 299 364 357 370
rect 299 330 311 364
rect 345 330 357 364
rect 299 324 357 330
rect 311 222 345 324
rect 299 216 357 222
rect 299 182 311 216
rect 345 182 357 216
rect 299 176 357 182
rect 0 54 550 60
rect 0 20 50 54
rect 84 20 186 54
rect 220 20 322 54
rect 356 20 458 54
rect 492 20 550 54
rect 0 0 550 20
<< labels >>
rlabel viali 54 570 54 570 1 S0
port 1 n
rlabel viali 68 48 68 48 1 vssd1
port 6 n
rlabel viali 476 840 476 840 1 vccd1
port 5 n
rlabel viali 329 348 329 348 1 Y
port 2 n
rlabel viali 415 422 415 422 1 A1
port 4 n
rlabel viali 253 494 253 494 1 A0
port 3 n
<< end >>
