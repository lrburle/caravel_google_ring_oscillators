magic
tech sky130A
magscale 1 2
timestamp 1709223702
<< obsli1 >>
rect 441400 176800 526832 491663
<< obsm1 >>
rect 441400 176800 580230 492652
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 444010 6559 580318 492969
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 444005 484836 583520 492965
rect 444005 484436 583440 484836
rect 444005 471644 583520 484436
rect 444005 471244 583440 471644
rect 444005 458316 583520 471244
rect 444005 457916 583440 458316
rect 444005 444988 583520 457916
rect 444005 444588 583440 444988
rect 444005 431796 583520 444588
rect 444005 431396 583440 431796
rect 444005 418468 583520 431396
rect 444005 418068 583440 418468
rect 444005 405140 583520 418068
rect 444005 404740 583440 405140
rect 444005 391948 583520 404740
rect 444005 391548 583440 391948
rect 444005 378620 583520 391548
rect 444005 378220 583440 378620
rect 444005 365292 583520 378220
rect 444005 364892 583440 365292
rect 444005 352100 583520 364892
rect 444005 351700 583440 352100
rect 444005 338772 583520 351700
rect 444005 338372 583440 338772
rect 444005 325444 583520 338372
rect 444005 325044 583440 325444
rect 444005 312252 583520 325044
rect 444005 311852 583440 312252
rect 444005 298924 583520 311852
rect 444005 298524 583440 298924
rect 444005 285596 583520 298524
rect 444005 285196 583440 285596
rect 444005 272404 583520 285196
rect 444005 272004 583440 272404
rect 444005 259076 583520 272004
rect 444005 258676 583440 259076
rect 444005 245748 583520 258676
rect 444005 245348 583440 245748
rect 444005 232556 583520 245348
rect 444005 232156 583440 232556
rect 444005 219228 583520 232156
rect 444005 218828 583440 219228
rect 444005 205900 583520 218828
rect 444005 205500 583440 205900
rect 444005 192708 583520 205500
rect 444005 192308 583440 192708
rect 444005 179380 583520 192308
rect 444005 178980 583440 179380
rect 444005 166052 583520 178980
rect 444005 165652 583440 166052
rect 444005 152860 583520 165652
rect 444005 152460 583440 152860
rect 444005 139532 583520 152460
rect 444005 139132 583440 139532
rect 444005 126204 583520 139132
rect 444005 125804 583440 126204
rect 444005 113012 583520 125804
rect 444005 112612 583440 113012
rect 444005 99684 583520 112612
rect 444005 99284 583440 99684
rect 444005 86356 583520 99284
rect 444005 85956 583440 86356
rect 444005 73164 583520 85956
rect 444005 72764 583440 73164
rect 444005 59836 583520 72764
rect 444005 59436 583440 59836
rect 444005 46508 583520 59436
rect 444005 46108 583440 46508
rect 444005 33316 583520 46108
rect 444005 32916 583440 33316
rect 444005 19988 583520 32916
rect 444005 19588 583440 19988
rect 444005 6796 583520 19588
rect 444005 6563 583440 6796
<< metal4 >>
rect -15462 -14390 -14050 718326
rect -13710 -12638 -12298 716574
rect -11958 -10886 -10546 714822
rect -10206 -9134 -8794 713070
rect -8454 -7382 -7042 711318
rect -6702 -5630 -5290 709566
rect -4950 -3878 -3538 707814
rect -3198 -2126 -1786 706062
rect 1144 -8054 1464 711990
rect 2876 -8054 3196 711990
rect 4608 -8054 4928 711990
rect 6340 -8054 6660 711990
rect 8072 -8054 8392 711990
rect 9804 -8054 10124 711990
rect 11536 -8054 11856 711990
rect 13268 -8054 13588 711990
rect 15144 -8054 15464 711990
rect 16876 -8054 17196 711990
rect 18608 -8054 18928 711990
rect 20340 -8054 20660 711990
rect 22072 -8054 22392 711990
rect 23804 -8054 24124 711990
rect 25536 -8054 25856 711990
rect 27268 -8054 27588 711990
rect 29144 -8054 29464 711990
rect 30876 -8054 31196 711990
rect 32608 -8054 32928 711990
rect 34340 -8054 34660 711990
rect 36072 -8054 36392 711990
rect 37804 -8054 38124 711990
rect 39536 -8054 39856 711990
rect 41268 -8054 41588 711990
rect 43144 -8054 43464 711990
rect 44876 -8054 45196 711990
rect 46608 -8054 46928 711990
rect 48340 -8054 48660 711990
rect 50072 -8054 50392 711990
rect 51804 -8054 52124 711990
rect 53536 -8054 53856 711990
rect 55268 -8054 55588 711990
rect 57144 -8054 57464 711990
rect 58876 -8054 59196 711990
rect 60608 -8054 60928 711990
rect 62340 -8054 62660 711990
rect 64072 -8054 64392 711990
rect 65804 -8054 66124 711990
rect 67536 -8054 67856 711990
rect 69268 -8054 69588 711990
rect 71144 -8054 71464 711990
rect 72876 -8054 73196 711990
rect 74608 -8054 74928 711990
rect 76340 -8054 76660 711990
rect 78072 -8054 78392 711990
rect 79804 -8054 80124 711990
rect 81536 -8054 81856 711990
rect 83268 -8054 83588 711990
rect 85144 -8054 85464 711990
rect 86876 -8054 87196 711990
rect 88608 -8054 88928 711990
rect 90340 -8054 90660 711990
rect 92072 -8054 92392 711990
rect 93804 -8054 94124 711990
rect 95536 -8054 95856 711990
rect 97268 -8054 97588 711990
rect 99144 -8054 99464 711990
rect 100876 -8054 101196 711990
rect 102608 -8054 102928 711990
rect 104340 -8054 104660 711990
rect 106072 -8054 106392 711990
rect 107804 -8054 108124 711990
rect 109536 -8054 109856 711990
rect 111268 -8054 111588 711990
rect 113144 -8054 113464 711990
rect 114876 -8054 115196 711990
rect 116608 -8054 116928 711990
rect 118340 -8054 118660 711990
rect 120072 -8054 120392 711990
rect 121804 -8054 122124 711990
rect 123536 -8054 123856 711990
rect 125268 -8054 125588 711990
rect 127144 -8054 127464 711990
rect 128876 -8054 129196 711990
rect 130608 -8054 130928 711990
rect 132340 -8054 132660 711990
rect 134072 -8054 134392 711990
rect 135804 -8054 136124 711990
rect 137536 -8054 137856 711990
rect 139268 -8054 139588 711990
rect 141144 -8054 141464 711990
rect 142876 -8054 143196 711990
rect 144608 -8054 144928 711990
rect 146340 -8054 146660 711990
rect 148072 -8054 148392 711990
rect 149804 -8054 150124 711990
rect 151536 -8054 151856 711990
rect 153268 -8054 153588 711990
rect 155144 -8054 155464 711990
rect 156876 -8054 157196 711990
rect 158608 -8054 158928 711990
rect 160340 -8054 160660 711990
rect 162072 -8054 162392 711990
rect 163804 -8054 164124 711990
rect 165536 -8054 165856 711990
rect 167268 -8054 167588 711990
rect 169144 -8054 169464 711990
rect 170876 -8054 171196 711990
rect 172608 -8054 172928 711990
rect 174340 -8054 174660 711990
rect 176072 -8054 176392 711990
rect 177804 -8054 178124 711990
rect 179536 -8054 179856 711990
rect 181268 -8054 181588 711990
rect 183144 -8054 183464 711990
rect 184876 -8054 185196 711990
rect 186608 -8054 186928 711990
rect 188340 -8054 188660 711990
rect 190072 -8054 190392 711990
rect 191804 -8054 192124 711990
rect 193536 -8054 193856 711990
rect 195268 -8054 195588 711990
rect 197144 -8054 197464 711990
rect 198876 -8054 199196 711990
rect 200608 -8054 200928 711990
rect 202340 -8054 202660 711990
rect 204072 -8054 204392 711990
rect 205804 -8054 206124 711990
rect 207536 -8054 207856 711990
rect 209268 -8054 209588 711990
rect 211144 -8054 211464 711990
rect 212876 -8054 213196 711990
rect 214608 -8054 214928 711990
rect 216340 -8054 216660 711990
rect 218072 -8054 218392 711990
rect 219804 -8054 220124 711990
rect 221536 -8054 221856 711990
rect 223268 -8054 223588 711990
rect 225144 -8054 225464 711990
rect 226876 -8054 227196 711990
rect 228608 -8054 228928 711990
rect 230340 -8054 230660 711990
rect 232072 -8054 232392 711990
rect 233804 -8054 234124 711990
rect 235536 -8054 235856 711990
rect 237268 -8054 237588 711990
rect 239144 -8054 239464 711990
rect 240876 -8054 241196 711990
rect 242608 -8054 242928 711990
rect 244340 -8054 244660 711990
rect 246072 -8054 246392 711990
rect 247804 -8054 248124 711990
rect 249536 -8054 249856 711990
rect 251268 -8054 251588 711990
rect 253144 -8054 253464 711990
rect 254876 -8054 255196 711990
rect 256608 -8054 256928 711990
rect 258340 -8054 258660 711990
rect 260072 -8054 260392 711990
rect 261804 -8054 262124 711990
rect 263536 -8054 263856 711990
rect 265268 -8054 265588 711990
rect 267144 -8054 267464 711990
rect 268876 -8054 269196 711990
rect 270608 -8054 270928 711990
rect 272340 -8054 272660 711990
rect 274072 -8054 274392 711990
rect 275804 -8054 276124 711990
rect 277536 -8054 277856 711990
rect 279268 -8054 279588 711990
rect 281144 -8054 281464 711990
rect 282876 -8054 283196 711990
rect 284608 -8054 284928 711990
rect 286340 -8054 286660 711990
rect 288072 -8054 288392 711990
rect 289804 -8054 290124 711990
rect 291536 -8054 291856 711990
rect 293268 -8054 293588 711990
rect 295144 -8054 295464 711990
rect 296876 -8054 297196 711990
rect 298608 -8054 298928 711990
rect 300340 -8054 300660 711990
rect 302072 -8054 302392 711990
rect 303804 -8054 304124 711990
rect 305536 -8054 305856 711990
rect 307268 -8054 307588 711990
rect 309144 -8054 309464 711990
rect 310876 -8054 311196 711990
rect 312608 -8054 312928 711990
rect 314340 -8054 314660 711990
rect 316072 -8054 316392 711990
rect 317804 -8054 318124 711990
rect 319536 -8054 319856 711990
rect 321268 -8054 321588 711990
rect 323144 -8054 323464 711990
rect 324876 -8054 325196 711990
rect 326608 -8054 326928 711990
rect 328340 -8054 328660 711990
rect 330072 -8054 330392 711990
rect 331804 -8054 332124 711990
rect 333536 -8054 333856 711990
rect 335268 -8054 335588 711990
rect 337144 -8054 337464 711990
rect 338876 -8054 339196 711990
rect 340608 -8054 340928 711990
rect 342340 -8054 342660 711990
rect 344072 -8054 344392 711990
rect 345804 -8054 346124 711990
rect 347536 -8054 347856 711990
rect 349268 -8054 349588 711990
rect 351144 -8054 351464 711990
rect 352876 -8054 353196 711990
rect 354608 -8054 354928 711990
rect 356340 -8054 356660 711990
rect 358072 -8054 358392 711990
rect 359804 -8054 360124 711990
rect 361536 -8054 361856 711990
rect 363268 -8054 363588 711990
rect 365144 -8054 365464 711990
rect 366876 -8054 367196 711990
rect 368608 -8054 368928 711990
rect 370340 -8054 370660 711990
rect 372072 -8054 372392 711990
rect 373804 -8054 374124 711990
rect 375536 -8054 375856 711990
rect 377268 -8054 377588 711990
rect 379144 -8054 379464 711990
rect 380876 -8054 381196 711990
rect 382608 -8054 382928 711990
rect 384340 -8054 384660 711990
rect 386072 -8054 386392 711990
rect 387804 -8054 388124 711990
rect 389536 -8054 389856 711990
rect 391268 -8054 391588 711990
rect 393144 -8054 393464 711990
rect 394876 -8054 395196 711990
rect 396608 -8054 396928 711990
rect 398340 -8054 398660 711990
rect 400072 -8054 400392 711990
rect 401804 -8054 402124 711990
rect 403536 -8054 403856 711990
rect 405268 -8054 405588 711990
rect 407144 -8054 407464 711990
rect 408876 -8054 409196 711990
rect 410608 -8054 410928 711990
rect 412340 -8054 412660 711990
rect 414072 -8054 414392 711990
rect 415804 -8054 416124 711990
rect 417536 -8054 417856 711990
rect 419268 -8054 419588 711990
rect 421144 -8054 421464 711990
rect 422876 -8054 423196 711990
rect 424608 -8054 424928 711990
rect 426340 -8054 426660 711990
rect 428072 -8054 428392 711990
rect 429804 -8054 430124 711990
rect 431536 -8054 431856 711990
rect 433268 -8054 433588 711990
rect 435144 -8054 435464 711990
rect 436876 -8054 437196 711990
rect 438608 -8054 438928 711990
rect 440340 -8054 440660 711990
rect 442072 -8054 442392 711990
rect 443804 -8054 444124 711990
rect 445536 368640 445856 711990
rect 447268 368640 447588 711990
rect 449144 368640 449464 711990
rect 450876 368640 451196 711990
rect 452608 368640 452928 711990
rect 454340 368640 454660 711990
rect 456072 368640 456392 711990
rect 457804 368640 458124 711990
rect 459536 368640 459856 711990
rect 461268 368640 461588 711990
rect 445536 200640 445856 364236
rect 447268 200640 447588 364236
rect 449144 200640 449464 364236
rect 450876 200640 451196 364236
rect 452608 200640 452928 364236
rect 454340 200640 454660 364236
rect 456072 200640 456392 364236
rect 457804 200640 458124 364236
rect 459536 200640 459856 364236
rect 461268 200640 461588 364236
rect 445536 -8054 445856 196236
rect 447268 -8054 447588 196236
rect 449144 -8054 449464 196236
rect 450876 -8054 451196 196236
rect 452608 -8054 452928 196236
rect 454340 -8054 454660 196236
rect 456072 -8054 456392 196236
rect 457804 -8054 458124 196236
rect 459536 -8054 459856 196236
rect 461268 -8054 461588 196236
rect 463144 -8054 463464 711990
rect 464876 -8054 465196 711990
rect 466608 -8054 466928 711990
rect 468340 -8054 468660 711990
rect 470072 -8054 470392 711990
rect 471804 -8054 472124 711990
rect 473536 -8054 473856 711990
rect 475268 -8054 475588 711990
rect 477144 -8054 477464 711990
rect 478876 -8054 479196 711990
rect 480608 -8054 480928 711990
rect 482340 -8054 482660 711990
rect 484072 -8054 484392 711990
rect 485804 -8054 486124 711990
rect 487536 -8054 487856 711990
rect 489268 -8054 489588 711990
rect 491144 -8054 491464 711990
rect 492876 -8054 493196 711990
rect 494608 -8054 494928 711990
rect 496340 -8054 496660 711990
rect 498072 -8054 498392 711990
rect 499804 -8054 500124 711990
rect 501536 -8054 501856 711990
rect 503268 -8054 503588 711990
rect 505144 -8054 505464 711990
rect 506876 -8054 507196 711990
rect 508608 -8054 508928 711990
rect 510340 -8054 510660 711990
rect 512072 -8054 512392 711990
rect 513804 -8054 514124 711990
rect 515536 -8054 515856 711990
rect 517268 -8054 517588 711990
rect 519144 -8054 519464 711990
rect 520876 421752 521196 711990
rect 522608 421752 522928 711990
rect 524340 421752 524660 711990
rect 526072 421752 526392 711990
rect 522608 381752 522928 400008
rect 524340 381752 524660 400008
rect 526072 381752 526392 400008
rect 526072 341752 526392 360008
rect 520876 -8054 521196 240008
rect 522608 -8054 522928 240008
rect 524340 -8054 524660 240008
rect 526072 -8054 526392 240008
rect 527804 -8054 528124 711990
rect 529536 -8054 529856 711990
rect 531268 -8054 531588 711990
rect 533144 -8054 533464 711990
rect 534876 -8054 535196 711990
rect 536608 -8054 536928 711990
rect 538340 -8054 538660 711990
rect 540072 -8054 540392 711990
rect 541804 -8054 542124 711990
rect 543536 -8054 543856 711990
rect 545268 -8054 545588 711990
rect 547144 -8054 547464 711990
rect 548876 -8054 549196 711990
rect 550608 -8054 550928 711990
rect 552340 -8054 552660 711990
rect 554072 -8054 554392 711990
rect 555804 -8054 556124 711990
rect 557536 -8054 557856 711990
rect 559268 -8054 559588 711990
rect 561144 -8054 561464 711990
rect 562876 -8054 563196 711990
rect 564608 -8054 564928 711990
rect 566340 -8054 566660 711990
rect 568072 -8054 568392 711990
rect 569804 -8054 570124 711990
rect 571536 -8054 571856 711990
rect 573268 -8054 573588 711990
rect 575144 -8054 575464 711990
rect 576876 -8054 577196 711990
rect 578608 -8054 578928 711990
rect 580340 -8054 580660 711990
rect 582072 -8054 582392 711990
rect 585710 -2126 587122 706062
rect 587462 -3878 588874 707814
rect 589214 -5630 590626 709566
rect 590966 -7382 592378 711318
rect 592718 -9134 594130 713070
rect 594470 -10886 595882 714822
rect 596222 -12638 597634 716574
rect 597974 -14390 599386 718326
<< obsm4 >>
rect 447668 368560 449064 419632
rect 449544 368560 450796 419632
rect 451276 368560 452528 419632
rect 453008 368560 454260 419632
rect 454740 368560 455992 419632
rect 456472 368560 457724 419632
rect 458204 368560 459456 419632
rect 459936 368560 461188 419632
rect 461668 368560 463064 419632
rect 447529 364316 463064 368560
rect 447668 200560 449064 364316
rect 449544 200560 450796 364316
rect 451276 200560 452528 364316
rect 453008 200560 454260 364316
rect 454740 200560 455992 364316
rect 456472 200560 457724 364316
rect 458204 200560 459456 364316
rect 459936 200560 461188 364316
rect 461668 200560 463064 364316
rect 447529 198356 463064 200560
rect 463544 198356 464796 419632
rect 465276 198356 466528 419632
rect 467008 198356 468260 419632
rect 468740 198356 469992 419632
rect 470472 198356 471724 419632
rect 472204 198356 473456 419632
rect 473936 198356 475188 419632
rect 475668 198356 477064 419632
rect 477544 198356 478796 419632
rect 479276 198356 480528 419632
rect 481008 198356 482260 419632
rect 482740 198356 483992 419632
rect 484472 198356 485724 419632
rect 486204 198356 487456 419632
rect 487936 198356 489188 419632
rect 489668 198356 491064 419632
rect 491544 198356 492796 419632
rect 493276 198356 494528 419632
rect 495008 198356 496260 419632
rect 496740 198356 497992 419632
rect 498472 198356 499724 419632
rect 500204 198356 501456 419632
rect 501936 198356 503188 419632
rect 503668 198356 505064 419632
rect 505544 198356 506796 419632
rect 507276 198356 508528 419632
rect 509008 198356 510260 419632
rect 510740 198356 511992 419632
rect 512472 198356 513724 419632
rect 514204 198356 515456 419632
rect 515936 198356 517188 419632
rect 517668 198356 519064 419632
rect 519544 400088 526992 419632
rect 519544 381672 522528 400088
rect 523008 381672 524260 400088
rect 524740 381672 525992 400088
rect 526472 381672 526992 400088
rect 519544 360088 526992 381672
rect 519544 341672 525992 360088
rect 526472 341672 526992 360088
rect 519544 240088 526992 341672
rect 519544 198356 520796 240088
rect 521276 198356 522528 240088
rect 523008 198356 524260 240088
rect 524740 198356 525992 240088
rect 526472 198356 526992 240088
<< metal5 >>
rect -9126 711370 593050 711990
rect -8166 710410 592090 711030
rect -7206 709450 591130 710070
rect -6246 708490 590170 709110
rect -5286 707530 589210 708150
rect -4326 706570 588250 707190
rect -3366 705610 587290 706230
rect -2406 704650 587122 705270
rect -15462 695685 599386 696005
rect -15462 694618 599386 694938
rect -15462 693551 599386 693871
rect -15462 692484 599386 692804
rect -15462 691417 599386 691737
rect -15462 690350 599386 690670
rect -15462 689283 599386 689603
rect -15462 688216 599386 688536
rect -15462 681685 599386 682005
rect -15462 680618 599386 680938
rect -15462 679551 599386 679871
rect -15462 678484 599386 678804
rect -15462 677417 599386 677737
rect -15462 676350 599386 676670
rect -15462 675283 599386 675603
rect -15462 674216 599386 674536
rect -15462 667685 599386 668005
rect -15462 666618 599386 666938
rect -15462 665551 599386 665871
rect -15462 664484 599386 664804
rect -15462 663417 599386 663737
rect -15462 662350 599386 662670
rect -15462 661283 599386 661603
rect -15462 660216 599386 660536
rect -15462 653685 599386 654005
rect -15462 652618 599386 652938
rect -15462 651551 599386 651871
rect -15462 650484 599386 650804
rect -15462 649417 599386 649737
rect -15462 648350 599386 648670
rect -15462 647283 599386 647603
rect -15462 646216 599386 646536
rect -15462 639685 599386 640005
rect -15462 638618 599386 638938
rect -15462 637551 599386 637871
rect -15462 636484 599386 636804
rect -15462 635417 599386 635737
rect -15462 634350 599386 634670
rect -15462 633283 599386 633603
rect -15462 632216 599386 632536
rect -15462 625685 599386 626005
rect -15462 624618 599386 624938
rect -15462 623551 599386 623871
rect -15462 622484 599386 622804
rect -15462 621417 599386 621737
rect -15462 620350 599386 620670
rect -15462 619283 599386 619603
rect -15462 618216 599386 618536
rect -15462 611685 599386 612005
rect -15462 610618 599386 610938
rect -15462 609551 599386 609871
rect -15462 608484 599386 608804
rect -15462 607417 599386 607737
rect -15462 606350 599386 606670
rect -15462 605283 599386 605603
rect -15462 604216 599386 604536
rect -15462 597685 599386 598005
rect -15462 596618 599386 596938
rect -15462 595551 599386 595871
rect -15462 594484 599386 594804
rect -15462 593417 599386 593737
rect -15462 592350 599386 592670
rect -15462 591283 599386 591603
rect -15462 590216 599386 590536
rect -15462 583685 599386 584005
rect -15462 582618 599386 582938
rect -15462 581551 599386 581871
rect -15462 580484 599386 580804
rect -15462 579417 599386 579737
rect -15462 578350 599386 578670
rect -15462 577283 599386 577603
rect -15462 576216 599386 576536
rect -15462 569685 599386 570005
rect -15462 568618 599386 568938
rect -15462 567551 599386 567871
rect -15462 566484 599386 566804
rect -15462 565417 599386 565737
rect -15462 564350 599386 564670
rect -15462 563283 599386 563603
rect -15462 562216 599386 562536
rect -15462 555685 599386 556005
rect -15462 554618 599386 554938
rect -15462 553551 599386 553871
rect -15462 552484 599386 552804
rect -15462 551417 599386 551737
rect -15462 550350 599386 550670
rect -15462 549283 599386 549603
rect -15462 548216 599386 548536
rect -15462 541685 599386 542005
rect -15462 540618 599386 540938
rect -15462 539551 599386 539871
rect -15462 538484 599386 538804
rect -15462 537417 599386 537737
rect -15462 536350 599386 536670
rect -15462 535283 599386 535603
rect -15462 534216 599386 534536
rect -15462 527685 599386 528005
rect -15462 526618 599386 526938
rect -15462 525551 599386 525871
rect -15462 524484 599386 524804
rect -15462 523417 599386 523737
rect -15462 522350 599386 522670
rect -15462 521283 599386 521603
rect -15462 520216 599386 520536
rect -15462 513685 599386 514005
rect -15462 512618 599386 512938
rect -15462 511551 599386 511871
rect -15462 510484 599386 510804
rect -15462 509417 599386 509737
rect -15462 508350 599386 508670
rect -15462 507283 599386 507603
rect -15462 506216 599386 506536
rect -15462 499685 599386 500005
rect -15462 498618 599386 498938
rect -15462 497551 599386 497871
rect -15462 496484 599386 496804
rect -15462 495417 599386 495737
rect -15462 494350 599386 494670
rect -15462 493283 599386 493603
rect -15462 492216 599386 492536
rect -15462 485685 599386 486005
rect -15462 484618 599386 484938
rect -15462 483551 599386 483871
rect -15462 482484 599386 482804
rect -15462 481417 599386 481737
rect -15462 480350 599386 480670
rect -15462 479283 599386 479603
rect -15462 478216 599386 478536
rect -15462 471685 599386 472005
rect -15462 470618 599386 470938
rect -15462 469551 599386 469871
rect -15462 468484 599386 468804
rect -15462 467417 599386 467737
rect -15462 466350 599386 466670
rect -15462 465283 599386 465603
rect -15462 464216 599386 464536
rect -15462 457685 599386 458005
rect -15462 456618 599386 456938
rect -15462 455551 599386 455871
rect -15462 454484 599386 454804
rect -15462 453417 599386 453737
rect -15462 452350 599386 452670
rect -15462 451283 599386 451603
rect -15462 450216 599386 450536
rect -15462 443685 599386 444005
rect -15462 442618 599386 442938
rect -15462 441551 599386 441871
rect -15462 440484 599386 440804
rect -15462 439417 599386 439737
rect -15462 438350 599386 438670
rect -15462 437283 599386 437603
rect -15462 436216 599386 436536
rect -15462 429685 599386 430005
rect -15462 428618 599386 428938
rect -15462 427551 599386 427871
rect -15462 426484 599386 426804
rect -15462 425417 599386 425737
rect -15462 424350 599386 424670
rect -15462 423283 599386 423603
rect -15462 422216 599386 422536
rect -15462 415685 599386 416005
rect -15462 414618 599386 414938
rect -15462 413551 599386 413871
rect -15462 412484 599386 412804
rect -15462 411417 599386 411737
rect -15462 410350 599386 410670
rect -15462 409283 599386 409603
rect -15462 408216 599386 408536
rect -15462 401685 599386 402005
rect -15462 400618 599386 400938
rect -15462 399551 599386 399871
rect -15462 398484 599386 398804
rect -15462 397417 599386 397737
rect -15462 396350 599386 396670
rect -15462 395283 599386 395603
rect -15462 394216 599386 394536
rect -15462 387685 599386 388005
rect -15462 386618 599386 386938
rect -15462 385551 599386 385871
rect -15462 384484 599386 384804
rect -15462 383417 599386 383737
rect -15462 382350 599386 382670
rect -15462 381283 599386 381603
rect -15462 380216 599386 380536
rect -15462 373685 599386 374005
rect -15462 372618 599386 372938
rect -15462 371551 599386 371871
rect -15462 370484 599386 370804
rect -15462 369417 599386 369737
rect -15462 368350 599386 368670
rect -15462 367283 599386 367603
rect -15462 366216 599386 366536
rect -15462 359685 599386 360005
rect -15462 358618 599386 358938
rect -15462 357551 599386 357871
rect -15462 356484 599386 356804
rect -15462 355417 599386 355737
rect -15462 354350 599386 354670
rect -15462 353283 599386 353603
rect -15462 352216 599386 352536
rect -15462 345685 599386 346005
rect -15462 344618 599386 344938
rect -15462 343551 599386 343871
rect -15462 342484 599386 342804
rect -15462 341417 599386 341737
rect -15462 340350 599386 340670
rect -15462 339283 599386 339603
rect -15462 338216 599386 338536
rect -15462 331685 599386 332005
rect -15462 330618 599386 330938
rect -15462 329551 599386 329871
rect -15462 328484 599386 328804
rect -15462 327417 599386 327737
rect -15462 326350 599386 326670
rect -15462 325283 599386 325603
rect -15462 324216 599386 324536
rect -15462 317685 599386 318005
rect -15462 316618 599386 316938
rect -15462 315551 599386 315871
rect -15462 314484 599386 314804
rect -15462 313417 599386 313737
rect -15462 312350 599386 312670
rect -15462 311283 599386 311603
rect -15462 310216 599386 310536
rect -15462 303685 599386 304005
rect -15462 302618 599386 302938
rect -15462 301551 599386 301871
rect -15462 300484 599386 300804
rect -15462 299417 599386 299737
rect -15462 298350 599386 298670
rect -15462 297283 599386 297603
rect -15462 296216 599386 296536
rect -15462 289685 599386 290005
rect -15462 288618 599386 288938
rect -15462 287551 599386 287871
rect -15462 286484 599386 286804
rect -15462 285417 599386 285737
rect -15462 284350 599386 284670
rect -15462 283283 599386 283603
rect -15462 282216 599386 282536
rect -15462 275685 599386 276005
rect -15462 274618 599386 274938
rect -15462 273551 599386 273871
rect -15462 272484 599386 272804
rect -15462 271417 599386 271737
rect -15462 270350 599386 270670
rect -15462 269283 599386 269603
rect -15462 268216 599386 268536
rect -15462 261685 599386 262005
rect -15462 260618 599386 260938
rect -15462 259551 599386 259871
rect -15462 258484 599386 258804
rect -15462 257417 599386 257737
rect -15462 256350 599386 256670
rect -15462 255283 599386 255603
rect -15462 254216 599386 254536
rect -15462 247685 599386 248005
rect -15462 246618 599386 246938
rect -15462 245551 599386 245871
rect -15462 244484 599386 244804
rect -15462 243417 599386 243737
rect -15462 242350 599386 242670
rect -15462 241283 599386 241603
rect -15462 240216 599386 240536
rect -15462 233685 599386 234005
rect -15462 232618 599386 232938
rect -15462 231551 599386 231871
rect -15462 230484 599386 230804
rect -15462 229417 599386 229737
rect -15462 228350 599386 228670
rect -15462 227283 599386 227603
rect -15462 226216 599386 226536
rect -15462 219685 599386 220005
rect -15462 218618 599386 218938
rect -15462 217551 599386 217871
rect -15462 216484 599386 216804
rect -15462 215417 599386 215737
rect -15462 214350 599386 214670
rect -15462 213283 599386 213603
rect -15462 212216 599386 212536
rect -15462 205685 599386 206005
rect -15462 204618 599386 204938
rect -15462 203551 599386 203871
rect -15462 202484 599386 202804
rect -15462 201417 599386 201737
rect -15462 200350 599386 200670
rect -15462 199283 599386 199603
rect -15462 198216 599386 198536
rect -15462 191685 599386 192005
rect -15462 190618 599386 190938
rect -15462 189551 599386 189871
rect -15462 188484 599386 188804
rect -15462 187417 599386 187737
rect -15462 186350 599386 186670
rect -15462 185283 599386 185603
rect -15462 184216 599386 184536
rect -15462 177685 599386 178005
rect -15462 176618 599386 176938
rect -15462 175551 599386 175871
rect -15462 174484 599386 174804
rect -15462 173417 599386 173737
rect -15462 172350 599386 172670
rect -15462 171283 599386 171603
rect -15462 170216 599386 170536
rect -15462 163685 599386 164005
rect -15462 162618 599386 162938
rect -15462 161551 599386 161871
rect -15462 160484 599386 160804
rect -15462 159417 599386 159737
rect -15462 158350 599386 158670
rect -15462 157283 599386 157603
rect -15462 156216 599386 156536
rect -15462 149685 599386 150005
rect -15462 148618 599386 148938
rect -15462 147551 599386 147871
rect -15462 146484 599386 146804
rect -15462 145417 599386 145737
rect -15462 144350 599386 144670
rect -15462 143283 599386 143603
rect -15462 142216 599386 142536
rect -15462 135685 599386 136005
rect -15462 134618 599386 134938
rect -15462 133551 599386 133871
rect -15462 132484 599386 132804
rect -15462 131417 599386 131737
rect -15462 130350 599386 130670
rect -15462 129283 599386 129603
rect -15462 128216 599386 128536
rect -15462 121685 599386 122005
rect -15462 120618 599386 120938
rect -15462 119551 599386 119871
rect -15462 118484 599386 118804
rect -15462 117417 599386 117737
rect -15462 116350 599386 116670
rect -15462 115283 599386 115603
rect -15462 114216 599386 114536
rect -15462 107685 599386 108005
rect -15462 106618 599386 106938
rect -15462 105551 599386 105871
rect -15462 104484 599386 104804
rect -15462 103417 599386 103737
rect -15462 102350 599386 102670
rect -15462 101283 599386 101603
rect -15462 100216 599386 100536
rect -15462 93685 599386 94005
rect -15462 92618 599386 92938
rect -15462 91551 599386 91871
rect -15462 90484 599386 90804
rect -15462 89417 599386 89737
rect -15462 88350 599386 88670
rect -15462 87283 599386 87603
rect -15462 86216 599386 86536
rect -15462 79685 599386 80005
rect -15462 78618 599386 78938
rect -15462 77551 599386 77871
rect -15462 76484 599386 76804
rect -15462 75417 599386 75737
rect -15462 74350 599386 74670
rect -15462 73283 599386 73603
rect -15462 72216 599386 72536
rect -15462 65685 599386 66005
rect -15462 64618 599386 64938
rect -15462 63551 599386 63871
rect -15462 62484 599386 62804
rect -15462 61417 599386 61737
rect -15462 60350 599386 60670
rect -15462 59283 599386 59603
rect -15462 58216 599386 58536
rect -15462 51685 599386 52005
rect -15462 50618 599386 50938
rect -15462 49551 599386 49871
rect -15462 48484 599386 48804
rect -15462 47417 599386 47737
rect -15462 46350 599386 46670
rect -15462 45283 599386 45603
rect -15462 44216 599386 44536
rect -15462 37685 599386 38005
rect -15462 36618 599386 36938
rect -15462 35551 599386 35871
rect -15462 34484 599386 34804
rect -15462 33417 599386 33737
rect -15462 32350 599386 32670
rect -15462 31283 599386 31603
rect -15462 30216 599386 30536
rect -15462 23685 599386 24005
rect -15462 22618 599386 22938
rect -15462 21551 599386 21871
rect -15462 20484 599386 20804
rect -15462 19417 599386 19737
rect -15462 18350 599386 18670
rect -15462 17283 599386 17603
rect -15462 16216 599386 16536
rect -15462 9685 599386 10005
rect -15462 8618 599386 8938
rect -15462 7551 599386 7871
rect -15462 6484 599386 6804
rect -15462 5417 599386 5737
rect -15462 4350 599386 4670
rect -15462 3283 599386 3603
rect -15462 2216 599386 2536
rect -2406 -1334 587122 -714
rect -3366 -2294 587290 -1674
rect -4326 -3254 588250 -2634
rect -5286 -4214 589210 -3594
rect -6246 -5174 590170 -4554
rect -7206 -6134 591130 -5514
rect -8166 -7094 592090 -6474
rect -9126 -8054 593050 -7434
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -3198 -2126 -1786 706062 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2406 -1334 587122 -714 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2406 704650 587122 705270 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585710 -2126 587122 706062 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 1144 -8054 1464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 15144 -8054 15464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 29144 -8054 29464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 43144 -8054 43464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 57144 -8054 57464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 71144 -8054 71464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 85144 -8054 85464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 99144 -8054 99464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 113144 -8054 113464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127144 -8054 127464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 141144 -8054 141464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 155144 -8054 155464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 169144 -8054 169464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 183144 -8054 183464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 197144 -8054 197464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 211144 -8054 211464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 225144 -8054 225464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 239144 -8054 239464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253144 -8054 253464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 267144 -8054 267464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 281144 -8054 281464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 295144 -8054 295464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 309144 -8054 309464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 323144 -8054 323464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 337144 -8054 337464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 351144 -8054 351464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 365144 -8054 365464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 379144 -8054 379464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 393144 -8054 393464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 407144 -8054 407464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 421144 -8054 421464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 435144 -8054 435464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 449144 -8054 449464 196236 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 449144 200640 449464 364236 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 449144 368640 449464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 463144 -8054 463464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 477144 -8054 477464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 491144 -8054 491464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505144 -8054 505464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 519144 -8054 519464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 533144 -8054 533464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 547144 -8054 547464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 561144 -8054 561464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 575144 -8054 575464 711990 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 2216 599386 2536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 16216 599386 16536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 30216 599386 30536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 44216 599386 44536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 58216 599386 58536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 72216 599386 72536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 86216 599386 86536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 100216 599386 100536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 114216 599386 114536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 128216 599386 128536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 142216 599386 142536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 156216 599386 156536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 170216 599386 170536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 184216 599386 184536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 198216 599386 198536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 212216 599386 212536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 226216 599386 226536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 240216 599386 240536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 254216 599386 254536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 268216 599386 268536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 282216 599386 282536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 296216 599386 296536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 310216 599386 310536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 324216 599386 324536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 338216 599386 338536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 352216 599386 352536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 366216 599386 366536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 380216 599386 380536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 394216 599386 394536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 408216 599386 408536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 422216 599386 422536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 436216 599386 436536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 450216 599386 450536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 464216 599386 464536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 478216 599386 478536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 492216 599386 492536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 506216 599386 506536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 520216 599386 520536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 534216 599386 534536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 548216 599386 548536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 562216 599386 562536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 576216 599386 576536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 590216 599386 590536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 604216 599386 604536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 618216 599386 618536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 632216 599386 632536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 646216 599386 646536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 660216 599386 660536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 674216 599386 674536 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -15462 688216 599386 688536 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -6702 -5630 -5290 709566 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4326 -3254 588250 -2634 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4326 706570 588250 707190 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 589214 -5630 590626 709566 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 4608 -8054 4928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 18608 -8054 18928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 32608 -8054 32928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 46608 -8054 46928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 60608 -8054 60928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 74608 -8054 74928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 88608 -8054 88928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 102608 -8054 102928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 116608 -8054 116928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 130608 -8054 130928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 144608 -8054 144928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 158608 -8054 158928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 172608 -8054 172928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 186608 -8054 186928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 200608 -8054 200928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 214608 -8054 214928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 228608 -8054 228928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 242608 -8054 242928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 256608 -8054 256928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 270608 -8054 270928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 284608 -8054 284928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 298608 -8054 298928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 312608 -8054 312928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 326608 -8054 326928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 340608 -8054 340928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 354608 -8054 354928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 368608 -8054 368928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 382608 -8054 382928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 396608 -8054 396928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 410608 -8054 410928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 424608 -8054 424928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 438608 -8054 438928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 452608 -8054 452928 196236 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 452608 200640 452928 364236 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 452608 368640 452928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 466608 -8054 466928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 480608 -8054 480928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 494608 -8054 494928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 508608 -8054 508928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 522608 -8054 522928 240008 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 522608 381752 522928 400008 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 522608 421752 522928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 536608 -8054 536928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 550608 -8054 550928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 564608 -8054 564928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 578608 -8054 578928 711990 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 4350 599386 4670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 18350 599386 18670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 32350 599386 32670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 46350 599386 46670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 60350 599386 60670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 74350 599386 74670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 88350 599386 88670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 102350 599386 102670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 116350 599386 116670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 130350 599386 130670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 144350 599386 144670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 158350 599386 158670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 172350 599386 172670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 186350 599386 186670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 200350 599386 200670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 214350 599386 214670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 228350 599386 228670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 242350 599386 242670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 256350 599386 256670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 270350 599386 270670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 284350 599386 284670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 298350 599386 298670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 312350 599386 312670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 326350 599386 326670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 340350 599386 340670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 354350 599386 354670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 368350 599386 368670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 382350 599386 382670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 396350 599386 396670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 410350 599386 410670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 424350 599386 424670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 438350 599386 438670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 452350 599386 452670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 466350 599386 466670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 480350 599386 480670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 494350 599386 494670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 508350 599386 508670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 522350 599386 522670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 536350 599386 536670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 550350 599386 550670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 564350 599386 564670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 578350 599386 578670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 592350 599386 592670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 606350 599386 606670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 620350 599386 620670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 634350 599386 634670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 648350 599386 648670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 662350 599386 662670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 676350 599386 676670 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -15462 690350 599386 690670 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -10206 -9134 -8794 713070 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -6246 -5174 590170 -4554 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -6246 708490 590170 709110 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 592718 -9134 594130 713070 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 8072 -8054 8392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 22072 -8054 22392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 36072 -8054 36392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 50072 -8054 50392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 64072 -8054 64392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 78072 -8054 78392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 92072 -8054 92392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 106072 -8054 106392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 120072 -8054 120392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 134072 -8054 134392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 148072 -8054 148392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 162072 -8054 162392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 176072 -8054 176392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 190072 -8054 190392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 204072 -8054 204392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 218072 -8054 218392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 232072 -8054 232392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 246072 -8054 246392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 260072 -8054 260392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 274072 -8054 274392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 288072 -8054 288392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 302072 -8054 302392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 316072 -8054 316392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 330072 -8054 330392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 344072 -8054 344392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 358072 -8054 358392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 372072 -8054 372392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 386072 -8054 386392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 400072 -8054 400392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 414072 -8054 414392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 428072 -8054 428392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 442072 -8054 442392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 456072 -8054 456392 196236 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 456072 200640 456392 364236 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 456072 368640 456392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 470072 -8054 470392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 484072 -8054 484392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 498072 -8054 498392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 512072 -8054 512392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526072 -8054 526392 240008 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526072 341752 526392 360008 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526072 381752 526392 400008 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526072 421752 526392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 540072 -8054 540392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 554072 -8054 554392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 568072 -8054 568392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 582072 -8054 582392 711990 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 6484 599386 6804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 20484 599386 20804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 34484 599386 34804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 48484 599386 48804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 62484 599386 62804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 76484 599386 76804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 90484 599386 90804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 104484 599386 104804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 118484 599386 118804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 132484 599386 132804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 146484 599386 146804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 160484 599386 160804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 174484 599386 174804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 188484 599386 188804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 202484 599386 202804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 216484 599386 216804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 230484 599386 230804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 244484 599386 244804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 258484 599386 258804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 272484 599386 272804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 286484 599386 286804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 300484 599386 300804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 314484 599386 314804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 328484 599386 328804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 342484 599386 342804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 356484 599386 356804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 370484 599386 370804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 384484 599386 384804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 398484 599386 398804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 412484 599386 412804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 426484 599386 426804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 440484 599386 440804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 454484 599386 454804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 468484 599386 468804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 482484 599386 482804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 496484 599386 496804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 510484 599386 510804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 524484 599386 524804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 538484 599386 538804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 552484 599386 552804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 566484 599386 566804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 580484 599386 580804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 594484 599386 594804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 608484 599386 608804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 622484 599386 622804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 636484 599386 636804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 650484 599386 650804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 664484 599386 664804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 678484 599386 678804 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -15462 692484 599386 692804 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -13710 -12638 -12298 716574 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8166 -7094 592090 -6474 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8166 710410 592090 711030 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 596222 -12638 597634 716574 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 11536 -8054 11856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 25536 -8054 25856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 39536 -8054 39856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 53536 -8054 53856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 67536 -8054 67856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 81536 -8054 81856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 95536 -8054 95856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 109536 -8054 109856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 123536 -8054 123856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 137536 -8054 137856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 151536 -8054 151856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 165536 -8054 165856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 179536 -8054 179856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 193536 -8054 193856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 207536 -8054 207856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 221536 -8054 221856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 235536 -8054 235856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 249536 -8054 249856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 263536 -8054 263856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 277536 -8054 277856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 291536 -8054 291856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 305536 -8054 305856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 319536 -8054 319856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 333536 -8054 333856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 347536 -8054 347856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 361536 -8054 361856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 375536 -8054 375856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 389536 -8054 389856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 403536 -8054 403856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 417536 -8054 417856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 431536 -8054 431856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 445536 -8054 445856 196236 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 445536 200640 445856 364236 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 445536 368640 445856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 459536 -8054 459856 196236 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 459536 200640 459856 364236 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 459536 368640 459856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 473536 -8054 473856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 487536 -8054 487856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 501536 -8054 501856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 515536 -8054 515856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 529536 -8054 529856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 543536 -8054 543856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 557536 -8054 557856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 571536 -8054 571856 711990 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 8618 599386 8938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 22618 599386 22938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 36618 599386 36938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 50618 599386 50938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 64618 599386 64938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 78618 599386 78938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 92618 599386 92938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 106618 599386 106938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 120618 599386 120938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 134618 599386 134938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 148618 599386 148938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 162618 599386 162938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 176618 599386 176938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 190618 599386 190938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 204618 599386 204938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 218618 599386 218938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 232618 599386 232938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 246618 599386 246938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 260618 599386 260938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 274618 599386 274938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 288618 599386 288938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 302618 599386 302938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 316618 599386 316938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 330618 599386 330938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 344618 599386 344938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 358618 599386 358938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 372618 599386 372938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 386618 599386 386938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 400618 599386 400938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 414618 599386 414938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 428618 599386 428938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 442618 599386 442938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 456618 599386 456938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 470618 599386 470938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 484618 599386 484938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 498618 599386 498938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 512618 599386 512938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 526618 599386 526938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 540618 599386 540938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 554618 599386 554938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 568618 599386 568938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 582618 599386 582938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 596618 599386 596938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 610618 599386 610938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 624618 599386 624938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 638618 599386 638938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 652618 599386 652938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 666618 599386 666938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 680618 599386 680938 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -15462 694618 599386 694938 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -11958 -10886 -10546 714822 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -7206 -6134 591130 -5514 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -7206 709450 591130 710070 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 594470 -10886 595882 714822 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 9804 -8054 10124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 23804 -8054 24124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 37804 -8054 38124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 51804 -8054 52124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 65804 -8054 66124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 79804 -8054 80124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 93804 -8054 94124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 107804 -8054 108124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 121804 -8054 122124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 135804 -8054 136124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 149804 -8054 150124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 163804 -8054 164124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 177804 -8054 178124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 191804 -8054 192124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 205804 -8054 206124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 219804 -8054 220124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 233804 -8054 234124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 247804 -8054 248124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 261804 -8054 262124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 275804 -8054 276124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 289804 -8054 290124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 303804 -8054 304124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 317804 -8054 318124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 331804 -8054 332124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 345804 -8054 346124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 359804 -8054 360124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 373804 -8054 374124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 387804 -8054 388124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 401804 -8054 402124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 415804 -8054 416124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 429804 -8054 430124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 443804 -8054 444124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 457804 -8054 458124 196236 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 457804 200640 458124 364236 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 457804 368640 458124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 471804 -8054 472124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 485804 -8054 486124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 499804 -8054 500124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 513804 -8054 514124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 527804 -8054 528124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 541804 -8054 542124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 555804 -8054 556124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 569804 -8054 570124 711990 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 7551 599386 7871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 21551 599386 21871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 35551 599386 35871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 49551 599386 49871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 63551 599386 63871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 77551 599386 77871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 91551 599386 91871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 105551 599386 105871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 119551 599386 119871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 133551 599386 133871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 147551 599386 147871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 161551 599386 161871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 175551 599386 175871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 189551 599386 189871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 203551 599386 203871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 217551 599386 217871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 231551 599386 231871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 245551 599386 245871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 259551 599386 259871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 273551 599386 273871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 287551 599386 287871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 301551 599386 301871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 315551 599386 315871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 329551 599386 329871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 343551 599386 343871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 357551 599386 357871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 371551 599386 371871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 385551 599386 385871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 399551 599386 399871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 413551 599386 413871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 427551 599386 427871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 441551 599386 441871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 455551 599386 455871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 469551 599386 469871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 483551 599386 483871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 497551 599386 497871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 511551 599386 511871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 525551 599386 525871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 539551 599386 539871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 553551 599386 553871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 567551 599386 567871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 581551 599386 581871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 595551 599386 595871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 609551 599386 609871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 623551 599386 623871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 637551 599386 637871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 651551 599386 651871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 665551 599386 665871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 679551 599386 679871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -15462 693551 599386 693871 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -15462 -14390 -14050 718326 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9126 -8054 593050 -7434 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9126 711370 593050 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 597974 -14390 599386 718326 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 13268 -8054 13588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 27268 -8054 27588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 41268 -8054 41588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 55268 -8054 55588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 69268 -8054 69588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 83268 -8054 83588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 97268 -8054 97588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 111268 -8054 111588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 125268 -8054 125588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 139268 -8054 139588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 153268 -8054 153588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 167268 -8054 167588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 181268 -8054 181588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 195268 -8054 195588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 209268 -8054 209588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 223268 -8054 223588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 237268 -8054 237588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 251268 -8054 251588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 265268 -8054 265588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 279268 -8054 279588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 293268 -8054 293588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 307268 -8054 307588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 321268 -8054 321588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 335268 -8054 335588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 349268 -8054 349588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 363268 -8054 363588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 377268 -8054 377588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 391268 -8054 391588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 405268 -8054 405588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 419268 -8054 419588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 433268 -8054 433588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 447268 -8054 447588 196236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 447268 200640 447588 364236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 447268 368640 447588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 461268 -8054 461588 196236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 461268 200640 461588 364236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 461268 368640 461588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 475268 -8054 475588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 489268 -8054 489588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 503268 -8054 503588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 517268 -8054 517588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 531268 -8054 531588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 545268 -8054 545588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 559268 -8054 559588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 573268 -8054 573588 711990 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 9685 599386 10005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 23685 599386 24005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 37685 599386 38005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 51685 599386 52005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 65685 599386 66005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 79685 599386 80005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 93685 599386 94005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 107685 599386 108005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 121685 599386 122005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 135685 599386 136005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 149685 599386 150005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 163685 599386 164005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 177685 599386 178005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 191685 599386 192005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 205685 599386 206005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 219685 599386 220005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 233685 599386 234005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 247685 599386 248005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 261685 599386 262005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 275685 599386 276005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 289685 599386 290005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 303685 599386 304005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 317685 599386 318005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 331685 599386 332005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 345685 599386 346005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 359685 599386 360005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 373685 599386 374005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 387685 599386 388005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 401685 599386 402005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 415685 599386 416005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 429685 599386 430005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 443685 599386 444005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 457685 599386 458005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 471685 599386 472005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 485685 599386 486005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 499685 599386 500005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 513685 599386 514005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 527685 599386 528005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 541685 599386 542005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 555685 599386 556005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 569685 599386 570005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 583685 599386 584005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 597685 599386 598005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 611685 599386 612005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 625685 599386 626005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 639685 599386 640005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 653685 599386 654005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 667685 599386 668005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 681685 599386 682005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -15462 695685 599386 696005 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -4950 -3878 -3538 707814 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -3366 -2294 587290 -1674 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -3366 705610 587290 706230 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 587462 -3878 588874 707814 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 2876 -8054 3196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 16876 -8054 17196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 30876 -8054 31196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 44876 -8054 45196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 58876 -8054 59196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 72876 -8054 73196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 86876 -8054 87196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 100876 -8054 101196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 114876 -8054 115196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 128876 -8054 129196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 142876 -8054 143196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 156876 -8054 157196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 170876 -8054 171196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 184876 -8054 185196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 198876 -8054 199196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 212876 -8054 213196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 226876 -8054 227196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 240876 -8054 241196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 254876 -8054 255196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 268876 -8054 269196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 282876 -8054 283196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 296876 -8054 297196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 310876 -8054 311196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 324876 -8054 325196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 338876 -8054 339196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 352876 -8054 353196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 366876 -8054 367196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 380876 -8054 381196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 394876 -8054 395196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 408876 -8054 409196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 422876 -8054 423196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 436876 -8054 437196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 450876 -8054 451196 196236 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 450876 200640 451196 364236 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 450876 368640 451196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 464876 -8054 465196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 478876 -8054 479196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 492876 -8054 493196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 506876 -8054 507196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 520876 -8054 521196 240008 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 520876 421752 521196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 534876 -8054 535196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 548876 -8054 549196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 562876 -8054 563196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 576876 -8054 577196 711990 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 3283 599386 3603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 17283 599386 17603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 31283 599386 31603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 45283 599386 45603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 59283 599386 59603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 73283 599386 73603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 87283 599386 87603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 101283 599386 101603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 115283 599386 115603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 129283 599386 129603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 143283 599386 143603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 157283 599386 157603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 171283 599386 171603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 185283 599386 185603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 199283 599386 199603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 213283 599386 213603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 227283 599386 227603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 241283 599386 241603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 255283 599386 255603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 269283 599386 269603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 283283 599386 283603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 297283 599386 297603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 311283 599386 311603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 325283 599386 325603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 339283 599386 339603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 353283 599386 353603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 367283 599386 367603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 381283 599386 381603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 395283 599386 395603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 409283 599386 409603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 423283 599386 423603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 437283 599386 437603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 451283 599386 451603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 465283 599386 465603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 479283 599386 479603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 493283 599386 493603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 507283 599386 507603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 521283 599386 521603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 535283 599386 535603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 549283 599386 549603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 563283 599386 563603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 577283 599386 577603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 591283 599386 591603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 605283 599386 605603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 619283 599386 619603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 633283 599386 633603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 647283 599386 647603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 661283 599386 661603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 675283 599386 675603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -15462 689283 599386 689603 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -8454 -7382 -7042 711318 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5286 -4214 589210 -3594 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5286 707530 589210 708150 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 590966 -7382 592378 711318 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 6340 -8054 6660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 20340 -8054 20660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 34340 -8054 34660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 48340 -8054 48660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 62340 -8054 62660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 76340 -8054 76660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 90340 -8054 90660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 104340 -8054 104660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 118340 -8054 118660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 132340 -8054 132660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 146340 -8054 146660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 160340 -8054 160660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 174340 -8054 174660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 188340 -8054 188660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 202340 -8054 202660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 216340 -8054 216660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 230340 -8054 230660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 244340 -8054 244660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 258340 -8054 258660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 272340 -8054 272660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 286340 -8054 286660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 300340 -8054 300660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 314340 -8054 314660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 328340 -8054 328660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 342340 -8054 342660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 356340 -8054 356660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 370340 -8054 370660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 384340 -8054 384660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 398340 -8054 398660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 412340 -8054 412660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 426340 -8054 426660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 440340 -8054 440660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 454340 -8054 454660 196236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 454340 200640 454660 364236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 454340 368640 454660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 468340 -8054 468660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 482340 -8054 482660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 496340 -8054 496660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 510340 -8054 510660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 524340 -8054 524660 240008 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 524340 381752 524660 400008 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 524340 421752 524660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 538340 -8054 538660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 552340 -8054 552660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 566340 -8054 566660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 580340 -8054 580660 711990 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 5417 599386 5737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 19417 599386 19737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 33417 599386 33737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 47417 599386 47737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 61417 599386 61737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 75417 599386 75737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 89417 599386 89737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 103417 599386 103737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 117417 599386 117737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 131417 599386 131737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 145417 599386 145737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 159417 599386 159737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 173417 599386 173737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 187417 599386 187737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 201417 599386 201737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 215417 599386 215737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 229417 599386 229737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 243417 599386 243737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 257417 599386 257737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 271417 599386 271737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 285417 599386 285737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 299417 599386 299737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 313417 599386 313737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 327417 599386 327737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 341417 599386 341737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 355417 599386 355737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 369417 599386 369737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 383417 599386 383737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 397417 599386 397737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 411417 599386 411737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 425417 599386 425737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 439417 599386 439737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 453417 599386 453737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 467417 599386 467737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 481417 599386 481737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 495417 599386 495737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 509417 599386 509737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 523417 599386 523737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 537417 599386 537737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 551417 599386 551737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 565417 599386 565737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 579417 599386 579737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 593417 599386 593737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 607417 599386 607737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 621417 599386 621737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 635417 599386 635737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 649417 599386 649737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 663417 599386 663737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 677417 599386 677737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -15462 691417 599386 691737 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4379016
string GDS_FILE /import/yukari1/lrburle/google_ring_oscillator/caravel/openlane/user_project_wrapper/runs/24_02_29_10_18/results/signoff/user_project_wrapper.magic.gds
string GDS_START 2369216
<< end >>

