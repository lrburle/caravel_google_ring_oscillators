magic
tech sky130A
magscale 1 2
timestamp 1716047795
<< nwell >>
rect 4996 1462 7827 1749
rect 9578 1636 9636 1694
rect 10670 1641 10701 1649
rect 12630 1636 12688 1694
rect 13724 1641 13760 1653
rect 15682 1636 15740 1694
rect 16791 1641 16816 1647
rect 18734 1636 18792 1694
rect 19826 1641 19856 1649
rect 4996 1407 5392 1462
rect 5436 1407 7827 1462
rect 4996 1087 20809 1407
rect 4996 820 7827 1087
rect 8480 985 8538 1043
rect 11532 985 11590 1043
rect 14584 985 14642 1043
rect 17636 985 17694 1043
rect 20688 985 20746 1043
<< ndiff >>
rect 8491 441 8526 475
rect 11543 441 11578 475
rect 14595 441 14630 475
rect 17647 441 17682 475
rect 20699 441 20734 475
<< pdiff >>
rect 5035 1648 5069 1682
rect 5029 1641 5078 1647
rect 6528 1636 6584 1694
rect 9580 1636 9636 1694
rect 12630 1636 12688 1694
rect 15684 1636 15740 1694
rect 18736 1636 18792 1694
<< locali >>
rect 0 2173 20800 2493
rect 5396 1407 5430 1471
rect 0 1087 20809 1407
rect 0 0 20809 320
<< viali >>
rect 5035 1648 5069 1682
rect 8492 441 8526 475
rect 11544 441 11578 475
rect 14596 441 14630 475
rect 17648 441 17682 475
rect 20700 441 20734 475
<< metal1 >>
rect 0 2173 20800 2493
rect 20727 2011 20735 2013
rect 20695 1999 20747 2011
rect 20695 1983 20759 1999
rect 20695 1977 20765 1983
rect 5292 1864 5298 1922
rect 5356 1864 5362 1922
rect 20695 1919 20701 1977
rect 20759 1919 20765 1977
rect 20695 1913 20765 1919
rect 8491 1854 8561 1860
rect 6927 1843 6997 1849
rect 6927 1785 6933 1843
rect 6991 1785 6997 1843
rect 6927 1779 6997 1785
rect 8491 1796 8497 1854
rect 8555 1796 8561 1854
rect 11542 1854 11613 1861
rect 8491 1790 8561 1796
rect 9979 1845 10049 1851
rect 8491 1773 8550 1790
rect 9979 1787 9985 1845
rect 10043 1787 10049 1845
rect 9979 1781 10049 1787
rect 11542 1796 11549 1854
rect 11607 1796 11613 1854
rect 14586 1854 14656 1860
rect 11542 1790 11613 1796
rect 13031 1845 13101 1851
rect 5217 1715 5223 1773
rect 5281 1715 5287 1773
rect 11542 1772 11602 1790
rect 13031 1787 13037 1845
rect 13095 1787 13101 1845
rect 13031 1781 13101 1787
rect 14586 1796 14592 1854
rect 14650 1796 14656 1854
rect 17638 1854 17708 1860
rect 14586 1790 14656 1796
rect 16084 1845 16154 1851
rect 14586 1772 14654 1790
rect 16084 1787 16090 1845
rect 16148 1787 16154 1845
rect 16084 1781 16154 1787
rect 17638 1796 17644 1854
rect 17702 1796 17708 1854
rect 17638 1790 17708 1796
rect 19135 1845 19205 1851
rect 17638 1772 17706 1790
rect 19135 1787 19141 1845
rect 19199 1787 19205 1845
rect 19135 1781 19205 1787
rect 5024 1682 5082 1687
rect 5024 1647 5029 1682
rect 5075 1647 5082 1682
rect 5024 1641 5082 1647
rect 6526 1636 6584 1694
rect 7640 1641 7666 1648
rect 9578 1636 9636 1694
rect 10670 1641 10701 1649
rect 12630 1636 12688 1694
rect 13724 1641 13760 1653
rect 15682 1636 15740 1694
rect 16791 1641 16816 1647
rect 18734 1636 18792 1694
rect 19826 1641 19856 1649
rect 0 1087 20809 1407
rect 0 0 20809 320
<< via1 >>
rect 5298 1864 5356 1922
rect 20701 1919 20759 1977
rect 6933 1785 6991 1843
rect 8497 1796 8555 1854
rect 9985 1787 10043 1845
rect 11549 1796 11607 1854
rect 5223 1715 5281 1773
rect 13037 1787 13095 1845
rect 14592 1796 14650 1854
rect 16090 1787 16148 1845
rect 17644 1796 17702 1854
rect 19141 1787 19199 1845
<< metal2 >>
rect 5235 2138 20735 2172
rect 5235 1779 5269 2138
rect 20701 1983 20735 2138
rect 20695 1977 20765 1983
rect 5298 1922 5356 1928
rect 20695 1919 20701 1977
rect 20759 1919 20765 1977
rect 20695 1913 20765 1919
rect 5356 1905 5362 1906
rect 5356 1871 5542 1905
rect 5298 1858 5356 1864
rect 5508 1829 5542 1871
rect 8491 1854 8561 1860
rect 6927 1843 6997 1849
rect 6927 1829 6933 1843
rect 5508 1795 6933 1829
rect 6927 1785 6933 1795
rect 6991 1785 6997 1843
rect 8491 1796 8497 1854
rect 8555 1836 8561 1854
rect 11543 1854 11613 1860
rect 9979 1845 10049 1851
rect 9979 1836 9985 1845
rect 8555 1796 9985 1836
rect 8491 1790 8561 1796
rect 6927 1779 6997 1785
rect 9979 1787 9985 1796
rect 10043 1787 10049 1845
rect 11543 1796 11549 1854
rect 11607 1836 11613 1854
rect 14586 1854 14656 1860
rect 13031 1845 13101 1851
rect 13031 1836 13037 1845
rect 11607 1796 13037 1836
rect 11543 1790 11613 1796
rect 9979 1781 10049 1787
rect 13031 1787 13037 1796
rect 13095 1787 13101 1845
rect 14586 1796 14592 1854
rect 14650 1836 14656 1854
rect 17638 1854 17708 1860
rect 16084 1845 16154 1851
rect 16084 1836 16090 1845
rect 14650 1796 16090 1836
rect 14586 1790 14656 1796
rect 13031 1781 13101 1787
rect 16084 1787 16090 1796
rect 16148 1787 16154 1845
rect 17638 1796 17644 1854
rect 17702 1836 17708 1854
rect 19135 1845 19205 1851
rect 19135 1836 19141 1845
rect 17702 1796 19141 1836
rect 17638 1790 17708 1796
rect 16084 1781 16154 1787
rect 19135 1787 19141 1796
rect 19199 1787 19205 1845
rect 19135 1781 19205 1787
rect 5223 1773 5281 1779
rect 5223 1709 5281 1715
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1714057206
transform 1 0 4999 0 -1 2234
box -10 0 552 902
use sky130_osu_single_mpr2xa_8_b0r1  sky130_osu_single_mpr2xa_8_b0r1_0
timestamp 1716047795
transform 1 0 17757 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2xa_8_b0r1  sky130_osu_single_mpr2xa_8_b0r1_1
timestamp 1716047795
transform 1 0 5549 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2xa_8_b0r1  sky130_osu_single_mpr2xa_8_b0r1_2
timestamp 1716047795
transform 1 0 8601 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2xa_8_b0r1  sky130_osu_single_mpr2xa_8_b0r1_3
timestamp 1716047795
transform 1 0 11653 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2xa_8_b0r1  sky130_osu_single_mpr2xa_8_b0r1_4
timestamp 1716047795
transform 1 0 14705 0 1 0
box 0 0 3052 2493
<< labels >>
flabel metal1 s 5024 1641 5082 1687 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel viali s 6538 1648 6572 1682 0 FreeSans 100 0 0 0 s1
port 16 nw signal input
flabel viali s 9590 1648 9624 1682 0 FreeSans 100 0 0 0 s2
port 17 nw signal input
flabel viali s 12642 1648 12676 1682 0 FreeSans 100 0 0 0 s3
port 18 nw signal input
flabel viali s 15694 1648 15728 1682 0 FreeSans 100 0 0 0 s4
port 19 nw signal input
flabel viali s 18746 1648 18780 1682 0 FreeSans 100 0 0 0 s5
port 20 nw signal input
flabel viali s 8492 441 8526 475 0 FreeSans 100 0 0 0 X1_Y1
port 6 se signal output
flabel viali s 11544 441 11578 475 0 FreeSans 100 0 0 0 X2_Y1
port 7 se signal output
flabel viali s 14596 441 14630 475 0 FreeSans 100 0 0 0 X3_Y1
port 8 se signal output
flabel viali s 17648 441 17682 475 0 FreeSans 100 0 0 0 X4_Y1
port 9 se signal output
flabel viali s 20700 441 20734 475 0 FreeSans 100 0 0 0 X5_Y1
port 10 se signal output
flabel metal1 s 0 2173 20800 2493 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 0 1087 20809 1407 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 0 0 20809 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
<< end >>
