magic
tech sky130A
magscale 1 2
timestamp 1710282110
<< nwell >>
rect -38 630 1510 827
rect -43 462 1510 630
rect -38 261 1510 462
<< pwell >>
rect -25 1105 95 1148
rect -25 1067 154 1105
rect 580 1098 614 1105
rect 399 1076 614 1098
rect 557 1067 614 1076
rect 1042 1067 1076 1105
rect 1318 1099 1352 1105
rect 1318 1077 1432 1099
rect 1318 1067 1375 1077
rect -25 1028 367 1067
rect 97 885 367 1028
rect 557 885 1375 1067
rect 3 60 1463 203
rect -25 21 1463 60
rect -25 -17 247 21
rect 488 -17 616 21
rect 1409 -17 1443 21
rect -25 -60 95 -17
<< scnmos >>
rect 175 911 205 1041
rect 259 911 289 1041
rect 635 911 665 1041
rect 719 911 749 1041
rect 907 911 937 1041
rect 991 911 1021 1041
rect 1183 911 1213 1041
rect 1267 911 1297 1041
rect 81 47 111 177
rect 165 47 195 177
rect 359 47 389 177
rect 443 47 473 177
rect 631 47 661 177
rect 715 47 745 177
rect 919 47 949 177
rect 1103 47 1133 177
rect 1187 47 1217 177
rect 1271 47 1301 177
rect 1355 47 1385 177
<< scpmoshvt >>
rect 175 591 205 791
rect 259 591 289 791
rect 635 591 665 791
rect 719 591 749 791
rect 907 591 937 791
rect 991 591 1021 791
rect 1183 591 1213 791
rect 1267 591 1297 791
rect 81 297 111 497
rect 165 297 195 497
rect 371 297 401 497
rect 443 297 473 497
rect 631 297 661 497
rect 703 297 733 497
rect 915 297 945 497
rect 1103 297 1133 497
rect 1187 297 1217 497
rect 1271 297 1301 497
rect 1355 297 1385 497
<< ndiff >>
rect 123 1029 175 1041
rect 123 995 131 1029
rect 165 995 175 1029
rect 123 961 175 995
rect 123 927 131 961
rect 165 927 175 961
rect 123 911 175 927
rect 205 911 259 1041
rect 289 1029 341 1041
rect 289 995 299 1029
rect 333 995 341 1029
rect 289 961 341 995
rect 289 927 299 961
rect 333 927 341 961
rect 289 911 341 927
rect 583 1029 635 1041
rect 583 995 591 1029
rect 625 995 635 1029
rect 583 961 635 995
rect 583 927 591 961
rect 625 927 635 961
rect 583 911 635 927
rect 665 911 719 1041
rect 749 1029 801 1041
rect 749 995 759 1029
rect 793 995 801 1029
rect 749 961 801 995
rect 749 927 759 961
rect 793 927 801 961
rect 749 911 801 927
rect 855 1029 907 1041
rect 855 995 863 1029
rect 897 995 907 1029
rect 855 961 907 995
rect 855 927 863 961
rect 897 927 907 961
rect 855 911 907 927
rect 937 911 991 1041
rect 1021 1029 1073 1041
rect 1021 995 1031 1029
rect 1065 995 1073 1029
rect 1021 961 1073 995
rect 1021 927 1031 961
rect 1065 927 1073 961
rect 1021 911 1073 927
rect 1131 1029 1183 1041
rect 1131 995 1139 1029
rect 1173 995 1183 1029
rect 1131 961 1183 995
rect 1131 927 1139 961
rect 1173 927 1183 961
rect 1131 911 1183 927
rect 1213 911 1267 1041
rect 1297 1029 1349 1041
rect 1297 995 1307 1029
rect 1341 995 1349 1029
rect 1297 961 1349 995
rect 1297 927 1307 961
rect 1341 927 1349 961
rect 1297 911 1349 927
rect 29 165 81 177
rect 29 131 37 165
rect 71 131 81 165
rect 29 93 81 131
rect 29 59 37 93
rect 71 59 81 93
rect 29 47 81 59
rect 111 165 165 177
rect 111 131 121 165
rect 155 131 165 165
rect 111 93 165 131
rect 111 59 121 93
rect 155 59 165 93
rect 111 47 165 59
rect 195 165 247 177
rect 195 131 205 165
rect 239 131 247 165
rect 195 93 247 131
rect 195 59 205 93
rect 239 59 247 93
rect 195 47 247 59
rect 307 163 359 177
rect 307 129 315 163
rect 349 129 359 163
rect 307 95 359 129
rect 307 61 315 95
rect 349 61 359 95
rect 307 47 359 61
rect 389 163 443 177
rect 389 129 399 163
rect 433 129 443 163
rect 389 95 443 129
rect 389 61 399 95
rect 433 61 443 95
rect 389 47 443 61
rect 473 163 525 177
rect 473 129 483 163
rect 517 129 525 163
rect 473 95 525 129
rect 473 61 483 95
rect 517 61 525 95
rect 473 47 525 61
rect 579 163 631 177
rect 579 129 587 163
rect 621 129 631 163
rect 579 95 631 129
rect 579 61 587 95
rect 621 61 631 95
rect 579 47 631 61
rect 661 163 715 177
rect 661 129 671 163
rect 705 129 715 163
rect 661 95 715 129
rect 661 61 671 95
rect 705 61 715 95
rect 661 47 715 61
rect 745 163 797 177
rect 745 129 755 163
rect 789 129 797 163
rect 745 95 797 129
rect 745 61 755 95
rect 789 61 797 95
rect 745 47 797 61
rect 855 168 919 177
rect 855 134 869 168
rect 903 134 919 168
rect 855 100 919 134
rect 855 66 869 100
rect 903 66 919 100
rect 855 47 919 66
rect 949 97 1103 177
rect 949 63 959 97
rect 993 63 1059 97
rect 1093 63 1103 97
rect 949 47 1103 63
rect 1133 47 1187 177
rect 1217 95 1271 177
rect 1217 61 1227 95
rect 1261 61 1271 95
rect 1217 47 1271 61
rect 1301 117 1355 177
rect 1301 83 1311 117
rect 1345 83 1355 117
rect 1301 47 1355 83
rect 1385 95 1437 177
rect 1385 61 1395 95
rect 1429 61 1437 95
rect 1385 47 1437 61
<< pdiff >>
rect 123 773 175 791
rect 123 739 131 773
rect 165 739 175 773
rect 123 705 175 739
rect 123 671 131 705
rect 165 671 175 705
rect 123 637 175 671
rect 123 603 131 637
rect 165 603 175 637
rect 123 591 175 603
rect 205 773 259 791
rect 205 739 215 773
rect 249 739 259 773
rect 205 705 259 739
rect 205 671 215 705
rect 249 671 259 705
rect 205 637 259 671
rect 205 603 215 637
rect 249 603 259 637
rect 205 591 259 603
rect 289 773 341 791
rect 289 739 299 773
rect 333 739 341 773
rect 289 705 341 739
rect 289 671 299 705
rect 333 671 341 705
rect 289 637 341 671
rect 289 603 299 637
rect 333 603 341 637
rect 289 591 341 603
rect 583 773 635 791
rect 583 739 591 773
rect 625 739 635 773
rect 583 705 635 739
rect 583 671 591 705
rect 625 671 635 705
rect 583 637 635 671
rect 583 603 591 637
rect 625 603 635 637
rect 583 591 635 603
rect 665 773 719 791
rect 665 739 675 773
rect 709 739 719 773
rect 665 705 719 739
rect 665 671 675 705
rect 709 671 719 705
rect 665 637 719 671
rect 665 603 675 637
rect 709 603 719 637
rect 665 591 719 603
rect 749 773 801 791
rect 749 739 759 773
rect 793 739 801 773
rect 749 705 801 739
rect 749 671 759 705
rect 793 671 801 705
rect 749 637 801 671
rect 749 603 759 637
rect 793 603 801 637
rect 749 591 801 603
rect 855 773 907 791
rect 855 739 863 773
rect 897 739 907 773
rect 855 705 907 739
rect 855 671 863 705
rect 897 671 907 705
rect 855 637 907 671
rect 855 603 863 637
rect 897 603 907 637
rect 855 591 907 603
rect 937 773 991 791
rect 937 739 947 773
rect 981 739 991 773
rect 937 705 991 739
rect 937 671 947 705
rect 981 671 991 705
rect 937 637 991 671
rect 937 603 947 637
rect 981 603 991 637
rect 937 591 991 603
rect 1021 773 1073 791
rect 1021 739 1031 773
rect 1065 739 1073 773
rect 1021 705 1073 739
rect 1021 671 1031 705
rect 1065 671 1073 705
rect 1021 637 1073 671
rect 1021 603 1031 637
rect 1065 603 1073 637
rect 1021 591 1073 603
rect 1131 773 1183 791
rect 1131 739 1139 773
rect 1173 739 1183 773
rect 1131 705 1183 739
rect 1131 671 1139 705
rect 1173 671 1183 705
rect 1131 637 1183 671
rect 1131 603 1139 637
rect 1173 603 1183 637
rect 1131 591 1183 603
rect 1213 773 1267 791
rect 1213 739 1223 773
rect 1257 739 1267 773
rect 1213 705 1267 739
rect 1213 671 1223 705
rect 1257 671 1267 705
rect 1213 637 1267 671
rect 1213 603 1223 637
rect 1257 603 1267 637
rect 1213 591 1267 603
rect 1297 773 1349 791
rect 1297 739 1307 773
rect 1341 739 1349 773
rect 1297 705 1349 739
rect 1297 671 1307 705
rect 1341 671 1349 705
rect 1297 637 1349 671
rect 1297 603 1307 637
rect 1341 603 1349 637
rect 1297 591 1349 603
rect 29 485 81 497
rect 29 451 37 485
rect 71 451 81 485
rect 29 417 81 451
rect 29 383 37 417
rect 71 383 81 417
rect 29 349 81 383
rect 29 315 37 349
rect 71 315 81 349
rect 29 297 81 315
rect 111 485 165 497
rect 111 451 121 485
rect 155 451 165 485
rect 111 417 165 451
rect 111 383 121 417
rect 155 383 165 417
rect 111 349 165 383
rect 111 315 121 349
rect 155 315 165 349
rect 111 297 165 315
rect 195 485 247 497
rect 195 451 205 485
rect 239 451 247 485
rect 195 417 247 451
rect 195 383 205 417
rect 239 383 247 417
rect 195 349 247 383
rect 195 315 205 349
rect 239 315 247 349
rect 195 297 247 315
rect 319 485 371 497
rect 319 451 327 485
rect 361 451 371 485
rect 319 417 371 451
rect 319 383 327 417
rect 361 383 371 417
rect 319 349 371 383
rect 319 315 327 349
rect 361 315 371 349
rect 319 297 371 315
rect 401 297 443 497
rect 473 485 525 497
rect 473 451 483 485
rect 517 451 525 485
rect 473 417 525 451
rect 473 383 483 417
rect 517 383 525 417
rect 473 349 525 383
rect 473 315 483 349
rect 517 315 525 349
rect 473 297 525 315
rect 579 485 631 497
rect 579 451 587 485
rect 621 451 631 485
rect 579 417 631 451
rect 579 383 587 417
rect 621 383 631 417
rect 579 349 631 383
rect 579 315 587 349
rect 621 315 631 349
rect 579 297 631 315
rect 661 297 703 497
rect 733 485 785 497
rect 733 451 743 485
rect 777 451 785 485
rect 733 417 785 451
rect 733 383 743 417
rect 777 383 785 417
rect 733 349 785 383
rect 733 315 743 349
rect 777 315 785 349
rect 733 297 785 315
rect 855 477 915 497
rect 855 443 871 477
rect 905 443 915 477
rect 855 409 915 443
rect 855 375 871 409
rect 905 375 915 409
rect 855 341 915 375
rect 855 307 871 341
rect 905 307 915 341
rect 855 297 915 307
rect 945 475 997 497
rect 945 441 955 475
rect 989 441 997 475
rect 945 407 997 441
rect 945 373 955 407
rect 989 373 997 407
rect 945 297 997 373
rect 1051 475 1103 497
rect 1051 441 1059 475
rect 1093 441 1103 475
rect 1051 297 1103 441
rect 1133 475 1187 497
rect 1133 441 1143 475
rect 1177 441 1187 475
rect 1133 407 1187 441
rect 1133 373 1143 407
rect 1177 373 1187 407
rect 1133 297 1187 373
rect 1217 475 1271 497
rect 1217 441 1227 475
rect 1261 441 1271 475
rect 1217 407 1271 441
rect 1217 373 1227 407
rect 1261 373 1271 407
rect 1217 297 1271 373
rect 1301 297 1355 497
rect 1385 485 1437 497
rect 1385 451 1395 485
rect 1429 451 1437 485
rect 1385 417 1437 451
rect 1385 383 1395 417
rect 1429 383 1437 417
rect 1385 297 1437 383
<< ndiffc >>
rect 131 995 165 1029
rect 131 927 165 961
rect 299 995 333 1029
rect 299 927 333 961
rect 591 995 625 1029
rect 591 927 625 961
rect 759 995 793 1029
rect 759 927 793 961
rect 863 995 897 1029
rect 863 927 897 961
rect 1031 995 1065 1029
rect 1031 927 1065 961
rect 1139 995 1173 1029
rect 1139 927 1173 961
rect 1307 995 1341 1029
rect 1307 927 1341 961
rect 37 131 71 165
rect 37 59 71 93
rect 121 131 155 165
rect 121 59 155 93
rect 205 131 239 165
rect 205 59 239 93
rect 315 129 349 163
rect 315 61 349 95
rect 399 129 433 163
rect 399 61 433 95
rect 483 129 517 163
rect 483 61 517 95
rect 587 129 621 163
rect 587 61 621 95
rect 671 129 705 163
rect 671 61 705 95
rect 755 129 789 163
rect 755 61 789 95
rect 869 134 903 168
rect 869 66 903 100
rect 959 63 993 97
rect 1059 63 1093 97
rect 1227 61 1261 95
rect 1311 83 1345 117
rect 1395 61 1429 95
<< pdiffc >>
rect 131 739 165 773
rect 131 671 165 705
rect 131 603 165 637
rect 215 739 249 773
rect 215 671 249 705
rect 215 603 249 637
rect 299 739 333 773
rect 299 671 333 705
rect 299 603 333 637
rect 591 739 625 773
rect 591 671 625 705
rect 591 603 625 637
rect 675 739 709 773
rect 675 671 709 705
rect 675 603 709 637
rect 759 739 793 773
rect 759 671 793 705
rect 759 603 793 637
rect 863 739 897 773
rect 863 671 897 705
rect 863 603 897 637
rect 947 739 981 773
rect 947 671 981 705
rect 947 603 981 637
rect 1031 739 1065 773
rect 1031 671 1065 705
rect 1031 603 1065 637
rect 1139 739 1173 773
rect 1139 671 1173 705
rect 1139 603 1173 637
rect 1223 739 1257 773
rect 1223 671 1257 705
rect 1223 603 1257 637
rect 1307 739 1341 773
rect 1307 671 1341 705
rect 1307 603 1341 637
rect 37 451 71 485
rect 37 383 71 417
rect 37 315 71 349
rect 121 451 155 485
rect 121 383 155 417
rect 121 315 155 349
rect 205 451 239 485
rect 205 383 239 417
rect 205 315 239 349
rect 327 451 361 485
rect 327 383 361 417
rect 327 315 361 349
rect 483 451 517 485
rect 483 383 517 417
rect 483 315 517 349
rect 587 451 621 485
rect 587 383 621 417
rect 587 315 621 349
rect 743 451 777 485
rect 743 383 777 417
rect 743 315 777 349
rect 871 443 905 477
rect 871 375 905 409
rect 871 307 905 341
rect 955 441 989 475
rect 955 373 989 407
rect 1059 441 1093 475
rect 1143 441 1177 475
rect 1143 373 1177 407
rect 1227 441 1261 475
rect 1227 373 1261 407
rect 1395 451 1429 485
rect 1395 383 1429 417
<< poly >>
rect 175 1041 205 1067
rect 259 1041 289 1067
rect 635 1041 665 1067
rect 719 1041 749 1067
rect 907 1041 937 1067
rect 991 1041 1021 1067
rect 1183 1041 1213 1067
rect 1267 1041 1297 1067
rect 175 889 205 911
rect 113 873 205 889
rect 113 839 128 873
rect 162 839 205 873
rect 113 823 205 839
rect 175 791 205 823
rect 259 889 289 911
rect 635 889 665 911
rect 259 873 347 889
rect 259 839 296 873
rect 330 839 347 873
rect 259 823 347 839
rect 573 873 665 889
rect 573 839 588 873
rect 622 839 665 873
rect 573 823 665 839
rect 259 791 289 823
rect 635 791 665 823
rect 719 889 749 911
rect 907 889 937 911
rect 719 873 807 889
rect 719 839 756 873
rect 790 839 807 873
rect 719 823 807 839
rect 849 873 937 889
rect 849 839 866 873
rect 900 839 937 873
rect 849 823 937 839
rect 719 791 749 823
rect 907 791 937 823
rect 991 889 1021 911
rect 1183 889 1213 911
rect 991 873 1083 889
rect 991 839 1034 873
rect 1068 839 1083 873
rect 991 823 1083 839
rect 1125 873 1213 889
rect 1125 839 1142 873
rect 1176 839 1213 873
rect 1125 823 1213 839
rect 991 791 1021 823
rect 1183 791 1213 823
rect 1267 889 1297 911
rect 1267 873 1359 889
rect 1267 839 1310 873
rect 1344 839 1359 873
rect 1267 823 1359 839
rect 1267 791 1297 823
rect 175 565 205 591
rect 259 565 289 591
rect 635 565 665 591
rect 719 565 749 591
rect 907 565 937 591
rect 991 565 1021 591
rect 1183 565 1213 591
rect 1267 565 1297 591
rect 81 497 111 523
rect 165 497 195 523
rect 371 497 401 523
rect 443 497 473 523
rect 631 497 661 523
rect 703 497 733 523
rect 915 497 945 523
rect 1103 497 1133 523
rect 1187 497 1217 523
rect 1271 497 1301 523
rect 1355 497 1385 523
rect 81 265 111 297
rect 165 265 195 297
rect 371 265 401 297
rect 81 249 255 265
rect 81 215 205 249
rect 239 215 255 249
rect 81 199 255 215
rect 297 249 401 265
rect 297 215 313 249
rect 347 235 401 249
rect 443 265 473 297
rect 631 265 661 297
rect 443 249 530 265
rect 347 215 389 235
rect 297 199 389 215
rect 81 177 111 199
rect 165 177 195 199
rect 359 177 389 199
rect 443 215 481 249
rect 515 215 530 249
rect 443 199 530 215
rect 574 249 661 265
rect 574 215 589 249
rect 623 215 661 249
rect 703 265 733 297
rect 915 265 945 297
rect 1103 265 1133 297
rect 1187 265 1217 297
rect 1271 265 1301 297
rect 1355 265 1385 297
rect 703 249 807 265
rect 703 235 757 249
rect 574 199 661 215
rect 443 177 473 199
rect 631 177 661 199
rect 715 215 757 235
rect 791 215 807 249
rect 915 249 1049 265
rect 915 232 1005 249
rect 715 199 807 215
rect 919 215 1005 232
rect 1039 215 1049 249
rect 919 199 1049 215
rect 1091 249 1145 265
rect 1091 215 1101 249
rect 1135 215 1145 249
rect 1091 199 1145 215
rect 1187 249 1301 265
rect 1187 215 1236 249
rect 1270 215 1301 249
rect 1187 199 1301 215
rect 1343 249 1397 265
rect 1343 215 1353 249
rect 1387 215 1397 249
rect 1343 199 1397 215
rect 715 177 745 199
rect 919 177 949 199
rect 1103 177 1133 199
rect 1187 177 1217 199
rect 1271 177 1301 199
rect 1355 177 1385 199
rect 81 21 111 47
rect 165 21 195 47
rect 359 21 389 47
rect 443 21 473 47
rect 631 21 661 47
rect 715 21 745 47
rect 919 21 949 47
rect 1103 21 1133 47
rect 1187 21 1217 47
rect 1271 21 1301 47
rect 1355 21 1385 47
<< polycont >>
rect 128 839 162 873
rect 296 839 330 873
rect 588 839 622 873
rect 756 839 790 873
rect 866 839 900 873
rect 1034 839 1068 873
rect 1142 839 1176 873
rect 1310 839 1344 873
rect 205 215 239 249
rect 313 215 347 249
rect 481 215 515 249
rect 589 215 623 249
rect 757 215 791 249
rect 1005 215 1039 249
rect 1101 215 1135 249
rect 1236 215 1270 249
rect 1353 215 1387 249
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1472 1105
rect 109 1029 171 1071
rect 109 995 131 1029
rect 165 995 171 1029
rect 109 961 171 995
rect 109 927 131 961
rect 165 927 171 961
rect 109 911 171 927
rect 212 1029 351 1037
rect 212 995 299 1029
rect 333 995 351 1029
rect 569 1029 631 1071
rect 212 961 351 995
rect 212 927 299 961
rect 333 927 351 961
rect 212 911 351 927
rect 111 873 178 877
rect 111 867 128 873
rect 51 839 128 867
rect 162 839 178 873
rect 51 833 178 839
rect 111 823 178 833
rect 212 791 246 911
rect 280 839 296 873
rect 330 867 347 873
rect 425 867 459 969
rect 569 995 591 1029
rect 625 995 631 1029
rect 569 961 631 995
rect 569 927 591 961
rect 625 927 631 961
rect 569 911 631 927
rect 672 1029 811 1037
rect 672 995 759 1029
rect 793 995 811 1029
rect 672 961 811 995
rect 672 927 759 961
rect 793 927 811 961
rect 672 911 811 927
rect 845 1029 984 1037
rect 845 995 863 1029
rect 897 1003 984 1029
rect 897 995 901 1003
rect 845 969 901 995
rect 935 969 984 1003
rect 845 961 984 969
rect 845 927 863 961
rect 897 927 984 961
rect 845 911 984 927
rect 1025 1029 1087 1071
rect 1025 995 1031 1029
rect 1065 995 1087 1029
rect 1025 961 1087 995
rect 1025 927 1031 961
rect 1065 927 1087 961
rect 1025 911 1087 927
rect 1121 1029 1260 1037
rect 1121 995 1139 1029
rect 1173 1003 1260 1029
rect 1121 969 1173 995
rect 1207 969 1260 1003
rect 1121 961 1260 969
rect 1121 927 1139 961
rect 1173 927 1260 961
rect 1121 911 1260 927
rect 1301 1029 1363 1071
rect 1301 995 1307 1029
rect 1341 995 1363 1029
rect 1301 961 1363 995
rect 1301 927 1307 961
rect 1341 927 1363 961
rect 1301 911 1363 927
rect 571 873 638 877
rect 571 867 588 873
rect 330 839 459 867
rect 280 833 459 839
rect 527 839 588 867
rect 622 839 638 873
rect 527 833 638 839
rect 280 823 347 833
rect 571 823 638 833
rect 672 791 706 911
rect 740 839 756 873
rect 790 867 807 873
rect 849 867 866 873
rect 797 839 866 867
rect 900 839 916 873
rect 740 833 763 839
rect 797 833 916 839
rect 740 823 807 833
rect 849 823 916 833
rect 950 791 984 911
rect 1018 873 1085 877
rect 1018 839 1034 873
rect 1068 867 1085 873
rect 1018 833 1037 839
rect 1071 833 1085 867
rect 1018 823 1085 833
rect 1125 867 1142 873
rect 1125 833 1139 867
rect 1176 839 1192 873
rect 1173 833 1192 839
rect 1125 823 1192 833
rect 1226 791 1260 911
rect 1294 873 1361 877
rect 1294 867 1310 873
rect 1294 833 1309 867
rect 1344 839 1361 873
rect 1343 833 1361 839
rect 1294 823 1361 833
rect 109 773 165 789
rect 109 739 131 773
rect 109 705 165 739
rect 109 671 131 705
rect 109 637 165 671
rect 109 603 131 637
rect 109 561 165 603
rect 199 773 265 791
rect 199 739 215 773
rect 249 739 265 773
rect 199 705 265 739
rect 199 671 215 705
rect 249 671 265 705
rect 199 663 265 671
rect 199 637 221 663
rect 199 603 215 637
rect 255 629 265 663
rect 249 603 265 629
rect 199 595 265 603
rect 299 773 351 789
rect 333 739 351 773
rect 299 705 351 739
rect 333 671 351 705
rect 299 637 351 671
rect 333 603 351 637
rect 299 561 351 603
rect 569 773 625 789
rect 569 739 591 773
rect 569 705 625 739
rect 569 671 591 705
rect 569 637 625 671
rect 569 603 591 637
rect 569 561 625 603
rect 659 773 725 791
rect 659 739 675 773
rect 709 739 725 773
rect 659 705 725 739
rect 659 671 675 705
rect 709 671 725 705
rect 659 663 725 671
rect 659 629 673 663
rect 707 637 725 663
rect 659 603 675 629
rect 709 603 725 637
rect 659 595 725 603
rect 759 773 811 789
rect 793 739 811 773
rect 759 705 811 739
rect 793 671 811 705
rect 759 637 811 671
rect 793 603 811 637
rect 759 561 811 603
rect 845 773 897 789
rect 845 739 863 773
rect 845 705 897 739
rect 845 671 863 705
rect 845 637 897 671
rect 845 603 863 637
rect 845 561 897 603
rect 931 773 997 791
rect 931 739 947 773
rect 981 739 997 773
rect 931 705 997 739
rect 931 671 947 705
rect 981 671 997 705
rect 931 637 997 671
rect 931 603 947 637
rect 981 603 997 637
rect 931 595 997 603
rect 1031 773 1087 789
rect 1065 739 1087 773
rect 1031 705 1087 739
rect 1065 671 1087 705
rect 1031 637 1087 671
rect 1065 603 1087 637
rect 1031 561 1087 603
rect 1121 773 1173 789
rect 1121 739 1139 773
rect 1121 705 1173 739
rect 1121 671 1139 705
rect 1121 637 1173 671
rect 1121 603 1139 637
rect 1121 561 1173 603
rect 1207 773 1273 791
rect 1207 739 1223 773
rect 1257 739 1273 773
rect 1207 705 1273 739
rect 1207 671 1223 705
rect 1257 671 1273 705
rect 1207 637 1273 671
rect 1207 603 1223 637
rect 1257 603 1273 637
rect 1207 595 1273 603
rect 1307 773 1363 789
rect 1341 739 1363 773
rect 1307 705 1363 739
rect 1341 671 1363 705
rect 1307 637 1363 671
rect 1341 603 1363 637
rect 1307 561 1363 603
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 29 485 71 527
rect 29 451 37 485
rect 29 417 71 451
rect 29 383 37 417
rect 29 349 71 383
rect 29 315 37 349
rect 29 299 71 315
rect 105 485 171 493
rect 105 451 121 485
rect 155 451 171 485
rect 105 417 171 451
rect 105 391 121 417
rect 105 357 119 391
rect 155 383 171 417
rect 153 357 171 383
rect 105 349 171 357
rect 105 315 121 349
rect 155 315 171 349
rect 105 297 171 315
rect 205 485 251 527
rect 239 451 251 485
rect 205 417 251 451
rect 239 383 251 417
rect 205 349 251 383
rect 239 315 251 349
rect 205 299 251 315
rect 295 485 361 527
rect 295 451 327 485
rect 295 417 361 451
rect 295 383 327 417
rect 295 349 361 383
rect 295 315 327 349
rect 467 485 533 490
rect 467 451 483 485
rect 517 459 533 485
rect 467 425 493 451
rect 527 425 533 459
rect 467 417 533 425
rect 467 383 483 417
rect 517 383 533 417
rect 467 349 533 383
rect 467 333 483 349
rect 295 299 361 315
rect 397 315 483 333
rect 517 315 533 349
rect 397 299 533 315
rect 571 485 637 490
rect 571 451 587 485
rect 621 451 637 485
rect 571 417 637 451
rect 571 383 587 417
rect 621 383 637 417
rect 571 349 637 383
rect 571 315 587 349
rect 621 333 637 349
rect 743 485 809 527
rect 777 451 809 485
rect 743 417 809 451
rect 777 383 809 417
rect 743 349 809 383
rect 621 315 707 333
rect 571 299 707 315
rect 777 315 809 349
rect 743 299 809 315
rect 845 477 909 493
rect 845 443 871 477
rect 905 443 909 477
rect 845 409 909 443
rect 845 375 871 409
rect 905 375 909 409
rect 845 341 909 375
rect 945 475 1025 493
rect 945 441 955 475
rect 989 441 1025 475
rect 945 407 1025 441
rect 1059 475 1093 527
rect 1059 425 1093 441
rect 1127 475 1193 493
rect 1127 441 1143 475
rect 1177 441 1193 475
rect 945 373 955 407
rect 989 391 1025 407
rect 1127 407 1193 441
rect 1127 391 1143 407
rect 989 373 1143 391
rect 1177 373 1193 407
rect 945 357 1193 373
rect 1227 475 1261 527
rect 1379 485 1455 493
rect 1227 407 1261 441
rect 1227 357 1261 373
rect 845 307 871 341
rect 905 323 909 341
rect 1309 323 1343 425
rect 1379 451 1395 485
rect 1429 451 1455 485
rect 1379 417 1455 451
rect 1379 383 1395 417
rect 1429 383 1455 417
rect 1379 357 1455 383
rect 29 165 71 181
rect 29 131 37 165
rect 29 93 71 131
rect 29 59 37 93
rect 29 17 71 59
rect 105 177 155 297
rect 189 255 255 265
rect 293 255 363 265
rect 189 249 221 255
rect 255 249 363 255
rect 189 215 205 249
rect 255 221 313 249
rect 239 215 255 221
rect 293 215 313 221
rect 347 215 363 249
rect 105 165 171 177
rect 105 131 121 165
rect 155 131 171 165
rect 105 93 171 131
rect 105 59 121 93
rect 155 59 171 93
rect 105 51 171 59
rect 205 165 251 181
rect 397 179 431 299
rect 465 256 535 265
rect 465 249 493 256
rect 465 215 481 249
rect 527 222 535 256
rect 515 215 535 222
rect 569 256 639 265
rect 569 249 595 256
rect 569 215 589 249
rect 629 222 639 256
rect 623 215 639 222
rect 673 179 707 299
rect 845 289 901 307
rect 935 289 971 307
rect 845 273 971 289
rect 741 255 811 265
rect 741 249 765 255
rect 741 215 757 249
rect 799 221 811 255
rect 791 215 811 221
rect 239 131 251 165
rect 205 93 251 131
rect 239 59 251 93
rect 205 17 251 59
rect 295 163 349 179
rect 295 129 315 163
rect 295 95 349 129
rect 295 61 315 95
rect 295 17 349 61
rect 383 163 449 179
rect 383 129 399 163
rect 433 129 449 163
rect 383 95 449 129
rect 383 61 399 95
rect 433 61 449 95
rect 383 51 449 61
rect 483 163 531 179
rect 517 129 531 163
rect 483 95 531 129
rect 517 61 531 95
rect 483 17 531 61
rect 573 163 621 179
rect 573 129 587 163
rect 573 95 621 129
rect 573 61 587 95
rect 573 17 621 61
rect 655 163 721 179
rect 655 153 671 163
rect 655 119 669 153
rect 705 129 721 163
rect 703 119 721 129
rect 655 95 721 119
rect 655 61 671 95
rect 705 61 721 95
rect 655 51 721 61
rect 755 163 809 179
rect 789 129 809 163
rect 755 95 809 129
rect 789 61 809 95
rect 755 17 809 61
rect 845 168 903 184
rect 845 134 869 168
rect 845 100 903 134
rect 845 66 869 100
rect 845 17 903 66
rect 937 97 971 273
rect 1126 289 1387 323
rect 1005 249 1051 265
rect 1126 249 1160 289
rect 1039 215 1051 249
rect 1085 215 1101 249
rect 1135 215 1160 249
rect 1194 249 1241 255
rect 1194 215 1236 249
rect 1275 221 1304 255
rect 1270 215 1304 221
rect 1338 249 1387 289
rect 1338 215 1353 249
rect 1005 165 1051 215
rect 1338 199 1387 215
rect 1421 165 1455 357
rect 1005 131 1455 165
rect 1311 117 1345 131
rect 937 63 959 97
rect 993 63 1059 97
rect 1093 63 1128 97
rect 1211 61 1227 95
rect 1261 61 1277 95
rect 1311 67 1345 83
rect 1211 17 1277 61
rect 1379 61 1395 95
rect 1429 61 1445 95
rect 1379 17 1445 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 425 969 459 1003
rect 17 833 51 867
rect 901 969 935 1003
rect 1173 969 1207 1003
rect 493 833 527 867
rect 763 839 790 867
rect 790 839 797 867
rect 763 833 797 839
rect 1037 839 1068 867
rect 1068 839 1071 867
rect 1037 833 1071 839
rect 1139 839 1142 867
rect 1142 839 1173 867
rect 1139 833 1173 839
rect 1309 839 1310 867
rect 1310 839 1343 867
rect 1309 833 1343 839
rect 221 637 255 663
rect 221 629 249 637
rect 249 629 255 637
rect 673 637 707 663
rect 673 629 675 637
rect 675 629 707 637
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 119 383 121 391
rect 121 383 153 391
rect 119 357 153 383
rect 493 451 517 459
rect 517 451 527 459
rect 493 425 527 451
rect 1309 425 1343 459
rect 901 307 905 323
rect 905 307 935 323
rect 221 249 255 255
rect 221 221 239 249
rect 239 221 255 249
rect 493 249 527 256
rect 493 222 515 249
rect 515 222 527 249
rect 595 249 629 256
rect 595 222 623 249
rect 623 222 629 249
rect 901 289 935 307
rect 765 249 799 255
rect 765 221 791 249
rect 791 221 799 249
rect 669 129 671 153
rect 671 129 703 153
rect 669 119 703 129
rect 1241 249 1275 255
rect 1241 221 1270 249
rect 1270 221 1275 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 1105 1472 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1472 1105
rect 0 1065 1472 1071
rect 413 1003 471 1009
rect 413 969 425 1003
rect 459 1000 471 1003
rect 614 1000 620 1006
rect 459 972 620 1000
rect 459 969 471 972
rect 413 963 471 969
rect 613 966 620 972
rect 614 954 620 966
rect 672 1000 678 1006
rect 672 972 796 1000
rect 672 966 679 972
rect 672 954 678 966
rect 768 929 796 972
rect 886 957 892 1009
rect 944 1000 950 1009
rect 1161 1003 1232 1009
rect 944 972 1005 1000
rect 944 957 950 972
rect 1161 969 1173 1003
rect 1207 969 1232 1003
rect 1161 960 1232 969
rect 1226 957 1232 960
rect 1284 957 1290 1009
rect 1226 954 1290 957
rect 768 901 1170 929
rect 5 867 63 873
rect 5 833 17 867
rect 51 864 63 867
rect 478 864 484 876
rect 51 836 484 864
rect 51 833 63 836
rect 5 827 63 833
rect 478 824 484 836
rect 536 824 542 876
rect 1142 873 1170 901
rect 751 867 822 873
rect 751 833 763 867
rect 797 833 822 867
rect 751 824 822 833
rect 816 821 822 824
rect 874 821 880 873
rect 1022 821 1028 873
rect 1080 821 1086 873
rect 1127 867 1185 873
rect 1127 833 1139 867
rect 1173 833 1185 867
rect 1127 827 1185 833
rect 1297 867 1355 873
rect 1297 833 1309 867
rect 1343 833 1355 867
rect 1297 827 1355 833
rect 1040 793 1068 821
rect 1312 793 1340 827
rect 1040 765 1340 793
rect 206 660 212 672
rect 151 632 212 660
rect 206 620 212 632
rect 264 620 270 672
rect 661 663 719 669
rect 661 629 673 663
rect 707 660 719 663
rect 1090 660 1096 672
rect 707 632 1096 660
rect 707 629 719 632
rect 661 623 719 629
rect 1090 620 1096 632
rect 1148 620 1154 672
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 481 459 539 465
rect 481 425 493 459
rect 527 456 539 459
rect 954 456 960 468
rect 527 428 960 456
rect 527 425 539 428
rect 481 419 539 425
rect 954 416 960 428
rect 1012 416 1018 468
rect 1090 416 1096 468
rect 1148 456 1154 468
rect 1297 459 1355 465
rect 1297 456 1309 459
rect 1148 428 1309 456
rect 1148 416 1154 428
rect 1297 425 1309 428
rect 1343 425 1355 459
rect 1297 419 1355 425
rect 107 391 165 397
rect 107 357 119 391
rect 153 388 165 391
rect 682 388 688 400
rect 153 360 688 388
rect 153 357 165 360
rect 107 351 165 357
rect 206 252 212 264
rect 151 224 212 252
rect 206 212 212 224
rect 264 212 270 264
rect 598 262 626 360
rect 682 348 688 360
rect 740 348 746 400
rect 886 320 892 332
rect 831 292 892 320
rect 886 280 892 292
rect 944 280 950 332
rect 481 256 539 262
rect 481 253 493 256
rect 360 225 493 253
rect 360 196 388 225
rect 481 222 493 225
rect 527 222 539 256
rect 481 216 539 222
rect 583 256 641 262
rect 583 222 595 256
rect 629 222 641 256
rect 750 252 756 264
rect 695 224 756 252
rect 583 216 641 222
rect 750 212 756 224
rect 808 212 814 264
rect 1226 252 1232 264
rect 1171 224 1232 252
rect 1226 212 1232 224
rect 1284 212 1290 264
rect 342 144 348 196
rect 400 144 406 196
rect 614 150 620 162
rect 672 159 678 162
rect 672 153 715 159
rect 596 122 620 150
rect 614 110 620 122
rect 703 119 715 153
rect 672 113 715 119
rect 672 110 678 113
rect 0 17 1472 23
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< via1 >>
rect 620 954 672 1006
rect 892 1003 944 1009
rect 892 969 901 1003
rect 901 969 935 1003
rect 935 969 944 1003
rect 892 957 944 969
rect 1232 957 1284 1009
rect 484 867 536 876
rect 484 833 493 867
rect 493 833 527 867
rect 527 833 536 867
rect 484 824 536 833
rect 822 821 874 873
rect 1028 867 1080 873
rect 1028 833 1037 867
rect 1037 833 1071 867
rect 1071 833 1080 867
rect 1028 821 1080 833
rect 212 663 264 672
rect 212 629 221 663
rect 221 629 255 663
rect 255 629 264 663
rect 212 620 264 629
rect 1096 620 1148 672
rect 960 416 1012 468
rect 1096 416 1148 468
rect 212 255 264 264
rect 212 221 221 255
rect 221 221 255 255
rect 255 221 264 255
rect 212 212 264 221
rect 688 348 740 400
rect 892 323 944 332
rect 892 289 901 323
rect 901 289 935 323
rect 935 289 944 323
rect 892 280 944 289
rect 756 255 808 264
rect 756 221 765 255
rect 765 221 799 255
rect 799 221 808 255
rect 756 212 808 221
rect 1232 255 1284 264
rect 1232 221 1241 255
rect 1241 221 1275 255
rect 1275 221 1284 255
rect 1232 212 1284 221
rect 348 144 400 196
rect 620 153 672 162
rect 620 119 669 153
rect 669 119 672 153
rect 620 110 672 119
<< metal2 >>
rect 618 1009 674 1018
rect 892 1009 944 1018
rect 1232 1009 1284 1018
rect 886 960 892 1009
rect 618 944 674 953
rect 944 960 950 1009
rect 892 951 944 957
rect 1232 951 1284 957
rect 482 877 538 886
rect 482 812 538 821
rect 820 877 876 886
rect 820 812 876 821
rect 904 728 932 951
rect 1028 877 1084 886
rect 1028 812 1084 821
rect 768 700 932 728
rect 212 672 264 678
rect 212 614 264 620
rect 224 270 252 614
rect 768 559 796 700
rect 1096 672 1148 678
rect 1096 614 1148 620
rect 346 550 402 559
rect 346 485 402 494
rect 754 550 810 559
rect 754 485 810 494
rect 212 264 264 270
rect 212 206 264 212
rect 360 202 388 485
rect 684 402 740 411
rect 684 337 740 346
rect 768 270 796 485
rect 958 470 1014 479
rect 1108 474 1136 614
rect 958 405 1014 414
rect 1096 468 1148 474
rect 1096 410 1148 416
rect 890 334 946 343
rect 756 264 808 270
rect 890 269 946 278
rect 1244 270 1272 951
rect 756 206 808 212
rect 1232 264 1284 270
rect 1232 206 1284 212
rect 348 196 400 202
rect 348 138 400 144
rect 618 164 674 173
rect 618 99 674 108
<< via2 >>
rect 618 1006 674 1009
rect 618 954 620 1006
rect 620 954 672 1006
rect 672 954 674 1006
rect 618 953 674 954
rect 482 876 538 877
rect 482 824 484 876
rect 484 824 536 876
rect 536 824 538 876
rect 482 821 538 824
rect 820 873 876 877
rect 820 821 822 873
rect 822 821 874 873
rect 874 821 876 873
rect 1028 873 1084 877
rect 1028 821 1080 873
rect 1080 821 1084 873
rect 346 494 402 550
rect 754 494 810 550
rect 684 400 740 402
rect 684 348 688 400
rect 688 348 740 400
rect 684 346 740 348
rect 958 468 1014 470
rect 958 416 960 468
rect 960 416 1012 468
rect 1012 416 1014 468
rect 958 414 1014 416
rect 890 332 946 334
rect 890 280 892 332
rect 892 280 944 332
rect 944 280 946 332
rect 890 278 946 280
rect 618 162 674 164
rect 618 110 620 162
rect 620 110 672 162
rect 672 110 674 162
rect 618 108 674 110
<< metal3 >>
rect 519 1009 679 1017
rect 519 957 618 1009
rect 595 953 618 957
rect 674 953 679 1009
rect 595 948 679 953
rect 595 943 655 948
rect 477 879 543 882
rect 815 879 881 882
rect 383 877 543 879
rect 383 821 482 877
rect 538 821 543 877
rect 383 819 543 821
rect 721 877 881 879
rect 721 821 820 877
rect 876 821 881 877
rect 721 819 881 821
rect 477 816 543 819
rect 815 816 881 819
rect 1023 879 1089 882
rect 1023 877 1183 879
rect 1023 821 1028 877
rect 1084 821 1183 877
rect 1023 819 1183 821
rect 1023 816 1094 819
rect 820 807 880 816
rect 1034 811 1094 816
rect 341 552 407 555
rect 749 552 815 555
rect 341 550 815 552
rect 341 494 346 550
rect 402 494 754 550
rect 810 494 815 550
rect 341 492 815 494
rect 341 489 407 492
rect 749 489 815 492
rect 953 472 1019 475
rect 953 470 1113 472
rect 953 414 958 470
rect 1014 414 1113 470
rect 953 412 1113 414
rect 953 409 1019 412
rect 679 404 745 407
rect 587 402 747 404
rect 956 403 1016 409
rect 587 346 684 402
rect 740 346 747 402
rect 587 344 747 346
rect 679 341 745 344
rect 885 336 951 339
rect 885 334 1045 336
rect 885 278 890 334
rect 946 278 1045 334
rect 885 276 1045 278
rect 885 273 962 276
rect 902 271 962 273
rect 613 166 679 169
rect 519 164 679 166
rect 519 108 618 164
rect 674 108 679 164
rect 519 106 679 108
rect 611 105 679 106
rect 613 103 679 105
<< labels >>
rlabel comment s 1472 0 1472 0 4 scs130hd_xor2_1
rlabel comment s 552 0 552 0 4 scs130hd_nor2_1
rlabel comment s 552 0 552 0 4 scs130hd_nor2_1
rlabel comment s 1104 1088 1104 1088 4 scs130hd_nand2_1
rlabel comment s 1380 1088 1380 1088 4 scs130hd_nand2_1
rlabel comment s 552 1088 552 1088 4 scs130hd_nand2_1
rlabel comment s 92 1088 92 1088 4 scs130hd_nand2_1
rlabel comment s 276 0 276 0 4 scs130hd_inv_2
rlabel comment s 368 1088 368 1088 4 scs130hd_fill_2
rlabel comment s 1380 1088 1380 1088 4 scs130hd_fill_1
rlabel comment s 0 1088 0 1088 4 scs130hd_fill_1
rlabel comment s 0 1088 0 1088 4 fill_T_1_1
rlabel metal3 s 815 816 881 882 4 A1
port 7 nsew
rlabel metal3 s 477 816 543 882 4 B0
port 15 nsew
rlabel metal3 s 1023 816 1089 882 4 B1
port 16 nsew
rlabel metal3 s 679 341 745 407 4 R0
port 17 nsew
rlabel metal3 s 885 273 951 339 4 R1
port 18 nsew
rlabel metal3 s 613 103 679 169 4 R2
port 19 nsew
rlabel metal3 s 953 409 1019 475 4 R3
port 20 nsew
rlabel pwell 82 -1 82 -1 1 VNB
port 21 n
rlabel metal1 136 0 136 0 1 vgnd
port 22 n
rlabel nwell 92 542 92 542 1 VPB
port 23 n
rlabel metal1 139 545 139 545 1 vpwr
port 24 n
rlabel pwell 46 1087 46 1087 1 VNB
port 21 n
rlabel viali 138 1089 138 1089 1 vgnd
port 22 n
rlabel metal3 s 613 948 679 1014 4 A0
port 14 nsew
<< properties >>
string FIXED_BBOX 0 0 1472 1088
string path 4.915 2.210 5.415 2.210 
<< end >>
