VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mux16x1_project
  CLASS BLOCK ;
  FOREIGN mux16x1_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 440.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 12.280 700.000 12.880 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 229.880 700.000 230.480 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 251.640 700.000 252.240 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 273.400 700.000 274.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 295.160 700.000 295.760 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 316.920 700.000 317.520 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 338.680 700.000 339.280 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 360.440 700.000 361.040 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 382.200 700.000 382.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 403.960 700.000 404.560 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 425.720 700.000 426.320 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 34.040 700.000 34.640 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 55.800 700.000 56.400 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 77.560 700.000 78.160 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 99.320 700.000 99.920 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 121.080 700.000 121.680 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 142.840 700.000 143.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 164.600 700.000 165.200 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 186.360 700.000 186.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 208.120 700.000 208.720 ;
    END
  END io_in[9]
  PIN io_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END io_out
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 427.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 427.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 694.140 427.125 ;
      LAYER met1 ;
        RECT 5.520 10.640 695.450 427.280 ;
      LAYER met2 ;
        RECT 7.910 10.695 695.430 427.225 ;
      LAYER met3 ;
        RECT 3.990 426.720 696.000 427.205 ;
        RECT 3.990 425.320 695.600 426.720 ;
        RECT 3.990 404.960 696.000 425.320 ;
        RECT 3.990 403.560 695.600 404.960 ;
        RECT 3.990 383.200 696.000 403.560 ;
        RECT 3.990 381.800 695.600 383.200 ;
        RECT 3.990 361.440 696.000 381.800 ;
        RECT 3.990 360.040 695.600 361.440 ;
        RECT 3.990 339.680 696.000 360.040 ;
        RECT 3.990 338.280 695.600 339.680 ;
        RECT 3.990 317.920 696.000 338.280 ;
        RECT 3.990 316.520 695.600 317.920 ;
        RECT 3.990 296.160 696.000 316.520 ;
        RECT 3.990 294.760 695.600 296.160 ;
        RECT 3.990 274.400 696.000 294.760 ;
        RECT 3.990 273.000 695.600 274.400 ;
        RECT 3.990 252.640 696.000 273.000 ;
        RECT 3.990 251.240 695.600 252.640 ;
        RECT 3.990 230.880 696.000 251.240 ;
        RECT 3.990 229.480 695.600 230.880 ;
        RECT 3.990 220.000 696.000 229.480 ;
        RECT 4.400 218.600 696.000 220.000 ;
        RECT 3.990 209.120 696.000 218.600 ;
        RECT 3.990 207.720 695.600 209.120 ;
        RECT 3.990 187.360 696.000 207.720 ;
        RECT 3.990 185.960 695.600 187.360 ;
        RECT 3.990 165.600 696.000 185.960 ;
        RECT 3.990 164.200 695.600 165.600 ;
        RECT 3.990 143.840 696.000 164.200 ;
        RECT 3.990 142.440 695.600 143.840 ;
        RECT 3.990 122.080 696.000 142.440 ;
        RECT 3.990 120.680 695.600 122.080 ;
        RECT 3.990 100.320 696.000 120.680 ;
        RECT 3.990 98.920 695.600 100.320 ;
        RECT 3.990 78.560 696.000 98.920 ;
        RECT 3.990 77.160 695.600 78.560 ;
        RECT 3.990 56.800 696.000 77.160 ;
        RECT 3.990 55.400 695.600 56.800 ;
        RECT 3.990 35.040 696.000 55.400 ;
        RECT 3.990 33.640 695.600 35.040 ;
        RECT 3.990 13.280 696.000 33.640 ;
        RECT 3.990 11.880 695.600 13.280 ;
        RECT 3.990 10.715 696.000 11.880 ;
  END
END mux16x1_project
END LIBRARY

