magic
tech sky130A
magscale 1 2
timestamp 1708010873
<< error_s >>
rect 1767 2133 1768 2144
rect 1957 2133 1958 2144
rect 2043 2133 2044 2144
rect 2719 2133 2720 2144
rect 2909 2133 2910 2144
rect 2995 2133 2996 2144
rect 3268 2133 3269 2144
rect 3466 2133 3467 2144
rect 1778 2093 1779 2133
rect 1968 2093 1969 2133
rect 2054 2093 2055 2133
rect 2730 2093 2731 2133
rect 2920 2093 2921 2133
rect 3006 2093 3007 2133
rect 3279 2093 3280 2133
rect 3477 2093 3478 2133
rect 2927 1966 2954 1973
rect 2927 1945 2995 1966
rect 2927 1939 2982 1945
rect 2966 1938 2967 1939
rect 2939 1932 2994 1938
rect 2966 1910 2967 1932
rect 1767 1703 1768 1714
rect 1957 1703 1958 1714
rect 2043 1703 2044 1714
rect 2719 1703 2720 1714
rect 2909 1703 2910 1714
rect 2995 1703 2996 1714
rect 3268 1703 3269 1714
rect 3466 1703 3467 1714
rect 1716 1671 1740 1677
rect 1744 1676 1768 1677
rect 1778 1507 1779 1703
rect 1968 1507 1969 1703
rect 2054 1507 2055 1703
rect 2730 1507 2731 1703
rect 2920 1507 2921 1703
rect 3006 1507 3007 1703
rect 3279 1507 3280 1703
rect 3477 1507 3478 1703
rect 2092 1403 2116 1437
rect 3044 1403 3068 1437
rect 3044 1085 3068 1119
rect 133 1057 142 1066
rect 180 1057 189 1066
rect 1444 1057 1453 1066
rect 1789 1057 1798 1066
rect 1836 1057 1845 1066
rect 1989 1057 1998 1066
rect 2036 1057 2045 1066
rect 124 1048 133 1057
rect 189 1048 198 1057
rect 1103 1038 1109 1044
rect 1149 1038 1155 1044
rect 1411 1043 1423 1051
rect 1433 1043 1445 1051
rect 1453 1048 1462 1057
rect 1512 1051 1528 1052
rect 1407 1040 1409 1043
rect 1447 1040 1449 1043
rect 1506 1039 1517 1051
rect 1780 1048 1789 1057
rect 1845 1051 1854 1057
rect 1786 1045 1789 1047
rect 1793 1045 1799 1051
rect 1839 1048 1854 1051
rect 1980 1048 1989 1057
rect 2045 1050 2054 1057
rect 1839 1045 1845 1048
rect 1097 1032 1103 1038
rect 1155 1032 1161 1038
rect 1388 1031 1394 1037
rect 1399 1031 1407 1039
rect 1410 1037 1445 1039
rect 1410 1036 1411 1037
rect 1409 1031 1410 1035
rect 1411 1031 1412 1036
rect 1443 1031 1445 1037
rect 130 1026 133 1030
rect 116 1023 155 1026
rect 1157 1023 1196 1028
rect 1382 1025 1388 1031
rect 1408 1026 1409 1031
rect 1407 1024 1408 1026
rect 113 1022 116 1023
rect 113 1015 125 1022
rect 130 1020 133 1023
rect 129 1016 130 1019
rect 113 1013 129 1015
rect 135 1013 147 1022
rect 155 1020 184 1023
rect 184 1014 188 1020
rect 924 1018 976 1020
rect 1196 1018 1210 1023
rect 1406 1020 1407 1023
rect 896 1016 976 1018
rect 896 1015 947 1016
rect 188 1013 189 1014
rect 871 1013 896 1015
rect 918 1014 924 1015
rect 947 1014 952 1015
rect 109 1011 113 1013
rect 125 1010 129 1013
rect 837 1011 867 1013
rect 913 1012 918 1014
rect 101 998 109 1010
rect 108 988 109 998
rect 113 1007 147 1010
rect 113 1003 115 1007
rect 113 996 114 1003
rect 125 1001 129 1007
rect 144 1005 147 1007
rect 150 1004 159 1010
rect 112 994 114 996
rect 111 988 117 994
rect 122 988 125 1001
rect 105 982 111 988
rect 108 976 109 982
rect 112 962 113 988
rect 145 982 147 1004
rect 151 998 159 1004
rect 189 1001 198 1010
rect 720 1005 734 1007
rect 746 1005 837 1011
rect 909 1007 913 1012
rect 720 1004 746 1005
rect 720 1003 734 1004
rect 714 1002 734 1003
rect 755 1002 760 1005
rect 905 1002 909 1007
rect 952 1005 969 1014
rect 969 1004 971 1005
rect 157 988 163 994
rect 180 992 189 1001
rect 705 997 729 1002
rect 760 997 766 1002
rect 904 1001 905 1002
rect 976 1001 993 1016
rect 1210 1015 1217 1018
rect 1405 1016 1406 1020
rect 1217 1014 1220 1015
rect 1220 1005 1242 1014
rect 1403 1012 1405 1016
rect 1443 1014 1447 1031
rect 1449 1027 1457 1039
rect 1715 1037 1727 1045
rect 1776 1041 1786 1045
rect 1787 1041 1793 1045
rect 1751 1037 1793 1041
rect 1845 1039 1851 1045
rect 1998 1044 2004 1050
rect 2044 1048 2054 1050
rect 2007 1044 2019 1048
rect 2029 1044 2041 1048
rect 2044 1044 2050 1048
rect 1992 1038 1998 1044
rect 2050 1038 2056 1044
rect 1496 1020 1506 1036
rect 1527 1034 1539 1037
rect 1721 1036 1727 1037
rect 1773 1036 1776 1037
rect 1521 1033 1541 1034
rect 1715 1033 1721 1036
rect 1757 1033 1787 1036
rect 1521 1031 1527 1033
rect 1541 1031 1571 1033
rect 1518 1025 1521 1031
rect 1515 1022 1521 1025
rect 1573 1024 1594 1031
rect 1621 1024 1627 1030
rect 1242 1004 1245 1005
rect 1102 1001 1103 1004
rect 163 982 169 988
rect 180 986 184 992
rect 692 989 705 997
rect 714 993 729 997
rect 178 974 179 979
rect 336 976 352 984
rect 519 976 535 989
rect 602 979 619 989
rect 678 981 692 989
rect 672 979 678 981
rect 619 978 672 979
rect 703 977 711 989
rect 715 987 720 989
rect 766 987 779 997
rect 336 974 393 976
rect 174 957 178 972
rect 336 968 381 974
rect 393 968 397 974
rect 112 944 119 957
rect 173 953 174 956
rect 172 949 173 952
rect 175 944 189 953
rect 320 952 336 968
rect 397 961 402 968
rect 584 952 590 958
rect 630 952 636 958
rect 703 956 711 967
rect 715 958 717 987
rect 965 984 967 1001
rect 971 999 993 1001
rect 971 989 979 999
rect 1097 992 1102 1001
rect 1245 996 1266 1004
rect 1400 1002 1403 1011
rect 1443 1007 1445 1014
rect 1434 1005 1445 1007
rect 1449 1010 1457 1017
rect 1449 1005 1462 1010
rect 1447 1004 1448 1005
rect 1453 1001 1462 1005
rect 1496 1002 1506 1018
rect 1515 1015 1518 1022
rect 1569 1018 1575 1024
rect 1627 1018 1633 1024
rect 1703 1021 1711 1033
rect 1715 1031 1749 1033
rect 1715 1030 1721 1031
rect 1715 1029 1718 1030
rect 1515 1014 1517 1015
rect 1515 1013 1519 1014
rect 1517 1001 1519 1013
rect 1155 995 1188 996
rect 1266 995 1268 996
rect 1190 993 1196 995
rect 1097 986 1103 992
rect 1155 987 1161 992
rect 1196 991 1200 993
rect 1268 991 1278 995
rect 1398 991 1400 997
rect 1440 993 1453 1001
rect 1515 998 1519 1001
rect 1703 999 1711 1011
rect 1715 1002 1717 1029
rect 1995 1024 1998 1036
rect 2050 1032 2053 1036
rect 2003 1018 2007 1031
rect 2050 1021 2066 1032
rect 2066 1018 2082 1021
rect 1792 1007 1793 1008
rect 1793 1005 1794 1006
rect 1715 1001 1718 1002
rect 1761 1001 1789 1002
rect 1715 999 1727 1001
rect 1761 1000 1787 1001
rect 1445 992 1453 993
rect 1506 991 1510 996
rect 1515 991 1520 998
rect 1715 997 1716 999
rect 1761 998 1783 1000
rect 1789 999 1793 1001
rect 1716 995 1719 997
rect 1761 996 1776 998
rect 1715 993 1721 995
rect 1761 994 1777 996
rect 1787 995 1793 999
rect 1796 997 1801 1003
rect 1845 1001 1854 1010
rect 1980 1001 1989 1010
rect 1989 1000 1995 1001
rect 824 981 840 984
rect 842 981 858 984
rect 818 978 838 981
rect 959 979 971 984
rect 1095 979 1096 983
rect 1103 980 1109 986
rect 1113 983 1181 987
rect 1200 986 1212 991
rect 862 974 863 978
rect 820 972 912 974
rect 959 972 979 979
rect 1094 974 1095 979
rect 1113 977 1139 983
rect 1149 980 1155 983
rect 1181 977 1194 983
rect 1212 978 1233 986
rect 1278 978 1312 991
rect 1444 988 1445 990
rect 1382 979 1388 985
rect 1398 983 1399 987
rect 1441 985 1444 986
rect 1093 972 1094 974
rect 1131 972 1139 977
rect 724 963 820 972
rect 862 969 863 972
rect 821 963 833 965
rect 724 960 821 963
rect 715 957 719 958
rect 724 957 820 960
rect 715 956 724 957
rect 698 955 722 956
rect 726 955 749 956
rect 698 953 717 955
rect 766 954 781 957
rect 691 952 698 953
rect 711 952 712 953
rect 327 944 336 952
rect 578 946 584 952
rect 636 946 642 952
rect 672 949 691 952
rect 759 951 766 954
rect 715 950 726 951
rect 757 950 759 951
rect 650 946 672 949
rect 642 945 664 946
rect 105 936 111 942
rect 111 930 117 936
rect 119 934 144 944
rect 159 936 175 944
rect 157 934 175 936
rect 323 935 327 944
rect 715 943 727 950
rect 330 940 336 941
rect 330 939 372 940
rect 376 939 382 941
rect 330 936 341 939
rect 330 935 336 936
rect 372 935 382 939
rect 323 934 330 935
rect 150 929 153 934
rect 157 930 163 934
rect 148 926 150 929
rect 146 923 148 926
rect 320 925 323 934
rect 324 929 330 934
rect 382 929 388 935
rect 389 933 401 941
rect 462 934 468 940
rect 508 934 514 940
rect 778 939 779 954
rect 808 952 818 957
rect 817 939 818 952
rect 863 952 874 968
rect 835 942 843 944
rect 825 940 835 942
rect 823 939 825 940
rect 403 932 405 933
rect 376 927 401 929
rect 318 924 320 925
rect 141 914 146 923
rect 234 922 264 924
rect 314 922 318 924
rect 139 907 141 914
rect 107 895 108 905
rect 137 896 139 907
rect 210 906 234 922
rect 264 916 314 922
rect 399 915 401 927
rect 405 917 413 929
rect 450 926 462 934
rect 514 928 520 934
rect 636 926 639 930
rect 765 927 823 939
rect 863 938 867 952
rect 904 947 905 968
rect 912 965 984 972
rect 908 963 984 965
rect 912 956 984 963
rect 993 962 994 968
rect 987 956 994 962
rect 1033 956 1039 962
rect 1088 956 1093 972
rect 955 955 996 956
rect 981 950 996 955
rect 1039 950 1045 956
rect 870 942 916 944
rect 916 940 924 942
rect 924 939 927 940
rect 835 930 847 938
rect 857 930 869 938
rect 760 926 765 927
rect 519 922 521 924
rect 399 906 402 915
rect 438 910 446 922
rect 450 920 468 922
rect 136 891 137 895
rect 135 888 136 891
rect 197 886 210 906
rect 399 902 401 906
rect 384 897 401 902
rect 376 896 401 897
rect 375 895 401 896
rect 405 895 413 907
rect 324 886 330 889
rect 372 886 401 895
rect 404 892 405 894
rect 438 888 446 900
rect 450 890 452 920
rect 521 916 528 922
rect 528 914 531 916
rect 639 914 653 926
rect 746 923 760 926
rect 769 924 778 927
rect 867 926 869 930
rect 927 927 974 939
rect 987 935 996 950
rect 1086 949 1088 956
rect 1104 952 1113 968
rect 1122 955 1131 972
rect 1194 968 1211 977
rect 1233 968 1272 978
rect 1085 946 1086 949
rect 989 934 994 935
rect 1039 933 1045 936
rect 974 926 979 927
rect 987 926 989 933
rect 1045 930 1052 933
rect 1062 930 1074 938
rect 1082 937 1084 942
rect 1104 937 1113 950
rect 1119 946 1122 955
rect 1164 954 1193 964
rect 1211 963 1272 968
rect 1211 957 1233 963
rect 1272 960 1282 963
rect 1157 945 1193 954
rect 1204 952 1213 954
rect 1116 937 1118 942
rect 1075 926 1082 937
rect 1104 934 1116 937
rect 1148 936 1157 945
rect 1164 944 1193 945
rect 1194 945 1213 952
rect 1233 950 1254 957
rect 1282 956 1292 960
rect 1312 956 1369 978
rect 1388 973 1394 979
rect 1399 977 1400 983
rect 1440 979 1446 985
rect 1400 972 1401 977
rect 1434 974 1440 979
rect 1441 974 1444 979
rect 1434 973 1441 974
rect 1440 972 1441 973
rect 1398 968 1401 972
rect 1449 971 1451 991
rect 1510 985 1516 991
rect 1521 988 1522 990
rect 1523 986 1526 987
rect 1526 985 1531 986
rect 1510 984 1566 985
rect 1715 984 1726 993
rect 1761 990 1773 994
rect 1787 993 1801 995
rect 1845 993 1851 999
rect 1989 998 1996 1000
rect 1998 998 2007 1018
rect 2082 1015 2095 1018
rect 2719 1015 2720 1026
rect 2909 1015 2910 1026
rect 2995 1015 2996 1026
rect 3268 1015 3269 1026
rect 3465 1015 3466 1026
rect 2095 1001 2159 1015
rect 2159 998 2169 1001
rect 1789 992 1799 993
rect 1836 992 1845 993
rect 1989 992 2007 998
rect 2050 992 2056 998
rect 2169 992 2214 998
rect 2309 994 2327 995
rect 2297 992 2309 994
rect 1761 986 1779 990
rect 1793 987 1799 992
rect 1839 987 1845 992
rect 1998 991 2004 992
rect 1998 989 2005 991
rect 2006 990 2007 992
rect 2036 991 2039 992
rect 1998 986 2004 989
rect 2006 987 2010 988
rect 2025 987 2036 991
rect 2041 986 2050 992
rect 2169 988 2297 992
rect 1510 983 1575 984
rect 1719 983 1727 984
rect 1527 981 1575 983
rect 1527 979 1539 981
rect 1721 978 1737 983
rect 1742 981 1743 984
rect 1569 972 1575 978
rect 1627 972 1633 978
rect 1398 967 1403 968
rect 1439 967 1440 971
rect 1389 958 1403 967
rect 1292 954 1297 956
rect 1369 955 1388 956
rect 1389 955 1401 958
rect 1297 951 1304 954
rect 1369 951 1401 955
rect 1403 951 1404 957
rect 1304 950 1306 951
rect 1194 944 1206 945
rect 1164 943 1171 944
rect 1213 943 1222 945
rect 1164 942 1169 943
rect 1164 941 1166 942
rect 1164 940 1210 941
rect 1211 940 1222 943
rect 1160 939 1165 940
rect 1172 939 1206 940
rect 1160 938 1206 939
rect 1160 937 1172 938
rect 1109 926 1116 934
rect 1159 931 1172 937
rect 1203 936 1206 938
rect 1210 937 1222 940
rect 1254 937 1356 950
rect 1369 949 1389 951
rect 1392 949 1408 950
rect 1382 948 1408 949
rect 1382 946 1389 948
rect 1392 945 1409 948
rect 1434 946 1439 967
rect 1451 951 1453 968
rect 1575 966 1581 972
rect 1584 967 1587 972
rect 1453 949 1458 950
rect 1204 931 1206 936
rect 1217 931 1223 937
rect 1254 934 1388 937
rect 1392 934 1408 945
rect 1409 943 1419 945
rect 1446 943 1458 949
rect 1587 948 1594 967
rect 1621 966 1633 972
rect 1726 968 1737 978
rect 1761 980 1780 986
rect 1761 973 1798 980
rect 1922 976 1938 984
rect 2000 982 2003 986
rect 1999 976 2000 981
rect 1743 968 1746 972
rect 1627 945 1633 966
rect 1737 953 1749 968
rect 1765 965 1798 973
rect 1882 968 1885 976
rect 1923 975 1938 976
rect 1998 970 1999 975
rect 2041 969 2044 986
rect 2053 972 2154 977
rect 2154 969 2165 972
rect 2196 969 2297 988
rect 2327 980 2349 994
rect 1743 951 1746 953
rect 1749 951 1751 953
rect 1419 934 1483 943
rect 1751 942 1771 951
rect 1780 948 1798 965
rect 1878 957 1882 968
rect 1873 955 1878 957
rect 1835 950 1836 953
rect 1584 936 1666 942
rect 1567 934 1584 936
rect 1160 930 1172 931
rect 737 921 746 923
rect 725 920 737 921
rect 764 920 769 924
rect 678 915 764 920
rect 666 914 678 915
rect 706 914 725 915
rect 823 914 831 926
rect 835 924 869 926
rect 531 913 661 914
rect 639 909 653 913
rect 695 911 706 914
rect 688 907 694 911
rect 578 900 584 906
rect 584 894 590 900
rect 612 892 625 900
rect 655 892 666 907
rect 680 900 685 904
rect 817 901 826 913
rect 835 901 837 924
rect 450 888 468 890
rect 612 889 621 892
rect 625 891 627 892
rect 667 889 669 891
rect 677 889 686 898
rect 826 892 837 901
rect 867 892 869 924
rect 873 914 881 926
rect 979 924 989 926
rect 1046 924 1074 926
rect 1075 924 1086 926
rect 979 923 987 924
rect 984 921 987 923
rect 1039 921 1040 924
rect 1072 921 1086 924
rect 905 907 919 921
rect 974 910 984 921
rect 1038 917 1039 921
rect 974 907 987 910
rect 1037 907 1038 916
rect 1072 915 1074 921
rect 1075 915 1086 921
rect 1109 924 1117 926
rect 1109 915 1116 924
rect 1117 921 1121 924
rect 1120 918 1126 921
rect 1121 916 1126 918
rect 1072 911 1075 915
rect 1077 914 1086 915
rect 1077 912 1078 914
rect 919 906 974 907
rect 981 904 987 907
rect 1036 904 1037 906
rect 1039 904 1045 910
rect 1072 906 1074 911
rect 1078 907 1080 912
rect 1080 906 1081 907
rect 1071 904 1074 906
rect 1081 904 1082 906
rect 987 898 993 904
rect 1029 902 1032 904
rect 1033 902 1039 904
rect 1028 898 1039 902
rect 1070 901 1071 904
rect 1028 892 1035 898
rect 1069 897 1070 900
rect 1067 894 1069 895
rect 1072 894 1074 904
rect 1040 892 1074 894
rect 1078 901 1086 904
rect 1078 892 1092 901
rect 1067 891 1069 892
rect 1092 890 1095 892
rect 193 879 197 885
rect 319 879 372 886
rect 382 883 388 886
rect 389 883 401 886
rect 456 884 462 888
rect 190 875 193 879
rect 289 875 319 879
rect 330 877 336 879
rect 135 871 136 875
rect 187 870 190 874
rect 251 870 289 875
rect 249 869 251 870
rect 186 868 187 869
rect 247 868 249 869
rect 338 868 340 879
rect 373 868 374 879
rect 376 877 382 883
rect 450 882 462 884
rect 514 882 520 888
rect 450 876 468 882
rect 508 876 514 882
rect 621 880 630 889
rect 667 888 677 889
rect 1065 888 1067 889
rect 668 887 677 888
rect 668 880 688 887
rect 870 885 871 888
rect 831 882 832 884
rect 1040 880 1052 888
rect 1062 882 1074 888
rect 1095 884 1097 890
rect 1099 885 1109 915
rect 1126 912 1139 916
rect 1139 907 1151 912
rect 1154 906 1156 907
rect 1165 906 1172 930
rect 1217 928 1218 931
rect 1340 919 1388 934
rect 1408 932 1483 934
rect 1500 933 1551 934
rect 1553 933 1564 934
rect 1500 932 1561 933
rect 1408 930 1500 932
rect 1156 904 1161 906
rect 1165 904 1217 906
rect 1161 901 1217 904
rect 1165 899 1217 901
rect 1148 889 1157 898
rect 1165 896 1234 899
rect 1165 891 1222 896
rect 1234 892 1259 896
rect 1356 894 1364 919
rect 1388 916 1395 919
rect 1408 918 1424 930
rect 1426 918 1442 930
rect 1547 929 1562 932
rect 1543 927 1547 929
rect 1527 922 1543 927
rect 1553 926 1562 929
rect 1596 926 1603 936
rect 1556 920 1561 922
rect 1374 900 1378 916
rect 1395 914 1426 916
rect 1427 914 1429 918
rect 1395 909 1427 914
rect 1418 907 1435 909
rect 1418 902 1427 907
rect 1435 906 1439 907
rect 1378 896 1379 899
rect 1398 898 1418 902
rect 1159 889 1223 891
rect 1259 890 1271 892
rect 1355 890 1356 893
rect 1157 885 1223 889
rect 1061 880 1074 882
rect 631 875 634 880
rect 675 879 688 880
rect 173 864 186 868
rect 241 864 247 868
rect 167 862 173 864
rect 238 862 241 864
rect 164 858 167 862
rect 231 857 238 862
rect 163 856 164 857
rect 230 856 231 857
rect 162 849 163 856
rect 227 849 230 856
rect 161 841 162 849
rect 229 838 238 842
rect 276 838 285 842
rect 288 838 304 854
rect 306 838 322 854
rect 340 838 344 867
rect 371 847 373 867
rect 634 860 641 875
rect 673 873 688 875
rect 384 849 398 854
rect 480 842 484 856
rect 157 804 161 838
rect 226 833 238 838
rect 272 833 288 838
rect 322 837 338 838
rect 329 834 338 837
rect 220 832 233 833
rect 272 832 294 833
rect 218 831 227 832
rect 218 811 220 831
rect 221 826 227 831
rect 217 810 220 811
rect 218 804 220 810
rect 226 820 227 826
rect 259 824 294 832
rect 259 823 288 824
rect 259 822 307 823
rect 333 822 338 834
rect 259 820 279 822
rect 288 820 307 822
rect 226 804 242 820
rect 272 804 288 820
rect 332 812 333 817
rect 161 799 174 804
rect 191 799 226 804
rect 174 797 191 799
rect 210 788 227 799
rect 288 797 291 803
rect 288 795 292 797
rect 288 788 298 795
rect 218 786 227 788
rect 292 786 298 788
rect 343 786 344 828
rect 368 822 381 838
rect 514 833 518 838
rect 536 837 548 845
rect 602 838 618 854
rect 641 842 650 860
rect 642 841 650 842
rect 654 845 655 862
rect 654 843 658 845
rect 686 844 688 873
rect 689 869 700 875
rect 692 863 700 869
rect 696 859 699 863
rect 832 860 836 879
rect 869 866 870 880
rect 951 867 957 873
rect 997 867 1003 873
rect 1061 870 1065 880
rect 1094 870 1099 884
rect 1157 880 1171 885
rect 1165 871 1171 880
rect 1207 880 1217 885
rect 1207 870 1208 880
rect 1211 879 1217 880
rect 1271 879 1338 890
rect 1354 885 1355 889
rect 1353 881 1354 885
rect 1339 875 1343 879
rect 1343 872 1346 875
rect 1350 871 1353 881
rect 1379 879 1383 896
rect 1393 891 1398 898
rect 1439 892 1496 906
rect 1496 891 1499 892
rect 1390 881 1392 889
rect 1499 888 1513 891
rect 1559 890 1561 920
rect 1565 910 1573 922
rect 1603 914 1608 926
rect 1608 902 1613 914
rect 1633 910 1640 936
rect 1666 934 1670 936
rect 1747 935 1748 942
rect 1771 936 1783 942
rect 1670 933 1671 934
rect 1671 927 1674 933
rect 1674 922 1677 927
rect 1677 919 1679 922
rect 1679 916 1680 919
rect 1530 888 1561 890
rect 1565 888 1573 900
rect 1613 899 1614 902
rect 1640 900 1642 910
rect 1680 902 1687 916
rect 1748 910 1752 935
rect 1783 934 1787 936
rect 1798 935 1799 942
rect 1785 933 1791 934
rect 1785 932 1793 933
rect 1799 932 1800 935
rect 1835 934 1850 950
rect 1873 948 1885 955
rect 1872 947 1885 948
rect 1895 947 1907 955
rect 1938 952 1954 968
rect 1869 945 1878 947
rect 1868 943 1869 945
rect 1872 943 1878 945
rect 1911 943 1912 945
rect 1918 943 1924 948
rect 1861 942 1868 943
rect 1872 942 1907 943
rect 1911 942 1924 943
rect 1861 937 1872 942
rect 1873 941 1907 942
rect 1859 934 1865 937
rect 1866 936 1872 937
rect 1906 936 1907 941
rect 1924 936 1930 942
rect 1938 934 1954 950
rect 1990 934 1998 968
rect 2044 956 2045 968
rect 2049 965 2050 969
rect 2165 968 2184 969
rect 2192 968 2196 969
rect 2156 964 2192 968
rect 2242 965 2246 969
rect 1855 932 1859 934
rect 1793 931 1834 932
rect 1799 918 1816 931
rect 1818 926 1834 931
rect 1852 930 1855 932
rect 1845 926 1852 930
rect 1937 927 1938 931
rect 1989 927 1990 932
rect 1818 918 1845 926
rect 1936 920 1938 927
rect 1988 922 1989 927
rect 1999 922 2007 934
rect 2011 922 2013 956
rect 2049 951 2050 964
rect 2156 960 2204 964
rect 2147 954 2156 960
rect 2044 945 2045 951
rect 2050 936 2051 945
rect 2136 936 2147 954
rect 2185 949 2204 960
rect 2204 948 2206 949
rect 2246 948 2251 965
rect 2349 961 2352 980
rect 2352 954 2353 960
rect 2206 945 2210 948
rect 2251 945 2252 948
rect 2131 934 2147 936
rect 2051 928 2057 934
rect 2052 922 2057 928
rect 2131 928 2143 934
rect 2153 928 2165 936
rect 2210 934 2225 945
rect 2252 934 2256 945
rect 2353 934 2356 954
rect 2225 932 2226 934
rect 2226 928 2227 930
rect 2256 929 2258 934
rect 2131 924 2136 928
rect 2169 926 2170 928
rect 2171 924 2174 925
rect 1935 919 1938 920
rect 1799 905 1800 918
rect 1827 916 1845 918
rect 1934 918 1938 919
rect 1934 916 1935 918
rect 1987 916 1988 919
rect 2007 916 2008 921
rect 1821 912 1827 916
rect 1930 909 1934 916
rect 1986 909 1987 916
rect 2008 912 2010 916
rect 2038 913 2045 922
rect 2052 916 2053 922
rect 2031 911 2038 913
rect 2049 911 2053 916
rect 2119 912 2127 924
rect 2131 922 2165 924
rect 2131 921 2134 922
rect 2011 910 2049 911
rect 1800 902 1801 904
rect 1687 899 1689 902
rect 1642 894 1643 899
rect 1689 896 1690 899
rect 1513 885 1524 888
rect 1527 885 1566 888
rect 1524 884 1566 885
rect 1383 872 1385 879
rect 1385 870 1386 872
rect 1387 871 1390 881
rect 1527 879 1566 884
rect 1615 881 1617 889
rect 1549 876 1561 879
rect 1566 874 1588 879
rect 1617 874 1618 881
rect 1602 872 1607 874
rect 1036 868 1037 869
rect 1060 867 1061 870
rect 945 861 951 867
rect 1003 861 1009 867
rect 1058 860 1060 867
rect 699 854 703 858
rect 699 853 714 854
rect 685 843 688 844
rect 654 841 688 843
rect 692 841 700 853
rect 703 850 714 853
rect 836 852 837 858
rect 870 854 871 858
rect 705 840 714 850
rect 471 831 548 833
rect 371 820 376 822
rect 368 804 381 820
rect 371 787 376 804
rect 384 788 400 799
rect 220 780 227 786
rect 285 785 298 786
rect 285 783 332 785
rect 260 780 307 783
rect 220 777 233 780
rect 273 777 279 780
rect 285 779 307 780
rect 285 777 294 779
rect 471 777 529 831
rect 546 799 548 831
rect 552 821 560 833
rect 618 822 634 838
rect 688 837 692 840
rect 712 838 714 840
rect 736 838 742 844
rect 782 839 788 844
rect 778 838 790 839
rect 837 838 840 850
rect 872 841 888 854
rect 943 852 951 858
rect 941 850 951 852
rect 1055 851 1058 860
rect 1004 848 1014 850
rect 1014 846 1020 848
rect 1053 847 1055 851
rect 931 844 945 846
rect 1020 844 1027 846
rect 871 840 888 841
rect 871 838 875 840
rect 654 829 666 837
rect 676 829 688 837
rect 714 832 794 838
rect 840 832 841 837
rect 654 828 655 829
rect 655 818 657 828
rect 714 822 730 832
rect 736 831 790 832
rect 736 827 788 831
rect 657 814 659 818
rect 659 809 660 812
rect 660 805 661 809
rect 661 799 662 803
rect 662 792 664 799
rect 736 793 756 827
rect 782 825 790 827
rect 788 794 790 825
rect 794 815 802 827
rect 782 793 790 794
rect 794 793 802 805
rect 818 804 826 820
rect 841 814 844 829
rect 856 822 875 838
rect 909 833 918 842
rect 931 841 951 844
rect 1027 843 1031 844
rect 1031 842 1036 843
rect 1052 842 1053 844
rect 1048 841 1059 842
rect 1084 841 1094 869
rect 1099 866 1100 869
rect 1100 854 1103 865
rect 1171 860 1176 870
rect 1347 869 1350 870
rect 1346 865 1350 869
rect 1347 860 1350 865
rect 1377 866 1387 870
rect 1607 866 1624 872
rect 1643 871 1647 890
rect 1690 888 1694 896
rect 1798 890 1801 896
rect 1807 891 1818 908
rect 1873 903 1885 909
rect 1985 908 1986 909
rect 1914 903 1930 908
rect 1984 903 1985 908
rect 2031 903 2038 910
rect 1885 902 1914 903
rect 1983 896 1984 899
rect 1866 890 1872 896
rect 1924 890 1930 896
rect 1694 874 1702 888
rect 1796 885 1798 889
rect 1804 886 1807 890
rect 1176 854 1177 860
rect 1346 854 1349 860
rect 1100 852 1106 854
rect 1103 841 1106 852
rect 1168 849 1184 854
rect 1167 848 1181 849
rect 1186 848 1202 854
rect 1159 841 1167 848
rect 1181 842 1204 848
rect 931 838 945 841
rect 1051 839 1052 841
rect 1059 840 1094 841
rect 1105 840 1106 841
rect 1157 840 1159 841
rect 1084 839 1132 840
rect 1155 838 1157 840
rect 1171 839 1183 842
rect 1264 841 1280 854
rect 1282 841 1298 854
rect 1344 847 1346 853
rect 1347 852 1349 854
rect 1377 852 1395 866
rect 1618 863 1633 866
rect 1204 840 1205 841
rect 1257 840 1258 841
rect 1176 838 1183 839
rect 925 834 939 838
rect 925 833 936 834
rect 900 824 909 833
rect 871 820 875 822
rect 856 814 875 820
rect 844 809 845 812
rect 845 799 847 808
rect 856 804 872 814
rect 931 812 939 824
rect 943 814 945 838
rect 1048 832 1051 838
rect 1003 815 1009 821
rect 1037 818 1055 832
rect 1043 815 1044 818
rect 997 814 1003 815
rect 1042 814 1043 815
rect 943 812 977 814
rect 986 812 1045 814
rect 1055 813 1061 818
rect 1056 812 1062 813
rect 875 808 876 812
rect 967 809 977 812
rect 981 810 986 812
rect 958 808 967 809
rect 970 808 976 809
rect 978 808 981 810
rect 997 809 1003 812
rect 876 804 877 808
rect 943 805 955 808
rect 958 805 977 808
rect 943 804 956 805
rect 872 794 880 804
rect 903 800 955 804
rect 965 800 977 805
rect 1033 800 1042 811
rect 1045 810 1053 812
rect 1056 810 1067 812
rect 1075 811 1084 838
rect 1106 822 1122 838
rect 1146 832 1154 838
rect 1053 809 1067 810
rect 1069 809 1075 810
rect 1053 808 1075 809
rect 1106 808 1122 820
rect 1175 811 1177 838
rect 1178 837 1183 838
rect 1180 836 1183 837
rect 1205 838 1206 840
rect 1256 838 1257 840
rect 1181 834 1185 836
rect 1186 832 1187 834
rect 1205 832 1218 838
rect 1179 828 1183 830
rect 1056 804 1122 808
rect 1065 800 1106 804
rect 1146 801 1147 804
rect 872 793 882 794
rect 736 792 788 793
rect 872 792 884 793
rect 664 789 670 792
rect 670 784 677 789
rect 730 788 810 792
rect 848 790 849 792
rect 872 789 893 792
rect 872 788 887 789
rect 730 786 794 788
rect 882 786 887 788
rect 893 787 898 789
rect 898 786 902 787
rect 903 786 954 800
rect 966 793 970 800
rect 1028 793 1033 799
rect 965 790 966 793
rect 1026 790 1028 793
rect 677 783 678 784
rect 713 783 714 785
rect 679 779 685 783
rect 710 779 713 783
rect 736 780 742 786
rect 778 781 790 786
rect 898 785 909 786
rect 900 783 909 785
rect 900 782 912 783
rect 782 780 788 781
rect 848 779 849 781
rect 685 777 690 779
rect 709 777 710 779
rect 107 755 108 775
rect 136 772 137 775
rect 227 774 266 777
rect 273 774 285 777
rect 137 759 145 772
rect 229 768 266 774
rect 276 768 285 774
rect 342 768 343 777
rect 137 755 148 759
rect 108 749 109 755
rect 145 753 148 755
rect 146 750 151 753
rect 120 747 149 748
rect 152 747 153 749
rect 102 713 109 725
rect 114 716 115 747
rect 143 745 148 747
rect 147 716 148 745
rect 149 738 160 747
rect 376 740 380 777
rect 685 776 709 777
rect 846 775 848 779
rect 900 777 909 782
rect 915 779 918 781
rect 918 777 937 779
rect 965 777 974 786
rect 996 782 1002 788
rect 1023 786 1026 790
rect 1042 782 1048 788
rect 1060 786 1069 800
rect 1072 788 1088 800
rect 1090 796 1126 800
rect 1147 798 1149 801
rect 1174 800 1175 810
rect 1181 798 1183 828
rect 1187 818 1195 830
rect 1204 822 1218 832
rect 1248 836 1256 838
rect 1310 837 1314 841
rect 1342 839 1344 847
rect 1377 838 1387 852
rect 1395 848 1398 852
rect 1525 842 1531 844
rect 1525 838 1539 842
rect 1571 838 1577 844
rect 1578 838 1594 854
rect 1618 838 1624 863
rect 1633 853 1636 863
rect 1636 838 1641 852
rect 1248 822 1255 836
rect 1272 826 1284 832
rect 1269 825 1328 826
rect 1332 825 1342 838
rect 1269 823 1277 825
rect 1328 823 1342 825
rect 1349 823 1352 838
rect 1204 820 1207 822
rect 1268 821 1269 823
rect 1147 796 1183 798
rect 1187 796 1195 808
rect 1204 804 1218 820
rect 1260 816 1268 820
rect 1272 818 1279 820
rect 1260 808 1266 816
rect 1272 814 1273 818
rect 1332 816 1357 823
rect 1366 816 1377 837
rect 1398 822 1410 838
rect 1519 832 1525 838
rect 1523 830 1525 832
rect 1527 830 1560 838
rect 1577 832 1583 838
rect 1594 832 1610 838
rect 1624 832 1625 838
rect 1577 830 1610 832
rect 1641 830 1644 838
rect 1647 830 1659 870
rect 1702 863 1707 874
rect 1749 871 1752 885
rect 1786 881 1796 885
rect 1872 884 1878 890
rect 1882 887 1883 890
rect 1892 886 1899 890
rect 1883 883 1886 885
rect 1889 884 1891 885
rect 1918 884 1924 890
rect 1981 888 1983 896
rect 1883 882 1888 883
rect 1784 874 1802 881
rect 1767 870 1784 874
rect 1786 870 1796 874
rect 1707 859 1709 863
rect 1733 838 1749 870
rect 1767 866 1786 870
rect 1765 863 1767 866
rect 1763 859 1765 863
rect 1779 859 1786 866
rect 1761 856 1763 859
rect 1759 854 1761 856
rect 1752 851 1761 854
rect 1752 839 1759 851
rect 1752 838 1753 839
rect 1709 830 1710 838
rect 1733 830 1752 838
rect 1766 830 1779 859
rect 1796 846 1803 858
rect 1808 848 1809 880
rect 1875 876 1881 879
rect 1872 874 1875 876
rect 1863 869 1872 874
rect 1883 870 1886 882
rect 1920 870 1923 884
rect 1980 881 1981 888
rect 1979 874 1980 881
rect 1856 860 1857 863
rect 1886 860 1888 870
rect 1920 862 1934 870
rect 1976 863 1979 874
rect 1851 848 1856 860
rect 1808 847 1813 848
rect 1808 846 1842 847
rect 1849 846 1854 848
rect 1803 844 1804 846
rect 1848 844 1849 846
rect 1845 842 1847 843
rect 1808 834 1820 841
rect 1830 834 1842 841
rect 1888 830 1899 859
rect 1923 830 1934 862
rect 1975 856 1976 859
rect 2013 856 2031 903
rect 2119 890 2127 902
rect 2131 890 2133 921
rect 2164 920 2165 922
rect 2171 912 2177 924
rect 2227 913 2229 925
rect 2258 924 2274 928
rect 2344 925 2353 934
rect 2336 924 2344 925
rect 2258 913 2336 924
rect 2171 911 2174 912
rect 2174 903 2179 910
rect 2212 905 2274 913
rect 2206 903 2212 905
rect 2165 890 2206 903
rect 2174 888 2179 890
rect 2229 889 2231 905
rect 2127 886 2130 888
rect 2179 886 2180 888
rect 2231 885 2232 888
rect 2130 884 2132 885
rect 2131 883 2133 884
rect 2131 879 2134 883
rect 2180 880 2181 882
rect 2131 878 2135 879
rect 2134 876 2135 878
rect 2181 876 2182 880
rect 2232 876 2233 879
rect 2258 878 2274 905
rect 2135 869 2138 874
rect 2138 863 2140 869
rect 2073 861 2074 862
rect 2140 860 2141 863
rect 1952 851 1968 854
rect 1972 851 1975 856
rect 2011 851 2013 856
rect 2054 854 2066 855
rect 1952 843 1972 851
rect 2008 843 2011 851
rect 2048 849 2066 854
rect 2076 849 2088 855
rect 2048 843 2139 849
rect 2141 848 2145 860
rect 2145 844 2146 847
rect 2162 843 2178 854
rect 1950 839 1953 843
rect 2006 839 2008 843
rect 2042 842 2047 843
rect 2042 840 2046 842
rect 2048 841 2088 843
rect 2035 839 2045 840
rect 2048 839 2054 841
rect 2029 838 2034 839
rect 2048 838 2049 839
rect 1936 830 1950 838
rect 2003 836 2006 838
rect 2025 837 2029 838
rect 2016 836 2022 837
rect 2003 834 2016 836
rect 1993 833 1997 834
rect 1987 832 1993 833
rect 1974 830 1987 832
rect 2003 831 2006 834
rect 1515 827 1523 830
rect 1527 828 1530 830
rect 1514 821 1524 827
rect 1203 802 1204 804
rect 1205 800 1207 804
rect 1332 801 1342 816
rect 1344 812 1352 816
rect 1344 804 1353 812
rect 1357 807 1389 816
rect 1398 807 1410 820
rect 1490 807 1514 821
rect 1515 818 1523 821
rect 1353 801 1354 803
rect 1366 801 1377 807
rect 1389 804 1410 807
rect 1090 788 1106 796
rect 1126 795 1131 796
rect 1131 793 1142 795
rect 1149 794 1156 796
rect 1156 793 1162 794
rect 1173 793 1174 796
rect 1142 792 1147 793
rect 1162 792 1182 793
rect 1185 792 1187 795
rect 1202 794 1203 796
rect 1162 786 1183 792
rect 1199 789 1202 793
rect 1184 788 1202 789
rect 1184 786 1199 788
rect 1255 786 1256 788
rect 1260 786 1266 798
rect 1314 789 1315 801
rect 1329 790 1332 800
rect 1354 797 1382 801
rect 1389 797 1408 804
rect 1478 800 1490 807
rect 1476 799 1478 800
rect 1354 796 1408 797
rect 1469 796 1476 799
rect 1515 796 1523 808
rect 1527 796 1529 828
rect 1595 822 1824 830
rect 1595 820 1597 822
rect 1598 820 1824 822
rect 1595 814 1824 820
rect 1852 814 1974 830
rect 1997 818 2003 831
rect 2032 822 2048 838
rect 1995 815 2002 818
rect 1595 812 1852 814
rect 1597 804 1610 812
rect 1627 807 1629 812
rect 1597 803 1598 804
rect 1598 801 1599 802
rect 1595 796 1598 801
rect 1628 800 1629 807
rect 1640 804 1652 812
rect 1652 803 1653 804
rect 1657 803 1659 808
rect 1676 803 1755 812
rect 1653 802 1755 803
rect 1656 799 1672 802
rect 1273 787 1274 788
rect 1272 786 1278 787
rect 1054 782 1060 786
rect 1171 784 1183 786
rect 845 772 846 774
rect 909 772 937 777
rect 838 759 845 772
rect 909 768 918 772
rect 956 768 965 777
rect 990 776 996 782
rect 1048 776 1060 782
rect 1172 776 1173 781
rect 1048 766 1052 773
rect 1204 772 1205 786
rect 1256 783 1257 786
rect 1267 784 1269 785
rect 1313 784 1314 788
rect 1328 787 1329 790
rect 1354 789 1398 796
rect 1408 795 1410 796
rect 1410 792 1417 795
rect 1467 793 1469 796
rect 1566 795 1594 796
rect 1417 789 1421 792
rect 1354 788 1376 789
rect 1378 788 1394 789
rect 1421 788 1423 789
rect 1463 788 1467 793
rect 1578 792 1594 795
rect 1624 793 1628 799
rect 1335 787 1342 788
rect 1350 787 1364 788
rect 1423 787 1426 788
rect 1327 786 1335 787
rect 1322 785 1335 786
rect 1354 785 1364 787
rect 1519 786 1525 792
rect 1577 791 1594 792
rect 1621 791 1624 793
rect 1577 789 1633 791
rect 1654 789 1672 799
rect 1577 788 1594 789
rect 1621 788 1624 789
rect 1633 788 1672 789
rect 1674 788 1755 802
rect 1766 800 1779 812
rect 1842 804 1843 807
rect 1577 786 1583 788
rect 1620 786 1621 788
rect 1319 784 1328 785
rect 1257 780 1269 783
rect 1272 780 1273 781
rect 1281 780 1319 784
rect 1257 779 1316 780
rect 1272 774 1284 779
rect 1203 763 1205 772
rect 1322 763 1328 784
rect 1354 784 1368 785
rect 828 756 845 759
rect 1169 756 1172 763
rect 828 755 838 756
rect 828 754 835 755
rect 1168 754 1169 756
rect 828 753 832 754
rect 817 749 859 753
rect 817 748 844 749
rect 815 747 817 748
rect 859 747 862 749
rect 801 745 815 747
rect 333 738 339 740
rect 376 739 385 740
rect 153 735 171 738
rect 160 725 171 735
rect 333 734 345 738
rect 379 734 385 739
rect 768 738 801 745
rect 762 737 767 738
rect 327 728 333 734
rect 385 729 391 734
rect 739 733 762 737
rect 816 735 824 747
rect 828 746 833 747
rect 733 731 739 733
rect 727 729 729 731
rect 349 728 480 729
rect 333 726 349 728
rect 385 727 688 728
rect 715 727 721 729
rect 726 728 727 729
rect 480 726 481 727
rect 688 726 721 727
rect 724 726 726 728
rect 114 714 118 716
rect 145 714 148 716
rect 114 713 148 714
rect 153 713 171 725
rect 321 714 329 726
rect 333 724 339 726
rect 109 711 110 713
rect 110 708 115 711
rect 148 708 153 711
rect 114 707 126 708
rect 113 701 126 707
rect 136 701 148 708
rect 160 707 171 713
rect 113 694 115 701
rect 171 690 178 707
rect 321 692 329 704
rect 333 694 335 724
rect 482 719 486 726
rect 688 723 723 726
rect 761 723 767 729
rect 486 708 493 719
rect 709 717 715 723
rect 716 719 723 723
rect 767 719 773 723
rect 816 719 824 725
rect 828 719 830 746
rect 1157 744 1163 750
rect 1165 744 1168 754
rect 1203 750 1204 763
rect 1309 757 1315 762
rect 1321 757 1322 762
rect 1354 758 1364 784
rect 1368 783 1372 784
rect 1427 783 1433 786
rect 1462 783 1463 786
rect 1525 784 1539 786
rect 1525 783 1531 784
rect 1563 783 1567 784
rect 1434 781 1436 782
rect 1436 780 1439 781
rect 1452 780 1462 783
rect 1381 775 1387 779
rect 1387 772 1392 775
rect 1439 772 1462 780
rect 1393 766 1417 772
rect 1452 769 1484 772
rect 1490 769 1563 783
rect 1571 780 1577 786
rect 1578 784 1579 785
rect 1619 784 1620 786
rect 1654 783 1657 788
rect 1663 787 1755 788
rect 1727 786 1755 787
rect 1704 785 1755 786
rect 1763 785 1766 799
rect 1841 797 1842 801
rect 1888 800 1899 814
rect 1923 804 1934 814
rect 1936 804 1952 814
rect 1989 807 2002 815
rect 1986 805 2002 807
rect 2032 805 2048 820
rect 2086 811 2088 841
rect 2092 831 2100 843
rect 2139 838 2179 843
rect 2182 842 2189 874
rect 2224 840 2232 852
rect 2236 842 2238 874
rect 2268 857 2273 874
rect 2268 842 2270 857
rect 2273 852 2274 856
rect 2236 840 2270 842
rect 2274 840 2282 852
rect 2189 838 2190 840
rect 2276 838 2278 840
rect 2179 837 2194 838
rect 2236 837 2237 838
rect 2188 836 2194 837
rect 2233 836 2235 837
rect 2070 809 2088 811
rect 2092 809 2100 821
rect 2149 805 2159 836
rect 2188 832 2203 836
rect 2191 808 2203 832
rect 2236 828 2248 836
rect 2258 828 2270 836
rect 2276 828 2290 838
rect 2237 820 2239 828
rect 2190 807 2203 808
rect 1975 804 2088 805
rect 1952 803 2088 804
rect 1840 791 1841 796
rect 1839 788 1840 791
rect 1899 789 1902 799
rect 1934 794 1942 800
rect 1952 795 1968 803
rect 1970 799 2088 803
rect 2159 801 2163 805
rect 2189 804 2203 807
rect 2224 815 2239 820
rect 2278 822 2290 828
rect 2278 820 2280 822
rect 2224 804 2240 815
rect 2278 805 2290 820
rect 2730 819 2731 1015
rect 2920 819 2921 1015
rect 3006 819 3007 1015
rect 3279 819 3280 1015
rect 3476 819 3477 1015
rect 2280 804 2290 805
rect 2188 803 2189 804
rect 2187 801 2188 802
rect 2135 799 2178 801
rect 1970 796 2135 799
rect 1970 795 2076 796
rect 2159 795 2178 799
rect 1952 794 1986 795
rect 1934 792 1968 794
rect 1913 789 1942 792
rect 1828 785 1839 788
rect 1888 787 1913 789
rect 1875 786 1888 787
rect 1871 785 1875 786
rect 1730 784 1733 785
rect 1751 784 1839 785
rect 1751 783 1828 784
rect 1844 783 1871 785
rect 1899 784 1902 787
rect 1573 779 1574 780
rect 1611 769 1619 783
rect 1653 778 1654 783
rect 1729 781 1730 783
rect 1752 782 1754 783
rect 1728 778 1729 781
rect 1754 780 1757 782
rect 1762 781 1763 783
rect 1820 782 1844 783
rect 1809 779 1820 782
rect 1757 778 1760 779
rect 1309 756 1327 757
rect 1355 756 1361 758
rect 1303 750 1367 756
rect 1392 753 1422 766
rect 1452 763 1490 769
rect 1608 763 1611 769
rect 1452 759 1484 763
rect 1451 756 1452 758
rect 1392 750 1428 753
rect 1449 752 1451 756
rect 1453 755 1484 759
rect 1481 754 1483 755
rect 1484 754 1487 755
rect 1603 754 1608 763
rect 1480 752 1481 754
rect 1487 751 1492 754
rect 1602 752 1603 754
rect 1203 744 1209 750
rect 1309 745 1361 750
rect 1113 742 1157 744
rect 962 741 996 742
rect 1113 741 1119 742
rect 925 740 962 741
rect 902 739 925 740
rect 899 737 902 739
rect 1151 738 1157 742
rect 1209 738 1215 744
rect 874 723 899 737
rect 990 730 996 736
rect 1048 731 1054 736
rect 1303 733 1315 745
rect 1349 735 1354 745
rect 1079 731 1115 733
rect 996 724 1002 730
rect 1020 729 1079 731
rect 1115 729 1121 731
rect 1018 726 1020 729
rect 869 720 874 723
rect 767 717 849 719
rect 770 716 849 717
rect 866 716 874 720
rect 816 713 824 716
rect 828 715 830 716
rect 849 715 878 716
rect 828 713 862 715
rect 859 709 862 713
rect 866 713 874 715
rect 878 714 906 715
rect 866 711 869 713
rect 863 709 866 711
rect 906 710 920 714
rect 1012 713 1018 726
rect 1042 724 1048 729
rect 1121 726 1132 729
rect 1309 726 1315 733
rect 1111 722 1113 723
rect 1132 722 1143 726
rect 1308 723 1315 726
rect 1143 721 1145 722
rect 1145 720 1149 721
rect 493 707 494 708
rect 715 707 716 708
rect 828 701 840 709
rect 850 701 862 709
rect 920 705 926 710
rect 1010 708 1012 713
rect 1009 707 1010 708
rect 926 703 937 705
rect 554 697 688 700
rect 854 698 858 701
rect 937 699 950 703
rect 950 698 955 699
rect 430 695 554 697
rect 688 695 694 697
rect 333 692 339 694
rect 408 692 430 695
rect 694 692 700 695
rect 115 688 116 690
rect 329 688 331 691
rect 332 688 333 690
rect 385 689 408 692
rect 700 689 706 692
rect 838 690 854 698
rect 955 694 971 698
rect 971 692 987 694
rect 987 691 996 692
rect 1002 691 1009 706
rect 1103 693 1111 698
rect 1115 693 1117 720
rect 1303 711 1315 723
rect 1354 711 1356 726
rect 1392 723 1422 750
rect 1448 749 1449 751
rect 1492 750 1494 751
rect 1432 746 1434 747
rect 1446 745 1448 749
rect 1435 737 1449 745
rect 1477 744 1479 749
rect 1497 747 1500 749
rect 1500 746 1502 747
rect 1502 743 1506 746
rect 1526 743 1538 749
rect 1597 744 1600 749
rect 1632 744 1653 778
rect 1719 756 1728 778
rect 1757 776 1762 778
rect 1763 776 1809 779
rect 1902 778 1903 781
rect 1757 775 1809 776
rect 1757 756 1762 775
rect 1903 772 1907 778
rect 1903 756 1910 772
rect 1934 756 1942 789
rect 1952 788 1968 792
rect 1970 788 1986 794
rect 2048 788 2064 795
rect 2162 788 2178 795
rect 2165 787 2166 788
rect 2166 783 2167 785
rect 2168 772 2171 779
rect 2191 778 2203 804
rect 2240 799 2241 802
rect 2240 796 2242 799
rect 2278 796 2280 800
rect 2240 791 2248 796
rect 2275 791 2278 796
rect 2240 788 2256 791
rect 2258 788 2274 791
rect 1714 745 1719 756
rect 1754 744 1757 756
rect 1907 750 1910 756
rect 1907 744 1914 750
rect 1942 744 1944 756
rect 1972 751 1984 759
rect 1994 751 2006 759
rect 2171 755 2176 772
rect 2203 770 2207 778
rect 1954 747 1960 750
rect 2008 749 2010 750
rect 1963 747 1967 749
rect 1954 746 1963 747
rect 1953 744 1961 746
rect 1972 745 2008 747
rect 2010 745 2018 747
rect 1475 738 1477 743
rect 1506 741 1538 743
rect 1534 740 1539 741
rect 1541 737 1544 739
rect 1594 738 1597 744
rect 1629 739 1632 744
rect 1712 740 1714 744
rect 1729 740 1741 742
rect 1442 734 1443 737
rect 1449 734 1453 737
rect 1441 732 1442 734
rect 1453 732 1457 734
rect 1473 732 1475 737
rect 1503 736 1504 737
rect 1533 734 1543 737
rect 1544 734 1550 737
rect 1556 734 1562 737
rect 1538 732 1543 734
rect 1438 725 1441 731
rect 1457 729 1461 732
rect 1471 729 1473 731
rect 1437 722 1438 724
rect 1433 711 1437 721
rect 1461 712 1489 729
rect 1502 726 1503 731
rect 1543 727 1547 732
rect 1549 731 1562 734
rect 1587 732 1591 734
rect 1585 731 1587 732
rect 1602 731 1608 737
rect 1692 734 1698 740
rect 1710 734 1711 736
rect 1729 734 1744 740
rect 1753 738 1754 742
rect 1902 738 1908 744
rect 1960 738 1966 744
rect 1972 743 1974 745
rect 1752 734 1753 737
rect 1625 732 1626 734
rect 1686 732 1750 734
rect 1547 726 1549 727
rect 1550 726 1556 731
rect 1304 710 1308 711
rect 1309 710 1361 711
rect 1303 706 1367 710
rect 1298 704 1367 706
rect 1430 704 1433 711
rect 1157 698 1163 699
rect 1171 698 1209 699
rect 1151 695 1163 698
rect 1167 695 1215 698
rect 1151 693 1157 695
rect 1167 693 1205 695
rect 1209 693 1215 695
rect 1103 692 1215 693
rect 1103 691 1197 692
rect 706 688 709 689
rect 713 688 715 690
rect 116 669 126 688
rect 327 682 333 688
rect 385 682 391 688
rect 709 686 715 688
rect 332 680 345 682
rect 332 676 339 680
rect 379 676 385 682
rect 713 677 715 686
rect 815 681 838 690
rect 996 689 1018 691
rect 1103 689 1193 691
rect 815 679 885 681
rect 126 658 136 669
rect 128 656 142 658
rect 178 656 194 672
rect 332 668 333 676
rect 709 671 715 677
rect 767 678 838 679
rect 767 676 831 678
rect 885 676 894 679
rect 767 671 773 676
rect 332 656 344 668
rect 712 665 721 671
rect 761 665 767 671
rect 712 662 715 665
rect 796 662 815 676
rect 894 675 898 676
rect 898 672 900 675
rect 902 667 903 669
rect 712 658 714 662
rect 792 659 796 662
rect 903 660 918 667
rect 1002 662 1008 689
rect 1018 686 1053 689
rect 1103 686 1187 689
rect 1203 686 1209 692
rect 1298 690 1303 704
rect 1309 699 1327 704
rect 1309 698 1315 699
rect 1355 698 1361 704
rect 1428 699 1430 704
rect 1356 696 1357 698
rect 1426 695 1428 698
rect 1462 695 1470 712
rect 1490 709 1493 711
rect 1498 709 1502 726
rect 1549 717 1559 726
rect 1608 725 1614 731
rect 1621 725 1625 732
rect 1686 730 1744 732
rect 1745 730 1750 732
rect 1751 730 1752 732
rect 1686 728 1742 730
rect 1619 722 1620 724
rect 1559 709 1561 717
rect 1613 711 1619 721
rect 1493 708 1495 709
rect 1492 707 1496 708
rect 1492 703 1498 707
rect 1504 705 1505 707
rect 1504 703 1521 705
rect 1423 694 1426 695
rect 1419 692 1423 694
rect 1417 691 1419 692
rect 1053 684 1072 686
rect 1111 684 1175 686
rect 1072 683 1080 684
rect 1080 681 1101 683
rect 1111 681 1170 684
rect 1101 679 1170 681
rect 1294 679 1298 689
rect 1357 686 1359 690
rect 1413 689 1417 691
rect 1409 688 1413 689
rect 1459 688 1462 695
rect 1495 690 1498 703
rect 1501 699 1503 700
rect 1504 696 1528 699
rect 1504 691 1516 696
rect 1528 693 1542 696
rect 1561 693 1563 706
rect 1608 702 1613 711
rect 1692 696 1707 728
rect 1739 726 1742 728
rect 1745 726 1753 730
rect 1739 724 1741 726
rect 1740 700 1741 724
rect 1742 718 1753 726
rect 1742 714 1746 718
rect 1742 710 1745 714
rect 1748 712 1750 718
rect 2004 715 2006 745
rect 2008 742 2018 745
rect 2178 743 2180 749
rect 2188 743 2194 749
rect 2207 746 2230 770
rect 2234 743 2240 749
rect 2182 742 2188 743
rect 2010 738 2018 742
rect 2010 735 2028 738
rect 2018 731 2028 735
rect 2180 731 2188 742
rect 2193 738 2194 742
rect 2226 739 2232 742
rect 2191 731 2193 738
rect 2227 737 2232 739
rect 2240 737 2246 743
rect 1978 714 2006 715
rect 1973 713 2006 714
rect 2010 713 2018 725
rect 2028 721 2034 731
rect 2180 721 2191 731
rect 2172 720 2191 721
rect 2172 712 2181 720
rect 1747 710 1748 711
rect 1745 707 1749 710
rect 2007 709 2010 711
rect 1981 708 1984 709
rect 1744 702 1749 707
rect 1969 706 1979 708
rect 1960 704 1969 706
rect 1739 696 1741 699
rect 1542 692 1608 693
rect 1548 691 1608 692
rect 1382 686 1409 688
rect 1458 686 1459 688
rect 1357 684 1389 686
rect 1347 683 1389 684
rect 1320 681 1389 683
rect 1302 679 1389 681
rect 1455 679 1458 684
rect 1111 678 1170 679
rect 1114 677 1149 678
rect 1275 677 1389 679
rect 1114 676 1146 677
rect 1148 676 1149 677
rect 1115 674 1127 676
rect 1129 675 1148 676
rect 1253 675 1275 677
rect 1281 676 1389 677
rect 1294 675 1298 676
rect 1129 671 1156 675
rect 1205 671 1253 675
rect 1129 670 1167 671
rect 1194 670 1237 671
rect 1129 664 1237 670
rect 1131 662 1141 664
rect 1294 662 1295 675
rect 1359 672 1361 675
rect 1452 673 1455 679
rect 1008 660 1009 662
rect 790 658 792 659
rect 492 656 494 657
rect 712 656 713 658
rect 788 656 790 658
rect 144 640 160 656
rect 162 640 178 656
rect 345 653 347 656
rect 485 653 491 656
rect 714 653 717 656
rect 784 653 788 656
rect 347 651 349 653
rect 484 652 485 653
rect 782 652 784 653
rect 918 652 1030 660
rect 1122 658 1131 662
rect 1359 659 1362 672
rect 1491 666 1495 689
rect 1554 685 1608 691
rect 1692 688 1744 696
rect 1745 692 1749 702
rect 1902 693 1908 698
rect 1960 693 1966 698
rect 1902 692 1966 693
rect 1749 688 1751 690
rect 1550 679 1614 685
rect 1686 682 1751 688
rect 1908 686 1914 692
rect 1954 686 1960 692
rect 1972 690 1973 706
rect 1994 701 2006 709
rect 2185 707 2191 720
rect 2228 717 2232 737
rect 2184 706 2185 707
rect 2180 697 2184 706
rect 2232 697 2234 717
rect 2995 703 3017 722
rect 2966 697 2989 698
rect 2994 697 3017 703
rect 2180 693 2188 697
rect 2240 693 2246 697
rect 2180 691 2246 693
rect 2180 690 2184 691
rect 1973 686 1975 690
rect 1554 673 1562 679
rect 1602 673 1608 679
rect 1692 676 1698 682
rect 1738 676 1744 682
rect 1554 666 1561 673
rect 1694 672 1697 676
rect 1118 656 1122 658
rect 1295 656 1296 658
rect 1360 657 1362 659
rect 1358 656 1362 657
rect 1113 653 1118 656
rect 1296 653 1299 656
rect 1357 653 1358 656
rect 1392 654 1422 663
rect 1426 654 1439 660
rect 1491 659 1493 666
rect 1554 665 1562 666
rect 1108 652 1109 653
rect 1356 652 1357 653
rect 1389 652 1426 654
rect 1493 653 1495 659
rect 1551 656 1562 665
rect 1688 660 1697 672
rect 1750 672 1751 682
rect 1688 656 1694 660
rect 1750 656 1754 672
rect 1966 660 1975 686
rect 2174 674 2180 690
rect 2188 685 2194 691
rect 2234 685 2240 691
rect 2234 674 2237 685
rect 1550 653 1551 655
rect 1693 654 1694 656
rect 482 651 484 652
rect 349 649 425 651
rect 477 649 482 651
rect 717 649 721 652
rect 780 650 782 652
rect 770 649 780 650
rect 432 648 476 649
rect 728 640 744 649
rect 745 648 746 649
rect 1010 647 1012 651
rect 1030 647 1142 652
rect 1024 644 1142 647
rect 1240 644 1389 652
rect 1024 640 1040 644
rect 1142 641 1153 644
rect 1193 641 1240 644
rect 1153 640 1193 641
rect 1330 640 1346 644
rect 1392 636 1422 652
rect 1530 640 1546 653
rect 1693 644 1703 654
rect 1966 652 1979 660
rect 2034 656 2050 672
rect 2172 665 2181 674
rect 2234 667 2246 674
rect 2237 665 2246 667
rect 2174 656 2175 665
rect 2181 656 2190 665
rect 2228 656 2242 665
rect 2001 652 2034 656
rect 2234 652 2237 656
rect 1981 651 2000 652
rect 1749 645 1750 651
rect 1704 640 1720 644
rect 1722 640 1738 644
rect 2018 640 2034 652
rect 2175 645 2185 652
rect 2229 646 2234 652
rect 2223 645 2229 646
rect 2185 644 2226 645
rect 2210 640 2226 644
rect 1723 639 1724 640
rect 2939 623 2966 629
rect 2967 623 2994 624
rect 3510 481 3511 487
rect 3476 441 3511 475
rect 3522 463 3523 475
rect 3522 441 3523 453
rect 2719 429 2720 440
rect 2909 429 2910 440
rect 2995 429 2996 440
rect 3268 429 3269 440
rect 3465 429 3466 440
rect 3499 429 3511 435
rect 2730 389 2731 429
rect 2920 389 2921 429
rect 3006 389 3007 429
rect 3279 389 3280 429
rect 3476 389 3477 429
<< nwell >>
rect 3473 1778 3519 1779
rect 0 1120 3586 1778
rect 0 1116 606 1120
rect 0 1115 489 1116
rect 0 850 112 1115
rect 2394 1086 2620 1120
rect 2396 850 2610 1086
rect 2398 744 2610 850
rect 2631 800 2701 870
rect 3392 772 3422 807
rect 3541 744 3586 1120
<< ndiff >>
rect 3477 441 3511 475
<< locali >>
rect 2 2202 3587 2522
rect 1 1116 3586 1436
rect 2394 1086 2620 1116
rect 3550 1086 3586 1116
rect 444 886 484 922
rect 443 879 445 886
rect 442 875 444 879
rect 438 870 442 875
rect 437 869 438 870
rect 432 868 437 869
rect 471 868 484 886
rect 418 864 484 868
rect 415 862 484 864
rect 409 857 415 862
rect 408 856 409 857
rect 398 849 408 856
rect 418 849 484 862
rect 756 853 814 858
rect 756 852 818 853
rect 812 849 818 852
rect 381 842 484 849
rect 381 799 475 842
rect 514 833 587 838
rect 517 815 587 833
rect 817 813 818 832
rect 816 805 818 813
rect 530 799 618 805
rect 514 795 618 799
rect 530 783 618 795
rect 756 792 818 805
rect 75 320 2457 595
rect 1 0 3586 320
<< viali >>
rect 3477 1751 3511 1785
rect 3478 1491 3512 1525
rect 3477 997 3511 1031
rect 3477 441 3511 475
<< metal1 >>
rect 2 2202 3587 2522
rect 1815 1784 1849 2202
rect 1947 1963 2022 1972
rect 1947 1907 1957 1963
rect 2013 1907 2022 1963
rect 2955 1938 3239 1945
rect 2967 1932 3239 1938
rect 1947 1898 2022 1907
rect 2921 1911 3239 1932
rect 2921 1898 2967 1911
rect 3000 1876 3065 1883
rect 3000 1858 3007 1876
rect 2066 1824 3007 1858
rect 3059 1824 3065 1876
rect 3000 1818 3065 1824
rect 1815 1750 1886 1784
rect 2840 1738 2846 1796
rect 2898 1738 2904 1796
rect 2840 1732 2904 1738
rect 2629 1719 2699 1725
rect 2629 1710 2635 1719
rect 1744 1676 2635 1710
rect 2629 1661 2635 1676
rect 2693 1661 2699 1719
rect 3205 1675 3239 1911
rect 3314 1752 3437 1784
rect 3314 1751 3346 1752
rect 3404 1717 3437 1752
rect 3404 1716 3438 1717
rect 3406 1676 3438 1716
rect 2629 1655 2699 1661
rect 3458 1537 3533 1546
rect 3458 1479 3466 1537
rect 3524 1479 3533 1537
rect 3458 1470 3533 1479
rect 1 1116 3586 1436
rect 2394 1086 2620 1116
rect 3550 1086 3586 1116
rect 3456 1044 3532 1053
rect 2516 1009 2586 1015
rect 2516 951 2522 1009
rect 2580 951 2586 1009
rect 3456 986 3465 1044
rect 3523 986 3532 1044
rect 3456 977 3532 986
rect 2516 945 2586 951
rect 446 884 491 926
rect 506 833 517 837
rect 550 835 552 837
rect 486 831 517 833
rect 452 830 517 831
rect 452 829 490 830
rect 415 827 453 829
rect 378 825 416 827
rect 354 823 378 825
rect 288 822 354 823
rect 288 785 340 822
rect 462 804 535 807
rect 419 803 552 804
rect 401 799 564 803
rect 357 788 564 799
rect 750 788 794 831
rect 344 787 564 788
rect 342 785 564 787
rect 288 783 344 785
rect 288 782 342 783
rect 288 779 340 782
rect 401 775 564 785
rect 2534 699 2568 945
rect 2631 864 2701 870
rect 2631 806 2637 864
rect 2695 806 2701 864
rect 3206 819 3240 846
rect 3206 812 3241 819
rect 3207 809 3241 812
rect 2631 800 2701 806
rect 3206 806 3241 809
rect 2840 790 2904 796
rect 2840 772 2846 790
rect 2826 738 2846 772
rect 2898 738 2904 790
rect 2840 732 2904 738
rect 2995 716 3065 722
rect 2534 698 2858 699
rect 2534 664 2989 698
rect 2995 658 3001 716
rect 3059 658 3065 716
rect 2995 652 3065 658
rect 3206 624 3239 806
rect 3384 805 3449 852
rect 3384 772 3422 805
rect 3313 738 3422 772
rect 2921 623 2955 624
rect 2967 623 3239 624
rect 75 563 2457 595
rect 2921 590 3239 623
rect 75 510 476 563
rect 75 454 224 510
rect 280 506 476 510
rect 532 516 2457 563
rect 532 506 618 516
rect 280 460 618 506
rect 674 460 905 516
rect 961 460 2457 516
rect 2513 552 2588 561
rect 2513 496 2523 552
rect 2579 496 2588 552
rect 2513 487 2588 496
rect 280 454 2457 460
rect 75 320 2457 454
rect 1 0 3586 320
<< via1 >>
rect 1957 1907 2013 1963
rect 3007 1824 3059 1876
rect 2846 1738 2898 1796
rect 2635 1661 2693 1719
rect 3466 1525 3524 1537
rect 3466 1491 3478 1525
rect 3478 1491 3512 1525
rect 3512 1491 3524 1525
rect 3466 1479 3524 1491
rect 2522 951 2580 1009
rect 3465 1031 3523 1044
rect 3465 997 3477 1031
rect 3477 997 3511 1031
rect 3511 997 3523 1031
rect 3465 986 3523 997
rect 2637 806 2695 864
rect 2846 738 2898 790
rect 3001 658 3059 716
rect 476 506 532 563
rect 2523 496 2579 552
<< metal2 >>
rect 1947 1963 2022 1972
rect 1947 1907 1957 1963
rect 2013 1907 2022 1963
rect 1947 1898 2022 1907
rect 3000 1876 3065 1883
rect 3000 1870 3007 1876
rect 2777 1836 3007 1870
rect 2629 1719 2699 1725
rect 2629 1661 2635 1719
rect 2693 1661 2699 1719
rect 2629 1655 2699 1661
rect 1394 1131 2568 1165
rect 1394 1020 1432 1131
rect 1797 1022 1831 1045
rect 2534 1015 2568 1131
rect 2516 1009 2586 1015
rect 2516 951 2522 1009
rect 2580 951 2586 1009
rect 2516 945 2586 951
rect 2534 944 2568 945
rect 468 833 495 886
rect 514 870 518 883
rect 2644 870 2679 1655
rect 517 867 519 870
rect 519 851 524 867
rect 2631 864 2701 870
rect 524 847 529 851
rect 529 845 544 847
rect 543 841 549 845
rect 543 840 553 841
rect 546 833 553 840
rect 462 777 471 833
rect 527 825 560 833
rect 527 790 739 825
rect 2631 806 2637 864
rect 2695 806 2701 864
rect 2631 800 2701 806
rect 527 782 744 790
rect 527 777 560 782
rect 489 569 523 777
rect 2777 772 2809 1836
rect 3000 1824 3007 1836
rect 3059 1824 3065 1876
rect 3000 1818 3065 1824
rect 2840 1738 2846 1796
rect 2898 1738 2904 1796
rect 2840 1732 2904 1738
rect 2846 1696 2880 1732
rect 2846 1661 2881 1696
rect 2846 1626 3041 1661
rect 2840 790 2904 796
rect 2840 772 2846 790
rect 2777 738 2846 772
rect 2898 738 2904 790
rect 2840 732 2904 738
rect 3006 722 3041 1626
rect 3458 1537 3533 1546
rect 3458 1479 3466 1537
rect 3524 1479 3533 1537
rect 3458 1470 3533 1479
rect 3456 1044 3532 1053
rect 3456 986 3465 1044
rect 3523 986 3532 1044
rect 3456 977 3532 986
rect 2995 716 3065 722
rect 2995 658 3001 716
rect 3059 658 3065 716
rect 2995 652 3065 658
rect 470 563 539 569
rect 214 510 289 519
rect 214 454 224 510
rect 280 454 289 510
rect 470 506 476 563
rect 532 506 539 563
rect 2513 552 2588 561
rect 470 500 539 506
rect 608 516 683 525
rect 214 445 289 454
rect 608 459 618 516
rect 674 509 683 516
rect 895 516 970 525
rect 895 509 905 516
rect 674 475 905 509
rect 674 459 683 475
rect 608 451 683 459
rect 895 460 905 475
rect 961 509 970 516
rect 2513 509 2523 552
rect 961 496 2523 509
rect 2579 496 2588 552
rect 961 487 2588 496
rect 961 475 2574 487
rect 961 460 970 475
rect 895 451 970 460
<< via2 >>
rect 1957 1907 2013 1963
rect 471 777 527 833
rect 3466 1479 3524 1537
rect 3465 986 3523 1044
rect 224 454 280 510
rect 618 459 674 516
rect 905 460 961 516
rect 2523 496 2579 552
<< metal3 >>
rect 1947 1963 2022 1972
rect 1947 1907 1957 1963
rect 2013 1907 2022 1963
rect 1947 1898 2022 1907
rect 1954 1534 2016 1898
rect 3458 1537 3533 2522
rect 1954 1472 2573 1534
rect 223 519 283 834
rect 401 833 547 838
rect 334 779 336 782
rect 401 777 471 833
rect 527 777 547 833
rect 401 772 547 777
rect 617 525 677 921
rect 904 525 964 1041
rect 2511 561 2573 1472
rect 3458 1479 3466 1537
rect 3524 1479 3533 1537
rect 3458 1470 3533 1479
rect 3456 1044 3532 1053
rect 3456 986 3465 1044
rect 3523 986 3532 1044
rect 2513 552 2588 561
rect 214 513 289 519
rect 608 516 683 525
rect 608 513 618 516
rect 214 510 618 513
rect 214 454 224 510
rect 280 459 618 510
rect 674 459 683 516
rect 280 454 683 459
rect 214 453 683 454
rect 214 445 289 453
rect 608 451 683 453
rect 895 516 970 525
rect 895 460 905 516
rect 961 460 970 516
rect 2513 496 2523 552
rect 2579 496 2588 552
rect 2513 487 2588 496
rect 2513 484 2575 487
rect 895 451 970 460
rect 3456 0 3532 986
use scs130hd_mpr2at_8  scs130hd_mpr2at_8_0
timestamp 1696005323
transform 1 0 78 0 1 588
box -48 -47 2440 593
use sky130_osu_sc_12T_hs__fill_2  sky130_osu_sc_12T_hs__fill_2_0
timestamp 1604095901
transform 1 0 2047 0 -1 2263
box -7 0 161 1341
use sky130_osu_sc_12T_hs__fill_8  sky130_osu_sc_12T_hs__fill_8_0
timestamp 1604095905
transform 1 0 2218 0 -1 2263
box -9 0 179 897
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1706264206
transform 1 0 3159 0 1 259
box -10 0 198 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1706264206
transform 1 0 3356 0 1 259
box -10 0 198 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1706264206
transform 1 0 3357 0 -1 2263
box -10 0 198 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1706264206
transform 1 0 3159 0 -1 2263
box -10 0 198 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1698882961
transform 1 0 2610 0 1 259
box -8 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1698882961
transform 1 0 1658 0 -1 2263
box -8 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1698882961
transform 1 0 2610 0 -1 2263
box -8 0 552 902
<< labels >>
rlabel metal1 47 1157 47 1157 1 vccd1
port 6 n
rlabel metal1 47 287 47 287 1 vssd1
port 5 n
rlabel metal2 2664 837 2664 837 1 sel
port 8 n
rlabel metal1 50 2230 50 2230 1 vssd1
port 5 n
rlabel metal1 2066 1824 2089 1858 1 in
port 12 n
rlabel viali 3477 1751 3511 1785 1 Y0
port 10 n
rlabel viali 3477 441 3511 475 1 Y1
port 11 n
<< end >>
