* NGSPICE file created from sky130_osu_sc_12T_hs__fill_32.ext - technology: sky130A


* Top level circuit sky130_osu_sc_12T_hs__fill_32

.end

