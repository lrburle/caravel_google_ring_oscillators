magic
tech sky130A
magscale 1 2
timestamp 1713287902
<< error_p >>
rect 0 827 44 888
rect 50 485 161 897
rect 0 0 44 61
<< nwell >>
rect -7 485 50 897
<< locali >>
rect 0 827 44 888
rect 0 0 44 61
<< metal1 >>
rect 0 827 44 888
rect 0 0 44 61
<< labels >>
rlabel metal1 22 856 22 856 1 vccd1
rlabel metal1 23 28 23 28 1 vssd1
<< end >>
